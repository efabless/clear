magic
tech sky130A
magscale 1 2
timestamp 1656406099
<< viali >>
rect 1869 20553 1903 20587
rect 3893 20553 3927 20587
rect 10333 20553 10367 20587
rect 11897 20553 11931 20587
rect 12265 20553 12299 20587
rect 12633 20553 12667 20587
rect 12909 20553 12943 20587
rect 13369 20553 13403 20587
rect 13645 20553 13679 20587
rect 14197 20553 14231 20587
rect 14933 20553 14967 20587
rect 15301 20553 15335 20587
rect 15669 20553 15703 20587
rect 16037 20553 16071 20587
rect 17141 20553 17175 20587
rect 18337 20553 18371 20587
rect 19073 20553 19107 20587
rect 19533 20553 19567 20587
rect 19993 20553 20027 20587
rect 21465 20553 21499 20587
rect 2881 20485 2915 20519
rect 3617 20485 3651 20519
rect 7665 20485 7699 20519
rect 9045 20485 9079 20519
rect 1685 20417 1719 20451
rect 2053 20417 2087 20451
rect 2329 20417 2363 20451
rect 2697 20417 2731 20451
rect 3065 20417 3099 20451
rect 3433 20417 3467 20451
rect 4252 20417 4286 20451
rect 5825 20417 5859 20451
rect 7205 20417 7239 20451
rect 7481 20417 7515 20451
rect 8769 20417 8803 20451
rect 9137 20417 9171 20451
rect 10149 20417 10183 20451
rect 10517 20417 10551 20451
rect 11713 20417 11747 20451
rect 12081 20417 12115 20451
rect 12449 20417 12483 20451
rect 13093 20417 13127 20451
rect 13185 20417 13219 20451
rect 13829 20417 13863 20451
rect 14381 20417 14415 20451
rect 14749 20417 14783 20451
rect 15117 20417 15151 20451
rect 15485 20417 15519 20451
rect 15853 20417 15887 20451
rect 16221 20417 16255 20451
rect 16497 20417 16531 20451
rect 16681 20417 16715 20451
rect 17325 20417 17359 20451
rect 17417 20417 17451 20451
rect 17785 20417 17819 20451
rect 18153 20417 18187 20451
rect 18521 20417 18555 20451
rect 18889 20417 18923 20451
rect 19349 20417 19383 20451
rect 19717 20417 19751 20451
rect 19809 20417 19843 20451
rect 20177 20417 20211 20451
rect 20545 20417 20579 20451
rect 20913 20417 20947 20451
rect 21281 20417 21315 20451
rect 3985 20349 4019 20383
rect 5917 20349 5951 20383
rect 6009 20349 6043 20383
rect 6929 20349 6963 20383
rect 8493 20349 8527 20383
rect 9413 20349 9447 20383
rect 10793 20349 10827 20383
rect 3249 20281 3283 20315
rect 5457 20281 5491 20315
rect 11529 20281 11563 20315
rect 14565 20281 14599 20315
rect 16865 20281 16899 20315
rect 17601 20281 17635 20315
rect 18705 20281 18739 20315
rect 20729 20281 20763 20315
rect 1501 20213 1535 20247
rect 2421 20213 2455 20247
rect 5365 20213 5399 20247
rect 7297 20213 7331 20247
rect 7757 20213 7791 20247
rect 16313 20213 16347 20247
rect 17969 20213 18003 20247
rect 20361 20213 20395 20247
rect 21097 20213 21131 20247
rect 2237 20009 2271 20043
rect 2605 20009 2639 20043
rect 6377 20009 6411 20043
rect 11529 20009 11563 20043
rect 12265 20009 12299 20043
rect 15485 20009 15519 20043
rect 16865 20009 16899 20043
rect 17141 20009 17175 20043
rect 17601 20009 17635 20043
rect 17693 20009 17727 20043
rect 18429 20009 18463 20043
rect 15209 19941 15243 19975
rect 16589 19941 16623 19975
rect 17969 19941 18003 19975
rect 18889 19941 18923 19975
rect 3065 19873 3099 19907
rect 8953 19873 8987 19907
rect 13737 19873 13771 19907
rect 19625 19873 19659 19907
rect 20269 19873 20303 19907
rect 1685 19805 1719 19839
rect 2053 19805 2087 19839
rect 2421 19805 2455 19839
rect 2789 19805 2823 19839
rect 3249 19805 3283 19839
rect 4353 19805 4387 19839
rect 4629 19805 4663 19839
rect 4721 19805 4755 19839
rect 4997 19805 5031 19839
rect 6837 19805 6871 19839
rect 7093 19805 7127 19839
rect 10517 19805 10551 19839
rect 10885 19805 10919 19839
rect 11345 19805 11379 19839
rect 12081 19805 12115 19839
rect 14197 19805 14231 19839
rect 14565 19805 14599 19839
rect 15117 19805 15151 19839
rect 15393 19821 15427 19855
rect 15669 19805 15703 19839
rect 15945 19805 15979 19839
rect 16221 19805 16255 19839
rect 16497 19805 16531 19839
rect 16773 19805 16807 19839
rect 17049 19805 17083 19839
rect 17325 19805 17359 19839
rect 17417 19805 17451 19839
rect 17877 19805 17911 19839
rect 18153 19805 18187 19839
rect 18613 19805 18647 19839
rect 19073 19805 19107 19839
rect 19349 19805 19383 19839
rect 20545 19805 20579 19839
rect 20729 19805 20763 19839
rect 21281 19805 21315 19839
rect 5242 19737 5276 19771
rect 6469 19737 6503 19771
rect 6653 19737 6687 19771
rect 8677 19737 8711 19771
rect 9198 19737 9232 19771
rect 11805 19737 11839 19771
rect 13470 19737 13504 19771
rect 21005 19737 21039 19771
rect 1501 19669 1535 19703
rect 1869 19669 1903 19703
rect 3157 19669 3191 19703
rect 3617 19669 3651 19703
rect 4905 19669 4939 19703
rect 8217 19669 8251 19703
rect 8309 19669 8343 19703
rect 8585 19669 8619 19703
rect 10333 19669 10367 19703
rect 11897 19669 11931 19703
rect 12357 19669 12391 19703
rect 13829 19669 13863 19703
rect 14933 19669 14967 19703
rect 15761 19669 15795 19703
rect 16037 19669 16071 19703
rect 16313 19669 16347 19703
rect 21465 19669 21499 19703
rect 1869 19465 1903 19499
rect 3433 19465 3467 19499
rect 4261 19465 4295 19499
rect 4721 19465 4755 19499
rect 6193 19465 6227 19499
rect 8493 19465 8527 19499
rect 8953 19465 8987 19499
rect 9321 19465 9355 19499
rect 9597 19465 9631 19499
rect 11345 19465 11379 19499
rect 13001 19465 13035 19499
rect 13829 19465 13863 19499
rect 15669 19465 15703 19499
rect 16129 19465 16163 19499
rect 16405 19465 16439 19499
rect 17969 19465 18003 19499
rect 18797 19465 18831 19499
rect 19073 19465 19107 19499
rect 19533 19465 19567 19499
rect 19809 19465 19843 19499
rect 20545 19465 20579 19499
rect 21465 19465 21499 19499
rect 2697 19397 2731 19431
rect 5080 19397 5114 19431
rect 6745 19397 6779 19431
rect 8033 19397 8067 19431
rect 10824 19397 10858 19431
rect 11774 19397 11808 19431
rect 14464 19397 14498 19431
rect 1685 19329 1719 19363
rect 2053 19329 2087 19363
rect 3525 19329 3559 19363
rect 4353 19329 4387 19363
rect 4813 19329 4847 19363
rect 7297 19329 7331 19363
rect 7389 19329 7423 19363
rect 8125 19329 8159 19363
rect 8861 19329 8895 19363
rect 9413 19329 9447 19363
rect 11069 19329 11103 19363
rect 11161 19329 11195 19363
rect 11529 19329 11563 19363
rect 13369 19329 13403 19363
rect 14013 19329 14047 19363
rect 15853 19329 15887 19363
rect 15945 19353 15979 19387
rect 16221 19329 16255 19363
rect 16865 19329 16899 19363
rect 16957 19329 16991 19363
rect 17785 19329 17819 19363
rect 18429 19329 18463 19363
rect 18705 19329 18739 19363
rect 18981 19329 19015 19363
rect 19257 19329 19291 19363
rect 19349 19329 19383 19363
rect 19625 19329 19659 19363
rect 19993 19329 20027 19363
rect 20361 19329 20395 19363
rect 20729 19329 20763 19363
rect 21005 19329 21039 19363
rect 21281 19329 21315 19363
rect 2513 19261 2547 19295
rect 2605 19261 2639 19295
rect 3341 19261 3375 19295
rect 4169 19261 4203 19295
rect 7573 19261 7607 19295
rect 7849 19261 7883 19295
rect 8769 19261 8803 19295
rect 13461 19261 13495 19295
rect 13553 19261 13587 19295
rect 14197 19261 14231 19295
rect 18061 19261 18095 19295
rect 16681 19193 16715 19227
rect 17141 19193 17175 19227
rect 17325 19193 17359 19227
rect 18245 19193 18279 19227
rect 20177 19193 20211 19227
rect 1501 19125 1535 19159
rect 2237 19125 2271 19159
rect 3065 19125 3099 19159
rect 3893 19125 3927 19159
rect 6469 19125 6503 19159
rect 6653 19125 6687 19159
rect 6929 19125 6963 19159
rect 9689 19125 9723 19159
rect 12909 19125 12943 19159
rect 15577 19125 15611 19159
rect 17417 19125 17451 19159
rect 17693 19125 17727 19159
rect 18521 19125 18555 19159
rect 3801 18921 3835 18955
rect 6469 18921 6503 18955
rect 7665 18921 7699 18955
rect 8493 18921 8527 18955
rect 8953 18921 8987 18955
rect 10977 18921 11011 18955
rect 11253 18921 11287 18955
rect 12081 18921 12115 18955
rect 13737 18921 13771 18955
rect 15485 18921 15519 18955
rect 15761 18921 15795 18955
rect 17969 18921 18003 18955
rect 18521 18921 18555 18955
rect 18797 18921 18831 18955
rect 20453 18921 20487 18955
rect 1869 18853 1903 18887
rect 5365 18853 5399 18887
rect 9781 18853 9815 18887
rect 15209 18853 15243 18887
rect 18245 18853 18279 18887
rect 20177 18853 20211 18887
rect 3341 18785 3375 18819
rect 3433 18785 3467 18819
rect 4261 18785 4295 18819
rect 4445 18785 4479 18819
rect 4721 18785 4755 18819
rect 6009 18785 6043 18819
rect 7113 18785 7147 18819
rect 7205 18785 7239 18819
rect 7941 18785 7975 18819
rect 9505 18785 9539 18819
rect 10333 18785 10367 18819
rect 11529 18785 11563 18819
rect 11621 18785 11655 18819
rect 12265 18785 12299 18819
rect 12449 18785 12483 18819
rect 13185 18785 13219 18819
rect 14381 18785 14415 18819
rect 1685 18717 1719 18751
rect 2053 18717 2087 18751
rect 2329 18717 2363 18751
rect 2789 18717 2823 18751
rect 6285 18717 6319 18751
rect 8585 18717 8619 18751
rect 10241 18717 10275 18751
rect 10609 18717 10643 18751
rect 10793 18717 10827 18751
rect 11069 18717 11103 18751
rect 14565 18717 14599 18751
rect 15025 18717 15059 18751
rect 15301 18717 15335 18751
rect 15577 18717 15611 18751
rect 16129 18717 16163 18751
rect 18061 18717 18095 18751
rect 18337 18717 18371 18751
rect 18613 18717 18647 18751
rect 18889 18717 18923 18751
rect 19625 18693 19659 18727
rect 19717 18717 19751 18751
rect 19993 18717 20027 18751
rect 20269 18717 20303 18751
rect 20637 18717 20671 18751
rect 21281 18717 21315 18751
rect 2421 18649 2455 18683
rect 6653 18649 6687 18683
rect 7297 18649 7331 18683
rect 13369 18649 13403 18683
rect 14473 18649 14507 18683
rect 15853 18649 15887 18683
rect 17785 18649 17819 18683
rect 20913 18649 20947 18683
rect 1501 18581 1535 18615
rect 2145 18581 2179 18615
rect 2605 18581 2639 18615
rect 2881 18581 2915 18615
rect 3249 18581 3283 18615
rect 4169 18581 4203 18615
rect 4905 18581 4939 18615
rect 4997 18581 5031 18615
rect 5457 18581 5491 18615
rect 5825 18581 5859 18615
rect 5917 18581 5951 18615
rect 6745 18581 6779 18615
rect 8033 18581 8067 18615
rect 8125 18581 8159 18615
rect 8769 18581 8803 18615
rect 9321 18581 9355 18615
rect 9413 18581 9447 18615
rect 10149 18581 10183 18615
rect 11713 18581 11747 18615
rect 12541 18581 12575 18615
rect 12909 18581 12943 18615
rect 13277 18581 13311 18615
rect 13829 18581 13863 18615
rect 14933 18581 14967 18615
rect 16221 18581 16255 18615
rect 16405 18581 16439 18615
rect 17233 18581 17267 18615
rect 19073 18581 19107 18615
rect 19257 18581 19291 18615
rect 19441 18581 19475 18615
rect 19901 18581 19935 18615
rect 21465 18581 21499 18615
rect 2513 18377 2547 18411
rect 3065 18377 3099 18411
rect 3157 18377 3191 18411
rect 3617 18377 3651 18411
rect 5733 18377 5767 18411
rect 6193 18377 6227 18411
rect 6377 18377 6411 18411
rect 7757 18377 7791 18411
rect 8125 18377 8159 18411
rect 8953 18377 8987 18411
rect 9321 18377 9355 18411
rect 10149 18377 10183 18411
rect 10609 18377 10643 18411
rect 10977 18377 11011 18411
rect 11253 18377 11287 18411
rect 11897 18377 11931 18411
rect 13553 18377 13587 18411
rect 14197 18377 14231 18411
rect 14657 18377 14691 18411
rect 15393 18377 15427 18411
rect 18889 18377 18923 18411
rect 19349 18377 19383 18411
rect 19809 18377 19843 18411
rect 20821 18377 20855 18411
rect 6837 18309 6871 18343
rect 7481 18309 7515 18343
rect 12265 18309 12299 18343
rect 14013 18309 14047 18343
rect 18797 18309 18831 18343
rect 1685 18241 1719 18275
rect 2053 18241 2087 18275
rect 2237 18241 2271 18275
rect 2697 18241 2731 18275
rect 4730 18241 4764 18275
rect 5273 18241 5307 18275
rect 5825 18241 5859 18275
rect 6745 18241 6779 18275
rect 9597 18241 9631 18275
rect 9873 18241 9907 18275
rect 10333 18241 10367 18275
rect 10425 18241 10459 18275
rect 10793 18241 10827 18275
rect 11069 18241 11103 18275
rect 13093 18241 13127 18275
rect 14749 18241 14783 18275
rect 19257 18241 19291 18275
rect 19533 18241 19567 18275
rect 19625 18241 19659 18275
rect 19901 18241 19935 18275
rect 20361 18241 20395 18275
rect 20637 18265 20671 18299
rect 20913 18241 20947 18275
rect 21281 18241 21315 18275
rect 2973 18173 3007 18207
rect 4997 18173 5031 18207
rect 5549 18173 5583 18207
rect 6929 18173 6963 18207
rect 8217 18173 8251 18207
rect 8309 18173 8343 18207
rect 8677 18173 8711 18207
rect 8861 18173 8895 18207
rect 12357 18173 12391 18207
rect 12541 18173 12575 18207
rect 13185 18173 13219 18207
rect 13277 18173 13311 18207
rect 14565 18173 14599 18207
rect 20269 18173 20303 18207
rect 1869 18105 1903 18139
rect 3525 18105 3559 18139
rect 7297 18105 7331 18139
rect 10057 18105 10091 18139
rect 11621 18105 11655 18139
rect 12725 18105 12759 18139
rect 15117 18105 15151 18139
rect 19073 18105 19107 18139
rect 20545 18105 20579 18139
rect 21097 18105 21131 18139
rect 1501 18037 1535 18071
rect 2421 18037 2455 18071
rect 5089 18037 5123 18071
rect 9689 18037 9723 18071
rect 11713 18037 11747 18071
rect 13829 18037 13863 18071
rect 15301 18037 15335 18071
rect 15577 18037 15611 18071
rect 20085 18037 20119 18071
rect 21465 18037 21499 18071
rect 2421 17833 2455 17867
rect 2789 17833 2823 17867
rect 6469 17833 6503 17867
rect 8033 17833 8067 17867
rect 8953 17833 8987 17867
rect 9965 17833 9999 17867
rect 13001 17833 13035 17867
rect 14933 17833 14967 17867
rect 16957 17833 16991 17867
rect 19441 17833 19475 17867
rect 21005 17833 21039 17867
rect 3617 17765 3651 17799
rect 6193 17765 6227 17799
rect 7481 17765 7515 17799
rect 11529 17765 11563 17799
rect 19901 17765 19935 17799
rect 20361 17765 20395 17799
rect 20637 17765 20671 17799
rect 21465 17765 21499 17799
rect 3065 17697 3099 17731
rect 5917 17697 5951 17731
rect 6929 17697 6963 17731
rect 8585 17697 8619 17731
rect 9505 17697 9539 17731
rect 12357 17697 12391 17731
rect 13277 17697 13311 17731
rect 14289 17697 14323 17731
rect 16497 17697 16531 17731
rect 19625 17697 19659 17731
rect 1685 17629 1719 17663
rect 2053 17629 2087 17663
rect 2329 17629 2363 17663
rect 2605 17629 2639 17663
rect 3985 17629 4019 17663
rect 4445 17629 4479 17663
rect 6009 17629 6043 17663
rect 6377 17629 6411 17663
rect 10057 17629 10091 17663
rect 11713 17629 11747 17663
rect 12541 17629 12575 17663
rect 13093 17629 13127 17663
rect 13553 17629 13587 17663
rect 16230 17629 16264 17663
rect 20085 17629 20119 17663
rect 20177 17629 20211 17663
rect 20453 17629 20487 17663
rect 20729 17629 20763 17663
rect 21189 17629 21223 17663
rect 21281 17629 21315 17663
rect 5650 17561 5684 17595
rect 7113 17561 7147 17595
rect 7941 17561 7975 17595
rect 8401 17561 8435 17595
rect 9413 17561 9447 17595
rect 10324 17561 10358 17595
rect 11805 17561 11839 17595
rect 13829 17561 13863 17595
rect 14473 17561 14507 17595
rect 16773 17561 16807 17595
rect 19717 17561 19751 17595
rect 1501 17493 1535 17527
rect 1869 17493 1903 17527
rect 2145 17493 2179 17527
rect 3157 17493 3191 17527
rect 3249 17493 3283 17527
rect 3801 17493 3835 17527
rect 4169 17493 4203 17527
rect 4261 17493 4295 17527
rect 4537 17493 4571 17527
rect 7021 17493 7055 17527
rect 7573 17493 7607 17527
rect 8493 17493 8527 17527
rect 9321 17493 9355 17527
rect 11437 17493 11471 17527
rect 12173 17493 12207 17527
rect 12633 17493 12667 17527
rect 13737 17493 13771 17527
rect 14565 17493 14599 17527
rect 15117 17493 15151 17527
rect 20913 17493 20947 17527
rect 4629 17289 4663 17323
rect 5089 17289 5123 17323
rect 5457 17289 5491 17323
rect 5825 17289 5859 17323
rect 5917 17289 5951 17323
rect 6377 17289 6411 17323
rect 8033 17289 8067 17323
rect 8861 17289 8895 17323
rect 14933 17289 14967 17323
rect 16129 17289 16163 17323
rect 16681 17289 16715 17323
rect 17049 17289 17083 17323
rect 19809 17289 19843 17323
rect 20269 17289 20303 17323
rect 21005 17289 21039 17323
rect 3402 17221 3436 17255
rect 11796 17221 11830 17255
rect 20729 17221 20763 17255
rect 1593 17153 1627 17187
rect 2809 17153 2843 17187
rect 4997 17153 5031 17187
rect 6561 17153 6595 17187
rect 7021 17153 7055 17187
rect 7113 17153 7147 17187
rect 7665 17153 7699 17187
rect 7757 17153 7791 17187
rect 8401 17153 8435 17187
rect 10158 17153 10192 17187
rect 10609 17153 10643 17187
rect 10977 17153 11011 17187
rect 11529 17153 11563 17187
rect 13461 17153 13495 17187
rect 13728 17153 13762 17187
rect 15301 17153 15335 17187
rect 19993 17153 20027 17187
rect 20821 17153 20855 17187
rect 21281 17153 21315 17187
rect 3065 17085 3099 17119
rect 3157 17085 3191 17119
rect 5273 17085 5307 17119
rect 6101 17085 6135 17119
rect 7297 17085 7331 17119
rect 8493 17085 8527 17119
rect 8677 17085 8711 17119
rect 10425 17085 10459 17119
rect 15393 17085 15427 17119
rect 15577 17085 15611 17119
rect 16221 17085 16255 17119
rect 16313 17085 16347 17119
rect 17141 17085 17175 17119
rect 17233 17085 17267 17119
rect 7481 17017 7515 17051
rect 9045 17017 9079 17051
rect 13001 17017 13035 17051
rect 14841 17017 14875 17051
rect 15761 17017 15795 17051
rect 20177 17017 20211 17051
rect 21189 17017 21223 17051
rect 1409 16949 1443 16983
rect 1685 16949 1719 16983
rect 4537 16949 4571 16983
rect 6653 16949 6687 16983
rect 7941 16949 7975 16983
rect 12909 16949 12943 16983
rect 13185 16949 13219 16983
rect 17509 16949 17543 16983
rect 20453 16949 20487 16983
rect 21465 16949 21499 16983
rect 3801 16745 3835 16779
rect 4813 16745 4847 16779
rect 6561 16745 6595 16779
rect 7757 16745 7791 16779
rect 9413 16745 9447 16779
rect 12357 16745 12391 16779
rect 13461 16745 13495 16779
rect 14105 16745 14139 16779
rect 16405 16745 16439 16779
rect 17233 16745 17267 16779
rect 20545 16745 20579 16779
rect 20821 16745 20855 16779
rect 3617 16677 3651 16711
rect 21097 16677 21131 16711
rect 2237 16609 2271 16643
rect 4353 16609 4387 16643
rect 5365 16609 5399 16643
rect 5457 16609 5491 16643
rect 6285 16609 6319 16643
rect 7021 16609 7055 16643
rect 7205 16609 7239 16643
rect 7941 16609 7975 16643
rect 8217 16609 8251 16643
rect 8309 16609 8343 16643
rect 9965 16609 9999 16643
rect 10149 16609 10183 16643
rect 10701 16609 10735 16643
rect 11345 16609 11379 16643
rect 11713 16609 11747 16643
rect 11805 16609 11839 16643
rect 12909 16609 12943 16643
rect 13645 16609 13679 16643
rect 15485 16609 15519 16643
rect 16221 16609 16255 16643
rect 17049 16609 17083 16643
rect 17693 16609 17727 16643
rect 17785 16609 17819 16643
rect 18153 16609 18187 16643
rect 19901 16609 19935 16643
rect 1409 16541 1443 16575
rect 2053 16541 2087 16575
rect 2504 16541 2538 16575
rect 4261 16541 4295 16575
rect 4629 16541 4663 16575
rect 6101 16541 6135 16575
rect 7573 16541 7607 16575
rect 9137 16541 9171 16575
rect 10793 16541 10827 16575
rect 12817 16541 12851 16575
rect 13369 16541 13403 16575
rect 15218 16541 15252 16575
rect 16865 16541 16899 16575
rect 20177 16541 20211 16575
rect 20361 16541 20395 16575
rect 20637 16541 20671 16575
rect 20913 16541 20947 16575
rect 21281 16541 21315 16575
rect 5273 16473 5307 16507
rect 8401 16473 8435 16507
rect 10885 16473 10919 16507
rect 16773 16473 16807 16507
rect 1593 16405 1627 16439
rect 1869 16405 1903 16439
rect 4169 16405 4203 16439
rect 4905 16405 4939 16439
rect 5733 16405 5767 16439
rect 6193 16405 6227 16439
rect 6929 16405 6963 16439
rect 7389 16405 7423 16439
rect 8769 16405 8803 16439
rect 8953 16405 8987 16439
rect 9505 16405 9539 16439
rect 9873 16405 9907 16439
rect 10425 16405 10459 16439
rect 11253 16405 11287 16439
rect 11897 16405 11931 16439
rect 12265 16405 12299 16439
rect 12725 16405 12759 16439
rect 13185 16405 13219 16439
rect 15577 16405 15611 16439
rect 15945 16405 15979 16439
rect 16037 16405 16071 16439
rect 17601 16405 17635 16439
rect 20085 16405 20119 16439
rect 21465 16405 21499 16439
rect 1869 16201 1903 16235
rect 2513 16201 2547 16235
rect 2973 16201 3007 16235
rect 5733 16201 5767 16235
rect 6101 16201 6135 16235
rect 8033 16201 8067 16235
rect 9505 16201 9539 16235
rect 10425 16201 10459 16235
rect 10885 16201 10919 16235
rect 12173 16201 12207 16235
rect 12449 16201 12483 16235
rect 15485 16201 15519 16235
rect 19625 16201 19659 16235
rect 20177 16201 20211 16235
rect 20729 16201 20763 16235
rect 21005 16201 21039 16235
rect 4620 16133 4654 16167
rect 6920 16133 6954 16167
rect 8370 16133 8404 16167
rect 10057 16133 10091 16167
rect 11989 16133 12023 16167
rect 13584 16133 13618 16167
rect 14197 16133 14231 16167
rect 16405 16133 16439 16167
rect 19533 16133 19567 16167
rect 1685 16065 1719 16099
rect 2053 16065 2087 16099
rect 3341 16065 3375 16099
rect 3801 16065 3835 16099
rect 4261 16065 4295 16099
rect 4353 16065 4387 16099
rect 5825 16065 5859 16099
rect 8125 16065 8159 16099
rect 11713 16065 11747 16099
rect 13829 16065 13863 16099
rect 14565 16065 14599 16099
rect 15117 16065 15151 16099
rect 17417 16065 17451 16099
rect 18797 16065 18831 16099
rect 19993 16065 20027 16099
rect 20269 16065 20303 16099
rect 20545 16065 20579 16099
rect 20821 16065 20855 16099
rect 21281 16065 21315 16099
rect 2237 15997 2271 16031
rect 2421 15997 2455 16031
rect 3433 15997 3467 16031
rect 3617 15997 3651 16031
rect 6377 15997 6411 16031
rect 6653 15997 6687 16031
rect 9781 15997 9815 16031
rect 9965 15997 9999 16031
rect 10977 15997 11011 16031
rect 11069 15997 11103 16031
rect 11529 15997 11563 16031
rect 14933 15997 14967 16031
rect 15025 15997 15059 16031
rect 17141 15997 17175 16031
rect 19073 15997 19107 16031
rect 19349 15997 19383 16031
rect 2881 15929 2915 15963
rect 4077 15929 4111 15963
rect 20453 15929 20487 15963
rect 1501 15861 1535 15895
rect 6009 15861 6043 15895
rect 10517 15861 10551 15895
rect 12265 15861 12299 15895
rect 16221 15861 16255 15895
rect 18981 15861 19015 15895
rect 19809 15861 19843 15895
rect 21097 15861 21131 15895
rect 21465 15861 21499 15895
rect 2145 15657 2179 15691
rect 3617 15657 3651 15691
rect 4353 15657 4387 15691
rect 5641 15657 5675 15691
rect 6745 15657 6779 15691
rect 6929 15657 6963 15691
rect 8677 15657 8711 15691
rect 9965 15657 9999 15691
rect 10793 15657 10827 15691
rect 13093 15657 13127 15691
rect 20453 15657 20487 15691
rect 2053 15589 2087 15623
rect 2421 15589 2455 15623
rect 3801 15589 3835 15623
rect 5549 15589 5583 15623
rect 8585 15589 8619 15623
rect 14473 15589 14507 15623
rect 16037 15589 16071 15623
rect 18153 15589 18187 15623
rect 18613 15589 18647 15623
rect 19533 15589 19567 15623
rect 19901 15589 19935 15623
rect 2973 15521 3007 15555
rect 5089 15521 5123 15555
rect 6193 15521 6227 15555
rect 7481 15521 7515 15555
rect 7849 15521 7883 15555
rect 8953 15521 8987 15555
rect 9321 15521 9355 15555
rect 10517 15521 10551 15555
rect 11345 15521 11379 15555
rect 12541 15521 12575 15555
rect 15485 15521 15519 15555
rect 16221 15521 16255 15555
rect 17141 15521 17175 15555
rect 17233 15521 17267 15555
rect 21097 15521 21131 15555
rect 1685 15453 1719 15487
rect 1869 15453 1903 15487
rect 2329 15453 2363 15487
rect 2605 15453 2639 15487
rect 2789 15453 2823 15487
rect 3985 15469 4019 15503
rect 4261 15453 4295 15487
rect 4997 15453 5031 15487
rect 5365 15453 5399 15487
rect 6101 15453 6135 15487
rect 7389 15453 7423 15487
rect 8309 15453 8343 15487
rect 9413 15453 9447 15487
rect 10425 15453 10459 15487
rect 11161 15453 11195 15487
rect 12173 15453 12207 15487
rect 16405 15453 16439 15487
rect 17969 15453 18003 15487
rect 18981 15453 19015 15487
rect 19717 15453 19751 15487
rect 20269 15453 20303 15487
rect 20545 15453 20579 15487
rect 20821 15453 20855 15487
rect 21281 15453 21315 15487
rect 3249 15385 3283 15419
rect 6009 15385 6043 15419
rect 7297 15385 7331 15419
rect 8033 15385 8067 15419
rect 10333 15385 10367 15419
rect 11621 15385 11655 15419
rect 12633 15385 12667 15419
rect 17325 15385 17359 15419
rect 1501 15317 1535 15351
rect 3157 15317 3191 15351
rect 4077 15317 4111 15351
rect 4537 15317 4571 15351
rect 4905 15317 4939 15351
rect 6469 15317 6503 15351
rect 8125 15317 8159 15351
rect 9505 15317 9539 15351
rect 9873 15317 9907 15351
rect 11253 15317 11287 15351
rect 11989 15317 12023 15351
rect 12725 15317 12759 15351
rect 13369 15317 13403 15351
rect 14565 15317 14599 15351
rect 15577 15317 15611 15351
rect 15669 15317 15703 15351
rect 16497 15317 16531 15351
rect 16865 15317 16899 15351
rect 17693 15317 17727 15351
rect 17785 15317 17819 15351
rect 18337 15317 18371 15351
rect 18521 15317 18555 15351
rect 18889 15317 18923 15351
rect 19349 15317 19383 15351
rect 20177 15317 20211 15351
rect 20729 15317 20763 15351
rect 21005 15317 21039 15351
rect 21465 15317 21499 15351
rect 3985 15113 4019 15147
rect 5273 15113 5307 15147
rect 6101 15113 6135 15147
rect 7849 15113 7883 15147
rect 8401 15113 8435 15147
rect 8953 15113 8987 15147
rect 10241 15113 10275 15147
rect 12725 15113 12759 15147
rect 13461 15113 13495 15147
rect 13921 15113 13955 15147
rect 16129 15113 16163 15147
rect 20361 15113 20395 15147
rect 4445 15045 4479 15079
rect 8677 15045 8711 15079
rect 9873 15045 9907 15079
rect 12081 15045 12115 15079
rect 13553 15045 13587 15079
rect 14381 15045 14415 15079
rect 20269 15045 20303 15079
rect 1685 14977 1719 15011
rect 2053 14977 2087 15011
rect 2329 14977 2363 15011
rect 2513 14977 2547 15011
rect 2780 14977 2814 15011
rect 4353 14977 4387 15011
rect 5089 14977 5123 15011
rect 5641 14977 5675 15011
rect 6561 14977 6595 15011
rect 7389 14977 7423 15011
rect 7757 14977 7791 15011
rect 8033 14977 8067 15011
rect 9137 14977 9171 15011
rect 9413 14977 9447 15011
rect 10701 14977 10735 15011
rect 11161 14977 11195 15011
rect 11989 14977 12023 15011
rect 12633 14977 12667 15011
rect 14289 14977 14323 15011
rect 15005 14977 15039 15011
rect 17049 14977 17083 15011
rect 17305 14977 17339 15011
rect 18777 14977 18811 15011
rect 20913 14977 20947 15011
rect 21281 14977 21315 15011
rect 4537 14909 4571 14943
rect 5733 14909 5767 14943
rect 5825 14909 5859 14943
rect 7021 14909 7055 14943
rect 9689 14909 9723 14943
rect 9781 14909 9815 14943
rect 10793 14909 10827 14943
rect 10977 14909 11011 14943
rect 11805 14909 11839 14943
rect 12817 14909 12851 14943
rect 13645 14909 13679 14943
rect 14473 14909 14507 14943
rect 14749 14909 14783 14943
rect 16865 14909 16899 14943
rect 18521 14909 18555 14943
rect 20085 14909 20119 14943
rect 1869 14841 1903 14875
rect 2145 14841 2179 14875
rect 3893 14841 3927 14875
rect 8217 14841 8251 14875
rect 8493 14841 8527 14875
rect 10333 14841 10367 14875
rect 11529 14841 11563 14875
rect 21097 14841 21131 14875
rect 1501 14773 1535 14807
rect 4997 14773 5031 14807
rect 6377 14773 6411 14807
rect 7573 14773 7607 14807
rect 12265 14773 12299 14807
rect 13093 14773 13127 14807
rect 18429 14773 18463 14807
rect 19901 14773 19935 14807
rect 20729 14773 20763 14807
rect 21465 14773 21499 14807
rect 1777 14569 1811 14603
rect 2145 14569 2179 14603
rect 3065 14569 3099 14603
rect 3341 14569 3375 14603
rect 11897 14569 11931 14603
rect 13369 14569 13403 14603
rect 17233 14569 17267 14603
rect 18521 14569 18555 14603
rect 2513 14501 2547 14535
rect 3617 14501 3651 14535
rect 15485 14501 15519 14535
rect 17141 14501 17175 14535
rect 18153 14501 18187 14535
rect 18889 14501 18923 14535
rect 5549 14433 5583 14467
rect 5641 14433 5675 14467
rect 8585 14433 8619 14467
rect 9505 14433 9539 14467
rect 10057 14433 10091 14467
rect 11989 14433 12023 14467
rect 17785 14433 17819 14467
rect 19441 14433 19475 14467
rect 20637 14433 20671 14467
rect 1685 14365 1719 14399
rect 1961 14365 1995 14399
rect 2421 14365 2455 14399
rect 2697 14365 2731 14399
rect 2881 14365 2915 14399
rect 3157 14365 3191 14399
rect 3433 14365 3467 14399
rect 3801 14365 3835 14399
rect 8329 14365 8363 14399
rect 10333 14365 10367 14399
rect 10517 14365 10551 14399
rect 12256 14365 12290 14399
rect 14105 14365 14139 14399
rect 14361 14365 14395 14399
rect 15761 14365 15795 14399
rect 17601 14365 17635 14399
rect 17693 14365 17727 14399
rect 18337 14365 18371 14399
rect 18797 14365 18831 14399
rect 20453 14365 20487 14399
rect 20913 14365 20947 14399
rect 21281 14365 21315 14399
rect 5304 14297 5338 14331
rect 5886 14297 5920 14331
rect 10784 14297 10818 14331
rect 16028 14297 16062 14331
rect 19625 14297 19659 14331
rect 20545 14297 20579 14331
rect 1501 14229 1535 14263
rect 2237 14229 2271 14263
rect 3985 14229 4019 14263
rect 4169 14229 4203 14263
rect 7021 14229 7055 14263
rect 7205 14229 7239 14263
rect 8769 14229 8803 14263
rect 8953 14229 8987 14263
rect 9321 14229 9355 14263
rect 9413 14229 9447 14263
rect 9873 14229 9907 14263
rect 10149 14229 10183 14263
rect 13461 14229 13495 14263
rect 18613 14229 18647 14263
rect 19533 14229 19567 14263
rect 19993 14229 20027 14263
rect 20085 14229 20119 14263
rect 21097 14229 21131 14263
rect 21465 14229 21499 14263
rect 2145 14025 2179 14059
rect 2605 14025 2639 14059
rect 4353 14025 4387 14059
rect 4721 14025 4755 14059
rect 5917 14025 5951 14059
rect 6377 14025 6411 14059
rect 6837 14025 6871 14059
rect 7205 14025 7239 14059
rect 7573 14025 7607 14059
rect 9505 14025 9539 14059
rect 10885 14025 10919 14059
rect 11069 14025 11103 14059
rect 11345 14025 11379 14059
rect 12357 14025 12391 14059
rect 12725 14025 12759 14059
rect 13553 14025 13587 14059
rect 15117 14025 15151 14059
rect 15945 14025 15979 14059
rect 16681 14025 16715 14059
rect 17049 14025 17083 14059
rect 18245 14025 18279 14059
rect 3801 13957 3835 13991
rect 5549 13957 5583 13991
rect 6745 13957 6779 13991
rect 8278 13957 8312 13991
rect 10425 13957 10459 13991
rect 14657 13957 14691 13991
rect 14749 13957 14783 13991
rect 19472 13957 19506 13991
rect 20076 13957 20110 13991
rect 1685 13889 1719 13923
rect 2053 13889 2087 13923
rect 2329 13889 2363 13923
rect 2973 13889 3007 13923
rect 8033 13889 8067 13923
rect 9873 13889 9907 13923
rect 13185 13889 13219 13923
rect 14105 13889 14139 13923
rect 14289 13889 14323 13923
rect 15853 13889 15887 13923
rect 17141 13889 17175 13923
rect 17877 13889 17911 13923
rect 19717 13889 19751 13923
rect 19809 13889 19843 13923
rect 21281 13889 21315 13923
rect 2421 13821 2455 13855
rect 3065 13821 3099 13855
rect 3157 13821 3191 13855
rect 3893 13821 3927 13855
rect 4077 13821 4111 13855
rect 4813 13821 4847 13855
rect 4905 13821 4939 13855
rect 5273 13821 5307 13855
rect 5457 13821 5491 13855
rect 6009 13821 6043 13855
rect 6929 13821 6963 13855
rect 7665 13821 7699 13855
rect 7757 13821 7791 13855
rect 9965 13821 9999 13855
rect 10057 13821 10091 13855
rect 10609 13821 10643 13855
rect 10701 13821 10735 13855
rect 11529 13821 11563 13855
rect 11713 13821 11747 13855
rect 12081 13821 12115 13855
rect 12265 13821 12299 13855
rect 12909 13821 12943 13855
rect 13093 13821 13127 13855
rect 13921 13821 13955 13855
rect 14565 13821 14599 13855
rect 16037 13821 16071 13855
rect 17233 13821 17267 13855
rect 17693 13821 17727 13855
rect 17785 13821 17819 13855
rect 15485 13753 15519 13787
rect 18337 13753 18371 13787
rect 1501 13685 1535 13719
rect 1869 13685 1903 13719
rect 3433 13685 3467 13719
rect 9413 13685 9447 13719
rect 13645 13685 13679 13719
rect 16313 13685 16347 13719
rect 21189 13685 21223 13719
rect 21465 13685 21499 13719
rect 1777 13481 1811 13515
rect 4169 13481 4203 13515
rect 5273 13481 5307 13515
rect 5365 13481 5399 13515
rect 6469 13481 6503 13515
rect 6929 13481 6963 13515
rect 7757 13481 7791 13515
rect 10517 13481 10551 13515
rect 11345 13481 11379 13515
rect 11621 13481 11655 13515
rect 11989 13481 12023 13515
rect 13093 13481 13127 13515
rect 13829 13481 13863 13515
rect 16497 13481 16531 13515
rect 18245 13481 18279 13515
rect 19717 13481 19751 13515
rect 20821 13481 20855 13515
rect 3617 13413 3651 13447
rect 6745 13413 6779 13447
rect 12081 13413 12115 13447
rect 16313 13413 16347 13447
rect 19625 13413 19659 13447
rect 3801 13345 3835 13379
rect 4445 13345 4479 13379
rect 4721 13345 4755 13379
rect 5917 13345 5951 13379
rect 7481 13345 7515 13379
rect 8309 13345 8343 13379
rect 9045 13345 9079 13379
rect 11069 13345 11103 13379
rect 12633 13345 12667 13379
rect 14473 13345 14507 13379
rect 17049 13345 17083 13379
rect 17601 13345 17635 13379
rect 18797 13345 18831 13379
rect 20177 13345 20211 13379
rect 20269 13345 20303 13379
rect 1685 13277 1719 13311
rect 3157 13277 3191 13311
rect 3433 13277 3467 13311
rect 4905 13277 4939 13311
rect 6285 13277 6319 13311
rect 8125 13277 8159 13311
rect 9301 13277 9335 13311
rect 10977 13277 11011 13311
rect 11805 13277 11839 13311
rect 14740 13277 14774 13311
rect 15945 13277 15979 13311
rect 18613 13277 18647 13311
rect 19257 13277 19291 13311
rect 19441 13277 19475 13311
rect 20085 13277 20119 13311
rect 20637 13277 20671 13311
rect 20913 13277 20947 13311
rect 21281 13277 21315 13311
rect 2912 13209 2946 13243
rect 4813 13209 4847 13243
rect 8585 13209 8619 13243
rect 13277 13209 13311 13243
rect 14381 13209 14415 13243
rect 16865 13209 16899 13243
rect 17785 13209 17819 13243
rect 1501 13141 1535 13175
rect 3249 13141 3283 13175
rect 5733 13141 5767 13175
rect 5825 13141 5859 13175
rect 6653 13141 6687 13175
rect 7297 13141 7331 13175
rect 7389 13141 7423 13175
rect 8217 13141 8251 13175
rect 10425 13141 10459 13175
rect 10885 13141 10919 13175
rect 12357 13141 12391 13175
rect 12817 13141 12851 13175
rect 13369 13141 13403 13175
rect 13553 13141 13587 13175
rect 14197 13141 14231 13175
rect 15853 13141 15887 13175
rect 16221 13141 16255 13175
rect 16957 13141 16991 13175
rect 17693 13141 17727 13175
rect 18153 13141 18187 13175
rect 18705 13141 18739 13175
rect 21097 13141 21131 13175
rect 21465 13141 21499 13175
rect 1501 12937 1535 12971
rect 4261 12937 4295 12971
rect 7849 12937 7883 12971
rect 8217 12937 8251 12971
rect 9597 12937 9631 12971
rect 10057 12937 10091 12971
rect 10793 12937 10827 12971
rect 11069 12937 11103 12971
rect 13369 12937 13403 12971
rect 13829 12937 13863 12971
rect 14105 12937 14139 12971
rect 15393 12937 15427 12971
rect 16681 12937 16715 12971
rect 18153 12937 18187 12971
rect 18521 12937 18555 12971
rect 18981 12937 19015 12971
rect 19901 12937 19935 12971
rect 20361 12937 20395 12971
rect 2513 12869 2547 12903
rect 4721 12869 4755 12903
rect 9137 12869 9171 12903
rect 13277 12869 13311 12903
rect 15025 12869 15059 12903
rect 18613 12869 18647 12903
rect 19349 12869 19383 12903
rect 21097 12869 21131 12903
rect 1685 12801 1719 12835
rect 1961 12801 1995 12835
rect 2789 12801 2823 12835
rect 3056 12801 3090 12835
rect 4629 12801 4663 12835
rect 5733 12801 5767 12835
rect 6644 12801 6678 12835
rect 8309 12801 8343 12835
rect 9965 12801 9999 12835
rect 11345 12801 11379 12835
rect 11529 12801 11563 12835
rect 11796 12801 11830 12835
rect 14381 12801 14415 12835
rect 15669 12801 15703 12835
rect 15853 12801 15887 12835
rect 16405 12801 16439 12835
rect 17794 12801 17828 12835
rect 20085 12801 20119 12835
rect 20177 12801 20211 12835
rect 20545 12801 20579 12835
rect 21281 12801 21315 12835
rect 4813 12733 4847 12767
rect 5181 12733 5215 12767
rect 5917 12733 5951 12767
rect 6377 12733 6411 12767
rect 8401 12733 8435 12767
rect 8953 12733 8987 12767
rect 9045 12733 9079 12767
rect 10241 12733 10275 12767
rect 13093 12733 13127 12767
rect 14749 12733 14783 12767
rect 14933 12733 14967 12767
rect 18061 12733 18095 12767
rect 18797 12733 18831 12767
rect 19441 12733 19475 12767
rect 19533 12733 19567 12767
rect 4169 12665 4203 12699
rect 7757 12665 7791 12699
rect 10609 12665 10643 12699
rect 14473 12665 14507 12699
rect 15485 12665 15519 12699
rect 6101 12597 6135 12631
rect 9505 12597 9539 12631
rect 10517 12597 10551 12631
rect 11161 12597 11195 12631
rect 12909 12597 12943 12631
rect 13737 12597 13771 12631
rect 21465 12597 21499 12631
rect 1593 12393 1627 12427
rect 3157 12393 3191 12427
rect 3433 12393 3467 12427
rect 4813 12393 4847 12427
rect 10057 12393 10091 12427
rect 13645 12393 13679 12427
rect 14473 12393 14507 12427
rect 15393 12393 15427 12427
rect 16865 12393 16899 12427
rect 17049 12393 17083 12427
rect 18705 12393 18739 12427
rect 3893 12325 3927 12359
rect 7481 12325 7515 12359
rect 10333 12325 10367 12359
rect 17877 12325 17911 12359
rect 4537 12257 4571 12291
rect 6193 12257 6227 12291
rect 6837 12257 6871 12291
rect 8401 12257 8435 12291
rect 9413 12257 9447 12291
rect 9505 12257 9539 12291
rect 12909 12257 12943 12291
rect 14749 12257 14783 12291
rect 14933 12257 14967 12291
rect 15485 12257 15519 12291
rect 18153 12257 18187 12291
rect 1409 12189 1443 12223
rect 1685 12189 1719 12223
rect 1952 12189 1986 12223
rect 3341 12189 3375 12223
rect 4353 12189 4387 12223
rect 4445 12189 4479 12223
rect 7665 12189 7699 12223
rect 8677 12189 8711 12223
rect 9965 12189 9999 12223
rect 11069 12189 11103 12223
rect 11336 12189 11370 12223
rect 13001 12189 13035 12223
rect 17509 12189 17543 12223
rect 17693 12189 17727 12223
rect 18337 12189 18371 12223
rect 18889 12189 18923 12223
rect 19257 12189 19291 12223
rect 19441 12189 19475 12223
rect 20177 12189 20211 12223
rect 20545 12189 20579 12223
rect 21281 12189 21315 12223
rect 5926 12121 5960 12155
rect 10793 12121 10827 12155
rect 12541 12121 12575 12155
rect 13093 12121 13127 12155
rect 14105 12121 14139 12155
rect 15752 12121 15786 12155
rect 17233 12121 17267 12155
rect 19901 12121 19935 12155
rect 20913 12121 20947 12155
rect 21097 12121 21131 12155
rect 3065 12053 3099 12087
rect 3985 12053 4019 12087
rect 6285 12053 6319 12087
rect 6653 12053 6687 12087
rect 6745 12053 6779 12087
rect 7113 12053 7147 12087
rect 7389 12053 7423 12087
rect 7941 12053 7975 12087
rect 8125 12053 8159 12087
rect 8493 12053 8527 12087
rect 8953 12053 8987 12087
rect 9321 12053 9355 12087
rect 9781 12053 9815 12087
rect 10425 12053 10459 12087
rect 10701 12053 10735 12087
rect 12449 12053 12483 12087
rect 13461 12053 13495 12087
rect 13921 12053 13955 12087
rect 14381 12053 14415 12087
rect 15025 12053 15059 12087
rect 18245 12053 18279 12087
rect 19073 12053 19107 12087
rect 19809 12053 19843 12087
rect 21465 12053 21499 12087
rect 3249 11849 3283 11883
rect 3617 11849 3651 11883
rect 3709 11849 3743 11883
rect 4353 11849 4387 11883
rect 5733 11849 5767 11883
rect 6469 11849 6503 11883
rect 6929 11849 6963 11883
rect 7297 11849 7331 11883
rect 7757 11849 7791 11883
rect 8125 11849 8159 11883
rect 8493 11849 8527 11883
rect 11345 11849 11379 11883
rect 11897 11849 11931 11883
rect 12725 11849 12759 11883
rect 13645 11849 13679 11883
rect 16221 11849 16255 11883
rect 16957 11849 16991 11883
rect 18061 11849 18095 11883
rect 18613 11849 18647 11883
rect 5181 11781 5215 11815
rect 6837 11781 6871 11815
rect 13553 11781 13587 11815
rect 14381 11781 14415 11815
rect 16681 11781 16715 11815
rect 18153 11781 18187 11815
rect 20002 11781 20036 11815
rect 1961 11713 1995 11747
rect 2237 11713 2271 11747
rect 2697 11713 2731 11747
rect 4077 11713 4111 11747
rect 5825 11713 5859 11747
rect 7665 11713 7699 11747
rect 8585 11713 8619 11747
rect 9413 11713 9447 11747
rect 9781 11713 9815 11747
rect 10221 11713 10255 11747
rect 14289 11713 14323 11747
rect 15761 11713 15795 11747
rect 15853 11713 15887 11747
rect 17877 11713 17911 11747
rect 18337 11713 18371 11747
rect 18797 11713 18831 11747
rect 20545 11713 20579 11747
rect 20729 11713 20763 11747
rect 21005 11713 21039 11747
rect 2513 11645 2547 11679
rect 2605 11645 2639 11679
rect 3893 11645 3927 11679
rect 5641 11645 5675 11679
rect 7113 11645 7147 11679
rect 7941 11645 7975 11679
rect 8677 11645 8711 11679
rect 9965 11645 9999 11679
rect 11713 11645 11747 11679
rect 11805 11645 11839 11679
rect 12817 11645 12851 11679
rect 13001 11645 13035 11679
rect 13737 11645 13771 11679
rect 14197 11645 14231 11679
rect 15669 11645 15703 11679
rect 20269 11645 20303 11679
rect 4445 11577 4479 11611
rect 6193 11577 6227 11611
rect 12265 11577 12299 11611
rect 14749 11577 14783 11611
rect 17693 11577 17727 11611
rect 18521 11577 18555 11611
rect 3065 11509 3099 11543
rect 4629 11509 4663 11543
rect 4813 11509 4847 11543
rect 5089 11509 5123 11543
rect 9045 11509 9079 11543
rect 12357 11509 12391 11543
rect 13185 11509 13219 11543
rect 14933 11509 14967 11543
rect 15209 11509 15243 11543
rect 15393 11509 15427 11543
rect 16405 11509 16439 11543
rect 17049 11509 17083 11543
rect 17325 11509 17359 11543
rect 17509 11509 17543 11543
rect 18889 11509 18923 11543
rect 20453 11509 20487 11543
rect 1501 11305 1535 11339
rect 2237 11305 2271 11339
rect 5641 11305 5675 11339
rect 6469 11305 6503 11339
rect 11161 11305 11195 11339
rect 13737 11305 13771 11339
rect 15761 11305 15795 11339
rect 19073 11305 19107 11339
rect 2053 11237 2087 11271
rect 3341 11237 3375 11271
rect 7481 11237 7515 11271
rect 8493 11237 8527 11271
rect 8677 11237 8711 11271
rect 9045 11237 9079 11271
rect 16589 11237 16623 11271
rect 17417 11237 17451 11271
rect 2513 11169 2547 11203
rect 5825 11169 5859 11203
rect 7113 11169 7147 11203
rect 7205 11169 7239 11203
rect 8033 11169 8067 11203
rect 10425 11169 10459 11203
rect 11437 11169 11471 11203
rect 12265 11169 12299 11203
rect 13369 11169 13403 11203
rect 13553 11169 13587 11203
rect 14289 11169 14323 11203
rect 16221 11169 16255 11203
rect 16313 11169 16347 11203
rect 17049 11169 17083 11203
rect 17233 11169 17267 11203
rect 21281 11169 21315 11203
rect 1685 11101 1719 11135
rect 1869 11101 1903 11135
rect 2973 11101 3007 11135
rect 3165 11101 3199 11135
rect 3617 11101 3651 11135
rect 4169 11101 4203 11135
rect 4261 11101 4295 11135
rect 6101 11101 6135 11135
rect 7941 11101 7975 11135
rect 8309 11101 8343 11135
rect 10158 11101 10192 11135
rect 11529 11101 11563 11135
rect 12449 11101 12483 11135
rect 14105 11101 14139 11135
rect 17693 11101 17727 11135
rect 19257 11101 19291 11135
rect 3801 11033 3835 11067
rect 4528 11033 4562 11067
rect 7849 11033 7883 11067
rect 10977 11033 11011 11067
rect 11621 11033 11655 11067
rect 14556 11033 14590 11067
rect 16129 11033 16163 11067
rect 17960 11033 17994 11067
rect 19524 11033 19558 11067
rect 21097 11033 21131 11067
rect 21189 11033 21223 11067
rect 3433 10965 3467 10999
rect 3985 10965 4019 10999
rect 6009 10965 6043 10999
rect 6653 10965 6687 10999
rect 7021 10965 7055 10999
rect 10517 10965 10551 10999
rect 11989 10965 12023 10999
rect 12357 10965 12391 10999
rect 12817 10965 12851 10999
rect 12909 10965 12943 10999
rect 13277 10965 13311 10999
rect 15669 10965 15703 10999
rect 16957 10965 16991 10999
rect 20637 10965 20671 10999
rect 20729 10965 20763 10999
rect 3157 10761 3191 10795
rect 6193 10761 6227 10795
rect 6377 10761 6411 10795
rect 9689 10761 9723 10795
rect 10057 10761 10091 10795
rect 10517 10761 10551 10795
rect 10977 10761 11011 10795
rect 11897 10761 11931 10795
rect 12357 10761 12391 10795
rect 14105 10761 14139 10795
rect 14933 10761 14967 10795
rect 15301 10761 15335 10795
rect 16129 10761 16163 10795
rect 16681 10761 16715 10795
rect 17509 10761 17543 10795
rect 17969 10761 18003 10795
rect 19165 10761 19199 10795
rect 19993 10761 20027 10795
rect 3494 10693 3528 10727
rect 8962 10693 8996 10727
rect 13562 10693 13596 10727
rect 15761 10693 15795 10727
rect 17141 10693 17175 10727
rect 21290 10693 21324 10727
rect 1501 10625 1535 10659
rect 1685 10625 1719 10659
rect 2044 10625 2078 10659
rect 3249 10625 3283 10659
rect 5365 10625 5399 10659
rect 5825 10625 5859 10659
rect 7490 10625 7524 10659
rect 9229 10625 9263 10659
rect 11253 10625 11287 10659
rect 11989 10625 12023 10659
rect 13829 10625 13863 10659
rect 13921 10625 13955 10659
rect 14381 10625 14415 10659
rect 16405 10625 16439 10659
rect 17049 10625 17083 10659
rect 17877 10625 17911 10659
rect 18705 10625 18739 10659
rect 19533 10625 19567 10659
rect 21557 10625 21591 10659
rect 1777 10557 1811 10591
rect 4813 10557 4847 10591
rect 5549 10557 5583 10591
rect 5733 10557 5767 10591
rect 7757 10557 7791 10591
rect 9413 10557 9447 10591
rect 9597 10557 9631 10591
rect 10609 10557 10643 10591
rect 10701 10557 10735 10591
rect 11713 10557 11747 10591
rect 14657 10557 14691 10591
rect 14841 10557 14875 10591
rect 15485 10557 15519 10591
rect 15669 10557 15703 10591
rect 17233 10557 17267 10591
rect 18153 10557 18187 10591
rect 18521 10557 18555 10591
rect 18613 10557 18647 10591
rect 19625 10557 19659 10591
rect 19809 10557 19843 10591
rect 4629 10489 4663 10523
rect 20177 10489 20211 10523
rect 5181 10421 5215 10455
rect 7849 10421 7883 10455
rect 10149 10421 10183 10455
rect 12449 10421 12483 10455
rect 14289 10421 14323 10455
rect 19073 10421 19107 10455
rect 3433 10217 3467 10251
rect 5181 10217 5215 10251
rect 6377 10217 6411 10251
rect 8769 10217 8803 10251
rect 11897 10217 11931 10251
rect 15669 10217 15703 10251
rect 18245 10217 18279 10251
rect 19257 10217 19291 10251
rect 1685 10149 1719 10183
rect 3341 10149 3375 10183
rect 5273 10149 5307 10183
rect 6193 10149 6227 10183
rect 9965 10149 9999 10183
rect 15485 10149 15519 10183
rect 16773 10149 16807 10183
rect 19073 10149 19107 10183
rect 1961 10081 1995 10115
rect 4629 10081 4663 10115
rect 5825 10081 5859 10115
rect 6561 10081 6595 10115
rect 7389 10081 7423 10115
rect 8217 10081 8251 10115
rect 9689 10081 9723 10115
rect 10517 10081 10551 10115
rect 11345 10081 11379 10115
rect 12081 10081 12115 10115
rect 12541 10081 12575 10115
rect 12725 10081 12759 10115
rect 13277 10081 13311 10115
rect 14105 10081 14139 10115
rect 16313 10081 16347 10115
rect 18429 10081 18463 10115
rect 19717 10081 19751 10115
rect 19809 10081 19843 10115
rect 21005 10081 21039 10115
rect 1501 10013 1535 10047
rect 3617 10013 3651 10047
rect 3801 10013 3835 10047
rect 4077 10013 4111 10047
rect 4813 10013 4847 10047
rect 9505 10013 9539 10047
rect 12265 10013 12299 10047
rect 12817 10013 12851 10047
rect 16865 10013 16899 10047
rect 18705 10013 18739 10047
rect 19625 10013 19659 10047
rect 20453 10013 20487 10047
rect 20729 10013 20763 10047
rect 2228 9945 2262 9979
rect 7113 9945 7147 9979
rect 9597 9945 9631 9979
rect 10609 9945 10643 9979
rect 10701 9945 10735 9979
rect 11529 9945 11563 9979
rect 13553 9945 13587 9979
rect 13829 9945 13863 9979
rect 14372 9945 14406 9979
rect 17110 9945 17144 9979
rect 20085 9945 20119 9979
rect 20269 9945 20303 9979
rect 1869 9877 1903 9911
rect 3985 9877 4019 9911
rect 4261 9877 4295 9911
rect 4721 9877 4755 9911
rect 5641 9877 5675 9911
rect 5733 9877 5767 9911
rect 6653 9877 6687 9911
rect 6929 9877 6963 9911
rect 7481 9877 7515 9911
rect 7573 9877 7607 9911
rect 7941 9877 7975 9911
rect 8309 9877 8343 9911
rect 8401 9877 8435 9911
rect 8953 9877 8987 9911
rect 9137 9877 9171 9911
rect 10149 9877 10183 9911
rect 11069 9877 11103 9911
rect 11437 9877 11471 9911
rect 13185 9877 13219 9911
rect 16037 9877 16071 9911
rect 16129 9877 16163 9911
rect 16497 9877 16531 9911
rect 18613 9877 18647 9911
rect 20637 9877 20671 9911
rect 7573 9673 7607 9707
rect 9781 9673 9815 9707
rect 9873 9673 9907 9707
rect 12909 9673 12943 9707
rect 19717 9673 19751 9707
rect 1501 9605 1535 9639
rect 7113 9605 7147 9639
rect 7941 9605 7975 9639
rect 10241 9605 10275 9639
rect 10885 9605 10919 9639
rect 12357 9605 12391 9639
rect 12817 9605 12851 9639
rect 15669 9605 15703 9639
rect 16129 9605 16163 9639
rect 16405 9605 16439 9639
rect 19257 9605 19291 9639
rect 21097 9605 21131 9639
rect 2237 9537 2271 9571
rect 2697 9537 2731 9571
rect 3801 9537 3835 9571
rect 3893 9537 3927 9571
rect 4721 9537 4755 9571
rect 5549 9537 5583 9571
rect 6193 9537 6227 9571
rect 6653 9537 6687 9571
rect 8401 9537 8435 9571
rect 8668 9537 8702 9571
rect 10333 9537 10367 9571
rect 10701 9537 10735 9571
rect 11897 9537 11931 9571
rect 13461 9537 13495 9571
rect 13829 9537 13863 9571
rect 14473 9537 14507 9571
rect 15025 9537 15059 9571
rect 15761 9537 15795 9571
rect 17141 9537 17175 9571
rect 17969 9537 18003 9571
rect 18797 9537 18831 9571
rect 19349 9537 19383 9571
rect 20177 9537 20211 9571
rect 21005 9537 21039 9571
rect 1961 9469 1995 9503
rect 2145 9469 2179 9503
rect 3525 9469 3559 9503
rect 4813 9469 4847 9503
rect 4905 9469 4939 9503
rect 5641 9469 5675 9503
rect 5733 9469 5767 9503
rect 6837 9469 6871 9503
rect 7021 9469 7055 9503
rect 8033 9469 8067 9503
rect 8125 9469 8159 9503
rect 10425 9469 10459 9503
rect 11161 9469 11195 9503
rect 11713 9469 11747 9503
rect 11805 9469 11839 9503
rect 12633 9469 12667 9503
rect 15945 9469 15979 9503
rect 16957 9469 16991 9503
rect 17049 9469 17083 9503
rect 18061 9469 18095 9503
rect 18153 9469 18187 9503
rect 19165 9469 19199 9503
rect 20269 9469 20303 9503
rect 20453 9469 20487 9503
rect 21281 9469 21315 9503
rect 1685 9401 1719 9435
rect 2605 9401 2639 9435
rect 4077 9401 4111 9435
rect 7481 9401 7515 9435
rect 11253 9401 11287 9435
rect 12265 9401 12299 9435
rect 15301 9401 15335 9435
rect 17601 9401 17635 9435
rect 18613 9401 18647 9435
rect 20637 9401 20671 9435
rect 2881 9333 2915 9367
rect 4353 9333 4387 9367
rect 5181 9333 5215 9367
rect 6009 9333 6043 9367
rect 6469 9333 6503 9367
rect 13277 9333 13311 9367
rect 14289 9333 14323 9367
rect 14657 9333 14691 9367
rect 14841 9333 14875 9367
rect 15209 9333 15243 9367
rect 17509 9333 17543 9367
rect 18521 9333 18555 9367
rect 19809 9333 19843 9367
rect 21465 9333 21499 9367
rect 2145 9129 2179 9163
rect 2237 9129 2271 9163
rect 3801 9129 3835 9163
rect 4629 9129 4663 9163
rect 5273 9129 5307 9163
rect 6101 9129 6135 9163
rect 8033 9129 8067 9163
rect 10333 9129 10367 9163
rect 10517 9129 10551 9163
rect 17141 9129 17175 9163
rect 20729 9129 20763 9163
rect 6929 9061 6963 9095
rect 7849 9061 7883 9095
rect 17049 9061 17083 9095
rect 1593 8993 1627 9027
rect 3617 8993 3651 9027
rect 4261 8993 4295 9027
rect 4353 8993 4387 9027
rect 5917 8993 5951 9027
rect 6745 8993 6779 9027
rect 7573 8993 7607 9027
rect 8493 8993 8527 9027
rect 8677 8993 8711 9027
rect 13093 8993 13127 9027
rect 15669 8993 15703 9027
rect 17785 8993 17819 9027
rect 18521 8993 18555 9027
rect 18797 8993 18831 9027
rect 21281 8993 21315 9027
rect 3350 8925 3384 8959
rect 4169 8925 4203 8959
rect 4813 8925 4847 8959
rect 4905 8925 4939 8959
rect 7297 8925 7331 8959
rect 8953 8925 8987 8959
rect 10977 8925 11011 8959
rect 12449 8925 12483 8959
rect 12909 8925 12943 8959
rect 14105 8925 14139 8959
rect 15936 8925 15970 8959
rect 19257 8925 19291 8959
rect 21097 8925 21131 8959
rect 1685 8857 1719 8891
rect 6561 8857 6595 8891
rect 9220 8857 9254 8891
rect 12182 8857 12216 8891
rect 13645 8857 13679 8891
rect 14350 8857 14384 8891
rect 17601 8857 17635 8891
rect 18429 8857 18463 8891
rect 18981 8857 19015 8891
rect 19502 8857 19536 8891
rect 1777 8789 1811 8823
rect 5089 8789 5123 8823
rect 5641 8789 5675 8823
rect 5733 8789 5767 8823
rect 6469 8789 6503 8823
rect 7389 8789 7423 8823
rect 8401 8789 8435 8823
rect 10609 8789 10643 8823
rect 10793 8789 10827 8823
rect 11069 8789 11103 8823
rect 12541 8789 12575 8823
rect 13001 8789 13035 8823
rect 13553 8789 13587 8823
rect 13921 8789 13955 8823
rect 15485 8789 15519 8823
rect 17509 8789 17543 8823
rect 17969 8789 18003 8823
rect 18337 8789 18371 8823
rect 20637 8789 20671 8823
rect 21189 8789 21223 8823
rect 1501 8585 1535 8619
rect 2329 8585 2363 8619
rect 2421 8585 2455 8619
rect 2881 8585 2915 8619
rect 3893 8585 3927 8619
rect 3985 8585 4019 8619
rect 4445 8585 4479 8619
rect 5273 8585 5307 8619
rect 5641 8585 5675 8619
rect 6193 8585 6227 8619
rect 7757 8585 7791 8619
rect 9229 8585 9263 8619
rect 9597 8585 9631 8619
rect 10149 8585 10183 8619
rect 10517 8585 10551 8619
rect 10977 8585 11011 8619
rect 11345 8585 11379 8619
rect 13001 8585 13035 8619
rect 14657 8585 14691 8619
rect 15393 8585 15427 8619
rect 15761 8585 15795 8619
rect 18337 8585 18371 8619
rect 18705 8585 18739 8619
rect 20269 8585 20303 8619
rect 20453 8585 20487 8619
rect 3525 8517 3559 8551
rect 6644 8517 6678 8551
rect 7849 8517 7883 8551
rect 8309 8517 8343 8551
rect 13461 8517 13495 8551
rect 15853 8517 15887 8551
rect 17794 8517 17828 8551
rect 20545 8517 20579 8551
rect 1961 8449 1995 8483
rect 2789 8449 2823 8483
rect 3341 8449 3375 8483
rect 4813 8449 4847 8483
rect 5733 8449 5767 8483
rect 8033 8449 8067 8483
rect 8677 8449 8711 8483
rect 9045 8449 9079 8483
rect 10885 8449 10919 8483
rect 12642 8449 12676 8483
rect 12909 8449 12943 8483
rect 13369 8449 13403 8483
rect 14105 8449 14139 8483
rect 16497 8449 16531 8483
rect 18429 8449 18463 8483
rect 19818 8449 19852 8483
rect 20729 8449 20763 8483
rect 1685 8381 1719 8415
rect 1869 8381 1903 8415
rect 3065 8381 3099 8415
rect 3709 8381 3743 8415
rect 4905 8381 4939 8415
rect 4997 8381 5031 8415
rect 5917 8381 5951 8415
rect 6377 8381 6411 8415
rect 9689 8381 9723 8415
rect 9873 8381 9907 8415
rect 10793 8381 10827 8415
rect 13553 8381 13587 8415
rect 13829 8381 13863 8415
rect 15209 8381 15243 8415
rect 15301 8381 15335 8415
rect 18061 8381 18095 8415
rect 20085 8381 20119 8415
rect 21005 8381 21039 8415
rect 10333 8313 10367 8347
rect 14289 8313 14323 8347
rect 14565 8313 14599 8347
rect 16037 8313 16071 8347
rect 16313 8313 16347 8347
rect 16681 8313 16715 8347
rect 18613 8313 18647 8347
rect 4353 8245 4387 8279
rect 11529 8245 11563 8279
rect 14933 8245 14967 8279
rect 1501 8041 1535 8075
rect 2329 8041 2363 8075
rect 3801 8041 3835 8075
rect 5181 8041 5215 8075
rect 6561 8041 6595 8075
rect 7573 8041 7607 8075
rect 10149 8041 10183 8075
rect 10609 8041 10643 8075
rect 15577 8041 15611 8075
rect 17233 8041 17267 8075
rect 18337 8041 18371 8075
rect 19257 8041 19291 8075
rect 20361 8041 20395 8075
rect 21281 8041 21315 8075
rect 9965 7973 9999 8007
rect 12909 7973 12943 8007
rect 16589 7973 16623 8007
rect 18245 7973 18279 8007
rect 1961 7905 1995 7939
rect 2145 7905 2179 7939
rect 2973 7905 3007 7939
rect 4261 7905 4295 7939
rect 4353 7905 4387 7939
rect 5733 7905 5767 7939
rect 6929 7905 6963 7939
rect 7113 7905 7147 7939
rect 8217 7905 8251 7939
rect 8401 7905 8435 7939
rect 9505 7905 9539 7939
rect 10885 7905 10919 7939
rect 13645 7905 13679 7939
rect 13921 7905 13955 7939
rect 15025 7905 15059 7939
rect 16221 7905 16255 7939
rect 16681 7905 16715 7939
rect 17693 7905 17727 7939
rect 18889 7905 18923 7939
rect 19809 7905 19843 7939
rect 20729 7905 20763 7939
rect 1869 7837 1903 7871
rect 4629 7837 4663 7871
rect 5089 7837 5123 7871
rect 6193 7837 6227 7871
rect 6469 7837 6503 7871
rect 6745 7837 6779 7871
rect 7205 7837 7239 7871
rect 9321 7837 9355 7871
rect 11529 7837 11563 7871
rect 13369 7837 13403 7871
rect 14289 7837 14323 7871
rect 16957 7837 16991 7871
rect 17417 7837 17451 7871
rect 19441 7837 19475 7871
rect 19901 7837 19935 7871
rect 19993 7837 20027 7871
rect 20913 7837 20947 7871
rect 2789 7769 2823 7803
rect 3249 7769 3283 7803
rect 3433 7769 3467 7803
rect 5549 7769 5583 7803
rect 9413 7769 9447 7803
rect 11069 7769 11103 7803
rect 11796 7769 11830 7803
rect 14381 7769 14415 7803
rect 14749 7769 14783 7803
rect 16037 7769 16071 7803
rect 16129 7769 16163 7803
rect 17785 7769 17819 7803
rect 18797 7769 18831 7803
rect 21373 7769 21407 7803
rect 2697 7701 2731 7735
rect 3617 7701 3651 7735
rect 4169 7701 4203 7735
rect 4905 7701 4939 7735
rect 5641 7701 5675 7735
rect 6009 7701 6043 7735
rect 6285 7701 6319 7735
rect 7757 7701 7791 7735
rect 8125 7701 8159 7735
rect 8585 7701 8619 7735
rect 8953 7701 8987 7735
rect 9781 7701 9815 7735
rect 10333 7701 10367 7735
rect 10977 7701 11011 7735
rect 11437 7701 11471 7735
rect 13001 7701 13035 7735
rect 13461 7701 13495 7735
rect 15117 7701 15151 7735
rect 15209 7701 15243 7735
rect 15669 7701 15703 7735
rect 17049 7701 17083 7735
rect 17877 7701 17911 7735
rect 18705 7701 18739 7735
rect 20821 7701 20855 7735
rect 1593 7497 1627 7531
rect 6193 7497 6227 7531
rect 7573 7497 7607 7531
rect 10149 7497 10183 7531
rect 11805 7497 11839 7531
rect 12265 7497 12299 7531
rect 13645 7497 13679 7531
rect 13737 7497 13771 7531
rect 15853 7497 15887 7531
rect 17141 7497 17175 7531
rect 17877 7497 17911 7531
rect 19717 7497 19751 7531
rect 20177 7497 20211 7531
rect 21189 7497 21223 7531
rect 2982 7429 3016 7463
rect 10057 7429 10091 7463
rect 12173 7429 12207 7463
rect 18604 7429 18638 7463
rect 20269 7429 20303 7463
rect 21465 7429 21499 7463
rect 1409 7361 1443 7395
rect 3249 7361 3283 7395
rect 3341 7361 3375 7395
rect 3597 7361 3631 7395
rect 5069 7361 5103 7395
rect 6745 7361 6779 7395
rect 7205 7361 7239 7395
rect 8686 7361 8720 7395
rect 8953 7361 8987 7395
rect 9045 7361 9079 7395
rect 11161 7361 11195 7395
rect 11529 7361 11563 7395
rect 12725 7361 12759 7395
rect 13277 7361 13311 7395
rect 14105 7361 14139 7395
rect 15025 7361 15059 7395
rect 15485 7361 15519 7395
rect 16313 7361 16347 7395
rect 17049 7361 17083 7395
rect 18337 7361 18371 7395
rect 19993 7361 20027 7395
rect 20821 7361 20855 7395
rect 4813 7293 4847 7327
rect 6469 7293 6503 7327
rect 6653 7293 6687 7327
rect 9321 7293 9355 7327
rect 10609 7293 10643 7327
rect 12357 7293 12391 7327
rect 13001 7293 13035 7327
rect 13185 7293 13219 7327
rect 14197 7293 14231 7327
rect 14289 7293 14323 7327
rect 14841 7293 14875 7327
rect 15209 7293 15243 7327
rect 15393 7293 15427 7327
rect 16037 7293 16071 7327
rect 17233 7293 17267 7327
rect 17969 7293 18003 7327
rect 18153 7293 18187 7327
rect 20637 7293 20671 7327
rect 20729 7293 20763 7327
rect 10701 7225 10735 7259
rect 11345 7225 11379 7259
rect 16681 7225 16715 7259
rect 1869 7157 1903 7191
rect 4721 7157 4755 7191
rect 7113 7157 7147 7191
rect 7389 7157 7423 7191
rect 10425 7157 10459 7191
rect 11069 7157 11103 7191
rect 11713 7157 11747 7191
rect 14657 7157 14691 7191
rect 16221 7157 16255 7191
rect 16497 7157 16531 7191
rect 17509 7157 17543 7191
rect 19809 7157 19843 7191
rect 21373 7157 21407 7191
rect 3617 6953 3651 6987
rect 3801 6953 3835 6987
rect 12173 6953 12207 6987
rect 13185 6953 13219 6987
rect 19993 6953 20027 6987
rect 4629 6885 4663 6919
rect 8769 6885 8803 6919
rect 11897 6885 11931 6919
rect 1961 6817 1995 6851
rect 2973 6817 3007 6851
rect 4261 6817 4295 6851
rect 4445 6817 4479 6851
rect 5273 6817 5307 6851
rect 6009 6817 6043 6851
rect 8217 6817 8251 6851
rect 9505 6817 9539 6851
rect 12633 6817 12667 6851
rect 13645 6817 13679 6851
rect 16221 6817 16255 6851
rect 17969 6817 18003 6851
rect 18429 6817 18463 6851
rect 19441 6817 19475 6851
rect 2237 6749 2271 6783
rect 3157 6749 3191 6783
rect 3249 6749 3283 6783
rect 5917 6749 5951 6783
rect 6469 6749 6503 6783
rect 6561 6749 6595 6783
rect 8585 6749 8619 6783
rect 9321 6749 9355 6783
rect 11253 6749 11287 6783
rect 11529 6749 11563 6783
rect 12725 6749 12759 6783
rect 14105 6749 14139 6783
rect 16405 6749 16439 6783
rect 17702 6749 17736 6783
rect 18245 6749 18279 6783
rect 20361 6749 20395 6783
rect 20545 6749 20579 6783
rect 20729 6749 20763 6783
rect 21005 6749 21039 6783
rect 2421 6681 2455 6715
rect 2605 6681 2639 6715
rect 4169 6681 4203 6715
rect 7950 6681 7984 6715
rect 8309 6681 8343 6715
rect 10986 6681 11020 6715
rect 11621 6681 11655 6715
rect 12081 6681 12115 6715
rect 14350 6681 14384 6715
rect 15945 6681 15979 6715
rect 19533 6681 19567 6715
rect 2697 6613 2731 6647
rect 4997 6613 5031 6647
rect 5089 6613 5123 6647
rect 5457 6613 5491 6647
rect 5825 6613 5859 6647
rect 6285 6613 6319 6647
rect 6745 6613 6779 6647
rect 6837 6613 6871 6647
rect 8953 6613 8987 6647
rect 9413 6613 9447 6647
rect 9873 6613 9907 6647
rect 11345 6613 11379 6647
rect 12817 6613 12851 6647
rect 13369 6613 13403 6647
rect 13461 6613 13495 6647
rect 13921 6613 13955 6647
rect 15485 6613 15519 6647
rect 15577 6613 15611 6647
rect 16037 6613 16071 6647
rect 16589 6613 16623 6647
rect 18061 6613 18095 6647
rect 18613 6613 18647 6647
rect 18705 6613 18739 6647
rect 19073 6613 19107 6647
rect 19625 6613 19659 6647
rect 20085 6613 20119 6647
rect 1869 6409 1903 6443
rect 2237 6409 2271 6443
rect 4721 6409 4755 6443
rect 5825 6409 5859 6443
rect 6377 6409 6411 6443
rect 6837 6409 6871 6443
rect 7573 6409 7607 6443
rect 8125 6409 8159 6443
rect 8493 6409 8527 6443
rect 8585 6409 8619 6443
rect 13369 6409 13403 6443
rect 16681 6409 16715 6443
rect 18705 6409 18739 6443
rect 19257 6409 19291 6443
rect 19717 6409 19751 6443
rect 19809 6409 19843 6443
rect 21005 6409 21039 6443
rect 21373 6409 21407 6443
rect 1501 6341 1535 6375
rect 1685 6341 1719 6375
rect 3157 6341 3191 6375
rect 7665 6341 7699 6375
rect 13001 6341 13035 6375
rect 2789 6273 2823 6307
rect 3249 6273 3283 6307
rect 3505 6273 3539 6307
rect 4905 6273 4939 6307
rect 4997 6273 5031 6307
rect 5733 6273 5767 6307
rect 6745 6273 6779 6307
rect 8953 6273 8987 6307
rect 10342 6273 10376 6307
rect 10701 6273 10735 6307
rect 11345 6273 11379 6307
rect 11897 6273 11931 6307
rect 14013 6273 14047 6307
rect 14473 6273 14507 6307
rect 14740 6273 14774 6307
rect 16129 6273 16163 6307
rect 16497 6273 16531 6307
rect 16865 6273 16899 6307
rect 17049 6273 17083 6307
rect 17325 6273 17359 6307
rect 17592 6273 17626 6307
rect 19349 6273 19383 6307
rect 20177 6273 20211 6307
rect 20913 6273 20947 6307
rect 2329 6205 2363 6239
rect 2513 6205 2547 6239
rect 5917 6205 5951 6239
rect 6929 6205 6963 6239
rect 7389 6205 7423 6239
rect 8769 6205 8803 6239
rect 10609 6205 10643 6239
rect 11069 6205 11103 6239
rect 11989 6205 12023 6239
rect 12081 6205 12115 6239
rect 12725 6205 12759 6239
rect 12909 6205 12943 6239
rect 13737 6205 13771 6239
rect 13921 6205 13955 6239
rect 19073 6205 19107 6239
rect 20269 6205 20303 6239
rect 20361 6205 20395 6239
rect 20821 6205 20855 6239
rect 2973 6137 3007 6171
rect 9137 6137 9171 6171
rect 11529 6137 11563 6171
rect 15853 6137 15887 6171
rect 17233 6137 17267 6171
rect 4629 6069 4663 6103
rect 5181 6069 5215 6103
rect 5365 6069 5399 6103
rect 8033 6069 8067 6103
rect 9229 6069 9263 6103
rect 10885 6069 10919 6103
rect 12449 6069 12483 6103
rect 13553 6069 13587 6103
rect 14381 6069 14415 6103
rect 15945 6069 15979 6103
rect 16313 6069 16347 6103
rect 18889 6069 18923 6103
rect 21557 6069 21591 6103
rect 3617 5865 3651 5899
rect 5917 5865 5951 5899
rect 6193 5865 6227 5899
rect 13921 5865 13955 5899
rect 15117 5865 15151 5899
rect 19533 5865 19567 5899
rect 20361 5865 20395 5899
rect 21373 5865 21407 5899
rect 6101 5797 6135 5831
rect 11345 5797 11379 5831
rect 16957 5797 16991 5831
rect 17325 5797 17359 5831
rect 19441 5797 19475 5831
rect 2789 5729 2823 5763
rect 3065 5729 3099 5763
rect 6745 5729 6779 5763
rect 7389 5729 7423 5763
rect 8217 5729 8251 5763
rect 9137 5729 9171 5763
rect 9873 5729 9907 5763
rect 10793 5729 10827 5763
rect 11529 5729 11563 5763
rect 13185 5729 13219 5763
rect 13369 5729 13403 5763
rect 14473 5729 14507 5763
rect 16589 5729 16623 5763
rect 18705 5729 18739 5763
rect 20177 5729 20211 5763
rect 20821 5729 20855 5763
rect 20913 5729 20947 5763
rect 3985 5661 4019 5695
rect 4261 5661 4295 5695
rect 5733 5661 5767 5695
rect 7573 5661 7607 5695
rect 9229 5661 9263 5695
rect 12449 5661 12483 5695
rect 13093 5661 13127 5695
rect 13737 5661 13771 5695
rect 14105 5661 14139 5695
rect 16773 5661 16807 5695
rect 17049 5661 17083 5695
rect 18981 5661 19015 5695
rect 19257 5661 19291 5695
rect 19901 5661 19935 5695
rect 2544 5593 2578 5627
rect 3249 5593 3283 5627
rect 4169 5593 4203 5627
rect 4528 5593 4562 5627
rect 8309 5593 8343 5627
rect 9321 5593 9355 5627
rect 10977 5593 11011 5627
rect 12265 5593 12299 5627
rect 14657 5593 14691 5627
rect 16322 5593 16356 5627
rect 18438 5593 18472 5627
rect 18797 5593 18831 5627
rect 19993 5593 20027 5627
rect 21465 5593 21499 5627
rect 1409 5525 1443 5559
rect 3157 5525 3191 5559
rect 5641 5525 5675 5559
rect 6561 5525 6595 5559
rect 6653 5525 6687 5559
rect 7021 5525 7055 5559
rect 7481 5525 7515 5559
rect 7941 5525 7975 5559
rect 8401 5525 8435 5559
rect 8769 5525 8803 5559
rect 9689 5525 9723 5559
rect 10057 5525 10091 5559
rect 10149 5525 10183 5559
rect 10517 5525 10551 5559
rect 10885 5525 10919 5559
rect 11713 5525 11747 5559
rect 11805 5525 11839 5559
rect 12173 5525 12207 5559
rect 12725 5525 12759 5559
rect 13553 5525 13587 5559
rect 14289 5525 14323 5559
rect 14749 5525 14783 5559
rect 15209 5525 15243 5559
rect 17233 5525 17267 5559
rect 20729 5525 20763 5559
rect 3341 5321 3375 5355
rect 4077 5321 4111 5355
rect 4169 5321 4203 5355
rect 5825 5321 5859 5355
rect 6837 5321 6871 5355
rect 7849 5321 7883 5355
rect 8309 5321 8343 5355
rect 8677 5321 8711 5355
rect 10425 5321 10459 5355
rect 10793 5321 10827 5355
rect 10885 5321 10919 5355
rect 11529 5321 11563 5355
rect 11989 5321 12023 5355
rect 17049 5321 17083 5355
rect 17141 5321 17175 5355
rect 17785 5321 17819 5355
rect 19533 5321 19567 5355
rect 21005 5321 21039 5355
rect 21373 5321 21407 5355
rect 2421 5253 2455 5287
rect 3249 5253 3283 5287
rect 9812 5253 9846 5287
rect 14688 5253 14722 5287
rect 16129 5253 16163 5287
rect 16313 5253 16347 5287
rect 19870 5253 19904 5287
rect 21465 5253 21499 5287
rect 1961 5185 1995 5219
rect 2789 5185 2823 5219
rect 4537 5185 4571 5219
rect 5917 5185 5951 5219
rect 6745 5185 6779 5219
rect 7481 5185 7515 5219
rect 7757 5185 7791 5219
rect 8217 5185 8251 5219
rect 10057 5185 10091 5219
rect 10149 5185 10183 5219
rect 11345 5185 11379 5219
rect 11897 5185 11931 5219
rect 12357 5185 12391 5219
rect 12909 5185 12943 5219
rect 13001 5185 13035 5219
rect 14933 5185 14967 5219
rect 15025 5185 15059 5219
rect 15669 5185 15703 5219
rect 17601 5185 17635 5219
rect 17877 5185 17911 5219
rect 18153 5185 18187 5219
rect 18420 5185 18454 5219
rect 21189 5185 21223 5219
rect 2237 5117 2271 5151
rect 3525 5117 3559 5151
rect 4353 5117 4387 5151
rect 4813 5117 4847 5151
rect 6101 5117 6135 5151
rect 6929 5117 6963 5151
rect 8493 5117 8527 5151
rect 10977 5117 11011 5151
rect 12081 5117 12115 5151
rect 12817 5117 12851 5151
rect 15393 5117 15427 5151
rect 15577 5117 15611 5151
rect 16957 5117 16991 5151
rect 19625 5117 19659 5151
rect 16037 5049 16071 5083
rect 17509 5049 17543 5083
rect 2513 4981 2547 5015
rect 2881 4981 2915 5015
rect 3709 4981 3743 5015
rect 5457 4981 5491 5015
rect 6377 4981 6411 5015
rect 7297 4981 7331 5015
rect 7573 4981 7607 5015
rect 10333 4981 10367 5015
rect 12541 4981 12575 5015
rect 13369 4981 13403 5015
rect 13553 4981 13587 5015
rect 15209 4981 15243 5015
rect 18061 4981 18095 5015
rect 4169 4777 4203 4811
rect 6285 4777 6319 4811
rect 7481 4777 7515 4811
rect 8953 4777 8987 4811
rect 9781 4777 9815 4811
rect 10609 4777 10643 4811
rect 8769 4709 8803 4743
rect 13093 4709 13127 4743
rect 14933 4709 14967 4743
rect 1961 4641 1995 4675
rect 2513 4641 2547 4675
rect 2605 4641 2639 4675
rect 3341 4641 3375 4675
rect 3525 4641 3559 4675
rect 4721 4641 4755 4675
rect 5733 4641 5767 4675
rect 5825 4641 5859 4675
rect 6469 4641 6503 4675
rect 7757 4641 7791 4675
rect 9597 4641 9631 4675
rect 10333 4641 10367 4675
rect 11161 4641 11195 4675
rect 11989 4641 12023 4675
rect 12541 4641 12575 4675
rect 13645 4641 13679 4675
rect 13737 4641 13771 4675
rect 14289 4641 14323 4675
rect 14473 4641 14507 4675
rect 15209 4641 15243 4675
rect 16497 4641 16531 4675
rect 17233 4641 17267 4675
rect 17693 4641 17727 4675
rect 17785 4641 17819 4675
rect 18797 4641 18831 4675
rect 18889 4641 18923 4675
rect 19441 4641 19475 4675
rect 20729 4641 20763 4675
rect 1501 4573 1535 4607
rect 2421 4573 2455 4607
rect 3985 4573 4019 4607
rect 4997 4573 5031 4607
rect 5641 4573 5675 4607
rect 6745 4573 6779 4607
rect 8585 4573 8619 4607
rect 10149 4573 10183 4607
rect 10241 4573 10275 4607
rect 10977 4573 11011 4607
rect 11805 4573 11839 4607
rect 13553 4573 13587 4607
rect 15301 4573 15335 4607
rect 15393 4573 15427 4607
rect 16221 4573 16255 4607
rect 20361 4573 20395 4607
rect 21005 4573 21039 4607
rect 1685 4505 1719 4539
rect 3249 4505 3283 4539
rect 4537 4505 4571 4539
rect 6193 4505 6227 4539
rect 9321 4505 9355 4539
rect 12633 4505 12667 4539
rect 12725 4505 12759 4539
rect 16313 4505 16347 4539
rect 17049 4505 17083 4539
rect 17877 4505 17911 4539
rect 18705 4505 18739 4539
rect 20545 4505 20579 4539
rect 2053 4437 2087 4471
rect 2881 4437 2915 4471
rect 4629 4437 4663 4471
rect 5181 4437 5215 4471
rect 5273 4437 5307 4471
rect 7849 4437 7883 4471
rect 7941 4437 7975 4471
rect 8309 4437 8343 4471
rect 9413 4437 9447 4471
rect 11069 4437 11103 4471
rect 11437 4437 11471 4471
rect 11897 4437 11931 4471
rect 13185 4437 13219 4471
rect 14565 4437 14599 4471
rect 15761 4437 15795 4471
rect 15853 4437 15887 4471
rect 16681 4437 16715 4471
rect 17141 4437 17175 4471
rect 18245 4437 18279 4471
rect 18337 4437 18371 4471
rect 19533 4437 19567 4471
rect 19625 4437 19659 4471
rect 19993 4437 20027 4471
rect 20085 4437 20119 4471
rect 2237 4233 2271 4267
rect 4169 4233 4203 4267
rect 5457 4233 5491 4267
rect 5825 4233 5859 4267
rect 5917 4233 5951 4267
rect 10977 4233 11011 4267
rect 11805 4233 11839 4267
rect 12541 4233 12575 4267
rect 13369 4233 13403 4267
rect 14289 4233 14323 4267
rect 14749 4233 14783 4267
rect 15209 4233 15243 4267
rect 15945 4233 15979 4267
rect 18337 4233 18371 4267
rect 18797 4233 18831 4267
rect 19257 4233 19291 4267
rect 19625 4233 19659 4267
rect 2329 4165 2363 4199
rect 8953 4165 8987 4199
rect 9045 4165 9079 4199
rect 1409 4097 1443 4131
rect 1869 4097 1903 4131
rect 2789 4097 2823 4131
rect 3056 4097 3090 4131
rect 4261 4097 4295 4131
rect 4997 4097 5031 4131
rect 6377 4097 6411 4131
rect 6653 4097 6687 4131
rect 6837 4097 6871 4131
rect 7288 4097 7322 4131
rect 9597 4097 9631 4131
rect 9873 4097 9907 4131
rect 11621 4097 11655 4131
rect 11897 4097 11931 4131
rect 12173 4097 12207 4131
rect 12633 4097 12667 4131
rect 13461 4097 13495 4131
rect 14197 4097 14231 4131
rect 15117 4097 15151 4131
rect 16681 4097 16715 4131
rect 16957 4097 16991 4131
rect 17224 4097 17258 4131
rect 20269 4097 20303 4131
rect 20545 4097 20579 4131
rect 21005 4097 21039 4131
rect 2145 4029 2179 4063
rect 5089 4029 5123 4063
rect 5273 4029 5307 4063
rect 6009 4029 6043 4063
rect 7021 4029 7055 4063
rect 9229 4029 9263 4063
rect 10241 4029 10275 4063
rect 11069 4029 11103 4063
rect 11161 4029 11195 4063
rect 13185 4029 13219 4063
rect 14105 4029 14139 4063
rect 15301 4029 15335 4063
rect 15761 4029 15795 4063
rect 15853 4029 15887 4063
rect 16405 4029 16439 4063
rect 18521 4029 18555 4063
rect 18705 4029 18739 4063
rect 19717 4029 19751 4063
rect 19809 4029 19843 4063
rect 20729 4029 20763 4063
rect 1685 3961 1719 3995
rect 2697 3961 2731 3995
rect 4445 3961 4479 3995
rect 8401 3961 8435 3995
rect 8585 3961 8619 3995
rect 12817 3961 12851 3995
rect 19165 3961 19199 3995
rect 1593 3893 1627 3927
rect 4629 3893 4663 3927
rect 6561 3893 6595 3927
rect 9505 3893 9539 3927
rect 10609 3893 10643 3927
rect 12081 3893 12115 3927
rect 12357 3893 12391 3927
rect 13001 3893 13035 3927
rect 13829 3893 13863 3927
rect 14657 3893 14691 3927
rect 16313 3893 16347 3927
rect 16865 3893 16899 3927
rect 20085 3893 20119 3927
rect 20361 3893 20395 3927
rect 1869 3689 1903 3723
rect 5181 3689 5215 3723
rect 6377 3689 6411 3723
rect 10517 3689 10551 3723
rect 14105 3689 14139 3723
rect 15577 3689 15611 3723
rect 17969 3689 18003 3723
rect 20453 3689 20487 3723
rect 3341 3621 3375 3655
rect 5549 3621 5583 3655
rect 10609 3621 10643 3655
rect 12265 3621 12299 3655
rect 15117 3621 15151 3655
rect 19349 3621 19383 3655
rect 19625 3621 19659 3655
rect 5825 3553 5859 3587
rect 8125 3553 8159 3587
rect 8309 3553 8343 3587
rect 11989 3553 12023 3587
rect 12173 3553 12207 3587
rect 14565 3553 14599 3587
rect 14657 3553 14691 3587
rect 17325 3553 17359 3587
rect 17509 3553 17543 3587
rect 18153 3553 18187 3587
rect 18337 3553 18371 3587
rect 21005 3553 21039 3587
rect 1409 3485 1443 3519
rect 1685 3485 1719 3519
rect 1961 3485 1995 3519
rect 3433 3485 3467 3519
rect 3801 3485 3835 3519
rect 7849 3485 7883 3519
rect 8953 3485 8987 3519
rect 9209 3485 9243 3519
rect 12449 3485 12483 3519
rect 12541 3485 12575 3519
rect 14933 3485 14967 3519
rect 17049 3485 17083 3519
rect 19073 3485 19107 3519
rect 19533 3485 19567 3519
rect 19809 3485 19843 3519
rect 20085 3485 20119 3519
rect 20361 3485 20395 3519
rect 21465 3485 21499 3519
rect 2228 3417 2262 3451
rect 4068 3417 4102 3451
rect 5365 3417 5399 3451
rect 7582 3417 7616 3451
rect 11744 3417 11778 3451
rect 12808 3417 12842 3451
rect 16804 3417 16838 3451
rect 20821 3417 20855 3451
rect 20913 3417 20947 3451
rect 1593 3349 1627 3383
rect 3617 3349 3651 3383
rect 5917 3349 5951 3383
rect 6009 3349 6043 3383
rect 6469 3349 6503 3383
rect 8401 3349 8435 3383
rect 8769 3349 8803 3383
rect 10333 3349 10367 3383
rect 13921 3349 13955 3383
rect 14473 3349 14507 3383
rect 15209 3349 15243 3383
rect 15669 3349 15703 3383
rect 17601 3349 17635 3383
rect 18429 3349 18463 3383
rect 18797 3349 18831 3383
rect 18889 3349 18923 3383
rect 19901 3349 19935 3383
rect 20177 3349 20211 3383
rect 21373 3349 21407 3383
rect 2421 3145 2455 3179
rect 2513 3145 2547 3179
rect 2973 3145 3007 3179
rect 3433 3145 3467 3179
rect 6469 3145 6503 3179
rect 6929 3145 6963 3179
rect 9413 3145 9447 3179
rect 9873 3145 9907 3179
rect 12817 3145 12851 3179
rect 14289 3145 14323 3179
rect 14749 3145 14783 3179
rect 17693 3145 17727 3179
rect 18153 3145 18187 3179
rect 18521 3145 18555 3179
rect 18981 3145 19015 3179
rect 19441 3145 19475 3179
rect 5080 3077 5114 3111
rect 9321 3077 9355 3111
rect 11989 3077 12023 3111
rect 19349 3077 19383 3111
rect 1593 3009 1627 3043
rect 1869 3009 1903 3043
rect 3341 3009 3375 3043
rect 4629 3009 4663 3043
rect 4813 3009 4847 3043
rect 6837 3009 6871 3043
rect 7665 3009 7699 3043
rect 8493 3009 8527 3043
rect 10221 3009 10255 3043
rect 11897 3009 11931 3043
rect 12357 3009 12391 3043
rect 13941 3009 13975 3043
rect 14657 3009 14691 3043
rect 15393 3009 15427 3043
rect 15577 3009 15611 3043
rect 16129 3009 16163 3043
rect 16405 3009 16439 3043
rect 16865 3009 16899 3043
rect 16957 3009 16991 3043
rect 17417 3009 17451 3043
rect 17509 3009 17543 3043
rect 17785 3009 17819 3043
rect 20085 3009 20119 3043
rect 20453 3009 20487 3043
rect 20545 3009 20579 3043
rect 20913 3009 20947 3043
rect 21281 3009 21315 3043
rect 2329 2941 2363 2975
rect 3617 2941 3651 2975
rect 4353 2941 4387 2975
rect 7113 2941 7147 2975
rect 7389 2941 7423 2975
rect 7573 2941 7607 2975
rect 8585 2941 8619 2975
rect 8769 2941 8803 2975
rect 9597 2941 9631 2975
rect 9965 2941 9999 2975
rect 12173 2941 12207 2975
rect 14197 2941 14231 2975
rect 14841 2941 14875 2975
rect 18613 2941 18647 2975
rect 18705 2941 18739 2975
rect 19533 2941 19567 2975
rect 1501 2873 1535 2907
rect 2881 2873 2915 2907
rect 6193 2873 6227 2907
rect 8033 2873 8067 2907
rect 11529 2873 11563 2907
rect 17141 2873 17175 2907
rect 20269 2873 20303 2907
rect 21097 2873 21131 2907
rect 1777 2805 1811 2839
rect 2053 2805 2087 2839
rect 8125 2805 8159 2839
rect 8953 2805 8987 2839
rect 11345 2805 11379 2839
rect 12541 2805 12575 2839
rect 15209 2805 15243 2839
rect 15761 2805 15795 2839
rect 15945 2805 15979 2839
rect 16221 2805 16255 2839
rect 16681 2805 16715 2839
rect 17233 2805 17267 2839
rect 17969 2805 18003 2839
rect 19901 2805 19935 2839
rect 20729 2805 20763 2839
rect 21465 2805 21499 2839
rect 5641 2601 5675 2635
rect 5825 2601 5859 2635
rect 7481 2601 7515 2635
rect 7665 2601 7699 2635
rect 11713 2601 11747 2635
rect 14841 2601 14875 2635
rect 16773 2601 16807 2635
rect 18705 2601 18739 2635
rect 20453 2601 20487 2635
rect 3617 2533 3651 2567
rect 4169 2533 4203 2567
rect 8677 2533 8711 2567
rect 12357 2533 12391 2567
rect 15025 2533 15059 2567
rect 16129 2533 16163 2567
rect 17141 2533 17175 2567
rect 18245 2533 18279 2567
rect 19257 2533 19291 2567
rect 20269 2533 20303 2567
rect 1961 2465 1995 2499
rect 6929 2465 6963 2499
rect 8033 2465 8067 2499
rect 8217 2465 8251 2499
rect 9505 2465 9539 2499
rect 9873 2465 9907 2499
rect 11161 2465 11195 2499
rect 14197 2465 14231 2499
rect 19809 2465 19843 2499
rect 21005 2465 21039 2499
rect 2237 2397 2271 2431
rect 3157 2397 3191 2431
rect 4261 2397 4295 2431
rect 7205 2397 7239 2431
rect 7297 2397 7331 2431
rect 8309 2397 8343 2431
rect 9413 2397 9447 2431
rect 10977 2397 11011 2431
rect 11621 2397 11655 2431
rect 11897 2397 11931 2431
rect 12541 2397 12575 2431
rect 12909 2397 12943 2431
rect 13001 2397 13035 2431
rect 13369 2397 13403 2431
rect 13921 2397 13955 2431
rect 14473 2397 14507 2431
rect 15209 2397 15243 2431
rect 15301 2397 15335 2431
rect 15669 2397 15703 2431
rect 16313 2397 16347 2431
rect 16957 2397 16991 2431
rect 17325 2397 17359 2431
rect 17693 2397 17727 2431
rect 18061 2397 18095 2431
rect 18429 2397 18463 2431
rect 18521 2397 18555 2431
rect 19073 2397 19107 2431
rect 20085 2397 20119 2431
rect 20637 2397 20671 2431
rect 20729 2397 20763 2431
rect 3433 2329 3467 2363
rect 3985 2329 4019 2363
rect 4506 2329 4540 2363
rect 5917 2329 5951 2363
rect 6101 2329 6135 2363
rect 7757 2329 7791 2363
rect 10149 2329 10183 2363
rect 11069 2329 11103 2363
rect 19625 2329 19659 2363
rect 2927 2261 2961 2295
rect 8953 2261 8987 2295
rect 9321 2261 9355 2295
rect 10057 2261 10091 2295
rect 10517 2261 10551 2295
rect 10609 2261 10643 2295
rect 12081 2261 12115 2295
rect 12725 2261 12759 2295
rect 13185 2261 13219 2295
rect 13553 2261 13587 2295
rect 13737 2261 13771 2295
rect 14381 2261 14415 2295
rect 15485 2261 15519 2295
rect 15853 2261 15887 2295
rect 16405 2261 16439 2295
rect 17509 2261 17543 2295
rect 17877 2261 17911 2295
rect 18889 2261 18923 2295
rect 19717 2261 19751 2295
<< metal1 >>
rect 1026 21224 1032 21276
rect 1084 21264 1090 21276
rect 14642 21264 14648 21276
rect 1084 21236 14648 21264
rect 1084 21224 1090 21236
rect 14642 21224 14648 21236
rect 14700 21224 14706 21276
rect 1210 21156 1216 21208
rect 1268 21196 1274 21208
rect 14274 21196 14280 21208
rect 1268 21168 14280 21196
rect 1268 21156 1274 21168
rect 14274 21156 14280 21168
rect 14332 21156 14338 21208
rect 1578 21088 1584 21140
rect 1636 21128 1642 21140
rect 2038 21128 2044 21140
rect 1636 21100 2044 21128
rect 1636 21088 1642 21100
rect 2038 21088 2044 21100
rect 2096 21088 2102 21140
rect 2406 21088 2412 21140
rect 2464 21128 2470 21140
rect 15930 21128 15936 21140
rect 2464 21100 15936 21128
rect 2464 21088 2470 21100
rect 15930 21088 15936 21100
rect 15988 21088 15994 21140
rect 2038 20952 2044 21004
rect 2096 20992 2102 21004
rect 16114 20992 16120 21004
rect 2096 20964 16120 20992
rect 2096 20952 2102 20964
rect 16114 20952 16120 20964
rect 16172 20952 16178 21004
rect 3878 20884 3884 20936
rect 3936 20924 3942 20936
rect 9122 20924 9128 20936
rect 3936 20896 9128 20924
rect 3936 20884 3942 20896
rect 9122 20884 9128 20896
rect 9180 20884 9186 20936
rect 2746 20828 12434 20856
rect 1946 20748 1952 20800
rect 2004 20788 2010 20800
rect 2746 20788 2774 20828
rect 2004 20760 2774 20788
rect 2004 20748 2010 20760
rect 4062 20748 4068 20800
rect 4120 20788 4126 20800
rect 7374 20788 7380 20800
rect 4120 20760 7380 20788
rect 4120 20748 4126 20760
rect 7374 20748 7380 20760
rect 7432 20748 7438 20800
rect 12406 20788 12434 20828
rect 17678 20788 17684 20800
rect 12406 20760 17684 20788
rect 17678 20748 17684 20760
rect 17736 20748 17742 20800
rect 18046 20748 18052 20800
rect 18104 20788 18110 20800
rect 19702 20788 19708 20800
rect 18104 20760 19708 20788
rect 18104 20748 18110 20760
rect 19702 20748 19708 20760
rect 19760 20748 19766 20800
rect 1104 20698 22056 20720
rect 1104 20646 6148 20698
rect 6200 20646 6212 20698
rect 6264 20646 6276 20698
rect 6328 20646 6340 20698
rect 6392 20646 6404 20698
rect 6456 20646 11346 20698
rect 11398 20646 11410 20698
rect 11462 20646 11474 20698
rect 11526 20646 11538 20698
rect 11590 20646 11602 20698
rect 11654 20646 16544 20698
rect 16596 20646 16608 20698
rect 16660 20646 16672 20698
rect 16724 20646 16736 20698
rect 16788 20646 16800 20698
rect 16852 20646 21742 20698
rect 21794 20646 21806 20698
rect 21858 20646 21870 20698
rect 21922 20646 21934 20698
rect 21986 20646 21998 20698
rect 22050 20646 22056 20698
rect 1104 20624 22056 20646
rect 1854 20584 1860 20596
rect 1815 20556 1860 20584
rect 1854 20544 1860 20556
rect 1912 20544 1918 20596
rect 3878 20584 3884 20596
rect 3839 20556 3884 20584
rect 3878 20544 3884 20556
rect 3936 20544 3942 20596
rect 9766 20584 9772 20596
rect 7668 20556 9772 20584
rect 2866 20516 2872 20528
rect 2827 20488 2872 20516
rect 2866 20476 2872 20488
rect 2924 20476 2930 20528
rect 3605 20519 3663 20525
rect 3605 20485 3617 20519
rect 3651 20516 3663 20519
rect 4154 20516 4160 20528
rect 3651 20488 4160 20516
rect 3651 20485 3663 20488
rect 3605 20479 3663 20485
rect 4154 20476 4160 20488
rect 4212 20476 4218 20528
rect 7668 20525 7696 20556
rect 9766 20544 9772 20556
rect 9824 20544 9830 20596
rect 10321 20587 10379 20593
rect 10321 20553 10333 20587
rect 10367 20584 10379 20587
rect 10870 20584 10876 20596
rect 10367 20556 10876 20584
rect 10367 20553 10379 20556
rect 10321 20547 10379 20553
rect 10870 20544 10876 20556
rect 10928 20544 10934 20596
rect 11698 20544 11704 20596
rect 11756 20584 11762 20596
rect 11885 20587 11943 20593
rect 11885 20584 11897 20587
rect 11756 20556 11897 20584
rect 11756 20544 11762 20556
rect 11885 20553 11897 20556
rect 11931 20553 11943 20587
rect 11885 20547 11943 20553
rect 11974 20544 11980 20596
rect 12032 20584 12038 20596
rect 12253 20587 12311 20593
rect 12253 20584 12265 20587
rect 12032 20556 12265 20584
rect 12032 20544 12038 20556
rect 12253 20553 12265 20556
rect 12299 20553 12311 20587
rect 12253 20547 12311 20553
rect 12434 20544 12440 20596
rect 12492 20584 12498 20596
rect 12621 20587 12679 20593
rect 12621 20584 12633 20587
rect 12492 20556 12633 20584
rect 12492 20544 12498 20556
rect 12621 20553 12633 20556
rect 12667 20553 12679 20587
rect 12621 20547 12679 20553
rect 12710 20544 12716 20596
rect 12768 20584 12774 20596
rect 12897 20587 12955 20593
rect 12897 20584 12909 20587
rect 12768 20556 12909 20584
rect 12768 20544 12774 20556
rect 12897 20553 12909 20556
rect 12943 20553 12955 20587
rect 12897 20547 12955 20553
rect 13078 20544 13084 20596
rect 13136 20584 13142 20596
rect 13357 20587 13415 20593
rect 13357 20584 13369 20587
rect 13136 20556 13369 20584
rect 13136 20544 13142 20556
rect 13357 20553 13369 20556
rect 13403 20553 13415 20587
rect 13357 20547 13415 20553
rect 13446 20544 13452 20596
rect 13504 20584 13510 20596
rect 13633 20587 13691 20593
rect 13633 20584 13645 20587
rect 13504 20556 13645 20584
rect 13504 20544 13510 20556
rect 13633 20553 13645 20556
rect 13679 20553 13691 20587
rect 13633 20547 13691 20553
rect 13814 20544 13820 20596
rect 13872 20584 13878 20596
rect 14185 20587 14243 20593
rect 14185 20584 14197 20587
rect 13872 20556 14197 20584
rect 13872 20544 13878 20556
rect 14185 20553 14197 20556
rect 14231 20553 14243 20587
rect 14185 20547 14243 20553
rect 14550 20544 14556 20596
rect 14608 20584 14614 20596
rect 14921 20587 14979 20593
rect 14921 20584 14933 20587
rect 14608 20556 14933 20584
rect 14608 20544 14614 20556
rect 14921 20553 14933 20556
rect 14967 20553 14979 20587
rect 14921 20547 14979 20553
rect 15194 20544 15200 20596
rect 15252 20584 15258 20596
rect 15289 20587 15347 20593
rect 15289 20584 15301 20587
rect 15252 20556 15301 20584
rect 15252 20544 15258 20556
rect 15289 20553 15301 20556
rect 15335 20553 15347 20587
rect 15289 20547 15347 20553
rect 15378 20544 15384 20596
rect 15436 20584 15442 20596
rect 15657 20587 15715 20593
rect 15657 20584 15669 20587
rect 15436 20556 15669 20584
rect 15436 20544 15442 20556
rect 15657 20553 15669 20556
rect 15703 20553 15715 20587
rect 15657 20547 15715 20553
rect 15746 20544 15752 20596
rect 15804 20584 15810 20596
rect 16025 20587 16083 20593
rect 16025 20584 16037 20587
rect 15804 20556 16037 20584
rect 15804 20544 15810 20556
rect 16025 20553 16037 20556
rect 16071 20553 16083 20587
rect 16025 20547 16083 20553
rect 16574 20544 16580 20596
rect 16632 20584 16638 20596
rect 17129 20587 17187 20593
rect 17129 20584 17141 20587
rect 16632 20556 17141 20584
rect 16632 20544 16638 20556
rect 17129 20553 17141 20556
rect 17175 20553 17187 20587
rect 17129 20547 17187 20553
rect 17494 20544 17500 20596
rect 17552 20584 17558 20596
rect 18325 20587 18383 20593
rect 18325 20584 18337 20587
rect 17552 20556 18337 20584
rect 17552 20544 17558 20556
rect 18325 20553 18337 20556
rect 18371 20553 18383 20587
rect 18325 20547 18383 20553
rect 19061 20587 19119 20593
rect 19061 20553 19073 20587
rect 19107 20553 19119 20587
rect 19518 20584 19524 20596
rect 19479 20556 19524 20584
rect 19061 20547 19119 20553
rect 7653 20519 7711 20525
rect 7392 20488 7604 20516
rect 1673 20451 1731 20457
rect 1673 20417 1685 20451
rect 1719 20448 1731 20451
rect 1946 20448 1952 20460
rect 1719 20420 1952 20448
rect 1719 20417 1731 20420
rect 1673 20411 1731 20417
rect 1946 20408 1952 20420
rect 2004 20408 2010 20460
rect 2038 20408 2044 20460
rect 2096 20448 2102 20460
rect 2317 20451 2375 20457
rect 2096 20420 2141 20448
rect 2096 20408 2102 20420
rect 2317 20417 2329 20451
rect 2363 20448 2375 20451
rect 2590 20448 2596 20460
rect 2363 20420 2596 20448
rect 2363 20417 2375 20420
rect 2317 20411 2375 20417
rect 2590 20408 2596 20420
rect 2648 20408 2654 20460
rect 2682 20408 2688 20460
rect 2740 20448 2746 20460
rect 2740 20420 2785 20448
rect 2740 20408 2746 20420
rect 2958 20408 2964 20460
rect 3016 20448 3022 20460
rect 3053 20451 3111 20457
rect 3053 20448 3065 20451
rect 3016 20420 3065 20448
rect 3016 20408 3022 20420
rect 3053 20417 3065 20420
rect 3099 20417 3111 20451
rect 3053 20411 3111 20417
rect 3326 20408 3332 20460
rect 3384 20448 3390 20460
rect 3421 20451 3479 20457
rect 3421 20448 3433 20451
rect 3384 20420 3433 20448
rect 3384 20408 3390 20420
rect 3421 20417 3433 20420
rect 3467 20417 3479 20451
rect 3421 20411 3479 20417
rect 4240 20451 4298 20457
rect 4240 20417 4252 20451
rect 4286 20448 4298 20451
rect 4706 20448 4712 20460
rect 4286 20420 4712 20448
rect 4286 20417 4298 20420
rect 4240 20411 4298 20417
rect 4706 20408 4712 20420
rect 4764 20408 4770 20460
rect 5813 20451 5871 20457
rect 5813 20417 5825 20451
rect 5859 20448 5871 20451
rect 7098 20448 7104 20460
rect 5859 20420 7104 20448
rect 5859 20417 5871 20420
rect 5813 20411 5871 20417
rect 7098 20408 7104 20420
rect 7156 20408 7162 20460
rect 7193 20451 7251 20457
rect 7193 20417 7205 20451
rect 7239 20448 7251 20451
rect 7282 20448 7288 20460
rect 7239 20420 7288 20448
rect 7239 20417 7251 20420
rect 7193 20411 7251 20417
rect 7282 20408 7288 20420
rect 7340 20408 7346 20460
rect 3970 20380 3976 20392
rect 3931 20352 3976 20380
rect 3970 20340 3976 20352
rect 4028 20340 4034 20392
rect 5902 20380 5908 20392
rect 5863 20352 5908 20380
rect 5902 20340 5908 20352
rect 5960 20340 5966 20392
rect 5997 20383 6055 20389
rect 5997 20349 6009 20383
rect 6043 20349 6055 20383
rect 5997 20343 6055 20349
rect 6917 20383 6975 20389
rect 6917 20349 6929 20383
rect 6963 20380 6975 20383
rect 7392 20380 7420 20488
rect 7469 20451 7527 20457
rect 7469 20417 7481 20451
rect 7515 20417 7527 20451
rect 7576 20448 7604 20488
rect 7653 20485 7665 20519
rect 7699 20485 7711 20519
rect 7653 20479 7711 20485
rect 9033 20519 9091 20525
rect 9033 20485 9045 20519
rect 9079 20516 9091 20519
rect 9079 20488 10548 20516
rect 9079 20485 9091 20488
rect 9033 20479 9091 20485
rect 10520 20460 10548 20488
rect 10594 20476 10600 20528
rect 10652 20516 10658 20528
rect 16298 20516 16304 20528
rect 10652 20488 12480 20516
rect 10652 20476 10658 20488
rect 7576 20420 8616 20448
rect 7469 20411 7527 20417
rect 6963 20352 7420 20380
rect 7484 20380 7512 20411
rect 8386 20380 8392 20392
rect 7484 20352 8392 20380
rect 6963 20349 6975 20352
rect 6917 20343 6975 20349
rect 3237 20315 3295 20321
rect 3237 20281 3249 20315
rect 3283 20312 3295 20315
rect 3418 20312 3424 20324
rect 3283 20284 3424 20312
rect 3283 20281 3295 20284
rect 3237 20275 3295 20281
rect 3418 20272 3424 20284
rect 3476 20272 3482 20324
rect 5445 20315 5503 20321
rect 5445 20312 5457 20315
rect 4908 20284 5457 20312
rect 1486 20244 1492 20256
rect 1447 20216 1492 20244
rect 1486 20204 1492 20216
rect 1544 20204 1550 20256
rect 2130 20204 2136 20256
rect 2188 20244 2194 20256
rect 2409 20247 2467 20253
rect 2409 20244 2421 20247
rect 2188 20216 2421 20244
rect 2188 20204 2194 20216
rect 2409 20213 2421 20216
rect 2455 20213 2467 20247
rect 2409 20207 2467 20213
rect 3878 20204 3884 20256
rect 3936 20244 3942 20256
rect 4908 20244 4936 20284
rect 5445 20281 5457 20284
rect 5491 20281 5503 20315
rect 6012 20312 6040 20343
rect 8386 20340 8392 20352
rect 8444 20340 8450 20392
rect 8481 20383 8539 20389
rect 8481 20349 8493 20383
rect 8527 20349 8539 20383
rect 8588 20380 8616 20420
rect 8662 20408 8668 20460
rect 8720 20448 8726 20460
rect 8757 20451 8815 20457
rect 8757 20448 8769 20451
rect 8720 20420 8769 20448
rect 8720 20408 8726 20420
rect 8757 20417 8769 20420
rect 8803 20417 8815 20451
rect 9122 20448 9128 20460
rect 9083 20420 9128 20448
rect 8757 20411 8815 20417
rect 9122 20408 9128 20420
rect 9180 20408 9186 20460
rect 10134 20448 10140 20460
rect 9324 20420 9996 20448
rect 10095 20420 10140 20448
rect 9324 20380 9352 20420
rect 8588 20352 9352 20380
rect 9401 20383 9459 20389
rect 8481 20343 8539 20349
rect 9401 20349 9413 20383
rect 9447 20380 9459 20383
rect 9490 20380 9496 20392
rect 9447 20352 9496 20380
rect 9447 20349 9459 20352
rect 9401 20343 9459 20349
rect 5445 20275 5503 20281
rect 5828 20284 6040 20312
rect 8496 20312 8524 20343
rect 9490 20340 9496 20352
rect 9548 20340 9554 20392
rect 9968 20380 9996 20420
rect 10134 20408 10140 20420
rect 10192 20408 10198 20460
rect 10502 20448 10508 20460
rect 10463 20420 10508 20448
rect 10502 20408 10508 20420
rect 10560 20408 10566 20460
rect 10686 20408 10692 20460
rect 10744 20448 10750 20460
rect 11701 20451 11759 20457
rect 11701 20448 11713 20451
rect 10744 20420 11713 20448
rect 10744 20408 10750 20420
rect 11701 20417 11713 20420
rect 11747 20417 11759 20451
rect 11701 20411 11759 20417
rect 11790 20408 11796 20460
rect 11848 20448 11854 20460
rect 12452 20457 12480 20488
rect 15120 20488 16304 20516
rect 12069 20451 12127 20457
rect 12069 20448 12081 20451
rect 11848 20420 12081 20448
rect 11848 20408 11854 20420
rect 12069 20417 12081 20420
rect 12115 20417 12127 20451
rect 12069 20411 12127 20417
rect 12437 20451 12495 20457
rect 12437 20417 12449 20451
rect 12483 20417 12495 20451
rect 13078 20448 13084 20460
rect 13039 20420 13084 20448
rect 12437 20411 12495 20417
rect 13078 20408 13084 20420
rect 13136 20408 13142 20460
rect 13173 20451 13231 20457
rect 13173 20417 13185 20451
rect 13219 20417 13231 20451
rect 13173 20411 13231 20417
rect 13817 20451 13875 20457
rect 13817 20417 13829 20451
rect 13863 20417 13875 20451
rect 14366 20448 14372 20460
rect 14327 20420 14372 20448
rect 13817 20411 13875 20417
rect 10410 20380 10416 20392
rect 9968 20352 10416 20380
rect 10410 20340 10416 20352
rect 10468 20340 10474 20392
rect 10778 20380 10784 20392
rect 10739 20352 10784 20380
rect 10778 20340 10784 20352
rect 10836 20340 10842 20392
rect 11882 20340 11888 20392
rect 11940 20380 11946 20392
rect 13188 20380 13216 20411
rect 11940 20352 13216 20380
rect 13832 20380 13860 20411
rect 14366 20408 14372 20420
rect 14424 20408 14430 20460
rect 14734 20448 14740 20460
rect 14695 20420 14740 20448
rect 14734 20408 14740 20420
rect 14792 20408 14798 20460
rect 15120 20457 15148 20488
rect 16298 20476 16304 20488
rect 16356 20476 16362 20528
rect 19076 20516 19104 20547
rect 19518 20544 19524 20556
rect 19576 20544 19582 20596
rect 19978 20584 19984 20596
rect 19939 20556 19984 20584
rect 19978 20544 19984 20556
rect 20036 20544 20042 20596
rect 21174 20544 21180 20596
rect 21232 20584 21238 20596
rect 21453 20587 21511 20593
rect 21453 20584 21465 20587
rect 21232 20556 21465 20584
rect 21232 20544 21238 20556
rect 21453 20553 21465 20556
rect 21499 20553 21511 20587
rect 21453 20547 21511 20553
rect 19076 20488 20208 20516
rect 15105 20451 15163 20457
rect 15105 20417 15117 20451
rect 15151 20417 15163 20451
rect 15470 20448 15476 20460
rect 15431 20420 15476 20448
rect 15105 20411 15163 20417
rect 15470 20408 15476 20420
rect 15528 20408 15534 20460
rect 15838 20448 15844 20460
rect 15799 20420 15844 20448
rect 15838 20408 15844 20420
rect 15896 20408 15902 20460
rect 16206 20448 16212 20460
rect 16167 20420 16212 20448
rect 16206 20408 16212 20420
rect 16264 20408 16270 20460
rect 16485 20451 16543 20457
rect 16485 20417 16497 20451
rect 16531 20417 16543 20451
rect 16485 20411 16543 20417
rect 16669 20451 16727 20457
rect 16669 20417 16681 20451
rect 16715 20448 16727 20451
rect 17034 20448 17040 20460
rect 16715 20420 17040 20448
rect 16715 20417 16727 20420
rect 16669 20411 16727 20417
rect 15562 20380 15568 20392
rect 13832 20352 15568 20380
rect 11940 20340 11946 20352
rect 15562 20340 15568 20352
rect 15620 20340 15626 20392
rect 16500 20380 16528 20411
rect 17034 20408 17040 20420
rect 17092 20408 17098 20460
rect 17126 20408 17132 20460
rect 17184 20448 17190 20460
rect 17313 20451 17371 20457
rect 17313 20448 17325 20451
rect 17184 20420 17325 20448
rect 17184 20408 17190 20420
rect 17313 20417 17325 20420
rect 17359 20417 17371 20451
rect 17313 20411 17371 20417
rect 17402 20408 17408 20460
rect 17460 20448 17466 20460
rect 17460 20420 17505 20448
rect 17460 20408 17466 20420
rect 17586 20408 17592 20460
rect 17644 20448 17650 20460
rect 17773 20451 17831 20457
rect 17773 20448 17785 20451
rect 17644 20420 17785 20448
rect 17644 20408 17650 20420
rect 17773 20417 17785 20420
rect 17819 20417 17831 20451
rect 18138 20448 18144 20460
rect 18099 20420 18144 20448
rect 17773 20411 17831 20417
rect 18138 20408 18144 20420
rect 18196 20408 18202 20460
rect 18322 20408 18328 20460
rect 18380 20448 18386 20460
rect 18509 20451 18567 20457
rect 18509 20448 18521 20451
rect 18380 20420 18521 20448
rect 18380 20408 18386 20420
rect 18509 20417 18521 20420
rect 18555 20417 18567 20451
rect 18509 20411 18567 20417
rect 18877 20451 18935 20457
rect 18877 20417 18889 20451
rect 18923 20417 18935 20451
rect 18877 20411 18935 20417
rect 16500 20352 17908 20380
rect 8496 20284 10180 20312
rect 5350 20244 5356 20256
rect 3936 20216 4936 20244
rect 5311 20216 5356 20244
rect 3936 20204 3942 20216
rect 5350 20204 5356 20216
rect 5408 20204 5414 20256
rect 5534 20204 5540 20256
rect 5592 20244 5598 20256
rect 5828 20244 5856 20284
rect 5592 20216 5856 20244
rect 5592 20204 5598 20216
rect 6822 20204 6828 20256
rect 6880 20244 6886 20256
rect 7285 20247 7343 20253
rect 7285 20244 7297 20247
rect 6880 20216 7297 20244
rect 6880 20204 6886 20216
rect 7285 20213 7297 20216
rect 7331 20213 7343 20247
rect 7742 20244 7748 20256
rect 7703 20216 7748 20244
rect 7285 20207 7343 20213
rect 7742 20204 7748 20216
rect 7800 20204 7806 20256
rect 8294 20204 8300 20256
rect 8352 20244 8358 20256
rect 9306 20244 9312 20256
rect 8352 20216 9312 20244
rect 8352 20204 8358 20216
rect 9306 20204 9312 20216
rect 9364 20204 9370 20256
rect 10152 20244 10180 20284
rect 10226 20272 10232 20324
rect 10284 20312 10290 20324
rect 10962 20312 10968 20324
rect 10284 20284 10968 20312
rect 10284 20272 10290 20284
rect 10962 20272 10968 20284
rect 11020 20312 11026 20324
rect 11517 20315 11575 20321
rect 11517 20312 11529 20315
rect 11020 20284 11529 20312
rect 11020 20272 11026 20284
rect 11517 20281 11529 20284
rect 11563 20281 11575 20315
rect 11517 20275 11575 20281
rect 14182 20272 14188 20324
rect 14240 20312 14246 20324
rect 14553 20315 14611 20321
rect 14553 20312 14565 20315
rect 14240 20284 14565 20312
rect 14240 20272 14246 20284
rect 14553 20281 14565 20284
rect 14599 20281 14611 20315
rect 14553 20275 14611 20281
rect 16022 20272 16028 20324
rect 16080 20312 16086 20324
rect 16853 20315 16911 20321
rect 16853 20312 16865 20315
rect 16080 20284 16865 20312
rect 16080 20272 16086 20284
rect 16853 20281 16865 20284
rect 16899 20281 16911 20315
rect 16853 20275 16911 20281
rect 16942 20272 16948 20324
rect 17000 20312 17006 20324
rect 17589 20315 17647 20321
rect 17589 20312 17601 20315
rect 17000 20284 17601 20312
rect 17000 20272 17006 20284
rect 17589 20281 17601 20284
rect 17635 20281 17647 20315
rect 17880 20312 17908 20352
rect 17954 20340 17960 20392
rect 18012 20380 18018 20392
rect 18892 20380 18920 20411
rect 18966 20408 18972 20460
rect 19024 20448 19030 20460
rect 19337 20451 19395 20457
rect 19337 20448 19349 20451
rect 19024 20420 19349 20448
rect 19024 20408 19030 20420
rect 19337 20417 19349 20420
rect 19383 20417 19395 20451
rect 19702 20448 19708 20460
rect 19663 20420 19708 20448
rect 19337 20411 19395 20417
rect 19702 20408 19708 20420
rect 19760 20408 19766 20460
rect 19794 20408 19800 20460
rect 19852 20448 19858 20460
rect 20180 20457 20208 20488
rect 20165 20451 20223 20457
rect 19852 20420 19897 20448
rect 19852 20408 19858 20420
rect 20165 20417 20177 20451
rect 20211 20417 20223 20451
rect 20165 20411 20223 20417
rect 20533 20451 20591 20457
rect 20533 20417 20545 20451
rect 20579 20417 20591 20451
rect 20533 20411 20591 20417
rect 19058 20380 19064 20392
rect 18012 20352 18736 20380
rect 18892 20352 19064 20380
rect 18012 20340 18018 20352
rect 18708 20321 18736 20352
rect 19058 20340 19064 20352
rect 19116 20340 19122 20392
rect 18693 20315 18751 20321
rect 17880 20284 18644 20312
rect 17589 20275 17647 20281
rect 11146 20244 11152 20256
rect 10152 20216 11152 20244
rect 11146 20204 11152 20216
rect 11204 20204 11210 20256
rect 13814 20204 13820 20256
rect 13872 20244 13878 20256
rect 15654 20244 15660 20256
rect 13872 20216 15660 20244
rect 13872 20204 13878 20216
rect 15654 20204 15660 20216
rect 15712 20204 15718 20256
rect 16114 20204 16120 20256
rect 16172 20244 16178 20256
rect 16301 20247 16359 20253
rect 16301 20244 16313 20247
rect 16172 20216 16313 20244
rect 16172 20204 16178 20216
rect 16301 20213 16313 20216
rect 16347 20213 16359 20247
rect 16301 20207 16359 20213
rect 17218 20204 17224 20256
rect 17276 20244 17282 20256
rect 17957 20247 18015 20253
rect 17957 20244 17969 20247
rect 17276 20216 17969 20244
rect 17276 20204 17282 20216
rect 17957 20213 17969 20216
rect 18003 20213 18015 20247
rect 18616 20244 18644 20284
rect 18693 20281 18705 20315
rect 18739 20281 18751 20315
rect 18693 20275 18751 20281
rect 18874 20272 18880 20324
rect 18932 20312 18938 20324
rect 20548 20312 20576 20411
rect 20714 20408 20720 20460
rect 20772 20448 20778 20460
rect 20901 20451 20959 20457
rect 20901 20448 20913 20451
rect 20772 20420 20913 20448
rect 20772 20408 20778 20420
rect 20901 20417 20913 20420
rect 20947 20417 20959 20451
rect 20901 20411 20959 20417
rect 21269 20451 21327 20457
rect 21269 20417 21281 20451
rect 21315 20448 21327 20451
rect 21358 20448 21364 20460
rect 21315 20420 21364 20448
rect 21315 20417 21327 20420
rect 21269 20411 21327 20417
rect 21358 20408 21364 20420
rect 21416 20408 21422 20460
rect 18932 20284 20576 20312
rect 20717 20315 20775 20321
rect 18932 20272 18938 20284
rect 20717 20281 20729 20315
rect 20763 20312 20775 20315
rect 21542 20312 21548 20324
rect 20763 20284 21548 20312
rect 20763 20281 20775 20284
rect 20717 20275 20775 20281
rect 21542 20272 21548 20284
rect 21600 20272 21606 20324
rect 20162 20244 20168 20256
rect 18616 20216 20168 20244
rect 17957 20207 18015 20213
rect 20162 20204 20168 20216
rect 20220 20204 20226 20256
rect 20346 20244 20352 20256
rect 20307 20216 20352 20244
rect 20346 20204 20352 20216
rect 20404 20204 20410 20256
rect 21082 20244 21088 20256
rect 21043 20216 21088 20244
rect 21082 20204 21088 20216
rect 21140 20204 21146 20256
rect 1104 20154 21896 20176
rect 1104 20102 3549 20154
rect 3601 20102 3613 20154
rect 3665 20102 3677 20154
rect 3729 20102 3741 20154
rect 3793 20102 3805 20154
rect 3857 20102 8747 20154
rect 8799 20102 8811 20154
rect 8863 20102 8875 20154
rect 8927 20102 8939 20154
rect 8991 20102 9003 20154
rect 9055 20102 13945 20154
rect 13997 20102 14009 20154
rect 14061 20102 14073 20154
rect 14125 20102 14137 20154
rect 14189 20102 14201 20154
rect 14253 20102 19143 20154
rect 19195 20102 19207 20154
rect 19259 20102 19271 20154
rect 19323 20102 19335 20154
rect 19387 20102 19399 20154
rect 19451 20102 21896 20154
rect 1104 20080 21896 20102
rect 2222 20040 2228 20052
rect 2183 20012 2228 20040
rect 2222 20000 2228 20012
rect 2280 20000 2286 20052
rect 2314 20000 2320 20052
rect 2372 20040 2378 20052
rect 2593 20043 2651 20049
rect 2593 20040 2605 20043
rect 2372 20012 2605 20040
rect 2372 20000 2378 20012
rect 2593 20009 2605 20012
rect 2639 20009 2651 20043
rect 6365 20043 6423 20049
rect 6365 20040 6377 20043
rect 2593 20003 2651 20009
rect 3068 20012 6377 20040
rect 3068 19913 3096 20012
rect 6365 20009 6377 20012
rect 6411 20009 6423 20043
rect 6365 20003 6423 20009
rect 3053 19907 3111 19913
rect 3053 19873 3065 19907
rect 3099 19873 3111 19907
rect 3053 19867 3111 19873
rect 4246 19864 4252 19916
rect 4304 19904 4310 19916
rect 4890 19904 4896 19916
rect 4304 19876 4896 19904
rect 4304 19864 4310 19876
rect 4890 19864 4896 19876
rect 4948 19864 4954 19916
rect 6380 19904 6408 20003
rect 6730 20000 6736 20052
rect 6788 20040 6794 20052
rect 7926 20040 7932 20052
rect 6788 20012 7932 20040
rect 6788 20000 6794 20012
rect 7926 20000 7932 20012
rect 7984 20040 7990 20052
rect 7984 20012 9904 20040
rect 7984 20000 7990 20012
rect 9876 19972 9904 20012
rect 11238 20000 11244 20052
rect 11296 20040 11302 20052
rect 11517 20043 11575 20049
rect 11517 20040 11529 20043
rect 11296 20012 11529 20040
rect 11296 20000 11302 20012
rect 11517 20009 11529 20012
rect 11563 20009 11575 20043
rect 11517 20003 11575 20009
rect 12253 20043 12311 20049
rect 12253 20009 12265 20043
rect 12299 20040 12311 20043
rect 15473 20043 15531 20049
rect 12299 20012 15424 20040
rect 12299 20009 12311 20012
rect 12253 20003 12311 20009
rect 12434 19972 12440 19984
rect 9876 19944 12440 19972
rect 12434 19932 12440 19944
rect 12492 19932 12498 19984
rect 14366 19932 14372 19984
rect 14424 19972 14430 19984
rect 15197 19975 15255 19981
rect 15197 19972 15209 19975
rect 14424 19944 15209 19972
rect 14424 19932 14430 19944
rect 15197 19941 15209 19944
rect 15243 19941 15255 19975
rect 15197 19935 15255 19941
rect 8294 19904 8300 19916
rect 6380 19876 6960 19904
rect 1673 19839 1731 19845
rect 1673 19805 1685 19839
rect 1719 19836 1731 19839
rect 1946 19836 1952 19848
rect 1719 19808 1952 19836
rect 1719 19805 1731 19808
rect 1673 19799 1731 19805
rect 1946 19796 1952 19808
rect 2004 19796 2010 19848
rect 2041 19839 2099 19845
rect 2041 19805 2053 19839
rect 2087 19836 2099 19839
rect 2314 19836 2320 19848
rect 2087 19808 2320 19836
rect 2087 19805 2099 19808
rect 2041 19799 2099 19805
rect 2314 19796 2320 19808
rect 2372 19796 2378 19848
rect 2406 19796 2412 19848
rect 2464 19836 2470 19848
rect 2777 19839 2835 19845
rect 2464 19808 2509 19836
rect 2464 19796 2470 19808
rect 2777 19805 2789 19839
rect 2823 19836 2835 19839
rect 3142 19836 3148 19848
rect 2823 19808 3148 19836
rect 2823 19805 2835 19808
rect 2777 19799 2835 19805
rect 3142 19796 3148 19808
rect 3200 19796 3206 19848
rect 3237 19839 3295 19845
rect 3237 19805 3249 19839
rect 3283 19836 3295 19839
rect 3878 19836 3884 19848
rect 3283 19808 3884 19836
rect 3283 19805 3295 19808
rect 3237 19799 3295 19805
rect 3878 19796 3884 19808
rect 3936 19796 3942 19848
rect 4341 19839 4399 19845
rect 4341 19805 4353 19839
rect 4387 19805 4399 19839
rect 4614 19836 4620 19848
rect 4575 19808 4620 19836
rect 4341 19799 4399 19805
rect 3050 19728 3056 19780
rect 3108 19768 3114 19780
rect 4246 19768 4252 19780
rect 3108 19740 4252 19768
rect 3108 19728 3114 19740
rect 4246 19728 4252 19740
rect 4304 19728 4310 19780
rect 1486 19700 1492 19712
rect 1447 19672 1492 19700
rect 1486 19660 1492 19672
rect 1544 19660 1550 19712
rect 1854 19700 1860 19712
rect 1815 19672 1860 19700
rect 1854 19660 1860 19672
rect 1912 19660 1918 19712
rect 3142 19700 3148 19712
rect 3103 19672 3148 19700
rect 3142 19660 3148 19672
rect 3200 19660 3206 19712
rect 3605 19703 3663 19709
rect 3605 19669 3617 19703
rect 3651 19700 3663 19703
rect 4062 19700 4068 19712
rect 3651 19672 4068 19700
rect 3651 19669 3663 19672
rect 3605 19663 3663 19669
rect 4062 19660 4068 19672
rect 4120 19660 4126 19712
rect 4356 19700 4384 19799
rect 4614 19796 4620 19808
rect 4672 19796 4678 19848
rect 4709 19839 4767 19845
rect 4709 19805 4721 19839
rect 4755 19805 4767 19839
rect 4709 19799 4767 19805
rect 4430 19728 4436 19780
rect 4488 19768 4494 19780
rect 4724 19768 4752 19799
rect 4798 19796 4804 19848
rect 4856 19836 4862 19848
rect 4985 19839 5043 19845
rect 4985 19836 4997 19839
rect 4856 19808 4997 19836
rect 4856 19796 4862 19808
rect 4985 19805 4997 19808
rect 5031 19836 5043 19839
rect 6822 19836 6828 19848
rect 5031 19808 6828 19836
rect 5031 19805 5043 19808
rect 4985 19799 5043 19805
rect 6822 19796 6828 19808
rect 6880 19796 6886 19848
rect 6932 19836 6960 19876
rect 7944 19876 8300 19904
rect 7081 19839 7139 19845
rect 7081 19836 7093 19839
rect 6932 19808 7093 19836
rect 7081 19805 7093 19808
rect 7127 19836 7139 19839
rect 7466 19836 7472 19848
rect 7127 19808 7472 19836
rect 7127 19805 7139 19808
rect 7081 19799 7139 19805
rect 7466 19796 7472 19808
rect 7524 19796 7530 19848
rect 5230 19771 5288 19777
rect 5230 19768 5242 19771
rect 4488 19740 5242 19768
rect 4488 19728 4494 19740
rect 5230 19737 5242 19740
rect 5276 19768 5288 19771
rect 5442 19768 5448 19780
rect 5276 19740 5448 19768
rect 5276 19737 5288 19740
rect 5230 19731 5288 19737
rect 5442 19728 5448 19740
rect 5500 19728 5506 19780
rect 5718 19728 5724 19780
rect 5776 19768 5782 19780
rect 6457 19771 6515 19777
rect 6457 19768 6469 19771
rect 5776 19740 6469 19768
rect 5776 19728 5782 19740
rect 6457 19737 6469 19740
rect 6503 19737 6515 19771
rect 6457 19731 6515 19737
rect 6641 19771 6699 19777
rect 6641 19737 6653 19771
rect 6687 19768 6699 19771
rect 7944 19768 7972 19876
rect 8294 19864 8300 19876
rect 8352 19864 8358 19916
rect 8386 19864 8392 19916
rect 8444 19904 8450 19916
rect 8941 19907 8999 19913
rect 8941 19904 8953 19907
rect 8444 19876 8953 19904
rect 8444 19864 8450 19876
rect 8941 19873 8953 19876
rect 8987 19873 8999 19907
rect 11054 19904 11060 19916
rect 8941 19867 8999 19873
rect 10244 19876 11060 19904
rect 8956 19836 8984 19867
rect 10244 19836 10272 19876
rect 11054 19864 11060 19876
rect 11112 19864 11118 19916
rect 13725 19907 13783 19913
rect 13725 19873 13737 19907
rect 13771 19904 13783 19907
rect 13771 19876 15056 19904
rect 13771 19873 13783 19876
rect 13725 19867 13783 19873
rect 10505 19839 10563 19845
rect 10505 19836 10517 19839
rect 6687 19740 7972 19768
rect 8220 19808 8800 19836
rect 8956 19808 10272 19836
rect 10336 19808 10517 19836
rect 6687 19737 6699 19740
rect 6641 19731 6699 19737
rect 4522 19700 4528 19712
rect 4356 19672 4528 19700
rect 4522 19660 4528 19672
rect 4580 19660 4586 19712
rect 4893 19703 4951 19709
rect 4893 19669 4905 19703
rect 4939 19700 4951 19703
rect 5074 19700 5080 19712
rect 4939 19672 5080 19700
rect 4939 19669 4951 19672
rect 4893 19663 4951 19669
rect 5074 19660 5080 19672
rect 5132 19660 5138 19712
rect 7742 19660 7748 19712
rect 7800 19700 7806 19712
rect 8220 19709 8248 19808
rect 8386 19728 8392 19780
rect 8444 19768 8450 19780
rect 8665 19771 8723 19777
rect 8665 19768 8677 19771
rect 8444 19740 8677 19768
rect 8444 19728 8450 19740
rect 8665 19737 8677 19740
rect 8711 19737 8723 19771
rect 8772 19768 8800 19808
rect 9186 19771 9244 19777
rect 9186 19768 9198 19771
rect 8772 19740 9198 19768
rect 8665 19731 8723 19737
rect 9186 19737 9198 19740
rect 9232 19737 9244 19771
rect 9186 19731 9244 19737
rect 8205 19703 8263 19709
rect 8205 19700 8217 19703
rect 7800 19672 8217 19700
rect 7800 19660 7806 19672
rect 8205 19669 8217 19672
rect 8251 19669 8263 19703
rect 8205 19663 8263 19669
rect 8294 19660 8300 19712
rect 8352 19700 8358 19712
rect 8570 19700 8576 19712
rect 8352 19672 8397 19700
rect 8531 19672 8576 19700
rect 8352 19660 8358 19672
rect 8570 19660 8576 19672
rect 8628 19660 8634 19712
rect 8754 19660 8760 19712
rect 8812 19700 8818 19712
rect 10336 19709 10364 19808
rect 10505 19805 10517 19808
rect 10551 19836 10563 19839
rect 10870 19836 10876 19848
rect 10551 19808 10876 19836
rect 10551 19805 10563 19808
rect 10505 19799 10563 19805
rect 10870 19796 10876 19808
rect 10928 19796 10934 19848
rect 11238 19796 11244 19848
rect 11296 19836 11302 19848
rect 11333 19839 11391 19845
rect 11333 19836 11345 19839
rect 11296 19808 11345 19836
rect 11296 19796 11302 19808
rect 11333 19805 11345 19808
rect 11379 19805 11391 19839
rect 11333 19799 11391 19805
rect 12069 19839 12127 19845
rect 12069 19805 12081 19839
rect 12115 19836 12127 19839
rect 12986 19836 12992 19848
rect 12115 19808 12992 19836
rect 12115 19805 12127 19808
rect 12069 19799 12127 19805
rect 12986 19796 12992 19808
rect 13044 19796 13050 19848
rect 14182 19836 14188 19848
rect 13556 19808 14188 19836
rect 10962 19728 10968 19780
rect 11020 19768 11026 19780
rect 11793 19771 11851 19777
rect 11793 19768 11805 19771
rect 11020 19740 11805 19768
rect 11020 19728 11026 19740
rect 11793 19737 11805 19740
rect 11839 19737 11851 19771
rect 11793 19731 11851 19737
rect 13170 19728 13176 19780
rect 13228 19768 13234 19780
rect 13458 19771 13516 19777
rect 13458 19768 13470 19771
rect 13228 19740 13470 19768
rect 13228 19728 13234 19740
rect 13458 19737 13470 19740
rect 13504 19737 13516 19771
rect 13458 19731 13516 19737
rect 13556 19712 13584 19808
rect 14182 19796 14188 19808
rect 14240 19836 14246 19848
rect 14553 19839 14611 19845
rect 14553 19836 14565 19839
rect 14240 19808 14565 19836
rect 14240 19796 14246 19808
rect 14553 19805 14565 19808
rect 14599 19805 14611 19839
rect 15028 19836 15056 19876
rect 15396 19861 15424 20012
rect 15473 20009 15485 20043
rect 15519 20040 15531 20043
rect 15562 20040 15568 20052
rect 15519 20012 15568 20040
rect 15519 20009 15531 20012
rect 15473 20003 15531 20009
rect 15562 20000 15568 20012
rect 15620 20000 15626 20052
rect 16206 20000 16212 20052
rect 16264 20040 16270 20052
rect 16853 20043 16911 20049
rect 16853 20040 16865 20043
rect 16264 20012 16865 20040
rect 16264 20000 16270 20012
rect 16853 20009 16865 20012
rect 16899 20009 16911 20043
rect 17126 20040 17132 20052
rect 17087 20012 17132 20040
rect 16853 20003 16911 20009
rect 17126 20000 17132 20012
rect 17184 20000 17190 20052
rect 17586 20040 17592 20052
rect 17547 20012 17592 20040
rect 17586 20000 17592 20012
rect 17644 20000 17650 20052
rect 17678 20000 17684 20052
rect 17736 20040 17742 20052
rect 17736 20012 17781 20040
rect 17736 20000 17742 20012
rect 18230 20000 18236 20052
rect 18288 20040 18294 20052
rect 18417 20043 18475 20049
rect 18417 20040 18429 20043
rect 18288 20012 18429 20040
rect 18288 20000 18294 20012
rect 18417 20009 18429 20012
rect 18463 20009 18475 20043
rect 18417 20003 18475 20009
rect 18690 20000 18696 20052
rect 18748 20040 18754 20052
rect 19334 20040 19340 20052
rect 18748 20012 19340 20040
rect 18748 20000 18754 20012
rect 19334 20000 19340 20012
rect 19392 20040 19398 20052
rect 20070 20040 20076 20052
rect 19392 20012 20076 20040
rect 19392 20000 19398 20012
rect 20070 20000 20076 20012
rect 20128 20000 20134 20052
rect 15838 19932 15844 19984
rect 15896 19972 15902 19984
rect 16577 19975 16635 19981
rect 16577 19972 16589 19975
rect 15896 19944 16589 19972
rect 15896 19932 15902 19944
rect 16577 19941 16589 19944
rect 16623 19941 16635 19975
rect 17954 19972 17960 19984
rect 17915 19944 17960 19972
rect 16577 19935 16635 19941
rect 17954 19932 17960 19944
rect 18012 19932 18018 19984
rect 18782 19932 18788 19984
rect 18840 19972 18846 19984
rect 18877 19975 18935 19981
rect 18877 19972 18889 19975
rect 18840 19944 18889 19972
rect 18840 19932 18846 19944
rect 18877 19941 18889 19944
rect 18923 19941 18935 19975
rect 18877 19935 18935 19941
rect 19058 19932 19064 19984
rect 19116 19932 19122 19984
rect 15746 19864 15752 19916
rect 15804 19904 15810 19916
rect 16390 19904 16396 19916
rect 15804 19876 16396 19904
rect 15804 19864 15810 19876
rect 15381 19855 15439 19861
rect 15105 19839 15163 19845
rect 15105 19836 15117 19839
rect 15028 19808 15117 19836
rect 14553 19799 14611 19805
rect 15105 19805 15117 19808
rect 15151 19805 15163 19839
rect 15381 19821 15393 19855
rect 15427 19821 15439 19855
rect 15654 19836 15660 19848
rect 15381 19815 15439 19821
rect 15615 19808 15660 19836
rect 15105 19799 15163 19805
rect 15120 19768 15148 19799
rect 15654 19796 15660 19808
rect 15712 19796 15718 19848
rect 16224 19845 16252 19876
rect 16390 19864 16396 19876
rect 16448 19864 16454 19916
rect 17678 19904 17684 19916
rect 17328 19876 17684 19904
rect 15933 19839 15991 19845
rect 15933 19805 15945 19839
rect 15979 19805 15991 19839
rect 15933 19799 15991 19805
rect 16209 19839 16267 19845
rect 16209 19805 16221 19839
rect 16255 19805 16267 19839
rect 16209 19799 16267 19805
rect 16485 19839 16543 19845
rect 16485 19805 16497 19839
rect 16531 19805 16543 19839
rect 16485 19799 16543 19805
rect 16761 19839 16819 19845
rect 16761 19805 16773 19839
rect 16807 19836 16819 19839
rect 16942 19836 16948 19848
rect 16807 19808 16948 19836
rect 16807 19805 16819 19808
rect 16761 19799 16819 19805
rect 15948 19768 15976 19799
rect 15120 19740 16068 19768
rect 10321 19703 10379 19709
rect 10321 19700 10333 19703
rect 8812 19672 10333 19700
rect 8812 19660 8818 19672
rect 10321 19669 10333 19672
rect 10367 19669 10379 19703
rect 10321 19663 10379 19669
rect 11698 19660 11704 19712
rect 11756 19700 11762 19712
rect 11885 19703 11943 19709
rect 11885 19700 11897 19703
rect 11756 19672 11897 19700
rect 11756 19660 11762 19672
rect 11885 19669 11897 19672
rect 11931 19669 11943 19703
rect 11885 19663 11943 19669
rect 12345 19703 12403 19709
rect 12345 19669 12357 19703
rect 12391 19700 12403 19703
rect 13538 19700 13544 19712
rect 12391 19672 13544 19700
rect 12391 19669 12403 19672
rect 12345 19663 12403 19669
rect 13538 19660 13544 19672
rect 13596 19660 13602 19712
rect 13814 19700 13820 19712
rect 13775 19672 13820 19700
rect 13814 19660 13820 19672
rect 13872 19660 13878 19712
rect 13906 19660 13912 19712
rect 13964 19700 13970 19712
rect 14921 19703 14979 19709
rect 14921 19700 14933 19703
rect 13964 19672 14933 19700
rect 13964 19660 13970 19672
rect 14921 19669 14933 19672
rect 14967 19669 14979 19703
rect 14921 19663 14979 19669
rect 15194 19660 15200 19712
rect 15252 19700 15258 19712
rect 16040 19709 16068 19740
rect 16390 19728 16396 19780
rect 16448 19768 16454 19780
rect 16500 19768 16528 19799
rect 16942 19796 16948 19808
rect 17000 19796 17006 19848
rect 17037 19839 17095 19845
rect 17037 19805 17049 19839
rect 17083 19836 17095 19839
rect 17218 19836 17224 19848
rect 17083 19808 17224 19836
rect 17083 19805 17095 19808
rect 17037 19799 17095 19805
rect 17218 19796 17224 19808
rect 17276 19796 17282 19848
rect 17328 19845 17356 19876
rect 17678 19864 17684 19876
rect 17736 19864 17742 19916
rect 19076 19904 19104 19932
rect 19610 19904 19616 19916
rect 17880 19876 19104 19904
rect 19571 19876 19616 19904
rect 17880 19845 17908 19876
rect 19610 19864 19616 19876
rect 19668 19904 19674 19916
rect 20254 19904 20260 19916
rect 19668 19876 20116 19904
rect 20215 19876 20260 19904
rect 19668 19864 19674 19876
rect 17313 19839 17371 19845
rect 17313 19805 17325 19839
rect 17359 19805 17371 19839
rect 17313 19799 17371 19805
rect 17405 19839 17463 19845
rect 17405 19805 17417 19839
rect 17451 19805 17463 19839
rect 17405 19799 17463 19805
rect 17865 19839 17923 19845
rect 17865 19805 17877 19839
rect 17911 19805 17923 19839
rect 17865 19799 17923 19805
rect 18141 19839 18199 19845
rect 18141 19805 18153 19839
rect 18187 19836 18199 19839
rect 18414 19836 18420 19848
rect 18187 19808 18420 19836
rect 18187 19805 18199 19808
rect 18141 19799 18199 19805
rect 16448 19740 16528 19768
rect 16448 19728 16454 19740
rect 17126 19728 17132 19780
rect 17184 19768 17190 19780
rect 17420 19768 17448 19799
rect 18414 19796 18420 19808
rect 18472 19796 18478 19848
rect 18601 19839 18659 19845
rect 18601 19805 18613 19839
rect 18647 19836 18659 19839
rect 18782 19836 18788 19848
rect 18647 19808 18788 19836
rect 18647 19805 18659 19808
rect 18601 19799 18659 19805
rect 18782 19796 18788 19808
rect 18840 19796 18846 19848
rect 19061 19839 19119 19845
rect 19061 19805 19073 19839
rect 19107 19805 19119 19839
rect 19061 19799 19119 19805
rect 19337 19839 19395 19845
rect 19337 19805 19349 19839
rect 19383 19836 19395 19839
rect 19518 19836 19524 19848
rect 19383 19808 19524 19836
rect 19383 19805 19395 19808
rect 19337 19799 19395 19805
rect 17184 19740 17448 19768
rect 19076 19768 19104 19799
rect 19518 19796 19524 19808
rect 19576 19796 19582 19848
rect 19610 19768 19616 19780
rect 19076 19740 19616 19768
rect 17184 19728 17190 19740
rect 19610 19728 19616 19740
rect 19668 19728 19674 19780
rect 20088 19768 20116 19876
rect 20254 19864 20260 19876
rect 20312 19864 20318 19916
rect 20438 19796 20444 19848
rect 20496 19836 20502 19848
rect 20533 19839 20591 19845
rect 20533 19836 20545 19839
rect 20496 19808 20545 19836
rect 20496 19796 20502 19808
rect 20533 19805 20545 19808
rect 20579 19836 20591 19839
rect 20717 19839 20775 19845
rect 20717 19836 20729 19839
rect 20579 19808 20729 19836
rect 20579 19805 20591 19808
rect 20533 19799 20591 19805
rect 20717 19805 20729 19808
rect 20763 19805 20775 19839
rect 20717 19799 20775 19805
rect 21174 19796 21180 19848
rect 21232 19836 21238 19848
rect 21269 19839 21327 19845
rect 21269 19836 21281 19839
rect 21232 19808 21281 19836
rect 21232 19796 21238 19808
rect 21269 19805 21281 19808
rect 21315 19805 21327 19839
rect 21269 19799 21327 19805
rect 20254 19768 20260 19780
rect 20088 19740 20260 19768
rect 20254 19728 20260 19740
rect 20312 19728 20318 19780
rect 20806 19728 20812 19780
rect 20864 19768 20870 19780
rect 20993 19771 21051 19777
rect 20993 19768 21005 19771
rect 20864 19740 21005 19768
rect 20864 19728 20870 19740
rect 20993 19737 21005 19740
rect 21039 19737 21051 19771
rect 20993 19731 21051 19737
rect 15749 19703 15807 19709
rect 15749 19700 15761 19703
rect 15252 19672 15761 19700
rect 15252 19660 15258 19672
rect 15749 19669 15761 19672
rect 15795 19669 15807 19703
rect 15749 19663 15807 19669
rect 16025 19703 16083 19709
rect 16025 19669 16037 19703
rect 16071 19669 16083 19703
rect 16298 19700 16304 19712
rect 16259 19672 16304 19700
rect 16025 19663 16083 19669
rect 16298 19660 16304 19672
rect 16356 19660 16362 19712
rect 21453 19703 21511 19709
rect 21453 19669 21465 19703
rect 21499 19700 21511 19703
rect 21542 19700 21548 19712
rect 21499 19672 21548 19700
rect 21499 19669 21511 19672
rect 21453 19663 21511 19669
rect 21542 19660 21548 19672
rect 21600 19660 21606 19712
rect 1104 19610 22056 19632
rect 1104 19558 6148 19610
rect 6200 19558 6212 19610
rect 6264 19558 6276 19610
rect 6328 19558 6340 19610
rect 6392 19558 6404 19610
rect 6456 19558 11346 19610
rect 11398 19558 11410 19610
rect 11462 19558 11474 19610
rect 11526 19558 11538 19610
rect 11590 19558 11602 19610
rect 11654 19558 16544 19610
rect 16596 19558 16608 19610
rect 16660 19558 16672 19610
rect 16724 19558 16736 19610
rect 16788 19558 16800 19610
rect 16852 19558 21742 19610
rect 21794 19558 21806 19610
rect 21858 19558 21870 19610
rect 21922 19558 21934 19610
rect 21986 19558 21998 19610
rect 22050 19558 22056 19610
rect 1104 19536 22056 19558
rect 1762 19456 1768 19508
rect 1820 19496 1826 19508
rect 1857 19499 1915 19505
rect 1857 19496 1869 19499
rect 1820 19468 1869 19496
rect 1820 19456 1826 19468
rect 1857 19465 1869 19468
rect 1903 19465 1915 19499
rect 3421 19499 3479 19505
rect 3421 19496 3433 19499
rect 1857 19459 1915 19465
rect 2608 19468 3433 19496
rect 14 19388 20 19440
rect 72 19428 78 19440
rect 934 19428 940 19440
rect 72 19400 940 19428
rect 72 19388 78 19400
rect 934 19388 940 19400
rect 992 19388 998 19440
rect 1394 19320 1400 19372
rect 1452 19360 1458 19372
rect 1673 19363 1731 19369
rect 1673 19360 1685 19363
rect 1452 19332 1685 19360
rect 1452 19320 1458 19332
rect 1673 19329 1685 19332
rect 1719 19329 1731 19363
rect 2038 19360 2044 19372
rect 1999 19332 2044 19360
rect 1673 19323 1731 19329
rect 2038 19320 2044 19332
rect 2096 19320 2102 19372
rect 2130 19320 2136 19372
rect 2188 19360 2194 19372
rect 2608 19360 2636 19468
rect 3421 19465 3433 19468
rect 3467 19496 3479 19499
rect 4249 19499 4307 19505
rect 4249 19496 4261 19499
rect 3467 19468 4261 19496
rect 3467 19465 3479 19468
rect 3421 19459 3479 19465
rect 4249 19465 4261 19468
rect 4295 19465 4307 19499
rect 4249 19459 4307 19465
rect 4709 19499 4767 19505
rect 4709 19465 4721 19499
rect 4755 19496 4767 19499
rect 4755 19468 5488 19496
rect 4755 19465 4767 19468
rect 4709 19459 4767 19465
rect 2685 19431 2743 19437
rect 2685 19397 2697 19431
rect 2731 19428 2743 19431
rect 3050 19428 3056 19440
rect 2731 19400 3056 19428
rect 2731 19397 2743 19400
rect 2685 19391 2743 19397
rect 3050 19388 3056 19400
rect 3108 19388 3114 19440
rect 5068 19431 5126 19437
rect 5068 19428 5080 19431
rect 3344 19400 5080 19428
rect 2188 19332 2636 19360
rect 2188 19320 2194 19332
rect 2608 19301 2636 19332
rect 3344 19301 3372 19400
rect 5068 19397 5080 19400
rect 5114 19428 5126 19431
rect 5350 19428 5356 19440
rect 5114 19400 5356 19428
rect 5114 19397 5126 19400
rect 5068 19391 5126 19397
rect 5350 19388 5356 19400
rect 5408 19388 5414 19440
rect 5460 19428 5488 19468
rect 5534 19456 5540 19508
rect 5592 19496 5598 19508
rect 6181 19499 6239 19505
rect 6181 19496 6193 19499
rect 5592 19468 6193 19496
rect 5592 19456 5598 19468
rect 6181 19465 6193 19468
rect 6227 19465 6239 19499
rect 8202 19496 8208 19508
rect 6181 19459 6239 19465
rect 6564 19468 8208 19496
rect 6564 19428 6592 19468
rect 8202 19456 8208 19468
rect 8260 19456 8266 19508
rect 8481 19499 8539 19505
rect 8481 19465 8493 19499
rect 8527 19496 8539 19499
rect 8941 19499 8999 19505
rect 8941 19496 8953 19499
rect 8527 19468 8953 19496
rect 8527 19465 8539 19468
rect 8481 19459 8539 19465
rect 8941 19465 8953 19468
rect 8987 19465 8999 19499
rect 8941 19459 8999 19465
rect 9309 19499 9367 19505
rect 9309 19465 9321 19499
rect 9355 19465 9367 19499
rect 9309 19459 9367 19465
rect 9585 19499 9643 19505
rect 9585 19465 9597 19499
rect 9631 19496 9643 19499
rect 10226 19496 10232 19508
rect 9631 19468 10232 19496
rect 9631 19465 9643 19468
rect 9585 19459 9643 19465
rect 6730 19428 6736 19440
rect 5460 19400 6592 19428
rect 6691 19400 6736 19428
rect 6730 19388 6736 19400
rect 6788 19388 6794 19440
rect 7926 19388 7932 19440
rect 7984 19388 7990 19440
rect 8021 19431 8079 19437
rect 8021 19397 8033 19431
rect 8067 19428 8079 19431
rect 8662 19428 8668 19440
rect 8067 19400 8668 19428
rect 8067 19397 8079 19400
rect 8021 19391 8079 19397
rect 8662 19388 8668 19400
rect 8720 19388 8726 19440
rect 9324 19428 9352 19459
rect 10226 19456 10232 19468
rect 10284 19456 10290 19508
rect 11333 19499 11391 19505
rect 11333 19465 11345 19499
rect 11379 19496 11391 19499
rect 11882 19496 11888 19508
rect 11379 19468 11888 19496
rect 11379 19465 11391 19468
rect 11333 19459 11391 19465
rect 11882 19456 11888 19468
rect 11940 19456 11946 19508
rect 12986 19496 12992 19508
rect 12947 19468 12992 19496
rect 12986 19456 12992 19468
rect 13044 19456 13050 19508
rect 13078 19456 13084 19508
rect 13136 19496 13142 19508
rect 13817 19499 13875 19505
rect 13817 19496 13829 19499
rect 13136 19468 13829 19496
rect 13136 19456 13142 19468
rect 13817 19465 13829 19468
rect 13863 19465 13875 19499
rect 13817 19459 13875 19465
rect 14182 19456 14188 19508
rect 14240 19496 14246 19508
rect 14240 19468 14504 19496
rect 14240 19456 14246 19468
rect 10410 19428 10416 19440
rect 9324 19400 10416 19428
rect 10410 19388 10416 19400
rect 10468 19388 10474 19440
rect 10870 19437 10876 19440
rect 10812 19431 10876 19437
rect 10812 19397 10824 19431
rect 10858 19397 10876 19431
rect 10812 19391 10876 19397
rect 10870 19388 10876 19391
rect 10928 19388 10934 19440
rect 11762 19431 11820 19437
rect 11072 19400 11560 19428
rect 3513 19363 3571 19369
rect 3513 19329 3525 19363
rect 3559 19329 3571 19363
rect 3513 19323 3571 19329
rect 2501 19295 2559 19301
rect 2501 19261 2513 19295
rect 2547 19261 2559 19295
rect 2501 19255 2559 19261
rect 2593 19295 2651 19301
rect 2593 19261 2605 19295
rect 2639 19292 2651 19295
rect 3329 19295 3387 19301
rect 2639 19264 2673 19292
rect 2639 19261 2651 19264
rect 2593 19255 2651 19261
rect 3329 19261 3341 19295
rect 3375 19261 3387 19295
rect 3329 19255 3387 19261
rect 2516 19224 2544 19255
rect 3418 19224 3424 19236
rect 2516 19196 3424 19224
rect 3418 19184 3424 19196
rect 3476 19184 3482 19236
rect 3528 19224 3556 19323
rect 3602 19320 3608 19372
rect 3660 19360 3666 19372
rect 4341 19363 4399 19369
rect 4341 19360 4353 19363
rect 3660 19332 4353 19360
rect 3660 19320 3666 19332
rect 4341 19329 4353 19332
rect 4387 19360 4399 19363
rect 4798 19360 4804 19372
rect 4387 19332 4660 19360
rect 4759 19332 4804 19360
rect 4387 19329 4399 19332
rect 4341 19323 4399 19329
rect 4157 19295 4215 19301
rect 4157 19261 4169 19295
rect 4203 19292 4215 19295
rect 4522 19292 4528 19304
rect 4203 19264 4528 19292
rect 4203 19261 4215 19264
rect 4157 19255 4215 19261
rect 4522 19252 4528 19264
rect 4580 19252 4586 19304
rect 4632 19292 4660 19332
rect 4798 19320 4804 19332
rect 4856 19320 4862 19372
rect 7098 19360 7104 19372
rect 4908 19332 7104 19360
rect 4908 19292 4936 19332
rect 7098 19320 7104 19332
rect 7156 19320 7162 19372
rect 7282 19360 7288 19372
rect 7243 19332 7288 19360
rect 7282 19320 7288 19332
rect 7340 19320 7346 19372
rect 7377 19363 7435 19369
rect 7377 19329 7389 19363
rect 7423 19360 7435 19363
rect 7944 19360 7972 19388
rect 11072 19372 11100 19400
rect 7423 19332 7972 19360
rect 8113 19363 8171 19369
rect 7423 19329 7435 19332
rect 7377 19323 7435 19329
rect 8113 19329 8125 19363
rect 8159 19360 8171 19363
rect 8478 19360 8484 19372
rect 8159 19332 8484 19360
rect 8159 19329 8171 19332
rect 8113 19323 8171 19329
rect 8478 19320 8484 19332
rect 8536 19320 8542 19372
rect 8849 19363 8907 19369
rect 8849 19360 8861 19363
rect 8588 19332 8861 19360
rect 4632 19264 4936 19292
rect 6270 19252 6276 19304
rect 6328 19292 6334 19304
rect 7006 19292 7012 19304
rect 6328 19264 7012 19292
rect 6328 19252 6334 19264
rect 7006 19252 7012 19264
rect 7064 19252 7070 19304
rect 7558 19292 7564 19304
rect 7519 19264 7564 19292
rect 7558 19252 7564 19264
rect 7616 19252 7622 19304
rect 7742 19252 7748 19304
rect 7800 19292 7806 19304
rect 7837 19295 7895 19301
rect 7837 19292 7849 19295
rect 7800 19264 7849 19292
rect 7800 19252 7806 19264
rect 7837 19261 7849 19264
rect 7883 19261 7895 19295
rect 7837 19255 7895 19261
rect 7926 19252 7932 19304
rect 7984 19292 7990 19304
rect 8588 19292 8616 19332
rect 8849 19329 8861 19332
rect 8895 19329 8907 19363
rect 8849 19323 8907 19329
rect 9122 19320 9128 19372
rect 9180 19360 9186 19372
rect 9401 19363 9459 19369
rect 9401 19360 9413 19363
rect 9180 19332 9413 19360
rect 9180 19320 9186 19332
rect 9401 19329 9413 19332
rect 9447 19329 9459 19363
rect 11054 19360 11060 19372
rect 11015 19332 11060 19360
rect 9401 19323 9459 19329
rect 11054 19320 11060 19332
rect 11112 19320 11118 19372
rect 11532 19369 11560 19400
rect 11762 19397 11774 19431
rect 11808 19428 11820 19431
rect 12158 19428 12164 19440
rect 11808 19400 12164 19428
rect 11808 19397 11820 19400
rect 11762 19391 11820 19397
rect 12158 19388 12164 19400
rect 12216 19388 12222 19440
rect 13906 19428 13912 19440
rect 12406 19400 13912 19428
rect 11149 19363 11207 19369
rect 11149 19329 11161 19363
rect 11195 19329 11207 19363
rect 11149 19323 11207 19329
rect 11517 19363 11575 19369
rect 11517 19329 11529 19363
rect 11563 19360 11575 19363
rect 12406 19360 12434 19400
rect 13906 19388 13912 19400
rect 13964 19388 13970 19440
rect 14476 19437 14504 19468
rect 14734 19456 14740 19508
rect 14792 19496 14798 19508
rect 15657 19499 15715 19505
rect 15657 19496 15669 19499
rect 14792 19468 15669 19496
rect 14792 19456 14798 19468
rect 15657 19465 15669 19468
rect 15703 19465 15715 19499
rect 15657 19459 15715 19465
rect 15838 19456 15844 19508
rect 15896 19496 15902 19508
rect 16117 19499 16175 19505
rect 15896 19468 15976 19496
rect 15896 19456 15902 19468
rect 14452 19431 14510 19437
rect 14452 19397 14464 19431
rect 14498 19397 14510 19431
rect 14452 19391 14510 19397
rect 15948 19393 15976 19468
rect 16117 19465 16129 19499
rect 16163 19465 16175 19499
rect 16117 19459 16175 19465
rect 16393 19499 16451 19505
rect 16393 19465 16405 19499
rect 16439 19496 16451 19499
rect 17402 19496 17408 19508
rect 16439 19468 17408 19496
rect 16439 19465 16451 19468
rect 16393 19459 16451 19465
rect 15933 19387 15991 19393
rect 13354 19360 13360 19372
rect 11563 19332 12434 19360
rect 13315 19332 13360 19360
rect 11563 19329 11575 19332
rect 11517 19323 11575 19329
rect 8754 19292 8760 19304
rect 7984 19264 8616 19292
rect 8715 19264 8760 19292
rect 7984 19252 7990 19264
rect 8754 19252 8760 19264
rect 8812 19252 8818 19304
rect 11164 19292 11192 19323
rect 13354 19320 13360 19332
rect 13412 19320 13418 19372
rect 14001 19363 14059 19369
rect 14001 19329 14013 19363
rect 14047 19360 14059 19363
rect 14090 19360 14096 19372
rect 14047 19332 14096 19360
rect 14047 19329 14059 19332
rect 14001 19323 14059 19329
rect 14090 19320 14096 19332
rect 14148 19320 14154 19372
rect 15746 19360 15752 19372
rect 14292 19332 15752 19360
rect 11072 19264 11192 19292
rect 11072 19236 11100 19264
rect 12894 19252 12900 19304
rect 12952 19292 12958 19304
rect 13449 19295 13507 19301
rect 13449 19292 13461 19295
rect 12952 19264 13461 19292
rect 12952 19252 12958 19264
rect 13449 19261 13461 19264
rect 13495 19261 13507 19295
rect 13449 19255 13507 19261
rect 13538 19252 13544 19304
rect 13596 19292 13602 19304
rect 14185 19295 14243 19301
rect 13596 19264 13641 19292
rect 13596 19252 13602 19264
rect 14185 19261 14197 19295
rect 14231 19292 14243 19295
rect 14292 19292 14320 19332
rect 15746 19320 15752 19332
rect 15804 19320 15810 19372
rect 15841 19363 15899 19369
rect 15841 19329 15853 19363
rect 15887 19329 15899 19363
rect 15933 19353 15945 19387
rect 15979 19353 15991 19387
rect 15933 19347 15991 19353
rect 16132 19360 16160 19459
rect 17402 19456 17408 19468
rect 17460 19456 17466 19508
rect 17957 19499 18015 19505
rect 17957 19465 17969 19499
rect 18003 19496 18015 19499
rect 18322 19496 18328 19508
rect 18003 19468 18328 19496
rect 18003 19465 18015 19468
rect 17957 19459 18015 19465
rect 18322 19456 18328 19468
rect 18380 19456 18386 19508
rect 18782 19496 18788 19508
rect 18743 19468 18788 19496
rect 18782 19456 18788 19468
rect 18840 19456 18846 19508
rect 18966 19456 18972 19508
rect 19024 19456 19030 19508
rect 19058 19456 19064 19508
rect 19116 19496 19122 19508
rect 19521 19499 19579 19505
rect 19116 19468 19161 19496
rect 19116 19456 19122 19468
rect 19521 19465 19533 19499
rect 19567 19465 19579 19499
rect 19521 19459 19579 19465
rect 19797 19499 19855 19505
rect 19797 19465 19809 19499
rect 19843 19496 19855 19499
rect 20070 19496 20076 19508
rect 19843 19468 20076 19496
rect 19843 19465 19855 19468
rect 19797 19459 19855 19465
rect 18138 19428 18144 19440
rect 17144 19400 18144 19428
rect 16209 19363 16267 19369
rect 16209 19360 16221 19363
rect 16132 19332 16221 19360
rect 15841 19323 15899 19329
rect 16209 19329 16221 19332
rect 16255 19329 16267 19363
rect 16850 19360 16856 19372
rect 16811 19332 16856 19360
rect 16209 19323 16267 19329
rect 14231 19264 14320 19292
rect 15856 19292 15884 19323
rect 16850 19320 16856 19332
rect 16908 19320 16914 19372
rect 16945 19363 17003 19369
rect 16945 19329 16957 19363
rect 16991 19329 17003 19363
rect 16945 19323 17003 19329
rect 16114 19292 16120 19304
rect 15856 19264 16120 19292
rect 14231 19261 14243 19264
rect 14185 19255 14243 19261
rect 16114 19252 16120 19264
rect 16172 19252 16178 19304
rect 8386 19224 8392 19236
rect 3528 19196 4844 19224
rect 1486 19156 1492 19168
rect 1447 19128 1492 19156
rect 1486 19116 1492 19128
rect 1544 19116 1550 19168
rect 2222 19156 2228 19168
rect 2183 19128 2228 19156
rect 2222 19116 2228 19128
rect 2280 19116 2286 19168
rect 3050 19156 3056 19168
rect 3011 19128 3056 19156
rect 3050 19116 3056 19128
rect 3108 19116 3114 19168
rect 3326 19116 3332 19168
rect 3384 19156 3390 19168
rect 3602 19156 3608 19168
rect 3384 19128 3608 19156
rect 3384 19116 3390 19128
rect 3602 19116 3608 19128
rect 3660 19116 3666 19168
rect 3878 19156 3884 19168
rect 3839 19128 3884 19156
rect 3878 19116 3884 19128
rect 3936 19116 3942 19168
rect 4816 19156 4844 19196
rect 6380 19196 8392 19224
rect 4982 19156 4988 19168
rect 4816 19128 4988 19156
rect 4982 19116 4988 19128
rect 5040 19116 5046 19168
rect 5074 19116 5080 19168
rect 5132 19156 5138 19168
rect 6380 19156 6408 19196
rect 8386 19184 8392 19196
rect 8444 19184 8450 19236
rect 8846 19184 8852 19236
rect 8904 19224 8910 19236
rect 8904 19196 9996 19224
rect 8904 19184 8910 19196
rect 5132 19128 6408 19156
rect 6457 19159 6515 19165
rect 5132 19116 5138 19128
rect 6457 19125 6469 19159
rect 6503 19156 6515 19159
rect 6546 19156 6552 19168
rect 6503 19128 6552 19156
rect 6503 19125 6515 19128
rect 6457 19119 6515 19125
rect 6546 19116 6552 19128
rect 6604 19116 6610 19168
rect 6641 19159 6699 19165
rect 6641 19125 6653 19159
rect 6687 19156 6699 19159
rect 6730 19156 6736 19168
rect 6687 19128 6736 19156
rect 6687 19125 6699 19128
rect 6641 19119 6699 19125
rect 6730 19116 6736 19128
rect 6788 19116 6794 19168
rect 6914 19156 6920 19168
rect 6875 19128 6920 19156
rect 6914 19116 6920 19128
rect 6972 19116 6978 19168
rect 7006 19116 7012 19168
rect 7064 19156 7070 19168
rect 7650 19156 7656 19168
rect 7064 19128 7656 19156
rect 7064 19116 7070 19128
rect 7650 19116 7656 19128
rect 7708 19116 7714 19168
rect 8404 19156 8432 19184
rect 9582 19156 9588 19168
rect 8404 19128 9588 19156
rect 9582 19116 9588 19128
rect 9640 19116 9646 19168
rect 9674 19116 9680 19168
rect 9732 19156 9738 19168
rect 9968 19156 9996 19196
rect 11054 19184 11060 19236
rect 11112 19184 11118 19236
rect 15930 19184 15936 19236
rect 15988 19224 15994 19236
rect 16669 19227 16727 19233
rect 16669 19224 16681 19227
rect 15988 19196 16681 19224
rect 15988 19184 15994 19196
rect 16669 19193 16681 19196
rect 16715 19193 16727 19227
rect 16669 19187 16727 19193
rect 12802 19156 12808 19168
rect 9732 19128 9777 19156
rect 9968 19128 12808 19156
rect 9732 19116 9738 19128
rect 12802 19116 12808 19128
rect 12860 19116 12866 19168
rect 12897 19159 12955 19165
rect 12897 19125 12909 19159
rect 12943 19156 12955 19159
rect 13170 19156 13176 19168
rect 12943 19128 13176 19156
rect 12943 19125 12955 19128
rect 12897 19119 12955 19125
rect 13170 19116 13176 19128
rect 13228 19116 13234 19168
rect 15565 19159 15623 19165
rect 15565 19125 15577 19159
rect 15611 19156 15623 19159
rect 15654 19156 15660 19168
rect 15611 19128 15660 19156
rect 15611 19125 15623 19128
rect 15565 19119 15623 19125
rect 15654 19116 15660 19128
rect 15712 19116 15718 19168
rect 16960 19156 16988 19323
rect 17144 19233 17172 19400
rect 18138 19388 18144 19400
rect 18196 19388 18202 19440
rect 18984 19428 19012 19456
rect 19536 19428 19564 19459
rect 20070 19456 20076 19468
rect 20128 19456 20134 19508
rect 20530 19496 20536 19508
rect 20491 19468 20536 19496
rect 20530 19456 20536 19468
rect 20588 19456 20594 19508
rect 21450 19496 21456 19508
rect 21411 19468 21456 19496
rect 21450 19456 21456 19468
rect 21508 19456 21514 19508
rect 20162 19428 20168 19440
rect 18984 19400 19380 19428
rect 19536 19400 20168 19428
rect 17770 19360 17776 19372
rect 17731 19332 17776 19360
rect 17770 19320 17776 19332
rect 17828 19320 17834 19372
rect 18230 19320 18236 19372
rect 18288 19320 18294 19372
rect 18417 19363 18475 19369
rect 18417 19329 18429 19363
rect 18463 19360 18475 19363
rect 18690 19360 18696 19372
rect 18463 19332 18552 19360
rect 18651 19332 18696 19360
rect 18463 19329 18475 19332
rect 18417 19323 18475 19329
rect 17788 19292 17816 19320
rect 18049 19295 18107 19301
rect 18049 19292 18061 19295
rect 17788 19264 18061 19292
rect 18049 19261 18061 19264
rect 18095 19261 18107 19295
rect 18049 19255 18107 19261
rect 17129 19227 17187 19233
rect 17129 19193 17141 19227
rect 17175 19193 17187 19227
rect 17310 19224 17316 19236
rect 17129 19187 17187 19193
rect 17236 19196 17316 19224
rect 17236 19156 17264 19196
rect 17310 19184 17316 19196
rect 17368 19184 17374 19236
rect 18248 19233 18276 19320
rect 18233 19227 18291 19233
rect 18233 19193 18245 19227
rect 18279 19193 18291 19227
rect 18233 19187 18291 19193
rect 17402 19156 17408 19168
rect 16960 19128 17264 19156
rect 17363 19128 17408 19156
rect 17402 19116 17408 19128
rect 17460 19116 17466 19168
rect 17678 19156 17684 19168
rect 17639 19128 17684 19156
rect 17678 19116 17684 19128
rect 17736 19116 17742 19168
rect 18524 19165 18552 19332
rect 18690 19320 18696 19332
rect 18748 19320 18754 19372
rect 18969 19363 19027 19369
rect 18969 19329 18981 19363
rect 19015 19360 19027 19363
rect 19150 19360 19156 19372
rect 19015 19332 19156 19360
rect 19015 19329 19027 19332
rect 18969 19323 19027 19329
rect 19150 19320 19156 19332
rect 19208 19320 19214 19372
rect 19352 19369 19380 19400
rect 20162 19388 20168 19400
rect 20220 19388 20226 19440
rect 20254 19388 20260 19440
rect 20312 19388 20318 19440
rect 19245 19363 19303 19369
rect 19245 19329 19257 19363
rect 19291 19329 19303 19363
rect 19245 19323 19303 19329
rect 19337 19363 19395 19369
rect 19337 19329 19349 19363
rect 19383 19329 19395 19363
rect 19337 19323 19395 19329
rect 18598 19252 18604 19304
rect 18656 19292 18662 19304
rect 19260 19292 19288 19323
rect 19426 19320 19432 19372
rect 19484 19360 19490 19372
rect 19613 19363 19671 19369
rect 19613 19360 19625 19363
rect 19484 19332 19625 19360
rect 19484 19320 19490 19332
rect 19613 19329 19625 19332
rect 19659 19360 19671 19363
rect 19886 19360 19892 19372
rect 19659 19332 19892 19360
rect 19659 19329 19671 19332
rect 19613 19323 19671 19329
rect 19886 19320 19892 19332
rect 19944 19320 19950 19372
rect 19981 19363 20039 19369
rect 19981 19329 19993 19363
rect 20027 19360 20039 19363
rect 20272 19360 20300 19388
rect 20027 19332 20300 19360
rect 20349 19363 20407 19369
rect 20027 19329 20039 19332
rect 19981 19323 20039 19329
rect 20349 19329 20361 19363
rect 20395 19329 20407 19363
rect 20349 19323 20407 19329
rect 18656 19264 19288 19292
rect 20364 19292 20392 19323
rect 20438 19320 20444 19372
rect 20496 19360 20502 19372
rect 20717 19363 20775 19369
rect 20717 19360 20729 19363
rect 20496 19332 20729 19360
rect 20496 19320 20502 19332
rect 20717 19329 20729 19332
rect 20763 19329 20775 19363
rect 20990 19360 20996 19372
rect 20951 19332 20996 19360
rect 20717 19323 20775 19329
rect 20990 19320 20996 19332
rect 21048 19320 21054 19372
rect 21266 19360 21272 19372
rect 21227 19332 21272 19360
rect 21266 19320 21272 19332
rect 21324 19320 21330 19372
rect 20622 19292 20628 19304
rect 20364 19264 20628 19292
rect 18656 19252 18662 19264
rect 20622 19252 20628 19264
rect 20680 19252 20686 19304
rect 20165 19227 20223 19233
rect 20165 19193 20177 19227
rect 20211 19224 20223 19227
rect 20254 19224 20260 19236
rect 20211 19196 20260 19224
rect 20211 19193 20223 19196
rect 20165 19187 20223 19193
rect 20254 19184 20260 19196
rect 20312 19184 20318 19236
rect 18509 19159 18567 19165
rect 18509 19125 18521 19159
rect 18555 19156 18567 19159
rect 18966 19156 18972 19168
rect 18555 19128 18972 19156
rect 18555 19125 18567 19128
rect 18509 19119 18567 19125
rect 18966 19116 18972 19128
rect 19024 19116 19030 19168
rect 1104 19066 21896 19088
rect 1104 19014 3549 19066
rect 3601 19014 3613 19066
rect 3665 19014 3677 19066
rect 3729 19014 3741 19066
rect 3793 19014 3805 19066
rect 3857 19014 8747 19066
rect 8799 19014 8811 19066
rect 8863 19014 8875 19066
rect 8927 19014 8939 19066
rect 8991 19014 9003 19066
rect 9055 19014 13945 19066
rect 13997 19014 14009 19066
rect 14061 19014 14073 19066
rect 14125 19014 14137 19066
rect 14189 19014 14201 19066
rect 14253 19014 19143 19066
rect 19195 19014 19207 19066
rect 19259 19014 19271 19066
rect 19323 19014 19335 19066
rect 19387 19014 19399 19066
rect 19451 19014 21896 19066
rect 1104 18992 21896 19014
rect 3142 18912 3148 18964
rect 3200 18952 3206 18964
rect 3789 18955 3847 18961
rect 3789 18952 3801 18955
rect 3200 18924 3801 18952
rect 3200 18912 3206 18924
rect 3789 18921 3801 18924
rect 3835 18921 3847 18955
rect 6270 18952 6276 18964
rect 3789 18915 3847 18921
rect 5276 18924 6276 18952
rect 1857 18887 1915 18893
rect 1857 18853 1869 18887
rect 1903 18853 1915 18887
rect 1857 18847 1915 18853
rect 1673 18751 1731 18757
rect 1673 18717 1685 18751
rect 1719 18748 1731 18751
rect 1872 18748 1900 18847
rect 2222 18844 2228 18896
rect 2280 18884 2286 18896
rect 5276 18884 5304 18924
rect 6270 18912 6276 18924
rect 6328 18912 6334 18964
rect 6457 18955 6515 18961
rect 6457 18921 6469 18955
rect 6503 18952 6515 18955
rect 6730 18952 6736 18964
rect 6503 18924 6736 18952
rect 6503 18921 6515 18924
rect 6457 18915 6515 18921
rect 6730 18912 6736 18924
rect 6788 18912 6794 18964
rect 7653 18955 7711 18961
rect 7653 18921 7665 18955
rect 7699 18952 7711 18955
rect 7926 18952 7932 18964
rect 7699 18924 7932 18952
rect 7699 18921 7711 18924
rect 7653 18915 7711 18921
rect 7926 18912 7932 18924
rect 7984 18912 7990 18964
rect 8478 18952 8484 18964
rect 8439 18924 8484 18952
rect 8478 18912 8484 18924
rect 8536 18912 8542 18964
rect 8662 18912 8668 18964
rect 8720 18952 8726 18964
rect 8941 18955 8999 18961
rect 8941 18952 8953 18955
rect 8720 18924 8953 18952
rect 8720 18912 8726 18924
rect 8941 18921 8953 18924
rect 8987 18921 8999 18955
rect 8941 18915 8999 18921
rect 10594 18912 10600 18964
rect 10652 18952 10658 18964
rect 10965 18955 11023 18961
rect 10965 18952 10977 18955
rect 10652 18924 10977 18952
rect 10652 18912 10658 18924
rect 10965 18921 10977 18924
rect 11011 18921 11023 18955
rect 10965 18915 11023 18921
rect 11241 18955 11299 18961
rect 11241 18921 11253 18955
rect 11287 18952 11299 18955
rect 11790 18952 11796 18964
rect 11287 18924 11796 18952
rect 11287 18921 11299 18924
rect 11241 18915 11299 18921
rect 11790 18912 11796 18924
rect 11848 18912 11854 18964
rect 12069 18955 12127 18961
rect 12069 18921 12081 18955
rect 12115 18952 12127 18955
rect 12894 18952 12900 18964
rect 12115 18924 12900 18952
rect 12115 18921 12127 18924
rect 12069 18915 12127 18921
rect 12894 18912 12900 18924
rect 12952 18912 12958 18964
rect 13354 18912 13360 18964
rect 13412 18952 13418 18964
rect 13725 18955 13783 18961
rect 13725 18952 13737 18955
rect 13412 18924 13737 18952
rect 13412 18912 13418 18924
rect 13725 18921 13737 18924
rect 13771 18921 13783 18955
rect 15470 18952 15476 18964
rect 15431 18924 15476 18952
rect 13725 18915 13783 18921
rect 15470 18912 15476 18924
rect 15528 18912 15534 18964
rect 15749 18955 15807 18961
rect 15749 18921 15761 18955
rect 15795 18952 15807 18955
rect 17034 18952 17040 18964
rect 15795 18924 17040 18952
rect 15795 18921 15807 18924
rect 15749 18915 15807 18921
rect 17034 18912 17040 18924
rect 17092 18912 17098 18964
rect 17957 18955 18015 18961
rect 17957 18921 17969 18955
rect 18003 18952 18015 18955
rect 18046 18952 18052 18964
rect 18003 18924 18052 18952
rect 18003 18921 18015 18924
rect 17957 18915 18015 18921
rect 18046 18912 18052 18924
rect 18104 18912 18110 18964
rect 18506 18952 18512 18964
rect 18467 18924 18512 18952
rect 18506 18912 18512 18924
rect 18564 18912 18570 18964
rect 18785 18955 18843 18961
rect 18785 18921 18797 18955
rect 18831 18952 18843 18955
rect 20441 18955 20499 18961
rect 18831 18924 20116 18952
rect 18831 18921 18843 18924
rect 18785 18915 18843 18921
rect 2280 18856 5304 18884
rect 2280 18844 2286 18856
rect 5350 18844 5356 18896
rect 5408 18884 5414 18896
rect 5408 18856 5453 18884
rect 5552 18856 7236 18884
rect 5408 18844 5414 18856
rect 3326 18816 3332 18828
rect 3287 18788 3332 18816
rect 3326 18776 3332 18788
rect 3384 18776 3390 18828
rect 3418 18776 3424 18828
rect 3476 18816 3482 18828
rect 3476 18788 3521 18816
rect 3476 18776 3482 18788
rect 3878 18776 3884 18828
rect 3936 18816 3942 18828
rect 4249 18819 4307 18825
rect 4249 18816 4261 18819
rect 3936 18788 4261 18816
rect 3936 18776 3942 18788
rect 4249 18785 4261 18788
rect 4295 18785 4307 18819
rect 4430 18816 4436 18828
rect 4391 18788 4436 18816
rect 4249 18779 4307 18785
rect 4430 18776 4436 18788
rect 4488 18776 4494 18828
rect 4706 18816 4712 18828
rect 4667 18788 4712 18816
rect 4706 18776 4712 18788
rect 4764 18776 4770 18828
rect 5552 18816 5580 18856
rect 5307 18788 5580 18816
rect 1719 18720 1900 18748
rect 2041 18751 2099 18757
rect 1719 18717 1731 18720
rect 1673 18711 1731 18717
rect 2041 18717 2053 18751
rect 2087 18748 2099 18751
rect 2222 18748 2228 18760
rect 2087 18720 2228 18748
rect 2087 18717 2099 18720
rect 2041 18711 2099 18717
rect 2222 18708 2228 18720
rect 2280 18708 2286 18760
rect 2317 18751 2375 18757
rect 2317 18717 2329 18751
rect 2363 18748 2375 18751
rect 2590 18748 2596 18760
rect 2363 18720 2596 18748
rect 2363 18717 2375 18720
rect 2317 18711 2375 18717
rect 2590 18708 2596 18720
rect 2648 18708 2654 18760
rect 2777 18751 2835 18757
rect 2777 18717 2789 18751
rect 2823 18748 2835 18751
rect 3970 18748 3976 18760
rect 2823 18720 3976 18748
rect 2823 18717 2835 18720
rect 2777 18711 2835 18717
rect 3970 18708 3976 18720
rect 4028 18708 4034 18760
rect 4062 18708 4068 18760
rect 4120 18748 4126 18760
rect 5307 18748 5335 18788
rect 5626 18776 5632 18828
rect 5684 18816 5690 18828
rect 7208 18825 7236 18856
rect 8110 18844 8116 18896
rect 8168 18884 8174 18896
rect 9769 18887 9827 18893
rect 9769 18884 9781 18887
rect 8168 18856 9781 18884
rect 8168 18844 8174 18856
rect 9769 18853 9781 18856
rect 9815 18853 9827 18887
rect 15197 18887 15255 18893
rect 9769 18847 9827 18853
rect 11532 18856 13216 18884
rect 5997 18819 6055 18825
rect 5997 18816 6009 18819
rect 5684 18788 6009 18816
rect 5684 18776 5690 18788
rect 5997 18785 6009 18788
rect 6043 18785 6055 18819
rect 5997 18779 6055 18785
rect 7101 18819 7159 18825
rect 7101 18785 7113 18819
rect 7147 18785 7159 18819
rect 7101 18779 7159 18785
rect 7193 18819 7251 18825
rect 7193 18785 7205 18819
rect 7239 18785 7251 18819
rect 7193 18779 7251 18785
rect 6270 18748 6276 18760
rect 4120 18720 5335 18748
rect 5368 18720 5672 18748
rect 6231 18720 6276 18748
rect 4120 18708 4126 18720
rect 2409 18683 2467 18689
rect 2409 18649 2421 18683
rect 2455 18680 2467 18683
rect 5368 18680 5396 18720
rect 2455 18652 5396 18680
rect 5644 18680 5672 18720
rect 6270 18708 6276 18720
rect 6328 18708 6334 18760
rect 7116 18744 7144 18779
rect 7558 18776 7564 18828
rect 7616 18816 7622 18828
rect 7929 18819 7987 18825
rect 7929 18816 7941 18819
rect 7616 18788 7941 18816
rect 7616 18776 7622 18788
rect 7929 18785 7941 18788
rect 7975 18816 7987 18819
rect 9493 18819 9551 18825
rect 9493 18816 9505 18819
rect 7975 18788 9505 18816
rect 7975 18785 7987 18788
rect 7929 18779 7987 18785
rect 9493 18785 9505 18788
rect 9539 18785 9551 18819
rect 9493 18779 9551 18785
rect 9582 18776 9588 18828
rect 9640 18816 9646 18828
rect 11532 18825 11560 18856
rect 13188 18828 13216 18856
rect 15197 18853 15209 18887
rect 15243 18884 15255 18887
rect 16942 18884 16948 18896
rect 15243 18856 16948 18884
rect 15243 18853 15255 18856
rect 15197 18847 15255 18853
rect 16942 18844 16948 18856
rect 17000 18844 17006 18896
rect 18233 18887 18291 18893
rect 18233 18853 18245 18887
rect 18279 18884 18291 18887
rect 18279 18856 19472 18884
rect 18279 18853 18291 18856
rect 18233 18847 18291 18853
rect 19444 18828 19472 18856
rect 10321 18819 10379 18825
rect 10321 18816 10333 18819
rect 9640 18788 10333 18816
rect 9640 18776 9646 18788
rect 10321 18785 10333 18788
rect 10367 18785 10379 18819
rect 11517 18819 11575 18825
rect 10321 18779 10379 18785
rect 10612 18788 11100 18816
rect 10612 18760 10640 18788
rect 7742 18748 7748 18760
rect 7208 18744 7748 18748
rect 7116 18720 7748 18744
rect 7116 18716 7236 18720
rect 7742 18708 7748 18720
rect 7800 18708 7806 18760
rect 8573 18751 8631 18757
rect 8573 18748 8585 18751
rect 7852 18720 8585 18748
rect 6638 18680 6644 18692
rect 5644 18652 6644 18680
rect 2455 18649 2467 18652
rect 2409 18643 2467 18649
rect 6638 18640 6644 18652
rect 6696 18640 6702 18692
rect 6914 18640 6920 18692
rect 6972 18680 6978 18692
rect 7285 18683 7343 18689
rect 7285 18680 7297 18683
rect 6972 18652 7297 18680
rect 6972 18640 6978 18652
rect 7285 18649 7297 18652
rect 7331 18649 7343 18683
rect 7285 18643 7343 18649
rect 1486 18612 1492 18624
rect 1447 18584 1492 18612
rect 1486 18572 1492 18584
rect 1544 18572 1550 18624
rect 2038 18572 2044 18624
rect 2096 18612 2102 18624
rect 2133 18615 2191 18621
rect 2133 18612 2145 18615
rect 2096 18584 2145 18612
rect 2096 18572 2102 18584
rect 2133 18581 2145 18584
rect 2179 18581 2191 18615
rect 2133 18575 2191 18581
rect 2498 18572 2504 18624
rect 2556 18612 2562 18624
rect 2593 18615 2651 18621
rect 2593 18612 2605 18615
rect 2556 18584 2605 18612
rect 2556 18572 2562 18584
rect 2593 18581 2605 18584
rect 2639 18612 2651 18615
rect 2682 18612 2688 18624
rect 2639 18584 2688 18612
rect 2639 18581 2651 18584
rect 2593 18575 2651 18581
rect 2682 18572 2688 18584
rect 2740 18572 2746 18624
rect 2869 18615 2927 18621
rect 2869 18581 2881 18615
rect 2915 18612 2927 18615
rect 3142 18612 3148 18624
rect 2915 18584 3148 18612
rect 2915 18581 2927 18584
rect 2869 18575 2927 18581
rect 3142 18572 3148 18584
rect 3200 18572 3206 18624
rect 3237 18615 3295 18621
rect 3237 18581 3249 18615
rect 3283 18612 3295 18615
rect 3326 18612 3332 18624
rect 3283 18584 3332 18612
rect 3283 18581 3295 18584
rect 3237 18575 3295 18581
rect 3326 18572 3332 18584
rect 3384 18572 3390 18624
rect 4157 18615 4215 18621
rect 4157 18581 4169 18615
rect 4203 18612 4215 18615
rect 4246 18612 4252 18624
rect 4203 18584 4252 18612
rect 4203 18581 4215 18584
rect 4157 18575 4215 18581
rect 4246 18572 4252 18584
rect 4304 18572 4310 18624
rect 4890 18612 4896 18624
rect 4851 18584 4896 18612
rect 4890 18572 4896 18584
rect 4948 18572 4954 18624
rect 4982 18572 4988 18624
rect 5040 18612 5046 18624
rect 5040 18584 5085 18612
rect 5040 18572 5046 18584
rect 5350 18572 5356 18624
rect 5408 18612 5414 18624
rect 5445 18615 5503 18621
rect 5445 18612 5457 18615
rect 5408 18584 5457 18612
rect 5408 18572 5414 18584
rect 5445 18581 5457 18584
rect 5491 18581 5503 18615
rect 5810 18612 5816 18624
rect 5771 18584 5816 18612
rect 5445 18575 5503 18581
rect 5810 18572 5816 18584
rect 5868 18572 5874 18624
rect 5902 18572 5908 18624
rect 5960 18612 5966 18624
rect 6733 18615 6791 18621
rect 5960 18584 6005 18612
rect 5960 18572 5966 18584
rect 6733 18581 6745 18615
rect 6779 18612 6791 18615
rect 7650 18612 7656 18624
rect 6779 18584 7656 18612
rect 6779 18581 6791 18584
rect 6733 18575 6791 18581
rect 7650 18572 7656 18584
rect 7708 18572 7714 18624
rect 7742 18572 7748 18624
rect 7800 18612 7806 18624
rect 7852 18612 7880 18720
rect 8573 18717 8585 18720
rect 8619 18717 8631 18751
rect 8573 18711 8631 18717
rect 9766 18708 9772 18760
rect 9824 18748 9830 18760
rect 10226 18748 10232 18760
rect 9824 18720 9996 18748
rect 10187 18720 10232 18748
rect 9824 18708 9830 18720
rect 8202 18640 8208 18692
rect 8260 18680 8266 18692
rect 9858 18680 9864 18692
rect 8260 18652 9864 18680
rect 8260 18640 8266 18652
rect 9858 18640 9864 18652
rect 9916 18640 9922 18692
rect 9968 18680 9996 18720
rect 10226 18708 10232 18720
rect 10284 18708 10290 18760
rect 10594 18748 10600 18760
rect 10555 18720 10600 18748
rect 10594 18708 10600 18720
rect 10652 18708 10658 18760
rect 10778 18748 10784 18760
rect 10739 18720 10784 18748
rect 10778 18708 10784 18720
rect 10836 18708 10842 18760
rect 11072 18757 11100 18788
rect 11517 18785 11529 18819
rect 11563 18785 11575 18819
rect 11517 18779 11575 18785
rect 11609 18819 11667 18825
rect 11609 18785 11621 18819
rect 11655 18816 11667 18819
rect 11882 18816 11888 18828
rect 11655 18788 11888 18816
rect 11655 18785 11667 18788
rect 11609 18779 11667 18785
rect 11882 18776 11888 18788
rect 11940 18776 11946 18828
rect 12158 18776 12164 18828
rect 12216 18816 12222 18828
rect 12253 18819 12311 18825
rect 12253 18816 12265 18819
rect 12216 18788 12265 18816
rect 12216 18776 12222 18788
rect 12253 18785 12265 18788
rect 12299 18785 12311 18819
rect 12253 18779 12311 18785
rect 12342 18776 12348 18828
rect 12400 18816 12406 18828
rect 12437 18819 12495 18825
rect 12437 18816 12449 18819
rect 12400 18788 12449 18816
rect 12400 18776 12406 18788
rect 12437 18785 12449 18788
rect 12483 18816 12495 18819
rect 12894 18816 12900 18828
rect 12483 18788 12900 18816
rect 12483 18785 12495 18788
rect 12437 18779 12495 18785
rect 12894 18776 12900 18788
rect 12952 18776 12958 18828
rect 13170 18816 13176 18828
rect 13131 18788 13176 18816
rect 13170 18776 13176 18788
rect 13228 18776 13234 18828
rect 14369 18819 14427 18825
rect 14369 18785 14381 18819
rect 14415 18816 14427 18819
rect 14415 18788 14872 18816
rect 14415 18785 14427 18788
rect 14369 18779 14427 18785
rect 11057 18751 11115 18757
rect 11057 18717 11069 18751
rect 11103 18717 11115 18751
rect 11974 18748 11980 18760
rect 11057 18711 11115 18717
rect 11164 18720 11980 18748
rect 11164 18680 11192 18720
rect 11974 18708 11980 18720
rect 12032 18708 12038 18760
rect 14553 18751 14611 18757
rect 14553 18748 14565 18751
rect 12406 18720 14565 18748
rect 12406 18680 12434 18720
rect 14553 18717 14565 18720
rect 14599 18717 14611 18751
rect 14553 18711 14611 18717
rect 13357 18683 13415 18689
rect 13357 18680 13369 18683
rect 9968 18652 11192 18680
rect 11624 18652 12434 18680
rect 12912 18652 13369 18680
rect 8018 18612 8024 18624
rect 7800 18584 7880 18612
rect 7979 18584 8024 18612
rect 7800 18572 7806 18584
rect 8018 18572 8024 18584
rect 8076 18572 8082 18624
rect 8110 18572 8116 18624
rect 8168 18612 8174 18624
rect 8168 18584 8213 18612
rect 8168 18572 8174 18584
rect 8294 18572 8300 18624
rect 8352 18612 8358 18624
rect 8478 18612 8484 18624
rect 8352 18584 8484 18612
rect 8352 18572 8358 18584
rect 8478 18572 8484 18584
rect 8536 18572 8542 18624
rect 8754 18612 8760 18624
rect 8715 18584 8760 18612
rect 8754 18572 8760 18584
rect 8812 18572 8818 18624
rect 9306 18612 9312 18624
rect 9267 18584 9312 18612
rect 9306 18572 9312 18584
rect 9364 18572 9370 18624
rect 9398 18572 9404 18624
rect 9456 18612 9462 18624
rect 9456 18584 9501 18612
rect 9456 18572 9462 18584
rect 9766 18572 9772 18624
rect 9824 18612 9830 18624
rect 10137 18615 10195 18621
rect 10137 18612 10149 18615
rect 9824 18584 10149 18612
rect 9824 18572 9830 18584
rect 10137 18581 10149 18584
rect 10183 18612 10195 18615
rect 11624 18612 11652 18652
rect 10183 18584 11652 18612
rect 11701 18615 11759 18621
rect 10183 18581 10195 18584
rect 10137 18575 10195 18581
rect 11701 18581 11713 18615
rect 11747 18612 11759 18615
rect 12066 18612 12072 18624
rect 11747 18584 12072 18612
rect 11747 18581 11759 18584
rect 11701 18575 11759 18581
rect 12066 18572 12072 18584
rect 12124 18572 12130 18624
rect 12526 18572 12532 18624
rect 12584 18612 12590 18624
rect 12912 18621 12940 18652
rect 13357 18649 13369 18652
rect 13403 18649 13415 18683
rect 13357 18643 13415 18649
rect 13446 18640 13452 18692
rect 13504 18680 13510 18692
rect 14461 18683 14519 18689
rect 14461 18680 14473 18683
rect 13504 18652 14473 18680
rect 13504 18640 13510 18652
rect 14461 18649 14473 18652
rect 14507 18649 14519 18683
rect 14844 18680 14872 18788
rect 16022 18776 16028 18828
rect 16080 18816 16086 18828
rect 17402 18816 17408 18828
rect 16080 18788 17408 18816
rect 16080 18776 16086 18788
rect 17402 18776 17408 18788
rect 17460 18776 17466 18828
rect 19288 18816 19294 18828
rect 18340 18788 19294 18816
rect 15010 18748 15016 18760
rect 14971 18720 15016 18748
rect 15010 18708 15016 18720
rect 15068 18708 15074 18760
rect 15102 18708 15108 18760
rect 15160 18748 15166 18760
rect 15289 18751 15347 18757
rect 15289 18748 15301 18751
rect 15160 18720 15301 18748
rect 15160 18708 15166 18720
rect 15289 18717 15301 18720
rect 15335 18717 15347 18751
rect 15562 18748 15568 18760
rect 15523 18720 15568 18748
rect 15289 18711 15347 18717
rect 15304 18680 15332 18711
rect 15562 18708 15568 18720
rect 15620 18748 15626 18760
rect 16117 18751 16175 18757
rect 16117 18748 16129 18751
rect 15620 18720 16129 18748
rect 15620 18708 15626 18720
rect 16117 18717 16129 18720
rect 16163 18717 16175 18751
rect 18046 18748 18052 18760
rect 18007 18720 18052 18748
rect 16117 18711 16175 18717
rect 18046 18708 18052 18720
rect 18104 18708 18110 18760
rect 18340 18757 18368 18788
rect 19288 18776 19294 18788
rect 19346 18776 19352 18828
rect 19426 18776 19432 18828
rect 19484 18776 19490 18828
rect 19527 18788 19748 18816
rect 18325 18751 18383 18757
rect 18325 18717 18337 18751
rect 18371 18717 18383 18751
rect 18325 18711 18383 18717
rect 18414 18708 18420 18760
rect 18472 18748 18478 18760
rect 18601 18751 18659 18757
rect 18601 18748 18613 18751
rect 18472 18720 18613 18748
rect 18472 18708 18478 18720
rect 18601 18717 18613 18720
rect 18647 18717 18659 18751
rect 18601 18711 18659 18717
rect 18782 18708 18788 18760
rect 18840 18748 18846 18760
rect 18877 18751 18935 18757
rect 18877 18748 18889 18751
rect 18840 18720 18889 18748
rect 18840 18708 18846 18720
rect 18877 18717 18889 18720
rect 18923 18717 18935 18751
rect 18877 18711 18935 18717
rect 18966 18708 18972 18760
rect 19024 18748 19030 18760
rect 19527 18748 19555 18788
rect 19720 18757 19748 18788
rect 19024 18720 19555 18748
rect 19705 18751 19763 18757
rect 19613 18727 19671 18733
rect 19024 18708 19030 18720
rect 19613 18693 19625 18727
rect 19659 18693 19671 18727
rect 19705 18717 19717 18751
rect 19751 18717 19763 18751
rect 19978 18748 19984 18760
rect 19939 18720 19984 18748
rect 19705 18711 19763 18717
rect 19978 18708 19984 18720
rect 20036 18708 20042 18760
rect 20088 18748 20116 18924
rect 20441 18921 20453 18955
rect 20487 18952 20499 18955
rect 22278 18952 22284 18964
rect 20487 18924 22284 18952
rect 20487 18921 20499 18924
rect 20441 18915 20499 18921
rect 22278 18912 22284 18924
rect 22336 18912 22342 18964
rect 20165 18887 20223 18893
rect 20165 18853 20177 18887
rect 20211 18884 20223 18887
rect 20714 18884 20720 18896
rect 20211 18856 20720 18884
rect 20211 18853 20223 18856
rect 20165 18847 20223 18853
rect 20714 18844 20720 18856
rect 20772 18844 20778 18896
rect 20530 18776 20536 18828
rect 20588 18776 20594 18828
rect 20257 18751 20315 18757
rect 20257 18748 20269 18751
rect 20088 18720 20269 18748
rect 20257 18717 20269 18720
rect 20303 18717 20315 18751
rect 20548 18748 20576 18776
rect 20625 18751 20683 18757
rect 20625 18748 20637 18751
rect 20548 18720 20637 18748
rect 20257 18711 20315 18717
rect 20625 18717 20637 18720
rect 20671 18717 20683 18751
rect 21269 18751 21327 18757
rect 21269 18748 21281 18751
rect 20625 18711 20683 18717
rect 20732 18720 21281 18748
rect 19613 18692 19671 18693
rect 15841 18683 15899 18689
rect 15841 18680 15853 18683
rect 14844 18652 15036 18680
rect 15304 18652 15853 18680
rect 14461 18643 14519 18649
rect 12897 18615 12955 18621
rect 12584 18584 12629 18612
rect 12584 18572 12590 18584
rect 12897 18581 12909 18615
rect 12943 18581 12955 18615
rect 13262 18612 13268 18624
rect 13223 18584 13268 18612
rect 12897 18575 12955 18581
rect 13262 18572 13268 18584
rect 13320 18572 13326 18624
rect 13722 18572 13728 18624
rect 13780 18612 13786 18624
rect 13817 18615 13875 18621
rect 13817 18612 13829 18615
rect 13780 18584 13829 18612
rect 13780 18572 13786 18584
rect 13817 18581 13829 18584
rect 13863 18612 13875 18615
rect 14274 18612 14280 18624
rect 13863 18584 14280 18612
rect 13863 18581 13875 18584
rect 13817 18575 13875 18581
rect 14274 18572 14280 18584
rect 14332 18572 14338 18624
rect 14642 18572 14648 18624
rect 14700 18612 14706 18624
rect 14921 18615 14979 18621
rect 14921 18612 14933 18615
rect 14700 18584 14933 18612
rect 14700 18572 14706 18584
rect 14921 18581 14933 18584
rect 14967 18581 14979 18615
rect 15008 18612 15036 18652
rect 15841 18649 15853 18652
rect 15887 18649 15899 18683
rect 15841 18643 15899 18649
rect 17773 18683 17831 18689
rect 17773 18649 17785 18683
rect 17819 18680 17831 18683
rect 17819 18652 19380 18680
rect 17819 18649 17831 18652
rect 17773 18643 17831 18649
rect 19352 18624 19380 18652
rect 19610 18640 19616 18692
rect 19668 18640 19674 18692
rect 20530 18640 20536 18692
rect 20588 18680 20594 18692
rect 20732 18680 20760 18720
rect 21269 18717 21281 18720
rect 21315 18717 21327 18751
rect 21269 18711 21327 18717
rect 20898 18680 20904 18692
rect 20588 18652 20760 18680
rect 20859 18652 20904 18680
rect 20588 18640 20594 18652
rect 20898 18640 20904 18652
rect 20956 18640 20962 18692
rect 15654 18612 15660 18624
rect 15008 18584 15660 18612
rect 14921 18575 14979 18581
rect 15654 18572 15660 18584
rect 15712 18572 15718 18624
rect 16114 18572 16120 18624
rect 16172 18612 16178 18624
rect 16209 18615 16267 18621
rect 16209 18612 16221 18615
rect 16172 18584 16221 18612
rect 16172 18572 16178 18584
rect 16209 18581 16221 18584
rect 16255 18581 16267 18615
rect 16390 18612 16396 18624
rect 16351 18584 16396 18612
rect 16209 18575 16267 18581
rect 16390 18572 16396 18584
rect 16448 18572 16454 18624
rect 17218 18612 17224 18624
rect 17179 18584 17224 18612
rect 17218 18572 17224 18584
rect 17276 18572 17282 18624
rect 18874 18572 18880 18624
rect 18932 18612 18938 18624
rect 19061 18615 19119 18621
rect 19061 18612 19073 18615
rect 18932 18584 19073 18612
rect 18932 18572 18938 18584
rect 19061 18581 19073 18584
rect 19107 18581 19119 18615
rect 19061 18575 19119 18581
rect 19150 18572 19156 18624
rect 19208 18612 19214 18624
rect 19245 18615 19303 18621
rect 19245 18612 19257 18615
rect 19208 18584 19257 18612
rect 19208 18572 19214 18584
rect 19245 18581 19257 18584
rect 19291 18581 19303 18615
rect 19245 18575 19303 18581
rect 19334 18572 19340 18624
rect 19392 18572 19398 18624
rect 19429 18615 19487 18621
rect 19429 18581 19441 18615
rect 19475 18612 19487 18615
rect 19518 18612 19524 18624
rect 19475 18584 19524 18612
rect 19475 18581 19487 18584
rect 19429 18575 19487 18581
rect 19518 18572 19524 18584
rect 19576 18572 19582 18624
rect 19889 18615 19947 18621
rect 19889 18581 19901 18615
rect 19935 18612 19947 18615
rect 20622 18612 20628 18624
rect 19935 18584 20628 18612
rect 19935 18581 19947 18584
rect 19889 18575 19947 18581
rect 20622 18572 20628 18584
rect 20680 18572 20686 18624
rect 21450 18612 21456 18624
rect 21411 18584 21456 18612
rect 21450 18572 21456 18584
rect 21508 18572 21514 18624
rect 1104 18522 22056 18544
rect 1104 18470 6148 18522
rect 6200 18470 6212 18522
rect 6264 18470 6276 18522
rect 6328 18470 6340 18522
rect 6392 18470 6404 18522
rect 6456 18470 11346 18522
rect 11398 18470 11410 18522
rect 11462 18470 11474 18522
rect 11526 18470 11538 18522
rect 11590 18470 11602 18522
rect 11654 18470 16544 18522
rect 16596 18470 16608 18522
rect 16660 18470 16672 18522
rect 16724 18470 16736 18522
rect 16788 18470 16800 18522
rect 16852 18470 21742 18522
rect 21794 18470 21806 18522
rect 21858 18470 21870 18522
rect 21922 18470 21934 18522
rect 21986 18470 21998 18522
rect 22050 18470 22056 18522
rect 1104 18448 22056 18470
rect 2501 18411 2559 18417
rect 2501 18377 2513 18411
rect 2547 18377 2559 18411
rect 3050 18408 3056 18420
rect 3011 18380 3056 18408
rect 2501 18371 2559 18377
rect 2516 18340 2544 18371
rect 3050 18368 3056 18380
rect 3108 18368 3114 18420
rect 3142 18368 3148 18420
rect 3200 18408 3206 18420
rect 3605 18411 3663 18417
rect 3200 18380 3245 18408
rect 3200 18368 3206 18380
rect 3605 18377 3617 18411
rect 3651 18408 3663 18411
rect 4062 18408 4068 18420
rect 3651 18380 4068 18408
rect 3651 18377 3663 18380
rect 3605 18371 3663 18377
rect 4062 18368 4068 18380
rect 4120 18368 4126 18420
rect 5074 18368 5080 18420
rect 5132 18408 5138 18420
rect 5721 18411 5779 18417
rect 5721 18408 5733 18411
rect 5132 18380 5733 18408
rect 5132 18368 5138 18380
rect 5721 18377 5733 18380
rect 5767 18377 5779 18411
rect 5721 18371 5779 18377
rect 1688 18312 2544 18340
rect 1688 18281 1716 18312
rect 3326 18300 3332 18352
rect 3384 18340 3390 18352
rect 3384 18312 5111 18340
rect 3384 18300 3390 18312
rect 1673 18275 1731 18281
rect 1673 18241 1685 18275
rect 1719 18241 1731 18275
rect 2038 18272 2044 18284
rect 1999 18244 2044 18272
rect 1673 18235 1731 18241
rect 2038 18232 2044 18244
rect 2096 18232 2102 18284
rect 2225 18275 2283 18281
rect 2225 18241 2237 18275
rect 2271 18272 2283 18275
rect 2406 18272 2412 18284
rect 2271 18244 2412 18272
rect 2271 18241 2283 18244
rect 2225 18235 2283 18241
rect 2406 18232 2412 18244
rect 2464 18232 2470 18284
rect 2498 18232 2504 18284
rect 2556 18272 2562 18284
rect 2685 18275 2743 18281
rect 2685 18272 2697 18275
rect 2556 18244 2697 18272
rect 2556 18232 2562 18244
rect 2685 18241 2697 18244
rect 2731 18241 2743 18275
rect 2685 18235 2743 18241
rect 3050 18232 3056 18284
rect 3108 18272 3114 18284
rect 3344 18272 3372 18300
rect 3108 18244 3372 18272
rect 3108 18232 3114 18244
rect 4706 18232 4712 18284
rect 4764 18281 4770 18284
rect 4764 18272 4776 18281
rect 4764 18244 4809 18272
rect 4764 18235 4776 18244
rect 4764 18232 4770 18235
rect 2958 18204 2964 18216
rect 2919 18176 2964 18204
rect 2958 18164 2964 18176
rect 3016 18164 3022 18216
rect 4985 18207 5043 18213
rect 4985 18173 4997 18207
rect 5031 18173 5043 18207
rect 4985 18167 5043 18173
rect 1854 18136 1860 18148
rect 1815 18108 1860 18136
rect 1854 18096 1860 18108
rect 1912 18096 1918 18148
rect 3513 18139 3571 18145
rect 3513 18105 3525 18139
rect 3559 18136 3571 18139
rect 3970 18136 3976 18148
rect 3559 18108 3976 18136
rect 3559 18105 3571 18108
rect 3513 18099 3571 18105
rect 3970 18096 3976 18108
rect 4028 18096 4034 18148
rect 1486 18068 1492 18080
rect 1447 18040 1492 18068
rect 1486 18028 1492 18040
rect 1544 18028 1550 18080
rect 2406 18068 2412 18080
rect 2367 18040 2412 18068
rect 2406 18028 2412 18040
rect 2464 18028 2470 18080
rect 4062 18028 4068 18080
rect 4120 18068 4126 18080
rect 5000 18068 5028 18167
rect 5083 18136 5111 18312
rect 5258 18232 5264 18284
rect 5316 18272 5322 18284
rect 5442 18272 5448 18284
rect 5316 18244 5448 18272
rect 5316 18232 5322 18244
rect 5442 18232 5448 18244
rect 5500 18232 5506 18284
rect 5534 18204 5540 18216
rect 5495 18176 5540 18204
rect 5534 18164 5540 18176
rect 5592 18164 5598 18216
rect 5736 18204 5764 18371
rect 5810 18368 5816 18420
rect 5868 18368 5874 18420
rect 5902 18368 5908 18420
rect 5960 18408 5966 18420
rect 6181 18411 6239 18417
rect 6181 18408 6193 18411
rect 5960 18380 6193 18408
rect 5960 18368 5966 18380
rect 6181 18377 6193 18380
rect 6227 18377 6239 18411
rect 6181 18371 6239 18377
rect 6365 18411 6423 18417
rect 6365 18377 6377 18411
rect 6411 18377 6423 18411
rect 6365 18371 6423 18377
rect 5828 18340 5856 18368
rect 6380 18340 6408 18371
rect 7282 18368 7288 18420
rect 7340 18408 7346 18420
rect 7745 18411 7803 18417
rect 7745 18408 7757 18411
rect 7340 18380 7757 18408
rect 7340 18368 7346 18380
rect 7745 18377 7757 18380
rect 7791 18377 7803 18411
rect 7745 18371 7803 18377
rect 7834 18368 7840 18420
rect 7892 18408 7898 18420
rect 8113 18411 8171 18417
rect 8113 18408 8125 18411
rect 7892 18380 8125 18408
rect 7892 18368 7898 18380
rect 8113 18377 8125 18380
rect 8159 18377 8171 18411
rect 8113 18371 8171 18377
rect 8294 18368 8300 18420
rect 8352 18408 8358 18420
rect 8941 18411 8999 18417
rect 8941 18408 8953 18411
rect 8352 18380 8953 18408
rect 8352 18368 8358 18380
rect 8941 18377 8953 18380
rect 8987 18377 8999 18411
rect 9306 18408 9312 18420
rect 9267 18380 9312 18408
rect 8941 18371 8999 18377
rect 9306 18368 9312 18380
rect 9364 18368 9370 18420
rect 10134 18408 10140 18420
rect 10095 18380 10140 18408
rect 10134 18368 10140 18380
rect 10192 18368 10198 18420
rect 10597 18411 10655 18417
rect 10597 18377 10609 18411
rect 10643 18377 10655 18411
rect 10597 18371 10655 18377
rect 5828 18312 6408 18340
rect 6825 18343 6883 18349
rect 6825 18309 6837 18343
rect 6871 18340 6883 18343
rect 6914 18340 6920 18352
rect 6871 18312 6920 18340
rect 6871 18309 6883 18312
rect 6825 18303 6883 18309
rect 6914 18300 6920 18312
rect 6972 18300 6978 18352
rect 7190 18300 7196 18352
rect 7248 18340 7254 18352
rect 7466 18340 7472 18352
rect 7248 18312 7472 18340
rect 7248 18300 7254 18312
rect 7466 18300 7472 18312
rect 7524 18300 7530 18352
rect 7650 18300 7656 18352
rect 7708 18340 7714 18352
rect 7708 18312 8708 18340
rect 7708 18300 7714 18312
rect 5810 18232 5816 18284
rect 5868 18272 5874 18284
rect 5868 18244 5913 18272
rect 5868 18232 5874 18244
rect 6546 18232 6552 18284
rect 6604 18272 6610 18284
rect 6733 18275 6791 18281
rect 6733 18272 6745 18275
rect 6604 18244 6745 18272
rect 6604 18232 6610 18244
rect 6733 18241 6745 18244
rect 6779 18272 6791 18275
rect 8680 18272 8708 18312
rect 8754 18300 8760 18352
rect 8812 18340 8818 18352
rect 8812 18312 10364 18340
rect 8812 18300 8818 18312
rect 6779 18244 7972 18272
rect 8680 18244 9444 18272
rect 6779 18241 6791 18244
rect 6733 18235 6791 18241
rect 6178 18204 6184 18216
rect 5736 18176 6184 18204
rect 6178 18164 6184 18176
rect 6236 18164 6242 18216
rect 6362 18164 6368 18216
rect 6420 18204 6426 18216
rect 6917 18207 6975 18213
rect 6917 18204 6929 18207
rect 6420 18176 6929 18204
rect 6420 18164 6426 18176
rect 6917 18173 6929 18176
rect 6963 18173 6975 18207
rect 7944 18204 7972 18244
rect 8205 18207 8263 18213
rect 8205 18204 8217 18207
rect 7944 18176 8217 18204
rect 6917 18167 6975 18173
rect 8205 18173 8217 18176
rect 8251 18173 8263 18207
rect 8205 18167 8263 18173
rect 6822 18136 6828 18148
rect 5083 18108 6828 18136
rect 6822 18096 6828 18108
rect 6880 18096 6886 18148
rect 7098 18096 7104 18148
rect 7156 18136 7162 18148
rect 7285 18139 7343 18145
rect 7285 18136 7297 18139
rect 7156 18108 7297 18136
rect 7156 18096 7162 18108
rect 7285 18105 7297 18108
rect 7331 18105 7343 18139
rect 7285 18099 7343 18105
rect 5077 18071 5135 18077
rect 5077 18068 5089 18071
rect 4120 18040 5089 18068
rect 4120 18028 4126 18040
rect 5077 18037 5089 18040
rect 5123 18037 5135 18071
rect 5077 18031 5135 18037
rect 5258 18028 5264 18080
rect 5316 18068 5322 18080
rect 5994 18068 6000 18080
rect 5316 18040 6000 18068
rect 5316 18028 5322 18040
rect 5994 18028 6000 18040
rect 6052 18028 6058 18080
rect 6270 18028 6276 18080
rect 6328 18068 6334 18080
rect 7742 18068 7748 18080
rect 6328 18040 7748 18068
rect 6328 18028 6334 18040
rect 7742 18028 7748 18040
rect 7800 18028 7806 18080
rect 8220 18068 8248 18167
rect 8294 18164 8300 18216
rect 8352 18204 8358 18216
rect 8352 18176 8397 18204
rect 8352 18164 8358 18176
rect 8570 18164 8576 18216
rect 8628 18204 8634 18216
rect 8665 18207 8723 18213
rect 8665 18204 8677 18207
rect 8628 18176 8677 18204
rect 8628 18164 8634 18176
rect 8665 18173 8677 18176
rect 8711 18173 8723 18207
rect 8665 18167 8723 18173
rect 8754 18164 8760 18216
rect 8812 18204 8818 18216
rect 8849 18207 8907 18213
rect 8849 18204 8861 18207
rect 8812 18176 8861 18204
rect 8812 18164 8818 18176
rect 8849 18173 8861 18176
rect 8895 18173 8907 18207
rect 9416 18204 9444 18244
rect 9490 18232 9496 18284
rect 9548 18272 9554 18284
rect 9585 18275 9643 18281
rect 9585 18272 9597 18275
rect 9548 18244 9597 18272
rect 9548 18232 9554 18244
rect 9585 18241 9597 18244
rect 9631 18241 9643 18275
rect 9858 18272 9864 18284
rect 9819 18244 9864 18272
rect 9585 18235 9643 18241
rect 9858 18232 9864 18244
rect 9916 18232 9922 18284
rect 10336 18281 10364 18312
rect 10321 18275 10379 18281
rect 10321 18241 10333 18275
rect 10367 18241 10379 18275
rect 10321 18235 10379 18241
rect 10410 18232 10416 18284
rect 10468 18272 10474 18284
rect 10612 18272 10640 18371
rect 10686 18368 10692 18420
rect 10744 18408 10750 18420
rect 10965 18411 11023 18417
rect 10965 18408 10977 18411
rect 10744 18380 10977 18408
rect 10744 18368 10750 18380
rect 10965 18377 10977 18380
rect 11011 18377 11023 18411
rect 11238 18408 11244 18420
rect 11199 18380 11244 18408
rect 10965 18371 11023 18377
rect 11238 18368 11244 18380
rect 11296 18368 11302 18420
rect 11882 18408 11888 18420
rect 11843 18380 11888 18408
rect 11882 18368 11888 18380
rect 11940 18368 11946 18420
rect 11974 18368 11980 18420
rect 12032 18408 12038 18420
rect 12032 18380 12480 18408
rect 12032 18368 12038 18380
rect 12253 18343 12311 18349
rect 12253 18309 12265 18343
rect 12299 18340 12311 18343
rect 12342 18340 12348 18352
rect 12299 18312 12348 18340
rect 12299 18309 12311 18312
rect 12253 18303 12311 18309
rect 12342 18300 12348 18312
rect 12400 18300 12406 18352
rect 12452 18340 12480 18380
rect 12526 18368 12532 18420
rect 12584 18408 12590 18420
rect 13541 18411 13599 18417
rect 13541 18408 13553 18411
rect 12584 18380 13553 18408
rect 12584 18368 12590 18380
rect 13541 18377 13553 18380
rect 13587 18377 13599 18411
rect 13541 18371 13599 18377
rect 13630 18368 13636 18420
rect 13688 18408 13694 18420
rect 14185 18411 14243 18417
rect 14185 18408 14197 18411
rect 13688 18380 14197 18408
rect 13688 18368 13694 18380
rect 14185 18377 14197 18380
rect 14231 18377 14243 18411
rect 14642 18408 14648 18420
rect 14603 18380 14648 18408
rect 14185 18371 14243 18377
rect 14642 18368 14648 18380
rect 14700 18368 14706 18420
rect 15378 18408 15384 18420
rect 15339 18380 15384 18408
rect 15378 18368 15384 18380
rect 15436 18368 15442 18420
rect 18598 18368 18604 18420
rect 18656 18408 18662 18420
rect 18877 18411 18935 18417
rect 18877 18408 18889 18411
rect 18656 18380 18889 18408
rect 18656 18368 18662 18380
rect 18877 18377 18889 18380
rect 18923 18377 18935 18411
rect 18877 18371 18935 18377
rect 19337 18411 19395 18417
rect 19337 18377 19349 18411
rect 19383 18408 19395 18411
rect 19610 18408 19616 18420
rect 19383 18380 19616 18408
rect 19383 18377 19395 18380
rect 19337 18371 19395 18377
rect 19610 18368 19616 18380
rect 19668 18368 19674 18420
rect 19794 18408 19800 18420
rect 19755 18380 19800 18408
rect 19794 18368 19800 18380
rect 19852 18368 19858 18420
rect 19886 18368 19892 18420
rect 19944 18368 19950 18420
rect 20622 18408 20628 18420
rect 20364 18380 20628 18408
rect 14001 18343 14059 18349
rect 14001 18340 14013 18343
rect 12452 18312 14013 18340
rect 14001 18309 14013 18312
rect 14047 18309 14059 18343
rect 14001 18303 14059 18309
rect 14274 18300 14280 18352
rect 14332 18340 14338 18352
rect 18506 18340 18512 18352
rect 14332 18312 18512 18340
rect 14332 18300 14338 18312
rect 18506 18300 18512 18312
rect 18564 18300 18570 18352
rect 18785 18343 18843 18349
rect 18785 18309 18797 18343
rect 18831 18340 18843 18343
rect 19904 18340 19932 18368
rect 18831 18312 19932 18340
rect 18831 18309 18843 18312
rect 18785 18303 18843 18309
rect 10781 18275 10839 18281
rect 10781 18272 10793 18275
rect 10468 18244 10513 18272
rect 10612 18244 10793 18272
rect 10468 18232 10474 18244
rect 10781 18241 10793 18244
rect 10827 18241 10839 18275
rect 10781 18235 10839 18241
rect 11057 18275 11115 18281
rect 11057 18241 11069 18275
rect 11103 18241 11115 18275
rect 11057 18235 11115 18241
rect 9950 18204 9956 18216
rect 9416 18176 9956 18204
rect 8849 18167 8907 18173
rect 9950 18164 9956 18176
rect 10008 18164 10014 18216
rect 11072 18204 11100 18235
rect 11698 18232 11704 18284
rect 11756 18272 11762 18284
rect 12158 18272 12164 18284
rect 11756 18244 12164 18272
rect 11756 18232 11762 18244
rect 12158 18232 12164 18244
rect 12216 18272 12222 18284
rect 13078 18272 13084 18284
rect 12216 18244 12572 18272
rect 13039 18244 13084 18272
rect 12216 18232 12222 18244
rect 10060 18176 11100 18204
rect 8386 18096 8392 18148
rect 8444 18136 8450 18148
rect 10060 18145 10088 18176
rect 11238 18164 11244 18216
rect 11296 18204 11302 18216
rect 12544 18213 12572 18244
rect 13078 18232 13084 18244
rect 13136 18232 13142 18284
rect 14737 18275 14795 18281
rect 14737 18241 14749 18275
rect 14783 18272 14795 18275
rect 15470 18272 15476 18284
rect 14783 18244 15476 18272
rect 14783 18241 14795 18244
rect 14737 18235 14795 18241
rect 15470 18232 15476 18244
rect 15528 18232 15534 18284
rect 19245 18275 19303 18281
rect 19245 18241 19257 18275
rect 19291 18241 19303 18275
rect 19245 18235 19303 18241
rect 12345 18207 12403 18213
rect 12345 18204 12357 18207
rect 11296 18176 12357 18204
rect 11296 18164 11302 18176
rect 12345 18173 12357 18176
rect 12391 18173 12403 18207
rect 12345 18167 12403 18173
rect 12529 18207 12587 18213
rect 12529 18173 12541 18207
rect 12575 18204 12587 18207
rect 13170 18204 13176 18216
rect 12575 18176 12848 18204
rect 13131 18176 13176 18204
rect 12575 18173 12587 18176
rect 12529 18167 12587 18173
rect 10045 18139 10103 18145
rect 8444 18108 9996 18136
rect 8444 18096 8450 18108
rect 9306 18068 9312 18080
rect 8220 18040 9312 18068
rect 9306 18028 9312 18040
rect 9364 18028 9370 18080
rect 9674 18028 9680 18080
rect 9732 18068 9738 18080
rect 9968 18068 9996 18108
rect 10045 18105 10057 18139
rect 10091 18105 10103 18139
rect 10045 18099 10103 18105
rect 10778 18096 10784 18148
rect 10836 18136 10842 18148
rect 11609 18139 11667 18145
rect 10836 18108 11560 18136
rect 10836 18096 10842 18108
rect 11238 18068 11244 18080
rect 9732 18040 9777 18068
rect 9968 18040 11244 18068
rect 9732 18028 9738 18040
rect 11238 18028 11244 18040
rect 11296 18028 11302 18080
rect 11532 18068 11560 18108
rect 11609 18105 11621 18139
rect 11655 18136 11667 18139
rect 11655 18108 12020 18136
rect 11655 18105 11667 18108
rect 11609 18099 11667 18105
rect 11701 18071 11759 18077
rect 11701 18068 11713 18071
rect 11532 18040 11713 18068
rect 11701 18037 11713 18040
rect 11747 18068 11759 18071
rect 11882 18068 11888 18080
rect 11747 18040 11888 18068
rect 11747 18037 11759 18040
rect 11701 18031 11759 18037
rect 11882 18028 11888 18040
rect 11940 18028 11946 18080
rect 11992 18068 12020 18108
rect 12066 18096 12072 18148
rect 12124 18136 12130 18148
rect 12713 18139 12771 18145
rect 12713 18136 12725 18139
rect 12124 18108 12725 18136
rect 12124 18096 12130 18108
rect 12713 18105 12725 18108
rect 12759 18105 12771 18139
rect 12820 18136 12848 18176
rect 13170 18164 13176 18176
rect 13228 18164 13234 18216
rect 13265 18207 13323 18213
rect 13265 18173 13277 18207
rect 13311 18173 13323 18207
rect 13265 18167 13323 18173
rect 14553 18207 14611 18213
rect 14553 18173 14565 18207
rect 14599 18204 14611 18207
rect 14918 18204 14924 18216
rect 14599 18176 14924 18204
rect 14599 18173 14611 18176
rect 14553 18167 14611 18173
rect 13280 18136 13308 18167
rect 14918 18164 14924 18176
rect 14976 18164 14982 18216
rect 16114 18204 16120 18216
rect 15028 18176 16120 18204
rect 12820 18108 13308 18136
rect 12713 18099 12771 18105
rect 13630 18096 13636 18148
rect 13688 18136 13694 18148
rect 15028 18136 15056 18176
rect 16114 18164 16120 18176
rect 16172 18164 16178 18216
rect 19260 18204 19288 18235
rect 19334 18232 19340 18284
rect 19392 18272 19398 18284
rect 19521 18275 19579 18281
rect 19521 18272 19533 18275
rect 19392 18244 19533 18272
rect 19392 18232 19398 18244
rect 19521 18241 19533 18244
rect 19567 18241 19579 18275
rect 19521 18235 19579 18241
rect 19613 18275 19671 18281
rect 19613 18241 19625 18275
rect 19659 18272 19671 18275
rect 19889 18275 19947 18281
rect 19889 18272 19901 18275
rect 19659 18244 19901 18272
rect 19659 18241 19671 18244
rect 19613 18235 19671 18241
rect 19889 18241 19901 18244
rect 19935 18272 19947 18275
rect 20162 18272 20168 18284
rect 19935 18244 20168 18272
rect 19935 18241 19947 18244
rect 19889 18235 19947 18241
rect 20162 18232 20168 18244
rect 20220 18232 20226 18284
rect 20364 18281 20392 18380
rect 20622 18368 20628 18380
rect 20680 18368 20686 18420
rect 20809 18411 20867 18417
rect 20809 18377 20821 18411
rect 20855 18408 20867 18411
rect 21266 18408 21272 18420
rect 20855 18380 21272 18408
rect 20855 18377 20867 18380
rect 20809 18371 20867 18377
rect 21266 18368 21272 18380
rect 21324 18368 21330 18420
rect 20625 18299 20683 18305
rect 20349 18275 20407 18281
rect 20349 18241 20361 18275
rect 20395 18241 20407 18275
rect 20625 18265 20637 18299
rect 20671 18296 20683 18299
rect 20671 18284 20852 18296
rect 20671 18268 20812 18284
rect 20671 18265 20683 18268
rect 20625 18259 20683 18265
rect 20349 18235 20407 18241
rect 20806 18232 20812 18268
rect 20864 18232 20870 18284
rect 20901 18275 20959 18281
rect 20901 18241 20913 18275
rect 20947 18272 20959 18275
rect 20990 18272 20996 18284
rect 20947 18244 20996 18272
rect 20947 18241 20959 18244
rect 20901 18235 20959 18241
rect 20990 18232 20996 18244
rect 21048 18232 21054 18284
rect 21082 18232 21088 18284
rect 21140 18232 21146 18284
rect 21266 18272 21272 18284
rect 21227 18244 21272 18272
rect 21266 18232 21272 18244
rect 21324 18232 21330 18284
rect 20257 18207 20315 18213
rect 20257 18204 20269 18207
rect 19260 18176 20269 18204
rect 20257 18173 20269 18176
rect 20303 18204 20315 18207
rect 21100 18204 21128 18232
rect 20303 18176 21128 18204
rect 20303 18173 20315 18176
rect 20257 18167 20315 18173
rect 13688 18108 15056 18136
rect 15105 18139 15163 18145
rect 13688 18096 13694 18108
rect 15105 18105 15117 18139
rect 15151 18136 15163 18139
rect 16206 18136 16212 18148
rect 15151 18108 16212 18136
rect 15151 18105 15163 18108
rect 15105 18099 15163 18105
rect 16206 18096 16212 18108
rect 16264 18096 16270 18148
rect 18414 18096 18420 18148
rect 18472 18136 18478 18148
rect 19061 18139 19119 18145
rect 19061 18136 19073 18139
rect 18472 18108 19073 18136
rect 18472 18096 18478 18108
rect 19061 18105 19073 18108
rect 19107 18136 19119 18139
rect 19242 18136 19248 18148
rect 19107 18108 19248 18136
rect 19107 18105 19119 18108
rect 19061 18099 19119 18105
rect 19242 18096 19248 18108
rect 19300 18136 19306 18148
rect 20162 18136 20168 18148
rect 19300 18108 20168 18136
rect 19300 18096 19306 18108
rect 20162 18096 20168 18108
rect 20220 18096 20226 18148
rect 20533 18139 20591 18145
rect 20533 18105 20545 18139
rect 20579 18136 20591 18139
rect 20622 18136 20628 18148
rect 20579 18108 20628 18136
rect 20579 18105 20591 18108
rect 20533 18099 20591 18105
rect 20622 18096 20628 18108
rect 20680 18096 20686 18148
rect 21082 18136 21088 18148
rect 21043 18108 21088 18136
rect 21082 18096 21088 18108
rect 21140 18096 21146 18148
rect 22186 18136 22192 18148
rect 21284 18108 22192 18136
rect 12250 18068 12256 18080
rect 11992 18040 12256 18068
rect 12250 18028 12256 18040
rect 12308 18028 12314 18080
rect 12434 18028 12440 18080
rect 12492 18068 12498 18080
rect 13817 18071 13875 18077
rect 13817 18068 13829 18071
rect 12492 18040 13829 18068
rect 12492 18028 12498 18040
rect 13817 18037 13829 18040
rect 13863 18037 13875 18071
rect 15286 18068 15292 18080
rect 15247 18040 15292 18068
rect 13817 18031 13875 18037
rect 15286 18028 15292 18040
rect 15344 18028 15350 18080
rect 15562 18068 15568 18080
rect 15523 18040 15568 18068
rect 15562 18028 15568 18040
rect 15620 18028 15626 18080
rect 20073 18071 20131 18077
rect 20073 18037 20085 18071
rect 20119 18068 20131 18071
rect 21284 18068 21312 18108
rect 22186 18096 22192 18108
rect 22244 18096 22250 18148
rect 21450 18068 21456 18080
rect 20119 18040 21312 18068
rect 21411 18040 21456 18068
rect 20119 18037 20131 18040
rect 20073 18031 20131 18037
rect 21450 18028 21456 18040
rect 21508 18028 21514 18080
rect 1104 17978 21896 18000
rect 1104 17926 3549 17978
rect 3601 17926 3613 17978
rect 3665 17926 3677 17978
rect 3729 17926 3741 17978
rect 3793 17926 3805 17978
rect 3857 17926 8747 17978
rect 8799 17926 8811 17978
rect 8863 17926 8875 17978
rect 8927 17926 8939 17978
rect 8991 17926 9003 17978
rect 9055 17926 13945 17978
rect 13997 17926 14009 17978
rect 14061 17926 14073 17978
rect 14125 17926 14137 17978
rect 14189 17926 14201 17978
rect 14253 17926 19143 17978
rect 19195 17926 19207 17978
rect 19259 17926 19271 17978
rect 19323 17926 19335 17978
rect 19387 17926 19399 17978
rect 19451 17926 21896 17978
rect 1104 17904 21896 17926
rect 1578 17824 1584 17876
rect 1636 17824 1642 17876
rect 2222 17824 2228 17876
rect 2280 17864 2286 17876
rect 2409 17867 2467 17873
rect 2409 17864 2421 17867
rect 2280 17836 2421 17864
rect 2280 17824 2286 17836
rect 2409 17833 2421 17836
rect 2455 17833 2467 17867
rect 2409 17827 2467 17833
rect 2777 17867 2835 17873
rect 2777 17833 2789 17867
rect 2823 17864 2835 17867
rect 5258 17864 5264 17876
rect 2823 17836 5264 17864
rect 2823 17833 2835 17836
rect 2777 17827 2835 17833
rect 5258 17824 5264 17836
rect 5316 17824 5322 17876
rect 5534 17824 5540 17876
rect 5592 17864 5598 17876
rect 6457 17867 6515 17873
rect 6457 17864 6469 17867
rect 5592 17836 6469 17864
rect 5592 17824 5598 17836
rect 6457 17833 6469 17836
rect 6503 17864 6515 17867
rect 7282 17864 7288 17876
rect 6503 17836 7288 17864
rect 6503 17833 6515 17836
rect 6457 17827 6515 17833
rect 7282 17824 7288 17836
rect 7340 17824 7346 17876
rect 8021 17867 8079 17873
rect 8021 17833 8033 17867
rect 8067 17864 8079 17867
rect 8110 17864 8116 17876
rect 8067 17836 8116 17864
rect 8067 17833 8079 17836
rect 8021 17827 8079 17833
rect 8110 17824 8116 17836
rect 8168 17824 8174 17876
rect 8941 17867 8999 17873
rect 8941 17833 8953 17867
rect 8987 17864 8999 17867
rect 9398 17864 9404 17876
rect 8987 17836 9404 17864
rect 8987 17833 8999 17836
rect 8941 17827 8999 17833
rect 9398 17824 9404 17836
rect 9456 17824 9462 17876
rect 9766 17824 9772 17876
rect 9824 17864 9830 17876
rect 9953 17867 10011 17873
rect 9953 17864 9965 17867
rect 9824 17836 9965 17864
rect 9824 17824 9830 17836
rect 9953 17833 9965 17836
rect 9999 17864 10011 17867
rect 10226 17864 10232 17876
rect 9999 17836 10232 17864
rect 9999 17833 10011 17836
rect 9953 17827 10011 17833
rect 10226 17824 10232 17836
rect 10284 17824 10290 17876
rect 10686 17824 10692 17876
rect 10744 17864 10750 17876
rect 12989 17867 13047 17873
rect 10744 17836 12434 17864
rect 10744 17824 10750 17836
rect 1596 17796 1624 17824
rect 3326 17796 3332 17808
rect 1596 17768 2728 17796
rect 1578 17688 1584 17740
rect 1636 17728 1642 17740
rect 1636 17700 2636 17728
rect 1636 17688 1642 17700
rect 1670 17660 1676 17672
rect 1631 17632 1676 17660
rect 1670 17620 1676 17632
rect 1728 17620 1734 17672
rect 2041 17663 2099 17669
rect 2041 17629 2053 17663
rect 2087 17660 2099 17663
rect 2087 17632 2176 17660
rect 2087 17629 2099 17632
rect 2041 17623 2099 17629
rect 1486 17524 1492 17536
rect 1447 17496 1492 17524
rect 1486 17484 1492 17496
rect 1544 17484 1550 17536
rect 1854 17524 1860 17536
rect 1815 17496 1860 17524
rect 1854 17484 1860 17496
rect 1912 17484 1918 17536
rect 2148 17533 2176 17632
rect 2222 17620 2228 17672
rect 2280 17660 2286 17672
rect 2608 17669 2636 17700
rect 2317 17663 2375 17669
rect 2317 17660 2329 17663
rect 2280 17632 2329 17660
rect 2280 17620 2286 17632
rect 2317 17629 2329 17632
rect 2363 17629 2375 17663
rect 2317 17623 2375 17629
rect 2593 17663 2651 17669
rect 2593 17629 2605 17663
rect 2639 17629 2651 17663
rect 2700 17660 2728 17768
rect 3068 17768 3332 17796
rect 3068 17737 3096 17768
rect 3326 17756 3332 17768
rect 3384 17756 3390 17808
rect 3605 17799 3663 17805
rect 3605 17765 3617 17799
rect 3651 17796 3663 17799
rect 3651 17768 4936 17796
rect 3651 17765 3663 17768
rect 3605 17759 3663 17765
rect 3053 17731 3111 17737
rect 3053 17697 3065 17731
rect 3099 17697 3111 17731
rect 3053 17691 3111 17697
rect 3234 17688 3240 17740
rect 3292 17728 3298 17740
rect 3694 17728 3700 17740
rect 3292 17700 3700 17728
rect 3292 17688 3298 17700
rect 3694 17688 3700 17700
rect 3752 17688 3758 17740
rect 3878 17660 3884 17672
rect 2700 17632 3884 17660
rect 2593 17623 2651 17629
rect 3878 17620 3884 17632
rect 3936 17620 3942 17672
rect 3973 17663 4031 17669
rect 3973 17629 3985 17663
rect 4019 17660 4031 17663
rect 4338 17660 4344 17672
rect 4019 17632 4344 17660
rect 4019 17629 4031 17632
rect 3973 17623 4031 17629
rect 4338 17620 4344 17632
rect 4396 17620 4402 17672
rect 4433 17663 4491 17669
rect 4433 17629 4445 17663
rect 4479 17660 4491 17663
rect 4798 17660 4804 17672
rect 4479 17632 4804 17660
rect 4479 17629 4491 17632
rect 4433 17623 4491 17629
rect 4798 17620 4804 17632
rect 4856 17620 4862 17672
rect 4908 17660 4936 17768
rect 5994 17756 6000 17808
rect 6052 17756 6058 17808
rect 6181 17799 6239 17805
rect 6181 17765 6193 17799
rect 6227 17796 6239 17799
rect 7469 17799 7527 17805
rect 6227 17768 7420 17796
rect 6227 17765 6239 17768
rect 6181 17759 6239 17765
rect 5902 17728 5908 17740
rect 5863 17700 5908 17728
rect 5902 17688 5908 17700
rect 5960 17688 5966 17740
rect 6012 17669 6040 17756
rect 6917 17731 6975 17737
rect 6917 17697 6929 17731
rect 6963 17697 6975 17731
rect 7392 17728 7420 17768
rect 7469 17765 7481 17799
rect 7515 17796 7527 17799
rect 8386 17796 8392 17808
rect 7515 17768 8392 17796
rect 7515 17765 7527 17768
rect 7469 17759 7527 17765
rect 8386 17756 8392 17768
rect 8444 17756 8450 17808
rect 11517 17799 11575 17805
rect 11517 17796 11529 17799
rect 11072 17768 11529 17796
rect 8110 17728 8116 17740
rect 7392 17700 8116 17728
rect 6917 17691 6975 17697
rect 5997 17663 6055 17669
rect 4908 17632 5957 17660
rect 3326 17552 3332 17604
rect 3384 17592 3390 17604
rect 3602 17592 3608 17604
rect 3384 17564 3608 17592
rect 3384 17552 3390 17564
rect 3602 17552 3608 17564
rect 3660 17552 3666 17604
rect 3694 17552 3700 17604
rect 3752 17592 3758 17604
rect 5258 17592 5264 17604
rect 3752 17564 5264 17592
rect 3752 17552 3758 17564
rect 5258 17552 5264 17564
rect 5316 17552 5322 17604
rect 5626 17552 5632 17604
rect 5684 17601 5690 17604
rect 5684 17592 5696 17601
rect 5929 17592 5957 17632
rect 5997 17629 6009 17663
rect 6043 17629 6055 17663
rect 5997 17623 6055 17629
rect 6086 17620 6092 17672
rect 6144 17660 6150 17672
rect 6362 17660 6368 17672
rect 6144 17632 6368 17660
rect 6144 17620 6150 17632
rect 6362 17620 6368 17632
rect 6420 17620 6426 17672
rect 6932 17660 6960 17691
rect 8110 17688 8116 17700
rect 8168 17688 8174 17740
rect 8570 17728 8576 17740
rect 8531 17700 8576 17728
rect 8570 17688 8576 17700
rect 8628 17728 8634 17740
rect 8938 17728 8944 17740
rect 8628 17700 8944 17728
rect 8628 17688 8634 17700
rect 8938 17688 8944 17700
rect 8996 17728 9002 17740
rect 9493 17731 9551 17737
rect 9493 17728 9505 17731
rect 8996 17700 9505 17728
rect 8996 17688 9002 17700
rect 9493 17697 9505 17700
rect 9539 17697 9551 17731
rect 9493 17691 9551 17697
rect 10045 17663 10103 17669
rect 6932 17632 9996 17660
rect 6270 17592 6276 17604
rect 5684 17564 5729 17592
rect 5929 17564 6276 17592
rect 5684 17555 5696 17564
rect 5684 17552 5690 17555
rect 6270 17552 6276 17564
rect 6328 17552 6334 17604
rect 6914 17552 6920 17604
rect 6972 17592 6978 17604
rect 7101 17595 7159 17601
rect 7101 17592 7113 17595
rect 6972 17564 7113 17592
rect 6972 17552 6978 17564
rect 7101 17561 7113 17564
rect 7147 17561 7159 17595
rect 7101 17555 7159 17561
rect 7929 17595 7987 17601
rect 7929 17561 7941 17595
rect 7975 17592 7987 17595
rect 8389 17595 8447 17601
rect 8389 17592 8401 17595
rect 7975 17564 8401 17592
rect 7975 17561 7987 17564
rect 7929 17555 7987 17561
rect 8389 17561 8401 17564
rect 8435 17561 8447 17595
rect 8389 17555 8447 17561
rect 9401 17595 9459 17601
rect 9401 17561 9413 17595
rect 9447 17592 9459 17595
rect 9766 17592 9772 17604
rect 9447 17564 9772 17592
rect 9447 17561 9459 17564
rect 9401 17555 9459 17561
rect 9766 17552 9772 17564
rect 9824 17552 9830 17604
rect 2133 17527 2191 17533
rect 2133 17493 2145 17527
rect 2179 17493 2191 17527
rect 3142 17524 3148 17536
rect 3103 17496 3148 17524
rect 2133 17487 2191 17493
rect 3142 17484 3148 17496
rect 3200 17484 3206 17536
rect 3234 17484 3240 17536
rect 3292 17524 3298 17536
rect 3786 17524 3792 17536
rect 3292 17496 3337 17524
rect 3747 17496 3792 17524
rect 3292 17484 3298 17496
rect 3786 17484 3792 17496
rect 3844 17484 3850 17536
rect 4062 17484 4068 17536
rect 4120 17524 4126 17536
rect 4157 17527 4215 17533
rect 4157 17524 4169 17527
rect 4120 17496 4169 17524
rect 4120 17484 4126 17496
rect 4157 17493 4169 17496
rect 4203 17493 4215 17527
rect 4157 17487 4215 17493
rect 4249 17527 4307 17533
rect 4249 17493 4261 17527
rect 4295 17524 4307 17527
rect 4430 17524 4436 17536
rect 4295 17496 4436 17524
rect 4295 17493 4307 17496
rect 4249 17487 4307 17493
rect 4430 17484 4436 17496
rect 4488 17484 4494 17536
rect 4525 17527 4583 17533
rect 4525 17493 4537 17527
rect 4571 17524 4583 17527
rect 4706 17524 4712 17536
rect 4571 17496 4712 17524
rect 4571 17493 4583 17496
rect 4525 17487 4583 17493
rect 4706 17484 4712 17496
rect 4764 17524 4770 17536
rect 5442 17524 5448 17536
rect 4764 17496 5448 17524
rect 4764 17484 4770 17496
rect 5442 17484 5448 17496
rect 5500 17484 5506 17536
rect 6178 17484 6184 17536
rect 6236 17524 6242 17536
rect 7009 17527 7067 17533
rect 7009 17524 7021 17527
rect 6236 17496 7021 17524
rect 6236 17484 6242 17496
rect 7009 17493 7021 17496
rect 7055 17524 7067 17527
rect 7190 17524 7196 17536
rect 7055 17496 7196 17524
rect 7055 17493 7067 17496
rect 7009 17487 7067 17493
rect 7190 17484 7196 17496
rect 7248 17484 7254 17536
rect 7558 17524 7564 17536
rect 7519 17496 7564 17524
rect 7558 17484 7564 17496
rect 7616 17524 7622 17536
rect 8202 17524 8208 17536
rect 7616 17496 8208 17524
rect 7616 17484 7622 17496
rect 8202 17484 8208 17496
rect 8260 17484 8266 17536
rect 8478 17524 8484 17536
rect 8439 17496 8484 17524
rect 8478 17484 8484 17496
rect 8536 17484 8542 17536
rect 8846 17484 8852 17536
rect 8904 17524 8910 17536
rect 9309 17527 9367 17533
rect 9309 17524 9321 17527
rect 8904 17496 9321 17524
rect 8904 17484 8910 17496
rect 9309 17493 9321 17496
rect 9355 17493 9367 17527
rect 9968 17524 9996 17632
rect 10045 17629 10057 17663
rect 10091 17660 10103 17663
rect 11072 17660 11100 17768
rect 11517 17765 11529 17768
rect 11563 17765 11575 17799
rect 12406 17796 12434 17836
rect 12989 17833 13001 17867
rect 13035 17864 13047 17867
rect 13170 17864 13176 17876
rect 13035 17836 13176 17864
rect 13035 17833 13047 17836
rect 12989 17827 13047 17833
rect 13170 17824 13176 17836
rect 13228 17824 13234 17876
rect 14921 17867 14979 17873
rect 14921 17833 14933 17867
rect 14967 17864 14979 17867
rect 15010 17864 15016 17876
rect 14967 17836 15016 17864
rect 14967 17833 14979 17836
rect 14921 17827 14979 17833
rect 15010 17824 15016 17836
rect 15068 17824 15074 17876
rect 15746 17824 15752 17876
rect 15804 17864 15810 17876
rect 16945 17867 17003 17873
rect 15804 17836 16528 17864
rect 15804 17824 15810 17836
rect 13446 17796 13452 17808
rect 12406 17768 13452 17796
rect 11517 17759 11575 17765
rect 13446 17756 13452 17768
rect 13504 17756 13510 17808
rect 11974 17728 11980 17740
rect 10091 17632 11100 17660
rect 11440 17700 11980 17728
rect 10091 17629 10103 17632
rect 10045 17623 10103 17629
rect 10428 17604 10456 17632
rect 10318 17601 10324 17604
rect 10312 17592 10324 17601
rect 10279 17564 10324 17592
rect 10312 17555 10324 17564
rect 10318 17552 10324 17555
rect 10376 17552 10382 17604
rect 10410 17552 10416 17604
rect 10468 17552 10474 17604
rect 11440 17533 11468 17700
rect 11974 17688 11980 17700
rect 12032 17728 12038 17740
rect 12345 17731 12403 17737
rect 12345 17728 12357 17731
rect 12032 17700 12357 17728
rect 12032 17688 12038 17700
rect 12345 17697 12357 17700
rect 12391 17697 12403 17731
rect 12345 17691 12403 17697
rect 12802 17688 12808 17740
rect 12860 17728 12866 17740
rect 13265 17731 13323 17737
rect 13265 17728 13277 17731
rect 12860 17700 13277 17728
rect 12860 17688 12866 17700
rect 13265 17697 13277 17700
rect 13311 17697 13323 17731
rect 14274 17728 14280 17740
rect 14235 17700 14280 17728
rect 13265 17691 13323 17697
rect 14274 17688 14280 17700
rect 14332 17688 14338 17740
rect 16500 17737 16528 17836
rect 16945 17833 16957 17867
rect 16991 17864 17003 17867
rect 17034 17864 17040 17876
rect 16991 17836 17040 17864
rect 16991 17833 17003 17836
rect 16945 17827 17003 17833
rect 17034 17824 17040 17836
rect 17092 17864 17098 17876
rect 17770 17864 17776 17876
rect 17092 17836 17776 17864
rect 17092 17824 17098 17836
rect 17770 17824 17776 17836
rect 17828 17864 17834 17876
rect 18782 17864 18788 17876
rect 17828 17836 18788 17864
rect 17828 17824 17834 17836
rect 18782 17824 18788 17836
rect 18840 17824 18846 17876
rect 19429 17867 19487 17873
rect 19429 17833 19441 17867
rect 19475 17864 19487 17867
rect 19610 17864 19616 17876
rect 19475 17836 19616 17864
rect 19475 17833 19487 17836
rect 19429 17827 19487 17833
rect 19610 17824 19616 17836
rect 19668 17864 19674 17876
rect 20438 17864 20444 17876
rect 19668 17836 20444 17864
rect 19668 17824 19674 17836
rect 20438 17824 20444 17836
rect 20496 17824 20502 17876
rect 20990 17864 20996 17876
rect 20951 17836 20996 17864
rect 20990 17824 20996 17836
rect 21048 17824 21054 17876
rect 19702 17756 19708 17808
rect 19760 17796 19766 17808
rect 19889 17799 19947 17805
rect 19889 17796 19901 17799
rect 19760 17768 19901 17796
rect 19760 17756 19766 17768
rect 19889 17765 19901 17768
rect 19935 17765 19947 17799
rect 19889 17759 19947 17765
rect 20349 17799 20407 17805
rect 20349 17765 20361 17799
rect 20395 17765 20407 17799
rect 20349 17759 20407 17765
rect 20625 17799 20683 17805
rect 20625 17765 20637 17799
rect 20671 17796 20683 17799
rect 21358 17796 21364 17808
rect 20671 17768 21364 17796
rect 20671 17765 20683 17768
rect 20625 17759 20683 17765
rect 16485 17731 16543 17737
rect 16485 17697 16497 17731
rect 16531 17697 16543 17731
rect 16485 17691 16543 17697
rect 19613 17731 19671 17737
rect 19613 17697 19625 17731
rect 19659 17728 19671 17731
rect 19978 17728 19984 17740
rect 19659 17700 19984 17728
rect 19659 17697 19671 17700
rect 19613 17691 19671 17697
rect 19978 17688 19984 17700
rect 20036 17688 20042 17740
rect 20364 17728 20392 17759
rect 21358 17756 21364 17768
rect 21416 17756 21422 17808
rect 21453 17799 21511 17805
rect 21453 17765 21465 17799
rect 21499 17796 21511 17799
rect 21542 17796 21548 17808
rect 21499 17768 21548 17796
rect 21499 17765 21511 17768
rect 21453 17759 21511 17765
rect 21542 17756 21548 17768
rect 21600 17756 21606 17808
rect 22278 17728 22284 17740
rect 20364 17700 22284 17728
rect 22278 17688 22284 17700
rect 22336 17688 22342 17740
rect 11701 17663 11759 17669
rect 11701 17629 11713 17663
rect 11747 17660 11759 17663
rect 11882 17660 11888 17672
rect 11747 17632 11888 17660
rect 11747 17629 11759 17632
rect 11701 17623 11759 17629
rect 11882 17620 11888 17632
rect 11940 17660 11946 17672
rect 12529 17663 12587 17669
rect 11940 17632 12480 17660
rect 11940 17620 11946 17632
rect 11514 17552 11520 17604
rect 11572 17592 11578 17604
rect 11793 17595 11851 17601
rect 11793 17592 11805 17595
rect 11572 17564 11805 17592
rect 11572 17552 11578 17564
rect 11793 17561 11805 17564
rect 11839 17561 11851 17595
rect 12452 17592 12480 17632
rect 12529 17629 12541 17663
rect 12575 17660 12587 17663
rect 12618 17660 12624 17672
rect 12575 17632 12624 17660
rect 12575 17629 12587 17632
rect 12529 17623 12587 17629
rect 12618 17620 12624 17632
rect 12676 17660 12682 17672
rect 13081 17663 13139 17669
rect 13081 17660 13093 17663
rect 12676 17632 13093 17660
rect 12676 17620 12682 17632
rect 13081 17629 13093 17632
rect 13127 17629 13139 17663
rect 13081 17623 13139 17629
rect 13446 17620 13452 17672
rect 13504 17660 13510 17672
rect 13541 17663 13599 17669
rect 13541 17660 13553 17663
rect 13504 17632 13553 17660
rect 13504 17620 13510 17632
rect 13541 17629 13553 17632
rect 13587 17660 13599 17663
rect 15194 17660 15200 17672
rect 13587 17632 15200 17660
rect 13587 17629 13599 17632
rect 13541 17623 13599 17629
rect 15194 17620 15200 17632
rect 15252 17620 15258 17672
rect 15654 17620 15660 17672
rect 15712 17660 15718 17672
rect 16218 17663 16276 17669
rect 16218 17660 16230 17663
rect 15712 17632 16230 17660
rect 15712 17620 15718 17632
rect 16218 17629 16230 17632
rect 16264 17629 16276 17663
rect 20070 17660 20076 17672
rect 20031 17632 20076 17660
rect 16218 17623 16276 17629
rect 20070 17620 20076 17632
rect 20128 17660 20134 17672
rect 20165 17663 20223 17669
rect 20165 17660 20177 17663
rect 20128 17632 20177 17660
rect 20128 17620 20134 17632
rect 20165 17629 20177 17632
rect 20211 17629 20223 17663
rect 20165 17623 20223 17629
rect 20254 17620 20260 17672
rect 20312 17660 20318 17672
rect 20441 17663 20499 17669
rect 20441 17660 20453 17663
rect 20312 17632 20453 17660
rect 20312 17620 20318 17632
rect 20441 17629 20453 17632
rect 20487 17629 20499 17663
rect 20714 17660 20720 17672
rect 20675 17632 20720 17660
rect 20441 17623 20499 17629
rect 20714 17620 20720 17632
rect 20772 17620 20778 17672
rect 21174 17660 21180 17672
rect 21135 17632 21180 17660
rect 21174 17620 21180 17632
rect 21232 17620 21238 17672
rect 21269 17663 21327 17669
rect 21269 17629 21281 17663
rect 21315 17629 21327 17663
rect 21269 17623 21327 17629
rect 13464 17592 13492 17620
rect 13814 17592 13820 17604
rect 12452 17564 13492 17592
rect 13775 17564 13820 17592
rect 11793 17555 11851 17561
rect 13814 17552 13820 17564
rect 13872 17552 13878 17604
rect 14461 17595 14519 17601
rect 14461 17561 14473 17595
rect 14507 17592 14519 17595
rect 15746 17592 15752 17604
rect 14507 17564 15752 17592
rect 14507 17561 14519 17564
rect 14461 17555 14519 17561
rect 15746 17552 15752 17564
rect 15804 17552 15810 17604
rect 16761 17595 16819 17601
rect 16761 17561 16773 17595
rect 16807 17592 16819 17595
rect 16942 17592 16948 17604
rect 16807 17564 16948 17592
rect 16807 17561 16819 17564
rect 16761 17555 16819 17561
rect 16942 17552 16948 17564
rect 17000 17552 17006 17604
rect 19702 17592 19708 17604
rect 19663 17564 19708 17592
rect 19702 17552 19708 17564
rect 19760 17552 19766 17604
rect 20530 17552 20536 17604
rect 20588 17592 20594 17604
rect 21284 17592 21312 17623
rect 22370 17592 22376 17604
rect 20588 17564 21312 17592
rect 21376 17564 22376 17592
rect 20588 17552 20594 17564
rect 11425 17527 11483 17533
rect 11425 17524 11437 17527
rect 9968 17496 11437 17524
rect 9309 17487 9367 17493
rect 11425 17493 11437 17496
rect 11471 17493 11483 17527
rect 11425 17487 11483 17493
rect 12161 17527 12219 17533
rect 12161 17493 12173 17527
rect 12207 17524 12219 17527
rect 12434 17524 12440 17536
rect 12207 17496 12440 17524
rect 12207 17493 12219 17496
rect 12161 17487 12219 17493
rect 12434 17484 12440 17496
rect 12492 17524 12498 17536
rect 12621 17527 12679 17533
rect 12621 17524 12633 17527
rect 12492 17496 12633 17524
rect 12492 17484 12498 17496
rect 12621 17493 12633 17496
rect 12667 17493 12679 17527
rect 12621 17487 12679 17493
rect 13354 17484 13360 17536
rect 13412 17524 13418 17536
rect 13725 17527 13783 17533
rect 13725 17524 13737 17527
rect 13412 17496 13737 17524
rect 13412 17484 13418 17496
rect 13725 17493 13737 17496
rect 13771 17493 13783 17527
rect 13725 17487 13783 17493
rect 14553 17527 14611 17533
rect 14553 17493 14565 17527
rect 14599 17524 14611 17527
rect 14918 17524 14924 17536
rect 14599 17496 14924 17524
rect 14599 17493 14611 17496
rect 14553 17487 14611 17493
rect 14918 17484 14924 17496
rect 14976 17484 14982 17536
rect 15102 17524 15108 17536
rect 15063 17496 15108 17524
rect 15102 17484 15108 17496
rect 15160 17484 15166 17536
rect 20162 17484 20168 17536
rect 20220 17524 20226 17536
rect 20714 17524 20720 17536
rect 20220 17496 20720 17524
rect 20220 17484 20226 17496
rect 20714 17484 20720 17496
rect 20772 17484 20778 17536
rect 20901 17527 20959 17533
rect 20901 17493 20913 17527
rect 20947 17524 20959 17527
rect 21376 17524 21404 17564
rect 22370 17552 22376 17564
rect 22428 17552 22434 17604
rect 20947 17496 21404 17524
rect 20947 17493 20959 17496
rect 20901 17487 20959 17493
rect 1104 17434 22056 17456
rect 1104 17382 6148 17434
rect 6200 17382 6212 17434
rect 6264 17382 6276 17434
rect 6328 17382 6340 17434
rect 6392 17382 6404 17434
rect 6456 17382 11346 17434
rect 11398 17382 11410 17434
rect 11462 17382 11474 17434
rect 11526 17382 11538 17434
rect 11590 17382 11602 17434
rect 11654 17382 16544 17434
rect 16596 17382 16608 17434
rect 16660 17382 16672 17434
rect 16724 17382 16736 17434
rect 16788 17382 16800 17434
rect 16852 17382 21742 17434
rect 21794 17382 21806 17434
rect 21858 17382 21870 17434
rect 21922 17382 21934 17434
rect 21986 17382 21998 17434
rect 22050 17382 22056 17434
rect 1104 17360 22056 17382
rect 1394 17280 1400 17332
rect 1452 17320 1458 17332
rect 4617 17323 4675 17329
rect 1452 17292 4568 17320
rect 1452 17280 1458 17292
rect 3418 17261 3424 17264
rect 3390 17255 3424 17261
rect 3390 17252 3402 17255
rect 1596 17224 3280 17252
rect 3331 17224 3402 17252
rect 1596 17193 1624 17224
rect 1581 17187 1639 17193
rect 1581 17153 1593 17187
rect 1627 17153 1639 17187
rect 1581 17147 1639 17153
rect 2797 17187 2855 17193
rect 2797 17153 2809 17187
rect 2843 17184 2855 17187
rect 2958 17184 2964 17196
rect 2843 17156 2964 17184
rect 2843 17153 2855 17156
rect 2797 17147 2855 17153
rect 2958 17144 2964 17156
rect 3016 17144 3022 17196
rect 3252 17184 3280 17224
rect 3390 17221 3402 17224
rect 3476 17252 3482 17264
rect 3602 17252 3608 17264
rect 3476 17224 3608 17252
rect 3390 17215 3424 17221
rect 3418 17212 3424 17215
rect 3476 17212 3482 17224
rect 3602 17212 3608 17224
rect 3660 17212 3666 17264
rect 4062 17212 4068 17264
rect 4120 17252 4126 17264
rect 4540 17252 4568 17292
rect 4617 17289 4629 17323
rect 4663 17320 4675 17323
rect 4982 17320 4988 17332
rect 4663 17292 4988 17320
rect 4663 17289 4675 17292
rect 4617 17283 4675 17289
rect 4982 17280 4988 17292
rect 5040 17280 5046 17332
rect 5077 17323 5135 17329
rect 5077 17289 5089 17323
rect 5123 17320 5135 17323
rect 5445 17323 5503 17329
rect 5445 17320 5457 17323
rect 5123 17292 5457 17320
rect 5123 17289 5135 17292
rect 5077 17283 5135 17289
rect 5445 17289 5457 17292
rect 5491 17289 5503 17323
rect 5445 17283 5503 17289
rect 5534 17280 5540 17332
rect 5592 17320 5598 17332
rect 5813 17323 5871 17329
rect 5813 17320 5825 17323
rect 5592 17292 5825 17320
rect 5592 17280 5598 17292
rect 5813 17289 5825 17292
rect 5859 17289 5871 17323
rect 5813 17283 5871 17289
rect 5905 17323 5963 17329
rect 5905 17289 5917 17323
rect 5951 17320 5963 17323
rect 6270 17320 6276 17332
rect 5951 17292 6276 17320
rect 5951 17289 5963 17292
rect 5905 17283 5963 17289
rect 6270 17280 6276 17292
rect 6328 17280 6334 17332
rect 6365 17323 6423 17329
rect 6365 17289 6377 17323
rect 6411 17289 6423 17323
rect 8018 17320 8024 17332
rect 6365 17283 6423 17289
rect 6472 17292 7788 17320
rect 7979 17292 8024 17320
rect 6380 17252 6408 17283
rect 4120 17224 4476 17252
rect 4540 17224 6408 17252
rect 4120 17212 4126 17224
rect 4448 17184 4476 17224
rect 4798 17184 4804 17196
rect 3252 17156 4200 17184
rect 4448 17156 4804 17184
rect 3053 17119 3111 17125
rect 3053 17085 3065 17119
rect 3099 17116 3111 17119
rect 3145 17119 3203 17125
rect 3145 17116 3157 17119
rect 3099 17088 3157 17116
rect 3099 17085 3111 17088
rect 3053 17079 3111 17085
rect 3145 17085 3157 17088
rect 3191 17085 3203 17119
rect 3145 17079 3203 17085
rect 1394 16980 1400 16992
rect 1355 16952 1400 16980
rect 1394 16940 1400 16952
rect 1452 16940 1458 16992
rect 1673 16983 1731 16989
rect 1673 16949 1685 16983
rect 1719 16980 1731 16983
rect 2130 16980 2136 16992
rect 1719 16952 2136 16980
rect 1719 16949 1731 16952
rect 1673 16943 1731 16949
rect 2130 16940 2136 16952
rect 2188 16940 2194 16992
rect 2682 16940 2688 16992
rect 2740 16980 2746 16992
rect 3068 16980 3096 17079
rect 4172 17048 4200 17156
rect 4798 17144 4804 17156
rect 4856 17144 4862 17196
rect 4982 17184 4988 17196
rect 4943 17156 4988 17184
rect 4982 17144 4988 17156
rect 5040 17144 5046 17196
rect 5083 17156 5681 17184
rect 4246 17076 4252 17128
rect 4304 17116 4310 17128
rect 5083 17116 5111 17156
rect 4304 17088 5111 17116
rect 5261 17119 5319 17125
rect 4304 17076 4310 17088
rect 5261 17085 5273 17119
rect 5307 17116 5319 17119
rect 5442 17116 5448 17128
rect 5307 17088 5448 17116
rect 5307 17085 5319 17088
rect 5261 17079 5319 17085
rect 5442 17076 5448 17088
rect 5500 17076 5506 17128
rect 5166 17048 5172 17060
rect 4172 17020 5172 17048
rect 5166 17008 5172 17020
rect 5224 17008 5230 17060
rect 5653 17048 5681 17156
rect 5902 17144 5908 17196
rect 5960 17184 5966 17196
rect 6472 17184 6500 17292
rect 6638 17212 6644 17264
rect 6696 17212 6702 17264
rect 6914 17212 6920 17264
rect 6972 17252 6978 17264
rect 7760 17252 7788 17292
rect 8018 17280 8024 17292
rect 8076 17280 8082 17332
rect 8202 17280 8208 17332
rect 8260 17320 8266 17332
rect 8846 17320 8852 17332
rect 8260 17292 8616 17320
rect 8807 17292 8852 17320
rect 8260 17280 8266 17292
rect 8478 17252 8484 17264
rect 6972 17224 7696 17252
rect 6972 17212 6978 17224
rect 5960 17156 6500 17184
rect 6549 17187 6607 17193
rect 5960 17144 5966 17156
rect 6549 17153 6561 17187
rect 6595 17184 6607 17187
rect 6656 17184 6684 17212
rect 6822 17184 6828 17196
rect 6595 17156 6828 17184
rect 6595 17153 6607 17156
rect 6549 17147 6607 17153
rect 6822 17144 6828 17156
rect 6880 17144 6886 17196
rect 7009 17187 7067 17193
rect 7009 17153 7021 17187
rect 7055 17153 7067 17187
rect 7009 17147 7067 17153
rect 7101 17187 7159 17193
rect 7101 17153 7113 17187
rect 7147 17184 7159 17187
rect 7466 17184 7472 17196
rect 7147 17156 7472 17184
rect 7147 17153 7159 17156
rect 7101 17147 7159 17153
rect 6089 17119 6147 17125
rect 6089 17085 6101 17119
rect 6135 17116 6147 17119
rect 6178 17116 6184 17128
rect 6135 17088 6184 17116
rect 6135 17085 6147 17088
rect 6089 17079 6147 17085
rect 6178 17076 6184 17088
rect 6236 17076 6242 17128
rect 6638 17076 6644 17128
rect 6696 17116 6702 17128
rect 7024 17116 7052 17147
rect 7466 17144 7472 17156
rect 7524 17144 7530 17196
rect 7668 17193 7696 17224
rect 7760 17224 8484 17252
rect 7760 17193 7788 17224
rect 8478 17212 8484 17224
rect 8536 17212 8542 17264
rect 7653 17187 7711 17193
rect 7653 17153 7665 17187
rect 7699 17153 7711 17187
rect 7653 17147 7711 17153
rect 7745 17187 7803 17193
rect 7745 17153 7757 17187
rect 7791 17153 7803 17187
rect 7745 17147 7803 17153
rect 7926 17144 7932 17196
rect 7984 17184 7990 17196
rect 8389 17187 8447 17193
rect 8389 17184 8401 17187
rect 7984 17156 8401 17184
rect 7984 17144 7990 17156
rect 8389 17153 8401 17156
rect 8435 17153 8447 17187
rect 8588 17184 8616 17292
rect 8846 17280 8852 17292
rect 8904 17280 8910 17332
rect 11054 17320 11060 17332
rect 8956 17292 11060 17320
rect 8662 17212 8668 17264
rect 8720 17252 8726 17264
rect 8956 17252 8984 17292
rect 11054 17280 11060 17292
rect 11112 17320 11118 17332
rect 11238 17320 11244 17332
rect 11112 17292 11244 17320
rect 11112 17280 11118 17292
rect 11238 17280 11244 17292
rect 11296 17280 11302 17332
rect 11882 17320 11888 17332
rect 11532 17292 11888 17320
rect 8720 17224 8984 17252
rect 8720 17212 8726 17224
rect 9030 17212 9036 17264
rect 9088 17252 9094 17264
rect 9950 17252 9956 17264
rect 9088 17224 9956 17252
rect 9088 17212 9094 17224
rect 9950 17212 9956 17224
rect 10008 17212 10014 17264
rect 9858 17184 9864 17196
rect 8588 17156 9864 17184
rect 8389 17147 8447 17153
rect 9858 17144 9864 17156
rect 9916 17144 9922 17196
rect 10134 17144 10140 17196
rect 10192 17193 10198 17196
rect 10192 17147 10204 17193
rect 10192 17144 10198 17147
rect 10594 17144 10600 17196
rect 10652 17184 10658 17196
rect 11532 17193 11560 17292
rect 11882 17280 11888 17292
rect 11940 17280 11946 17332
rect 12434 17280 12440 17332
rect 12492 17320 12498 17332
rect 13630 17320 13636 17332
rect 12492 17292 13636 17320
rect 12492 17280 12498 17292
rect 13630 17280 13636 17292
rect 13688 17280 13694 17332
rect 14918 17320 14924 17332
rect 14879 17292 14924 17320
rect 14918 17280 14924 17292
rect 14976 17280 14982 17332
rect 15010 17280 15016 17332
rect 15068 17320 15074 17332
rect 16117 17323 16175 17329
rect 15068 17292 15700 17320
rect 15068 17280 15074 17292
rect 11784 17255 11842 17261
rect 11784 17221 11796 17255
rect 11830 17252 11842 17255
rect 11974 17252 11980 17264
rect 11830 17224 11980 17252
rect 11830 17221 11842 17224
rect 11784 17215 11842 17221
rect 11974 17212 11980 17224
rect 12032 17252 12038 17264
rect 12894 17252 12900 17264
rect 12032 17224 12900 17252
rect 12032 17212 12038 17224
rect 12894 17212 12900 17224
rect 12952 17212 12958 17264
rect 15672 17252 15700 17292
rect 16117 17289 16129 17323
rect 16163 17320 16175 17323
rect 16669 17323 16727 17329
rect 16669 17320 16681 17323
rect 16163 17292 16681 17320
rect 16163 17289 16175 17292
rect 16117 17283 16175 17289
rect 16669 17289 16681 17292
rect 16715 17289 16727 17323
rect 17034 17320 17040 17332
rect 16995 17292 17040 17320
rect 16669 17283 16727 17289
rect 17034 17280 17040 17292
rect 17092 17280 17098 17332
rect 19610 17280 19616 17332
rect 19668 17320 19674 17332
rect 19797 17323 19855 17329
rect 19797 17320 19809 17323
rect 19668 17292 19809 17320
rect 19668 17280 19674 17292
rect 19797 17289 19809 17292
rect 19843 17320 19855 17323
rect 20257 17323 20315 17329
rect 20257 17320 20269 17323
rect 19843 17292 20269 17320
rect 19843 17289 19855 17292
rect 19797 17283 19855 17289
rect 20257 17289 20269 17292
rect 20303 17289 20315 17323
rect 20257 17283 20315 17289
rect 20993 17323 21051 17329
rect 20993 17289 21005 17323
rect 21039 17320 21051 17323
rect 21266 17320 21272 17332
rect 21039 17292 21272 17320
rect 21039 17289 21051 17292
rect 20993 17283 21051 17289
rect 21266 17280 21272 17292
rect 21324 17280 21330 17332
rect 20717 17255 20775 17261
rect 20717 17252 20729 17255
rect 15672 17224 20729 17252
rect 20717 17221 20729 17224
rect 20763 17252 20775 17255
rect 20763 17224 20852 17252
rect 20763 17221 20775 17224
rect 20717 17215 20775 17221
rect 10965 17187 11023 17193
rect 10965 17184 10977 17187
rect 10652 17156 10977 17184
rect 10652 17144 10658 17156
rect 10965 17153 10977 17156
rect 11011 17153 11023 17187
rect 10965 17147 11023 17153
rect 11517 17187 11575 17193
rect 11517 17153 11529 17187
rect 11563 17153 11575 17187
rect 13446 17184 13452 17196
rect 13407 17156 13452 17184
rect 11517 17147 11575 17153
rect 13446 17144 13452 17156
rect 13504 17144 13510 17196
rect 13716 17187 13774 17193
rect 13716 17153 13728 17187
rect 13762 17184 13774 17187
rect 15102 17184 15108 17196
rect 13762 17156 15108 17184
rect 13762 17153 13774 17156
rect 13716 17147 13774 17153
rect 15102 17144 15108 17156
rect 15160 17144 15166 17196
rect 15286 17184 15292 17196
rect 15247 17156 15292 17184
rect 15286 17144 15292 17156
rect 15344 17144 15350 17196
rect 15580 17156 16344 17184
rect 7282 17116 7288 17128
rect 6696 17088 7052 17116
rect 7243 17088 7288 17116
rect 6696 17076 6702 17088
rect 7282 17076 7288 17088
rect 7340 17076 7346 17128
rect 8294 17076 8300 17128
rect 8352 17116 8358 17128
rect 8481 17119 8539 17125
rect 8481 17116 8493 17119
rect 8352 17088 8493 17116
rect 8352 17076 8358 17088
rect 8481 17085 8493 17088
rect 8527 17085 8539 17119
rect 8481 17079 8539 17085
rect 8665 17119 8723 17125
rect 8665 17085 8677 17119
rect 8711 17116 8723 17119
rect 8938 17116 8944 17128
rect 8711 17088 8944 17116
rect 8711 17085 8723 17088
rect 8665 17079 8723 17085
rect 8938 17076 8944 17088
rect 8996 17076 9002 17128
rect 10410 17116 10416 17128
rect 10371 17088 10416 17116
rect 10410 17076 10416 17088
rect 10468 17076 10474 17128
rect 15010 17116 15016 17128
rect 14752 17088 15016 17116
rect 5653 17020 6776 17048
rect 2740 16952 3096 16980
rect 4525 16983 4583 16989
rect 2740 16940 2746 16952
rect 4525 16949 4537 16983
rect 4571 16980 4583 16983
rect 4614 16980 4620 16992
rect 4571 16952 4620 16980
rect 4571 16949 4583 16952
rect 4525 16943 4583 16949
rect 4614 16940 4620 16952
rect 4672 16980 4678 16992
rect 5994 16980 6000 16992
rect 4672 16952 6000 16980
rect 4672 16940 4678 16952
rect 5994 16940 6000 16952
rect 6052 16940 6058 16992
rect 6638 16980 6644 16992
rect 6599 16952 6644 16980
rect 6638 16940 6644 16952
rect 6696 16940 6702 16992
rect 6748 16980 6776 17020
rect 7006 17008 7012 17060
rect 7064 17048 7070 17060
rect 7469 17051 7527 17057
rect 7469 17048 7481 17051
rect 7064 17020 7481 17048
rect 7064 17008 7070 17020
rect 7469 17017 7481 17020
rect 7515 17017 7527 17051
rect 7469 17011 7527 17017
rect 8386 17008 8392 17060
rect 8444 17048 8450 17060
rect 9030 17048 9036 17060
rect 8444 17020 9036 17048
rect 8444 17008 8450 17020
rect 9030 17008 9036 17020
rect 9088 17008 9094 17060
rect 12526 17008 12532 17060
rect 12584 17048 12590 17060
rect 12989 17051 13047 17057
rect 12989 17048 13001 17051
rect 12584 17020 13001 17048
rect 12584 17008 12590 17020
rect 12989 17017 13001 17020
rect 13035 17017 13047 17051
rect 12989 17011 13047 17017
rect 7929 16983 7987 16989
rect 7929 16980 7941 16983
rect 6748 16952 7941 16980
rect 7929 16949 7941 16952
rect 7975 16980 7987 16983
rect 10686 16980 10692 16992
rect 7975 16952 10692 16980
rect 7975 16949 7987 16952
rect 7929 16943 7987 16949
rect 10686 16940 10692 16952
rect 10744 16940 10750 16992
rect 11698 16940 11704 16992
rect 11756 16980 11762 16992
rect 12897 16983 12955 16989
rect 12897 16980 12909 16983
rect 11756 16952 12909 16980
rect 11756 16940 11762 16952
rect 12897 16949 12909 16952
rect 12943 16949 12955 16983
rect 13170 16980 13176 16992
rect 13131 16952 13176 16980
rect 12897 16943 12955 16949
rect 13170 16940 13176 16952
rect 13228 16940 13234 16992
rect 13722 16940 13728 16992
rect 13780 16980 13786 16992
rect 14752 16980 14780 17088
rect 15010 17076 15016 17088
rect 15068 17076 15074 17128
rect 15378 17116 15384 17128
rect 15339 17088 15384 17116
rect 15378 17076 15384 17088
rect 15436 17076 15442 17128
rect 15580 17125 15608 17156
rect 15565 17119 15623 17125
rect 15565 17085 15577 17119
rect 15611 17085 15623 17119
rect 16206 17116 16212 17128
rect 16167 17088 16212 17116
rect 15565 17079 15623 17085
rect 14829 17051 14887 17057
rect 14829 17017 14841 17051
rect 14875 17048 14887 17051
rect 15194 17048 15200 17060
rect 14875 17020 15200 17048
rect 14875 17017 14887 17020
rect 14829 17011 14887 17017
rect 15194 17008 15200 17020
rect 15252 17048 15258 17060
rect 15580 17048 15608 17079
rect 16206 17076 16212 17088
rect 16264 17076 16270 17128
rect 16316 17125 16344 17156
rect 18966 17144 18972 17196
rect 19024 17184 19030 17196
rect 20824 17193 20852 17224
rect 19981 17187 20039 17193
rect 19981 17184 19993 17187
rect 19024 17156 19993 17184
rect 19024 17144 19030 17156
rect 19981 17153 19993 17156
rect 20027 17153 20039 17187
rect 19981 17147 20039 17153
rect 20809 17187 20867 17193
rect 20809 17153 20821 17187
rect 20855 17153 20867 17187
rect 21266 17184 21272 17196
rect 21227 17156 21272 17184
rect 20809 17147 20867 17153
rect 21266 17144 21272 17156
rect 21324 17144 21330 17196
rect 16301 17119 16359 17125
rect 16301 17085 16313 17119
rect 16347 17085 16359 17119
rect 17126 17116 17132 17128
rect 17087 17088 17132 17116
rect 16301 17079 16359 17085
rect 17126 17076 17132 17088
rect 17184 17076 17190 17128
rect 17218 17076 17224 17128
rect 17276 17116 17282 17128
rect 20622 17116 20628 17128
rect 17276 17088 17321 17116
rect 20180 17088 20628 17116
rect 17276 17076 17282 17088
rect 15746 17048 15752 17060
rect 15252 17020 15608 17048
rect 15707 17020 15752 17048
rect 15252 17008 15258 17020
rect 15746 17008 15752 17020
rect 15804 17008 15810 17060
rect 16390 17008 16396 17060
rect 16448 17048 16454 17060
rect 20180 17057 20208 17088
rect 20622 17076 20628 17088
rect 20680 17076 20686 17128
rect 20165 17051 20223 17057
rect 16448 17020 17540 17048
rect 16448 17008 16454 17020
rect 17512 16992 17540 17020
rect 20165 17017 20177 17051
rect 20211 17017 20223 17051
rect 21174 17048 21180 17060
rect 21087 17020 21180 17048
rect 20165 17011 20223 17017
rect 21174 17008 21180 17020
rect 21232 17048 21238 17060
rect 22922 17048 22928 17060
rect 21232 17020 22928 17048
rect 21232 17008 21238 17020
rect 22922 17008 22928 17020
rect 22980 17008 22986 17060
rect 13780 16952 14780 16980
rect 13780 16940 13786 16952
rect 15102 16940 15108 16992
rect 15160 16980 15166 16992
rect 17218 16980 17224 16992
rect 15160 16952 17224 16980
rect 15160 16940 15166 16952
rect 17218 16940 17224 16952
rect 17276 16940 17282 16992
rect 17494 16980 17500 16992
rect 17455 16952 17500 16980
rect 17494 16940 17500 16952
rect 17552 16940 17558 16992
rect 19610 16940 19616 16992
rect 19668 16980 19674 16992
rect 20441 16983 20499 16989
rect 20441 16980 20453 16983
rect 19668 16952 20453 16980
rect 19668 16940 19674 16952
rect 20441 16949 20453 16952
rect 20487 16980 20499 16983
rect 20806 16980 20812 16992
rect 20487 16952 20812 16980
rect 20487 16949 20499 16952
rect 20441 16943 20499 16949
rect 20806 16940 20812 16952
rect 20864 16940 20870 16992
rect 21450 16980 21456 16992
rect 21411 16952 21456 16980
rect 21450 16940 21456 16952
rect 21508 16940 21514 16992
rect 1104 16890 21896 16912
rect 1104 16838 3549 16890
rect 3601 16838 3613 16890
rect 3665 16838 3677 16890
rect 3729 16838 3741 16890
rect 3793 16838 3805 16890
rect 3857 16838 8747 16890
rect 8799 16838 8811 16890
rect 8863 16838 8875 16890
rect 8927 16838 8939 16890
rect 8991 16838 9003 16890
rect 9055 16838 13945 16890
rect 13997 16838 14009 16890
rect 14061 16838 14073 16890
rect 14125 16838 14137 16890
rect 14189 16838 14201 16890
rect 14253 16838 19143 16890
rect 19195 16838 19207 16890
rect 19259 16838 19271 16890
rect 19323 16838 19335 16890
rect 19387 16838 19399 16890
rect 19451 16838 21896 16890
rect 1104 16816 21896 16838
rect 2590 16776 2596 16788
rect 2240 16748 2596 16776
rect 1118 16668 1124 16720
rect 1176 16708 1182 16720
rect 1176 16680 1348 16708
rect 1176 16668 1182 16680
rect 1320 16652 1348 16680
rect 1302 16600 1308 16652
rect 1360 16600 1366 16652
rect 2240 16649 2268 16748
rect 2590 16736 2596 16748
rect 2648 16736 2654 16788
rect 3142 16736 3148 16788
rect 3200 16776 3206 16788
rect 3789 16779 3847 16785
rect 3789 16776 3801 16779
rect 3200 16748 3801 16776
rect 3200 16736 3206 16748
rect 3789 16745 3801 16748
rect 3835 16745 3847 16779
rect 3789 16739 3847 16745
rect 4801 16779 4859 16785
rect 4801 16745 4813 16779
rect 4847 16776 4859 16779
rect 5810 16776 5816 16788
rect 4847 16748 5816 16776
rect 4847 16745 4859 16748
rect 4801 16739 4859 16745
rect 5810 16736 5816 16748
rect 5868 16736 5874 16788
rect 6270 16736 6276 16788
rect 6328 16776 6334 16788
rect 6549 16779 6607 16785
rect 6549 16776 6561 16779
rect 6328 16748 6561 16776
rect 6328 16736 6334 16748
rect 6549 16745 6561 16748
rect 6595 16745 6607 16779
rect 7742 16776 7748 16788
rect 6549 16739 6607 16745
rect 7024 16748 7748 16776
rect 3418 16668 3424 16720
rect 3476 16708 3482 16720
rect 3605 16711 3663 16717
rect 3605 16708 3617 16711
rect 3476 16680 3617 16708
rect 3476 16668 3482 16680
rect 3605 16677 3617 16680
rect 3651 16677 3663 16711
rect 3605 16671 3663 16677
rect 3878 16668 3884 16720
rect 3936 16708 3942 16720
rect 5994 16708 6000 16720
rect 3936 16680 6000 16708
rect 3936 16668 3942 16680
rect 5994 16668 6000 16680
rect 6052 16708 6058 16720
rect 6914 16708 6920 16720
rect 6052 16680 6920 16708
rect 6052 16668 6058 16680
rect 6914 16668 6920 16680
rect 6972 16668 6978 16720
rect 2225 16643 2283 16649
rect 2225 16609 2237 16643
rect 2271 16609 2283 16643
rect 4341 16643 4399 16649
rect 4341 16640 4353 16643
rect 2225 16603 2283 16609
rect 3252 16612 4353 16640
rect 1394 16572 1400 16584
rect 1355 16544 1400 16572
rect 1394 16532 1400 16544
rect 1452 16532 1458 16584
rect 2038 16572 2044 16584
rect 1999 16544 2044 16572
rect 2038 16532 2044 16544
rect 2096 16532 2102 16584
rect 2492 16575 2550 16581
rect 2492 16572 2504 16575
rect 2240 16544 2504 16572
rect 2240 16516 2268 16544
rect 2492 16541 2504 16544
rect 2538 16572 2550 16575
rect 3252 16572 3280 16612
rect 4341 16609 4353 16612
rect 4387 16609 4399 16643
rect 5350 16640 5356 16652
rect 5311 16612 5356 16640
rect 4341 16603 4399 16609
rect 5350 16600 5356 16612
rect 5408 16600 5414 16652
rect 5442 16600 5448 16652
rect 5500 16640 5506 16652
rect 5500 16612 5545 16640
rect 5500 16600 5506 16612
rect 5626 16600 5632 16652
rect 5684 16640 5690 16652
rect 6178 16640 6184 16652
rect 5684 16612 6184 16640
rect 5684 16600 5690 16612
rect 6178 16600 6184 16612
rect 6236 16640 6242 16652
rect 7024 16649 7052 16748
rect 7742 16736 7748 16748
rect 7800 16736 7806 16788
rect 9401 16779 9459 16785
rect 9401 16745 9413 16779
rect 9447 16776 9459 16779
rect 9490 16776 9496 16788
rect 9447 16748 9496 16776
rect 9447 16745 9459 16748
rect 9401 16739 9459 16745
rect 9490 16736 9496 16748
rect 9548 16736 9554 16788
rect 9858 16736 9864 16788
rect 9916 16776 9922 16788
rect 10594 16776 10600 16788
rect 9916 16748 10600 16776
rect 9916 16736 9922 16748
rect 10594 16736 10600 16748
rect 10652 16736 10658 16788
rect 11146 16736 11152 16788
rect 11204 16776 11210 16788
rect 11790 16776 11796 16788
rect 11204 16748 11796 16776
rect 11204 16736 11210 16748
rect 11790 16736 11796 16748
rect 11848 16736 11854 16788
rect 12342 16776 12348 16788
rect 12303 16748 12348 16776
rect 12342 16736 12348 16748
rect 12400 16736 12406 16788
rect 12986 16736 12992 16788
rect 13044 16776 13050 16788
rect 13449 16779 13507 16785
rect 13449 16776 13461 16779
rect 13044 16748 13461 16776
rect 13044 16736 13050 16748
rect 13449 16745 13461 16748
rect 13495 16745 13507 16779
rect 13449 16739 13507 16745
rect 14093 16779 14151 16785
rect 14093 16745 14105 16779
rect 14139 16776 14151 16779
rect 14274 16776 14280 16788
rect 14139 16748 14280 16776
rect 14139 16745 14151 16748
rect 14093 16739 14151 16745
rect 14274 16736 14280 16748
rect 14332 16736 14338 16788
rect 15286 16736 15292 16788
rect 15344 16776 15350 16788
rect 16393 16779 16451 16785
rect 16393 16776 16405 16779
rect 15344 16748 16405 16776
rect 15344 16736 15350 16748
rect 16393 16745 16405 16748
rect 16439 16745 16451 16779
rect 16393 16739 16451 16745
rect 17126 16736 17132 16788
rect 17184 16776 17190 16788
rect 17221 16779 17279 16785
rect 17221 16776 17233 16779
rect 17184 16748 17233 16776
rect 17184 16736 17190 16748
rect 17221 16745 17233 16748
rect 17267 16745 17279 16779
rect 19518 16776 19524 16788
rect 17221 16739 17279 16745
rect 17604 16748 19524 16776
rect 8386 16708 8392 16720
rect 8220 16680 8392 16708
rect 6273 16643 6331 16649
rect 6273 16640 6285 16643
rect 6236 16612 6285 16640
rect 6236 16600 6242 16612
rect 6273 16609 6285 16612
rect 6319 16609 6331 16643
rect 6273 16603 6331 16609
rect 7009 16643 7067 16649
rect 7009 16609 7021 16643
rect 7055 16609 7067 16643
rect 7009 16603 7067 16609
rect 7193 16643 7251 16649
rect 7193 16609 7205 16643
rect 7239 16640 7251 16643
rect 7282 16640 7288 16652
rect 7239 16612 7288 16640
rect 7239 16609 7251 16612
rect 7193 16603 7251 16609
rect 7282 16600 7288 16612
rect 7340 16600 7346 16652
rect 7926 16640 7932 16652
rect 7887 16612 7932 16640
rect 7926 16600 7932 16612
rect 7984 16600 7990 16652
rect 8220 16649 8248 16680
rect 8386 16668 8392 16680
rect 8444 16668 8450 16720
rect 8662 16668 8668 16720
rect 8720 16708 8726 16720
rect 11054 16708 11060 16720
rect 8720 16680 11060 16708
rect 8720 16668 8726 16680
rect 11054 16668 11060 16680
rect 11112 16668 11118 16720
rect 11348 16680 11836 16708
rect 8205 16643 8263 16649
rect 8205 16609 8217 16643
rect 8251 16609 8263 16643
rect 8205 16603 8263 16609
rect 8297 16643 8355 16649
rect 8297 16609 8309 16643
rect 8343 16640 8355 16643
rect 9766 16640 9772 16652
rect 8343 16612 9772 16640
rect 8343 16609 8355 16612
rect 8297 16603 8355 16609
rect 9766 16600 9772 16612
rect 9824 16600 9830 16652
rect 9950 16640 9956 16652
rect 9911 16612 9956 16640
rect 9950 16600 9956 16612
rect 10008 16600 10014 16652
rect 10134 16640 10140 16652
rect 10095 16612 10140 16640
rect 10134 16600 10140 16612
rect 10192 16600 10198 16652
rect 10689 16643 10747 16649
rect 10689 16609 10701 16643
rect 10735 16640 10747 16643
rect 10735 16612 11008 16640
rect 10735 16609 10747 16612
rect 10689 16603 10747 16609
rect 2538 16544 3280 16572
rect 2538 16541 2550 16544
rect 2492 16535 2550 16541
rect 3970 16532 3976 16584
rect 4028 16572 4034 16584
rect 4249 16575 4307 16581
rect 4249 16572 4261 16575
rect 4028 16544 4261 16572
rect 4028 16532 4034 16544
rect 4249 16541 4261 16544
rect 4295 16541 4307 16575
rect 4617 16575 4675 16581
rect 4617 16572 4629 16575
rect 4249 16535 4307 16541
rect 4356 16544 4629 16572
rect 4356 16516 4384 16544
rect 4617 16541 4629 16544
rect 4663 16572 4675 16575
rect 4706 16572 4712 16584
rect 4663 16544 4712 16572
rect 4663 16541 4675 16544
rect 4617 16535 4675 16541
rect 4706 16532 4712 16544
rect 4764 16532 4770 16584
rect 6089 16575 6147 16581
rect 6089 16541 6101 16575
rect 6135 16572 6147 16575
rect 6638 16572 6644 16584
rect 6135 16544 6644 16572
rect 6135 16541 6147 16544
rect 6089 16535 6147 16541
rect 6638 16532 6644 16544
rect 6696 16532 6702 16584
rect 7561 16575 7619 16581
rect 7561 16541 7573 16575
rect 7607 16572 7619 16575
rect 7742 16572 7748 16584
rect 7607 16544 7748 16572
rect 7607 16541 7619 16544
rect 7561 16535 7619 16541
rect 7742 16532 7748 16544
rect 7800 16532 7806 16584
rect 8110 16532 8116 16584
rect 8168 16572 8174 16584
rect 9125 16575 9183 16581
rect 9125 16572 9137 16575
rect 8168 16544 9137 16572
rect 8168 16532 8174 16544
rect 9125 16541 9137 16544
rect 9171 16572 9183 16575
rect 10410 16572 10416 16584
rect 9171 16544 10416 16572
rect 9171 16541 9183 16544
rect 9125 16535 9183 16541
rect 10410 16532 10416 16544
rect 10468 16532 10474 16584
rect 10594 16532 10600 16584
rect 10652 16572 10658 16584
rect 10781 16575 10839 16581
rect 10781 16572 10793 16575
rect 10652 16544 10793 16572
rect 10652 16532 10658 16544
rect 10781 16541 10793 16544
rect 10827 16541 10839 16575
rect 10980 16572 11008 16612
rect 11146 16600 11152 16652
rect 11204 16640 11210 16652
rect 11348 16649 11376 16680
rect 11333 16643 11391 16649
rect 11333 16640 11345 16643
rect 11204 16612 11345 16640
rect 11204 16600 11210 16612
rect 11333 16609 11345 16612
rect 11379 16609 11391 16643
rect 11698 16640 11704 16652
rect 11659 16612 11704 16640
rect 11333 16603 11391 16609
rect 11698 16600 11704 16612
rect 11756 16600 11762 16652
rect 11808 16649 11836 16680
rect 12434 16668 12440 16720
rect 12492 16708 12498 16720
rect 12710 16708 12716 16720
rect 12492 16680 12716 16708
rect 12492 16668 12498 16680
rect 12710 16668 12716 16680
rect 12768 16668 12774 16720
rect 15654 16668 15660 16720
rect 15712 16708 15718 16720
rect 15712 16680 16252 16708
rect 15712 16668 15718 16680
rect 16224 16652 16252 16680
rect 11793 16643 11851 16649
rect 11793 16609 11805 16643
rect 11839 16609 11851 16643
rect 11793 16603 11851 16609
rect 12894 16600 12900 16652
rect 12952 16640 12958 16652
rect 13633 16643 13691 16649
rect 13633 16640 13645 16643
rect 12952 16612 12997 16640
rect 13096 16612 13645 16640
rect 12952 16600 12958 16612
rect 12710 16572 12716 16584
rect 10980 16544 12716 16572
rect 10781 16535 10839 16541
rect 12710 16532 12716 16544
rect 12768 16532 12774 16584
rect 12802 16532 12808 16584
rect 12860 16572 12866 16584
rect 13096 16572 13124 16612
rect 13633 16609 13645 16612
rect 13679 16609 13691 16643
rect 15473 16643 15531 16649
rect 15473 16640 15485 16643
rect 13633 16603 13691 16609
rect 15396 16612 15485 16640
rect 13354 16572 13360 16584
rect 12860 16544 13124 16572
rect 13315 16544 13360 16572
rect 12860 16532 12866 16544
rect 13354 16532 13360 16544
rect 13412 16532 13418 16584
rect 15194 16532 15200 16584
rect 15252 16581 15258 16584
rect 15252 16572 15264 16581
rect 15252 16544 15297 16572
rect 15252 16535 15264 16544
rect 15252 16532 15258 16535
rect 2222 16464 2228 16516
rect 2280 16464 2286 16516
rect 4338 16464 4344 16516
rect 4396 16464 4402 16516
rect 5261 16507 5319 16513
rect 5261 16473 5273 16507
rect 5307 16504 5319 16507
rect 5307 16476 5764 16504
rect 5307 16473 5319 16476
rect 5261 16467 5319 16473
rect 1578 16436 1584 16448
rect 1539 16408 1584 16436
rect 1578 16396 1584 16408
rect 1636 16396 1642 16448
rect 1854 16436 1860 16448
rect 1815 16408 1860 16436
rect 1854 16396 1860 16408
rect 1912 16396 1918 16448
rect 4154 16436 4160 16448
rect 4115 16408 4160 16436
rect 4154 16396 4160 16408
rect 4212 16396 4218 16448
rect 4890 16396 4896 16448
rect 4948 16436 4954 16448
rect 5736 16445 5764 16476
rect 5902 16464 5908 16516
rect 5960 16504 5966 16516
rect 7190 16504 7196 16516
rect 5960 16476 7196 16504
rect 5960 16464 5966 16476
rect 7190 16464 7196 16476
rect 7248 16464 7254 16516
rect 8389 16507 8447 16513
rect 8389 16473 8401 16507
rect 8435 16504 8447 16507
rect 8435 16476 9536 16504
rect 8435 16473 8447 16476
rect 8389 16467 8447 16473
rect 5721 16439 5779 16445
rect 4948 16408 4993 16436
rect 4948 16396 4954 16408
rect 5721 16405 5733 16439
rect 5767 16405 5779 16439
rect 5721 16399 5779 16405
rect 6181 16439 6239 16445
rect 6181 16405 6193 16439
rect 6227 16436 6239 16439
rect 6822 16436 6828 16448
rect 6227 16408 6828 16436
rect 6227 16405 6239 16408
rect 6181 16399 6239 16405
rect 6822 16396 6828 16408
rect 6880 16396 6886 16448
rect 6914 16396 6920 16448
rect 6972 16436 6978 16448
rect 7374 16436 7380 16448
rect 6972 16408 7017 16436
rect 7335 16408 7380 16436
rect 6972 16396 6978 16408
rect 7374 16396 7380 16408
rect 7432 16396 7438 16448
rect 8757 16439 8815 16445
rect 8757 16405 8769 16439
rect 8803 16436 8815 16439
rect 8846 16436 8852 16448
rect 8803 16408 8852 16436
rect 8803 16405 8815 16408
rect 8757 16399 8815 16405
rect 8846 16396 8852 16408
rect 8904 16396 8910 16448
rect 8938 16396 8944 16448
rect 8996 16436 9002 16448
rect 9508 16445 9536 16476
rect 9582 16464 9588 16516
rect 9640 16504 9646 16516
rect 10873 16507 10931 16513
rect 10873 16504 10885 16507
rect 9640 16476 10885 16504
rect 9640 16464 9646 16476
rect 10873 16473 10885 16476
rect 10919 16473 10931 16507
rect 10873 16467 10931 16473
rect 11054 16464 11060 16516
rect 11112 16504 11118 16516
rect 13262 16504 13268 16516
rect 11112 16476 11928 16504
rect 11112 16464 11118 16476
rect 9493 16439 9551 16445
rect 8996 16408 9041 16436
rect 8996 16396 9002 16408
rect 9493 16405 9505 16439
rect 9539 16405 9551 16439
rect 9858 16436 9864 16448
rect 9819 16408 9864 16436
rect 9493 16399 9551 16405
rect 9858 16396 9864 16408
rect 9916 16396 9922 16448
rect 10413 16439 10471 16445
rect 10413 16405 10425 16439
rect 10459 16436 10471 16439
rect 11072 16436 11100 16464
rect 11238 16436 11244 16448
rect 10459 16408 11100 16436
rect 11199 16408 11244 16436
rect 10459 16405 10471 16408
rect 10413 16399 10471 16405
rect 11238 16396 11244 16408
rect 11296 16396 11302 16448
rect 11900 16445 11928 16476
rect 12406 16476 13268 16504
rect 11885 16439 11943 16445
rect 11885 16405 11897 16439
rect 11931 16436 11943 16439
rect 11974 16436 11980 16448
rect 11931 16408 11980 16436
rect 11931 16405 11943 16408
rect 11885 16399 11943 16405
rect 11974 16396 11980 16408
rect 12032 16396 12038 16448
rect 12253 16439 12311 16445
rect 12253 16405 12265 16439
rect 12299 16436 12311 16439
rect 12406 16436 12434 16476
rect 13262 16464 13268 16476
rect 13320 16464 13326 16516
rect 13372 16504 13400 16532
rect 15396 16504 15424 16612
rect 15473 16609 15485 16612
rect 15519 16609 15531 16643
rect 16206 16640 16212 16652
rect 16167 16612 16212 16640
rect 15473 16603 15531 16609
rect 16206 16600 16212 16612
rect 16264 16600 16270 16652
rect 17037 16643 17095 16649
rect 17037 16609 17049 16643
rect 17083 16640 17095 16643
rect 17218 16640 17224 16652
rect 17083 16612 17224 16640
rect 17083 16609 17095 16612
rect 17037 16603 17095 16609
rect 17218 16600 17224 16612
rect 17276 16600 17282 16652
rect 16390 16532 16396 16584
rect 16448 16572 16454 16584
rect 16853 16575 16911 16581
rect 16853 16572 16865 16575
rect 16448 16544 16865 16572
rect 16448 16532 16454 16544
rect 16853 16541 16865 16544
rect 16899 16572 16911 16575
rect 17604 16572 17632 16748
rect 19518 16736 19524 16748
rect 19576 16776 19582 16788
rect 19978 16776 19984 16788
rect 19576 16748 19984 16776
rect 19576 16736 19582 16748
rect 19978 16736 19984 16748
rect 20036 16736 20042 16788
rect 20530 16776 20536 16788
rect 20491 16748 20536 16776
rect 20530 16736 20536 16748
rect 20588 16736 20594 16788
rect 20809 16779 20867 16785
rect 20809 16745 20821 16779
rect 20855 16776 20867 16779
rect 21266 16776 21272 16788
rect 20855 16748 21272 16776
rect 20855 16745 20867 16748
rect 20809 16739 20867 16745
rect 21266 16736 21272 16748
rect 21324 16736 21330 16788
rect 21085 16711 21143 16717
rect 17696 16680 20852 16708
rect 17696 16649 17724 16680
rect 20824 16652 20852 16680
rect 21085 16677 21097 16711
rect 21131 16677 21143 16711
rect 21085 16671 21143 16677
rect 17681 16643 17739 16649
rect 17681 16609 17693 16643
rect 17727 16609 17739 16643
rect 17681 16603 17739 16609
rect 17770 16600 17776 16652
rect 17828 16640 17834 16652
rect 18141 16643 18199 16649
rect 18141 16640 18153 16643
rect 17828 16612 17873 16640
rect 17963 16612 18153 16640
rect 17828 16600 17834 16612
rect 16899 16544 17632 16572
rect 16899 16541 16911 16544
rect 16853 16535 16911 16541
rect 13372 16476 15424 16504
rect 16761 16507 16819 16513
rect 16761 16473 16773 16507
rect 16807 16504 16819 16507
rect 16942 16504 16948 16516
rect 16807 16476 16948 16504
rect 16807 16473 16819 16476
rect 16761 16467 16819 16473
rect 16942 16464 16948 16476
rect 17000 16464 17006 16516
rect 17963 16504 17991 16612
rect 18141 16609 18153 16612
rect 18187 16640 18199 16643
rect 19794 16640 19800 16652
rect 18187 16612 19800 16640
rect 18187 16609 18199 16612
rect 18141 16603 18199 16609
rect 19794 16600 19800 16612
rect 19852 16600 19858 16652
rect 19889 16643 19947 16649
rect 19889 16609 19901 16643
rect 19935 16640 19947 16643
rect 20254 16640 20260 16652
rect 19935 16612 20260 16640
rect 19935 16609 19947 16612
rect 19889 16603 19947 16609
rect 20254 16600 20260 16612
rect 20312 16600 20318 16652
rect 20806 16600 20812 16652
rect 20864 16600 20870 16652
rect 21100 16584 21128 16671
rect 18046 16532 18052 16584
rect 18104 16572 18110 16584
rect 20165 16575 20223 16581
rect 20165 16572 20177 16575
rect 18104 16544 20177 16572
rect 18104 16532 18110 16544
rect 20165 16541 20177 16544
rect 20211 16572 20223 16575
rect 20349 16575 20407 16581
rect 20349 16572 20361 16575
rect 20211 16544 20361 16572
rect 20211 16541 20223 16544
rect 20165 16535 20223 16541
rect 20349 16541 20361 16544
rect 20395 16541 20407 16575
rect 20622 16572 20628 16584
rect 20583 16544 20628 16572
rect 20349 16535 20407 16541
rect 20622 16532 20628 16544
rect 20680 16532 20686 16584
rect 20901 16575 20959 16581
rect 20901 16541 20913 16575
rect 20947 16541 20959 16575
rect 20901 16535 20959 16541
rect 17052 16476 17991 16504
rect 12299 16408 12434 16436
rect 12299 16405 12311 16408
rect 12253 16399 12311 16405
rect 12526 16396 12532 16448
rect 12584 16436 12590 16448
rect 12713 16439 12771 16445
rect 12713 16436 12725 16439
rect 12584 16408 12725 16436
rect 12584 16396 12590 16408
rect 12713 16405 12725 16408
rect 12759 16436 12771 16439
rect 12986 16436 12992 16448
rect 12759 16408 12992 16436
rect 12759 16405 12771 16408
rect 12713 16399 12771 16405
rect 12986 16396 12992 16408
rect 13044 16396 13050 16448
rect 13170 16436 13176 16448
rect 13131 16408 13176 16436
rect 13170 16396 13176 16408
rect 13228 16396 13234 16448
rect 15470 16396 15476 16448
rect 15528 16436 15534 16448
rect 15565 16439 15623 16445
rect 15565 16436 15577 16439
rect 15528 16408 15577 16436
rect 15528 16396 15534 16408
rect 15565 16405 15577 16408
rect 15611 16405 15623 16439
rect 15930 16436 15936 16448
rect 15891 16408 15936 16436
rect 15565 16399 15623 16405
rect 15930 16396 15936 16408
rect 15988 16396 15994 16448
rect 16025 16439 16083 16445
rect 16025 16405 16037 16439
rect 16071 16436 16083 16439
rect 16114 16436 16120 16448
rect 16071 16408 16120 16436
rect 16071 16405 16083 16408
rect 16025 16399 16083 16405
rect 16114 16396 16120 16408
rect 16172 16436 16178 16448
rect 17052 16436 17080 16476
rect 20438 16464 20444 16516
rect 20496 16504 20502 16516
rect 20916 16504 20944 16535
rect 21082 16532 21088 16584
rect 21140 16532 21146 16584
rect 21269 16575 21327 16581
rect 21269 16541 21281 16575
rect 21315 16541 21327 16575
rect 21269 16535 21327 16541
rect 21284 16504 21312 16535
rect 20496 16476 20944 16504
rect 21008 16476 21312 16504
rect 20496 16464 20502 16476
rect 16172 16408 17080 16436
rect 16172 16396 16178 16408
rect 17494 16396 17500 16448
rect 17552 16436 17558 16448
rect 17589 16439 17647 16445
rect 17589 16436 17601 16439
rect 17552 16408 17601 16436
rect 17552 16396 17558 16408
rect 17589 16405 17601 16408
rect 17635 16405 17647 16439
rect 20070 16436 20076 16448
rect 20031 16408 20076 16436
rect 17589 16399 17647 16405
rect 20070 16396 20076 16408
rect 20128 16396 20134 16448
rect 20162 16396 20168 16448
rect 20220 16436 20226 16448
rect 21008 16436 21036 16476
rect 21450 16436 21456 16448
rect 20220 16408 21036 16436
rect 21411 16408 21456 16436
rect 20220 16396 20226 16408
rect 21450 16396 21456 16408
rect 21508 16396 21514 16448
rect 1104 16346 22056 16368
rect 14 16260 20 16312
rect 72 16300 78 16312
rect 934 16300 940 16312
rect 72 16272 940 16300
rect 72 16260 78 16272
rect 934 16260 940 16272
rect 992 16260 998 16312
rect 1104 16294 6148 16346
rect 6200 16294 6212 16346
rect 6264 16294 6276 16346
rect 6328 16294 6340 16346
rect 6392 16294 6404 16346
rect 6456 16294 11346 16346
rect 11398 16294 11410 16346
rect 11462 16294 11474 16346
rect 11526 16294 11538 16346
rect 11590 16294 11602 16346
rect 11654 16294 16544 16346
rect 16596 16294 16608 16346
rect 16660 16294 16672 16346
rect 16724 16294 16736 16346
rect 16788 16294 16800 16346
rect 16852 16294 21742 16346
rect 21794 16294 21806 16346
rect 21858 16294 21870 16346
rect 21922 16294 21934 16346
rect 21986 16294 21998 16346
rect 22050 16294 22056 16346
rect 1104 16272 22056 16294
rect 1857 16235 1915 16241
rect 1857 16201 1869 16235
rect 1903 16232 1915 16235
rect 2038 16232 2044 16244
rect 1903 16204 2044 16232
rect 1903 16201 1915 16204
rect 1857 16195 1915 16201
rect 2038 16192 2044 16204
rect 2096 16192 2102 16244
rect 2501 16235 2559 16241
rect 2501 16201 2513 16235
rect 2547 16232 2559 16235
rect 2961 16235 3019 16241
rect 2961 16232 2973 16235
rect 2547 16204 2973 16232
rect 2547 16201 2559 16204
rect 2501 16195 2559 16201
rect 2961 16201 2973 16204
rect 3007 16201 3019 16235
rect 2961 16195 3019 16201
rect 5626 16192 5632 16244
rect 5684 16232 5690 16244
rect 5721 16235 5779 16241
rect 5721 16232 5733 16235
rect 5684 16204 5733 16232
rect 5684 16192 5690 16204
rect 5721 16201 5733 16204
rect 5767 16201 5779 16235
rect 5721 16195 5779 16201
rect 4614 16173 4620 16176
rect 4608 16164 4620 16173
rect 1688 16136 4108 16164
rect 4575 16136 4620 16164
rect 1688 16105 1716 16136
rect 1673 16099 1731 16105
rect 1673 16065 1685 16099
rect 1719 16065 1731 16099
rect 1673 16059 1731 16065
rect 2041 16099 2099 16105
rect 2041 16065 2053 16099
rect 2087 16096 2099 16099
rect 2130 16096 2136 16108
rect 2087 16068 2136 16096
rect 2087 16065 2099 16068
rect 2041 16059 2099 16065
rect 2130 16056 2136 16068
rect 2188 16056 2194 16108
rect 3329 16099 3387 16105
rect 3329 16065 3341 16099
rect 3375 16096 3387 16099
rect 3789 16099 3847 16105
rect 3789 16096 3801 16099
rect 3375 16068 3801 16096
rect 3375 16065 3387 16068
rect 3329 16059 3387 16065
rect 3789 16065 3801 16068
rect 3835 16065 3847 16099
rect 3789 16059 3847 16065
rect 2222 16028 2228 16040
rect 2183 16000 2228 16028
rect 2222 15988 2228 16000
rect 2280 15988 2286 16040
rect 2406 16028 2412 16040
rect 2367 16000 2412 16028
rect 2406 15988 2412 16000
rect 2464 15988 2470 16040
rect 3234 15988 3240 16040
rect 3292 16028 3298 16040
rect 3421 16031 3479 16037
rect 3421 16028 3433 16031
rect 3292 16000 3433 16028
rect 3292 15988 3298 16000
rect 3421 15997 3433 16000
rect 3467 15997 3479 16031
rect 3421 15991 3479 15997
rect 3605 16031 3663 16037
rect 3605 15997 3617 16031
rect 3651 16028 3663 16031
rect 3878 16028 3884 16040
rect 3651 16000 3884 16028
rect 3651 15997 3663 16000
rect 3605 15991 3663 15997
rect 3878 15988 3884 16000
rect 3936 15988 3942 16040
rect 106 15920 112 15972
rect 164 15960 170 15972
rect 2869 15963 2927 15969
rect 164 15932 2840 15960
rect 164 15920 170 15932
rect 1486 15892 1492 15904
rect 1447 15864 1492 15892
rect 1486 15852 1492 15864
rect 1544 15852 1550 15904
rect 2812 15892 2840 15932
rect 2869 15929 2881 15963
rect 2915 15960 2927 15963
rect 3142 15960 3148 15972
rect 2915 15932 3148 15960
rect 2915 15929 2927 15932
rect 2869 15923 2927 15929
rect 3142 15920 3148 15932
rect 3200 15920 3206 15972
rect 4080 15969 4108 16136
rect 4608 16127 4620 16136
rect 4614 16124 4620 16127
rect 4672 16124 4678 16176
rect 5258 16124 5264 16176
rect 5316 16124 5322 16176
rect 5736 16164 5764 16195
rect 5994 16192 6000 16244
rect 6052 16232 6058 16244
rect 6089 16235 6147 16241
rect 6089 16232 6101 16235
rect 6052 16204 6101 16232
rect 6052 16192 6058 16204
rect 6089 16201 6101 16204
rect 6135 16201 6147 16235
rect 6089 16195 6147 16201
rect 8021 16235 8079 16241
rect 8021 16201 8033 16235
rect 8067 16201 8079 16235
rect 8021 16195 8079 16201
rect 9493 16235 9551 16241
rect 9493 16201 9505 16235
rect 9539 16232 9551 16235
rect 10134 16232 10140 16244
rect 9539 16204 10140 16232
rect 9539 16201 9551 16204
rect 9493 16195 9551 16201
rect 6178 16164 6184 16176
rect 5736 16136 6184 16164
rect 6178 16124 6184 16136
rect 6236 16124 6242 16176
rect 6908 16167 6966 16173
rect 6908 16133 6920 16167
rect 6954 16164 6966 16167
rect 7006 16164 7012 16176
rect 6954 16136 7012 16164
rect 6954 16133 6966 16136
rect 6908 16127 6966 16133
rect 7006 16124 7012 16136
rect 7064 16124 7070 16176
rect 8036 16164 8064 16195
rect 10134 16192 10140 16204
rect 10192 16192 10198 16244
rect 10413 16235 10471 16241
rect 10413 16201 10425 16235
rect 10459 16232 10471 16235
rect 10873 16235 10931 16241
rect 10873 16232 10885 16235
rect 10459 16204 10885 16232
rect 10459 16201 10471 16204
rect 10413 16195 10471 16201
rect 10873 16201 10885 16204
rect 10919 16201 10931 16235
rect 10873 16195 10931 16201
rect 11330 16192 11336 16244
rect 11388 16232 11394 16244
rect 12158 16232 12164 16244
rect 11388 16204 12020 16232
rect 12119 16204 12164 16232
rect 11388 16192 11394 16204
rect 11992 16173 12020 16204
rect 12158 16192 12164 16204
rect 12216 16192 12222 16244
rect 12437 16235 12495 16241
rect 12437 16201 12449 16235
rect 12483 16232 12495 16235
rect 12710 16232 12716 16244
rect 12483 16204 12716 16232
rect 12483 16201 12495 16204
rect 12437 16195 12495 16201
rect 12710 16192 12716 16204
rect 12768 16192 12774 16244
rect 15378 16192 15384 16244
rect 15436 16232 15442 16244
rect 15473 16235 15531 16241
rect 15473 16232 15485 16235
rect 15436 16204 15485 16232
rect 15436 16192 15442 16204
rect 15473 16201 15485 16204
rect 15519 16201 15531 16235
rect 15473 16195 15531 16201
rect 15746 16192 15752 16244
rect 15804 16232 15810 16244
rect 19613 16235 19671 16241
rect 19613 16232 19625 16235
rect 15804 16204 19625 16232
rect 15804 16192 15810 16204
rect 19613 16201 19625 16204
rect 19659 16232 19671 16235
rect 19659 16204 20107 16232
rect 19659 16201 19671 16204
rect 19613 16195 19671 16201
rect 8358 16167 8416 16173
rect 8358 16164 8370 16167
rect 8036 16136 8370 16164
rect 8358 16133 8370 16136
rect 8404 16164 8416 16167
rect 10045 16167 10103 16173
rect 8404 16136 9812 16164
rect 8404 16133 8416 16136
rect 8358 16127 8416 16133
rect 4249 16099 4307 16105
rect 4249 16065 4261 16099
rect 4295 16065 4307 16099
rect 4249 16059 4307 16065
rect 4341 16099 4399 16105
rect 4341 16065 4353 16099
rect 4387 16096 4399 16099
rect 4430 16096 4436 16108
rect 4387 16068 4436 16096
rect 4387 16065 4399 16068
rect 4341 16059 4399 16065
rect 4264 16028 4292 16059
rect 4430 16056 4436 16068
rect 4488 16056 4494 16108
rect 5276 16096 5304 16124
rect 5813 16099 5871 16105
rect 5813 16096 5825 16099
rect 5276 16068 5825 16096
rect 5813 16065 5825 16068
rect 5859 16096 5871 16099
rect 5994 16096 6000 16108
rect 5859 16068 6000 16096
rect 5859 16065 5871 16068
rect 5813 16059 5871 16065
rect 5994 16056 6000 16068
rect 6052 16056 6058 16108
rect 7190 16056 7196 16108
rect 7248 16096 7254 16108
rect 7834 16096 7840 16108
rect 7248 16068 7840 16096
rect 7248 16056 7254 16068
rect 7834 16056 7840 16068
rect 7892 16056 7898 16108
rect 8110 16096 8116 16108
rect 8071 16068 8116 16096
rect 8110 16056 8116 16068
rect 8168 16056 8174 16108
rect 8754 16056 8760 16108
rect 8812 16096 8818 16108
rect 9398 16096 9404 16108
rect 8812 16068 9404 16096
rect 8812 16056 8818 16068
rect 9398 16056 9404 16068
rect 9456 16056 9462 16108
rect 6362 16028 6368 16040
rect 4264 16000 4384 16028
rect 6323 16000 6368 16028
rect 4065 15963 4123 15969
rect 4065 15929 4077 15963
rect 4111 15929 4123 15963
rect 4065 15923 4123 15929
rect 4246 15892 4252 15904
rect 2812 15864 4252 15892
rect 4246 15852 4252 15864
rect 4304 15852 4310 15904
rect 4356 15892 4384 16000
rect 6362 15988 6368 16000
rect 6420 15988 6426 16040
rect 6641 16031 6699 16037
rect 6641 15997 6653 16031
rect 6687 15997 6699 16031
rect 6641 15991 6699 15997
rect 5442 15892 5448 15904
rect 4356 15864 5448 15892
rect 5442 15852 5448 15864
rect 5500 15852 5506 15904
rect 5997 15895 6055 15901
rect 5997 15861 6009 15895
rect 6043 15892 6055 15895
rect 6546 15892 6552 15904
rect 6043 15864 6552 15892
rect 6043 15861 6055 15864
rect 5997 15855 6055 15861
rect 6546 15852 6552 15864
rect 6604 15852 6610 15904
rect 6656 15892 6684 15991
rect 9674 15988 9680 16040
rect 9732 16028 9738 16040
rect 9784 16037 9812 16136
rect 10045 16133 10057 16167
rect 10091 16164 10103 16167
rect 11977 16167 12035 16173
rect 10091 16136 11560 16164
rect 10091 16133 10103 16136
rect 10045 16127 10103 16133
rect 10060 16096 10088 16127
rect 9876 16068 10088 16096
rect 9769 16031 9827 16037
rect 9769 16028 9781 16031
rect 9732 16000 9781 16028
rect 9732 15988 9738 16000
rect 9769 15997 9781 16000
rect 9815 15997 9827 16031
rect 9769 15991 9827 15997
rect 9582 15920 9588 15972
rect 9640 15960 9646 15972
rect 9876 15960 9904 16068
rect 10134 16056 10140 16108
rect 10192 16096 10198 16108
rect 10192 16068 11100 16096
rect 10192 16056 10198 16068
rect 9953 16031 10011 16037
rect 9953 15997 9965 16031
rect 9999 16028 10011 16031
rect 10778 16028 10784 16040
rect 9999 16000 10784 16028
rect 9999 15997 10011 16000
rect 9953 15991 10011 15997
rect 10778 15988 10784 16000
rect 10836 15988 10842 16040
rect 10962 16028 10968 16040
rect 10923 16000 10968 16028
rect 10962 15988 10968 16000
rect 11020 15988 11026 16040
rect 11072 16037 11100 16068
rect 11532 16040 11560 16136
rect 11977 16133 11989 16167
rect 12023 16164 12035 16167
rect 12066 16164 12072 16176
rect 12023 16136 12072 16164
rect 12023 16133 12035 16136
rect 11977 16127 12035 16133
rect 12066 16124 12072 16136
rect 12124 16124 12130 16176
rect 13354 16124 13360 16176
rect 13412 16124 13418 16176
rect 13572 16167 13630 16173
rect 13572 16133 13584 16167
rect 13618 16164 13630 16167
rect 14185 16167 14243 16173
rect 14185 16164 14197 16167
rect 13618 16136 14197 16164
rect 13618 16133 13630 16136
rect 13572 16127 13630 16133
rect 14185 16133 14197 16136
rect 14231 16164 14243 16167
rect 14274 16164 14280 16176
rect 14231 16136 14280 16164
rect 14231 16133 14243 16136
rect 14185 16127 14243 16133
rect 14274 16124 14280 16136
rect 14332 16164 14338 16176
rect 14332 16136 14596 16164
rect 14332 16124 14338 16136
rect 11606 16056 11612 16108
rect 11664 16096 11670 16108
rect 11701 16099 11759 16105
rect 11701 16096 11713 16099
rect 11664 16068 11713 16096
rect 11664 16056 11670 16068
rect 11701 16065 11713 16068
rect 11747 16065 11759 16099
rect 11701 16059 11759 16065
rect 11790 16056 11796 16108
rect 11848 16096 11854 16108
rect 13170 16096 13176 16108
rect 11848 16068 13176 16096
rect 11848 16056 11854 16068
rect 13170 16056 13176 16068
rect 13228 16056 13234 16108
rect 13372 16096 13400 16124
rect 14568 16105 14596 16136
rect 15930 16124 15936 16176
rect 15988 16164 15994 16176
rect 16393 16167 16451 16173
rect 16393 16164 16405 16167
rect 15988 16136 16405 16164
rect 15988 16124 15994 16136
rect 16393 16133 16405 16136
rect 16439 16164 16451 16167
rect 17862 16164 17868 16176
rect 16439 16136 17868 16164
rect 16439 16133 16451 16136
rect 16393 16127 16451 16133
rect 17862 16124 17868 16136
rect 17920 16124 17926 16176
rect 17954 16124 17960 16176
rect 18012 16164 18018 16176
rect 19521 16167 19579 16173
rect 19521 16164 19533 16167
rect 18012 16136 19533 16164
rect 18012 16124 18018 16136
rect 19521 16133 19533 16136
rect 19567 16164 19579 16167
rect 19702 16164 19708 16176
rect 19567 16136 19708 16164
rect 19567 16133 19579 16136
rect 19521 16127 19579 16133
rect 19702 16124 19708 16136
rect 19760 16124 19766 16176
rect 13817 16099 13875 16105
rect 13817 16096 13829 16099
rect 13372 16068 13829 16096
rect 13817 16065 13829 16068
rect 13863 16065 13875 16099
rect 13817 16059 13875 16065
rect 14553 16099 14611 16105
rect 14553 16065 14565 16099
rect 14599 16065 14611 16099
rect 15102 16096 15108 16108
rect 15015 16068 15108 16096
rect 14553 16059 14611 16065
rect 15102 16056 15108 16068
rect 15160 16096 15166 16108
rect 16114 16096 16120 16108
rect 15160 16068 16120 16096
rect 15160 16056 15166 16068
rect 16114 16056 16120 16068
rect 16172 16056 16178 16108
rect 17405 16099 17463 16105
rect 17405 16065 17417 16099
rect 17451 16065 17463 16099
rect 17405 16059 17463 16065
rect 11057 16031 11115 16037
rect 11057 15997 11069 16031
rect 11103 15997 11115 16031
rect 11514 16028 11520 16040
rect 11475 16000 11520 16028
rect 11057 15991 11115 15997
rect 11514 15988 11520 16000
rect 11572 15988 11578 16040
rect 14918 16028 14924 16040
rect 14879 16000 14924 16028
rect 14918 15988 14924 16000
rect 14976 15988 14982 16040
rect 15010 15988 15016 16040
rect 15068 16028 15074 16040
rect 15068 16000 15113 16028
rect 15068 15988 15074 16000
rect 15378 15988 15384 16040
rect 15436 16028 15442 16040
rect 17126 16028 17132 16040
rect 15436 16000 16988 16028
rect 17087 16000 17132 16028
rect 15436 15988 15442 16000
rect 9640 15932 9904 15960
rect 9640 15920 9646 15932
rect 10318 15920 10324 15972
rect 10376 15960 10382 15972
rect 16960 15960 16988 16000
rect 17126 15988 17132 16000
rect 17184 16028 17190 16040
rect 17420 16028 17448 16059
rect 17678 16056 17684 16108
rect 17736 16096 17742 16108
rect 18785 16099 18843 16105
rect 18785 16096 18797 16099
rect 17736 16068 18797 16096
rect 17736 16056 17742 16068
rect 18785 16065 18797 16068
rect 18831 16065 18843 16099
rect 18785 16059 18843 16065
rect 18892 16068 19288 16096
rect 17184 16000 17448 16028
rect 17184 15988 17190 16000
rect 18892 15960 18920 16068
rect 18966 15988 18972 16040
rect 19024 15988 19030 16040
rect 19058 15988 19064 16040
rect 19116 16028 19122 16040
rect 19116 16000 19161 16028
rect 19116 15988 19122 16000
rect 10376 15932 12940 15960
rect 16960 15932 18920 15960
rect 10376 15920 10382 15932
rect 12912 15904 12940 15932
rect 8294 15892 8300 15904
rect 6656 15864 8300 15892
rect 8294 15852 8300 15864
rect 8352 15892 8358 15904
rect 8846 15892 8852 15904
rect 8352 15864 8852 15892
rect 8352 15852 8358 15864
rect 8846 15852 8852 15864
rect 8904 15852 8910 15904
rect 9766 15852 9772 15904
rect 9824 15892 9830 15904
rect 10505 15895 10563 15901
rect 10505 15892 10517 15895
rect 9824 15864 10517 15892
rect 9824 15852 9830 15864
rect 10505 15861 10517 15864
rect 10551 15861 10563 15895
rect 10505 15855 10563 15861
rect 10870 15852 10876 15904
rect 10928 15892 10934 15904
rect 12253 15895 12311 15901
rect 12253 15892 12265 15895
rect 10928 15864 12265 15892
rect 10928 15852 10934 15864
rect 12253 15861 12265 15864
rect 12299 15861 12311 15895
rect 12253 15855 12311 15861
rect 12894 15852 12900 15904
rect 12952 15852 12958 15904
rect 13446 15852 13452 15904
rect 13504 15892 13510 15904
rect 16209 15895 16267 15901
rect 16209 15892 16221 15895
rect 13504 15864 16221 15892
rect 13504 15852 13510 15864
rect 16209 15861 16221 15864
rect 16255 15892 16267 15895
rect 16390 15892 16396 15904
rect 16255 15864 16396 15892
rect 16255 15861 16267 15864
rect 16209 15855 16267 15861
rect 16390 15852 16396 15864
rect 16448 15852 16454 15904
rect 17586 15852 17592 15904
rect 17644 15892 17650 15904
rect 18874 15892 18880 15904
rect 17644 15864 18880 15892
rect 17644 15852 17650 15864
rect 18874 15852 18880 15864
rect 18932 15852 18938 15904
rect 18984 15901 19012 15988
rect 19260 15960 19288 16068
rect 19794 16056 19800 16108
rect 19852 16096 19858 16108
rect 19904 16105 20033 16120
rect 19904 16099 20039 16105
rect 19904 16096 19993 16099
rect 19852 16092 19993 16096
rect 19852 16068 19932 16092
rect 19852 16056 19858 16068
rect 19981 16065 19993 16092
rect 20027 16065 20039 16099
rect 20079 16096 20107 16204
rect 20162 16192 20168 16244
rect 20220 16232 20226 16244
rect 20717 16235 20775 16241
rect 20220 16204 20265 16232
rect 20220 16192 20226 16204
rect 20717 16201 20729 16235
rect 20763 16201 20775 16235
rect 20990 16232 20996 16244
rect 20951 16204 20996 16232
rect 20717 16195 20775 16201
rect 20732 16164 20760 16195
rect 20990 16192 20996 16204
rect 21048 16192 21054 16244
rect 20364 16136 20692 16164
rect 20732 16136 21312 16164
rect 20257 16099 20315 16105
rect 20257 16096 20269 16099
rect 20079 16068 20269 16096
rect 19981 16059 20039 16065
rect 20257 16065 20269 16068
rect 20303 16065 20315 16099
rect 20257 16059 20315 16065
rect 19337 16031 19395 16037
rect 19337 15997 19349 16031
rect 19383 16028 19395 16031
rect 20364 16028 20392 16136
rect 20438 16056 20444 16108
rect 20496 16056 20502 16108
rect 20530 16056 20536 16108
rect 20588 16096 20594 16108
rect 20588 16068 20633 16096
rect 20588 16056 20594 16068
rect 19383 16000 20392 16028
rect 19383 15997 19395 16000
rect 19337 15991 19395 15997
rect 20456 15969 20484 16056
rect 20664 16028 20692 16136
rect 20806 16096 20812 16108
rect 20767 16068 20812 16096
rect 20806 16056 20812 16068
rect 20864 16056 20870 16108
rect 21284 16105 21312 16136
rect 21269 16099 21327 16105
rect 21269 16065 21281 16099
rect 21315 16065 21327 16099
rect 21269 16059 21327 16065
rect 22094 16028 22100 16040
rect 20664 16000 22100 16028
rect 22094 15988 22100 16000
rect 22152 15988 22158 16040
rect 20441 15963 20499 15969
rect 19260 15932 20116 15960
rect 18969 15895 19027 15901
rect 18969 15861 18981 15895
rect 19015 15861 19027 15895
rect 18969 15855 19027 15861
rect 19610 15852 19616 15904
rect 19668 15892 19674 15904
rect 19794 15892 19800 15904
rect 19668 15864 19800 15892
rect 19668 15852 19674 15864
rect 19794 15852 19800 15864
rect 19852 15852 19858 15904
rect 20088 15892 20116 15932
rect 20441 15929 20453 15963
rect 20487 15929 20499 15963
rect 20441 15923 20499 15929
rect 20530 15892 20536 15904
rect 20088 15864 20536 15892
rect 20530 15852 20536 15864
rect 20588 15892 20594 15904
rect 21085 15895 21143 15901
rect 21085 15892 21097 15895
rect 20588 15864 21097 15892
rect 20588 15852 20594 15864
rect 21085 15861 21097 15864
rect 21131 15861 21143 15895
rect 21450 15892 21456 15904
rect 21411 15864 21456 15892
rect 21085 15855 21143 15861
rect 21450 15852 21456 15864
rect 21508 15852 21514 15904
rect 1104 15802 21896 15824
rect 1104 15750 3549 15802
rect 3601 15750 3613 15802
rect 3665 15750 3677 15802
rect 3729 15750 3741 15802
rect 3793 15750 3805 15802
rect 3857 15750 8747 15802
rect 8799 15750 8811 15802
rect 8863 15750 8875 15802
rect 8927 15750 8939 15802
rect 8991 15750 9003 15802
rect 9055 15750 13945 15802
rect 13997 15750 14009 15802
rect 14061 15750 14073 15802
rect 14125 15750 14137 15802
rect 14189 15750 14201 15802
rect 14253 15750 19143 15802
rect 19195 15750 19207 15802
rect 19259 15750 19271 15802
rect 19323 15750 19335 15802
rect 19387 15750 19399 15802
rect 19451 15750 21896 15802
rect 1104 15728 21896 15750
rect 1670 15648 1676 15700
rect 1728 15688 1734 15700
rect 2133 15691 2191 15697
rect 2133 15688 2145 15691
rect 1728 15660 2145 15688
rect 1728 15648 1734 15660
rect 2133 15657 2145 15660
rect 2179 15657 2191 15691
rect 3605 15691 3663 15697
rect 2133 15651 2191 15657
rect 2332 15660 2636 15688
rect 2041 15623 2099 15629
rect 2041 15589 2053 15623
rect 2087 15620 2099 15623
rect 2332 15620 2360 15660
rect 2087 15592 2360 15620
rect 2409 15623 2467 15629
rect 2087 15589 2099 15592
rect 2041 15583 2099 15589
rect 2409 15589 2421 15623
rect 2455 15589 2467 15623
rect 2409 15583 2467 15589
rect 2424 15552 2452 15583
rect 1688 15524 2452 15552
rect 1688 15493 1716 15524
rect 1673 15487 1731 15493
rect 1673 15453 1685 15487
rect 1719 15453 1731 15487
rect 1673 15447 1731 15453
rect 1857 15487 1915 15493
rect 1857 15453 1869 15487
rect 1903 15484 1915 15487
rect 2314 15484 2320 15496
rect 1903 15456 2176 15484
rect 2275 15456 2320 15484
rect 1903 15453 1915 15456
rect 1857 15447 1915 15453
rect 1486 15348 1492 15360
rect 1447 15320 1492 15348
rect 1486 15308 1492 15320
rect 1544 15308 1550 15360
rect 2148 15348 2176 15456
rect 2314 15444 2320 15456
rect 2372 15444 2378 15496
rect 2608 15493 2636 15660
rect 3605 15657 3617 15691
rect 3651 15688 3663 15691
rect 4154 15688 4160 15700
rect 3651 15660 4160 15688
rect 3651 15657 3663 15660
rect 3605 15651 3663 15657
rect 4154 15648 4160 15660
rect 4212 15648 4218 15700
rect 4338 15688 4344 15700
rect 4299 15660 4344 15688
rect 4338 15648 4344 15660
rect 4396 15648 4402 15700
rect 4982 15648 4988 15700
rect 5040 15688 5046 15700
rect 5629 15691 5687 15697
rect 5629 15688 5641 15691
rect 5040 15660 5641 15688
rect 5040 15648 5046 15660
rect 5629 15657 5641 15660
rect 5675 15657 5687 15691
rect 5629 15651 5687 15657
rect 6638 15648 6644 15700
rect 6696 15688 6702 15700
rect 6733 15691 6791 15697
rect 6733 15688 6745 15691
rect 6696 15660 6745 15688
rect 6696 15648 6702 15660
rect 6733 15657 6745 15660
rect 6779 15657 6791 15691
rect 6733 15651 6791 15657
rect 6822 15648 6828 15700
rect 6880 15688 6886 15700
rect 6917 15691 6975 15697
rect 6917 15688 6929 15691
rect 6880 15660 6929 15688
rect 6880 15648 6886 15660
rect 6917 15657 6929 15660
rect 6963 15657 6975 15691
rect 6917 15651 6975 15657
rect 7466 15648 7472 15700
rect 7524 15648 7530 15700
rect 8665 15691 8723 15697
rect 8665 15688 8677 15691
rect 7852 15660 8677 15688
rect 3418 15580 3424 15632
rect 3476 15620 3482 15632
rect 3789 15623 3847 15629
rect 3789 15620 3801 15623
rect 3476 15592 3801 15620
rect 3476 15580 3482 15592
rect 3789 15589 3801 15592
rect 3835 15589 3847 15623
rect 5537 15623 5595 15629
rect 3789 15583 3847 15589
rect 4080 15592 5488 15620
rect 2958 15552 2964 15564
rect 2919 15524 2964 15552
rect 2958 15512 2964 15524
rect 3016 15552 3022 15564
rect 3878 15552 3884 15564
rect 3016 15524 3884 15552
rect 3016 15512 3022 15524
rect 3878 15512 3884 15524
rect 3936 15512 3942 15564
rect 3973 15503 4031 15509
rect 2593 15487 2651 15493
rect 2593 15453 2605 15487
rect 2639 15453 2651 15487
rect 2593 15447 2651 15453
rect 2777 15487 2835 15493
rect 2777 15453 2789 15487
rect 2823 15484 2835 15487
rect 3786 15484 3792 15496
rect 2823 15456 3792 15484
rect 2823 15453 2835 15456
rect 2777 15447 2835 15453
rect 3786 15444 3792 15456
rect 3844 15444 3850 15496
rect 3973 15469 3985 15503
rect 4019 15500 4031 15503
rect 4080 15500 4108 15592
rect 4614 15512 4620 15564
rect 4672 15552 4678 15564
rect 5077 15555 5135 15561
rect 5077 15552 5089 15555
rect 4672 15524 5089 15552
rect 4672 15512 4678 15524
rect 5077 15521 5089 15524
rect 5123 15521 5135 15555
rect 5460 15552 5488 15592
rect 5537 15589 5549 15623
rect 5583 15620 5595 15623
rect 5902 15620 5908 15632
rect 5583 15592 5908 15620
rect 5583 15589 5595 15592
rect 5537 15583 5595 15589
rect 5902 15580 5908 15592
rect 5960 15580 5966 15632
rect 7484 15620 7512 15648
rect 7852 15620 7880 15660
rect 8665 15657 8677 15660
rect 8711 15688 8723 15691
rect 9306 15688 9312 15700
rect 8711 15660 9312 15688
rect 8711 15657 8723 15660
rect 8665 15651 8723 15657
rect 9306 15648 9312 15660
rect 9364 15648 9370 15700
rect 9858 15648 9864 15700
rect 9916 15688 9922 15700
rect 9953 15691 10011 15697
rect 9953 15688 9965 15691
rect 9916 15660 9965 15688
rect 9916 15648 9922 15660
rect 9953 15657 9965 15660
rect 9999 15657 10011 15691
rect 10778 15688 10784 15700
rect 10739 15660 10784 15688
rect 9953 15651 10011 15657
rect 10778 15648 10784 15660
rect 10836 15648 10842 15700
rect 11238 15648 11244 15700
rect 11296 15688 11302 15700
rect 12894 15688 12900 15700
rect 11296 15660 12900 15688
rect 11296 15648 11302 15660
rect 12894 15648 12900 15660
rect 12952 15648 12958 15700
rect 13081 15691 13139 15697
rect 13081 15657 13093 15691
rect 13127 15688 13139 15691
rect 15838 15688 15844 15700
rect 13127 15660 15844 15688
rect 13127 15657 13139 15660
rect 13081 15651 13139 15657
rect 15838 15648 15844 15660
rect 15896 15648 15902 15700
rect 16114 15648 16120 15700
rect 16172 15688 16178 15700
rect 19610 15688 19616 15700
rect 16172 15660 19616 15688
rect 16172 15648 16178 15660
rect 19610 15648 19616 15660
rect 19668 15648 19674 15700
rect 20441 15691 20499 15697
rect 20441 15657 20453 15691
rect 20487 15688 20499 15691
rect 20806 15688 20812 15700
rect 20487 15660 20812 15688
rect 20487 15657 20499 15660
rect 20441 15651 20499 15657
rect 20806 15648 20812 15660
rect 20864 15648 20870 15700
rect 6012 15592 7880 15620
rect 6012 15552 6040 15592
rect 7926 15580 7932 15632
rect 7984 15620 7990 15632
rect 8570 15620 8576 15632
rect 7984 15592 8576 15620
rect 7984 15580 7990 15592
rect 8570 15580 8576 15592
rect 8628 15580 8634 15632
rect 8956 15592 10640 15620
rect 6178 15552 6184 15564
rect 5460 15524 6040 15552
rect 6139 15524 6184 15552
rect 5077 15515 5135 15521
rect 6178 15512 6184 15524
rect 6236 15512 6242 15564
rect 7282 15512 7288 15564
rect 7340 15552 7346 15564
rect 7469 15555 7527 15561
rect 7469 15552 7481 15555
rect 7340 15524 7481 15552
rect 7340 15512 7346 15524
rect 7469 15521 7481 15524
rect 7515 15521 7527 15555
rect 7834 15552 7840 15564
rect 7795 15524 7840 15552
rect 7469 15515 7527 15521
rect 7834 15512 7840 15524
rect 7892 15512 7898 15564
rect 8110 15512 8116 15564
rect 8168 15552 8174 15564
rect 8956 15561 8984 15592
rect 8941 15555 8999 15561
rect 8941 15552 8953 15555
rect 8168 15524 8953 15552
rect 8168 15512 8174 15524
rect 8941 15521 8953 15524
rect 8987 15521 8999 15555
rect 8941 15515 8999 15521
rect 9309 15555 9367 15561
rect 9309 15521 9321 15555
rect 9355 15552 9367 15555
rect 9674 15552 9680 15564
rect 9355 15524 9680 15552
rect 9355 15521 9367 15524
rect 9309 15515 9367 15521
rect 9674 15512 9680 15524
rect 9732 15552 9738 15564
rect 10505 15555 10563 15561
rect 10505 15552 10517 15555
rect 9732 15524 10517 15552
rect 9732 15512 9738 15524
rect 10505 15521 10517 15524
rect 10551 15521 10563 15555
rect 10505 15515 10563 15521
rect 4019 15472 4108 15500
rect 4246 15484 4252 15496
rect 4019 15469 4031 15472
rect 3973 15463 4031 15469
rect 4207 15456 4252 15484
rect 4246 15444 4252 15456
rect 4304 15444 4310 15496
rect 4982 15444 4988 15496
rect 5040 15484 5046 15496
rect 5040 15456 5085 15484
rect 5040 15444 5046 15456
rect 5258 15444 5264 15496
rect 5316 15484 5322 15496
rect 5353 15487 5411 15493
rect 5353 15484 5365 15487
rect 5316 15456 5365 15484
rect 5316 15444 5322 15456
rect 5353 15453 5365 15456
rect 5399 15453 5411 15487
rect 6089 15487 6147 15493
rect 6089 15484 6101 15487
rect 5353 15447 5411 15453
rect 5552 15456 6101 15484
rect 3237 15419 3295 15425
rect 3237 15385 3249 15419
rect 3283 15416 3295 15419
rect 3283 15388 4568 15416
rect 3283 15385 3295 15388
rect 3237 15379 3295 15385
rect 2958 15348 2964 15360
rect 2148 15320 2964 15348
rect 2958 15308 2964 15320
rect 3016 15308 3022 15360
rect 3142 15348 3148 15360
rect 3103 15320 3148 15348
rect 3142 15308 3148 15320
rect 3200 15308 3206 15360
rect 4062 15348 4068 15360
rect 4023 15320 4068 15348
rect 4062 15308 4068 15320
rect 4120 15308 4126 15360
rect 4540 15357 4568 15388
rect 4706 15376 4712 15428
rect 4764 15416 4770 15428
rect 5552 15416 5580 15456
rect 6089 15453 6101 15456
rect 6135 15453 6147 15487
rect 6089 15447 6147 15453
rect 7377 15487 7435 15493
rect 7377 15453 7389 15487
rect 7423 15484 7435 15487
rect 7852 15484 7880 15512
rect 10612 15496 10640 15592
rect 11054 15580 11060 15632
rect 11112 15580 11118 15632
rect 11974 15580 11980 15632
rect 12032 15620 12038 15632
rect 14461 15623 14519 15629
rect 12032 15592 13952 15620
rect 12032 15580 12038 15592
rect 10778 15512 10784 15564
rect 10836 15552 10842 15564
rect 11072 15552 11100 15580
rect 11333 15555 11391 15561
rect 11333 15552 11345 15555
rect 10836 15524 11345 15552
rect 10836 15512 10842 15524
rect 11333 15521 11345 15524
rect 11379 15521 11391 15555
rect 11333 15515 11391 15521
rect 12529 15555 12587 15561
rect 12529 15521 12541 15555
rect 12575 15552 12587 15555
rect 13262 15552 13268 15564
rect 12575 15524 13268 15552
rect 12575 15521 12587 15524
rect 12529 15515 12587 15521
rect 13262 15512 13268 15524
rect 13320 15512 13326 15564
rect 7423 15456 7880 15484
rect 8297 15487 8355 15493
rect 7423 15453 7435 15456
rect 7377 15447 7435 15453
rect 8297 15453 8309 15487
rect 8343 15484 8355 15487
rect 8478 15484 8484 15496
rect 8343 15456 8484 15484
rect 8343 15453 8355 15456
rect 8297 15447 8355 15453
rect 8478 15444 8484 15456
rect 8536 15444 8542 15496
rect 9398 15484 9404 15496
rect 9359 15456 9404 15484
rect 9398 15444 9404 15456
rect 9456 15444 9462 15496
rect 10413 15487 10471 15493
rect 10413 15453 10425 15487
rect 10459 15484 10471 15487
rect 10594 15484 10600 15496
rect 10459 15456 10600 15484
rect 10459 15453 10471 15456
rect 10413 15447 10471 15453
rect 10594 15444 10600 15456
rect 10652 15444 10658 15496
rect 11149 15487 11207 15493
rect 11149 15453 11161 15487
rect 11195 15484 11207 15487
rect 12161 15487 12219 15493
rect 12161 15484 12173 15487
rect 11195 15456 12173 15484
rect 11195 15453 11207 15456
rect 11149 15447 11207 15453
rect 12161 15453 12173 15456
rect 12207 15484 12219 15487
rect 13170 15484 13176 15496
rect 12207 15456 13176 15484
rect 12207 15453 12219 15456
rect 12161 15447 12219 15453
rect 13170 15444 13176 15456
rect 13228 15484 13234 15496
rect 13814 15484 13820 15496
rect 13228 15456 13820 15484
rect 13228 15444 13234 15456
rect 13814 15444 13820 15456
rect 13872 15444 13878 15496
rect 13924 15484 13952 15592
rect 14461 15589 14473 15623
rect 14507 15620 14519 15623
rect 14918 15620 14924 15632
rect 14507 15592 14924 15620
rect 14507 15589 14519 15592
rect 14461 15583 14519 15589
rect 14918 15580 14924 15592
rect 14976 15620 14982 15632
rect 15102 15620 15108 15632
rect 14976 15592 15108 15620
rect 14976 15580 14982 15592
rect 15102 15580 15108 15592
rect 15160 15580 15166 15632
rect 16025 15623 16083 15629
rect 16025 15589 16037 15623
rect 16071 15620 16083 15623
rect 18138 15620 18144 15632
rect 16071 15592 17264 15620
rect 18099 15592 18144 15620
rect 16071 15589 16083 15592
rect 16025 15583 16083 15589
rect 15473 15555 15531 15561
rect 15473 15521 15485 15555
rect 15519 15552 15531 15555
rect 16114 15552 16120 15564
rect 15519 15524 16120 15552
rect 15519 15521 15531 15524
rect 15473 15515 15531 15521
rect 16114 15512 16120 15524
rect 16172 15552 16178 15564
rect 16209 15555 16267 15561
rect 16209 15552 16221 15555
rect 16172 15524 16221 15552
rect 16172 15512 16178 15524
rect 16209 15521 16221 15524
rect 16255 15521 16267 15555
rect 17126 15552 17132 15564
rect 17087 15524 17132 15552
rect 16209 15515 16267 15521
rect 17126 15512 17132 15524
rect 17184 15512 17190 15564
rect 17236 15561 17264 15592
rect 18138 15580 18144 15592
rect 18196 15580 18202 15632
rect 18506 15580 18512 15632
rect 18564 15620 18570 15632
rect 18601 15623 18659 15629
rect 18601 15620 18613 15623
rect 18564 15592 18613 15620
rect 18564 15580 18570 15592
rect 18601 15589 18613 15592
rect 18647 15589 18659 15623
rect 19518 15620 19524 15632
rect 19479 15592 19524 15620
rect 18601 15583 18659 15589
rect 19518 15580 19524 15592
rect 19576 15580 19582 15632
rect 19889 15623 19947 15629
rect 19889 15589 19901 15623
rect 19935 15620 19947 15623
rect 20622 15620 20628 15632
rect 19935 15592 20628 15620
rect 19935 15589 19947 15592
rect 19889 15583 19947 15589
rect 20622 15580 20628 15592
rect 20680 15580 20686 15632
rect 17221 15555 17279 15561
rect 17221 15521 17233 15555
rect 17267 15521 17279 15555
rect 17221 15515 17279 15521
rect 19306 15524 20668 15552
rect 16298 15484 16304 15496
rect 13924 15456 16304 15484
rect 16298 15444 16304 15456
rect 16356 15444 16362 15496
rect 16393 15487 16451 15493
rect 16393 15453 16405 15487
rect 16439 15484 16451 15487
rect 16942 15484 16948 15496
rect 16439 15456 16948 15484
rect 16439 15453 16451 15456
rect 16393 15447 16451 15453
rect 16942 15444 16948 15456
rect 17000 15444 17006 15496
rect 17957 15487 18015 15493
rect 17957 15453 17969 15487
rect 18003 15484 18015 15487
rect 18506 15484 18512 15496
rect 18003 15456 18512 15484
rect 18003 15453 18015 15456
rect 17957 15447 18015 15453
rect 18506 15444 18512 15456
rect 18564 15444 18570 15496
rect 18598 15444 18604 15496
rect 18656 15484 18662 15496
rect 18969 15487 19027 15493
rect 18969 15484 18981 15487
rect 18656 15456 18981 15484
rect 18656 15444 18662 15456
rect 18969 15453 18981 15456
rect 19015 15484 19027 15487
rect 19306 15484 19334 15524
rect 19702 15484 19708 15496
rect 19015 15456 19334 15484
rect 19663 15456 19708 15484
rect 19015 15453 19027 15456
rect 18969 15447 19027 15453
rect 19702 15444 19708 15456
rect 19760 15444 19766 15496
rect 20257 15487 20315 15493
rect 20257 15453 20269 15487
rect 20303 15453 20315 15487
rect 20530 15484 20536 15496
rect 20491 15456 20536 15484
rect 20257 15447 20315 15453
rect 4764 15388 5580 15416
rect 5997 15419 6055 15425
rect 4764 15376 4770 15388
rect 5997 15385 6009 15419
rect 6043 15416 6055 15419
rect 6362 15416 6368 15428
rect 6043 15388 6368 15416
rect 6043 15385 6055 15388
rect 5997 15379 6055 15385
rect 6362 15376 6368 15388
rect 6420 15376 6426 15428
rect 7285 15419 7343 15425
rect 7285 15385 7297 15419
rect 7331 15416 7343 15419
rect 8021 15419 8079 15425
rect 8021 15416 8033 15419
rect 7331 15388 8033 15416
rect 7331 15385 7343 15388
rect 7285 15379 7343 15385
rect 8021 15385 8033 15388
rect 8067 15416 8079 15419
rect 8067 15388 8340 15416
rect 8067 15385 8079 15388
rect 8021 15379 8079 15385
rect 4525 15351 4583 15357
rect 4525 15317 4537 15351
rect 4571 15317 4583 15351
rect 4525 15311 4583 15317
rect 4893 15351 4951 15357
rect 4893 15317 4905 15351
rect 4939 15348 4951 15351
rect 5902 15348 5908 15360
rect 4939 15320 5908 15348
rect 4939 15317 4951 15320
rect 4893 15311 4951 15317
rect 5902 15308 5908 15320
rect 5960 15348 5966 15360
rect 6457 15351 6515 15357
rect 6457 15348 6469 15351
rect 5960 15320 6469 15348
rect 5960 15308 5966 15320
rect 6457 15317 6469 15320
rect 6503 15348 6515 15351
rect 6638 15348 6644 15360
rect 6503 15320 6644 15348
rect 6503 15317 6515 15320
rect 6457 15311 6515 15317
rect 6638 15308 6644 15320
rect 6696 15308 6702 15360
rect 7374 15308 7380 15360
rect 7432 15348 7438 15360
rect 8113 15351 8171 15357
rect 8113 15348 8125 15351
rect 7432 15320 8125 15348
rect 7432 15308 7438 15320
rect 8113 15317 8125 15320
rect 8159 15348 8171 15351
rect 8202 15348 8208 15360
rect 8159 15320 8208 15348
rect 8159 15317 8171 15320
rect 8113 15311 8171 15317
rect 8202 15308 8208 15320
rect 8260 15308 8266 15360
rect 8312 15348 8340 15388
rect 8386 15376 8392 15428
rect 8444 15416 8450 15428
rect 9766 15416 9772 15428
rect 8444 15388 9772 15416
rect 8444 15376 8450 15388
rect 9766 15376 9772 15388
rect 9824 15376 9830 15428
rect 10321 15419 10379 15425
rect 10321 15385 10333 15419
rect 10367 15416 10379 15419
rect 11609 15419 11667 15425
rect 11609 15416 11621 15419
rect 10367 15388 11621 15416
rect 10367 15385 10379 15388
rect 10321 15379 10379 15385
rect 11609 15385 11621 15388
rect 11655 15385 11667 15419
rect 11609 15379 11667 15385
rect 12621 15419 12679 15425
rect 12621 15385 12633 15419
rect 12667 15416 12679 15419
rect 13906 15416 13912 15428
rect 12667 15388 13912 15416
rect 12667 15385 12679 15388
rect 12621 15379 12679 15385
rect 13906 15376 13912 15388
rect 13964 15376 13970 15428
rect 17313 15419 17371 15425
rect 17313 15416 17325 15419
rect 16868 15388 17325 15416
rect 8570 15348 8576 15360
rect 8312 15320 8576 15348
rect 8570 15308 8576 15320
rect 8628 15308 8634 15360
rect 9490 15308 9496 15360
rect 9548 15348 9554 15360
rect 9861 15351 9919 15357
rect 9548 15320 9593 15348
rect 9548 15308 9554 15320
rect 9861 15317 9873 15351
rect 9907 15348 9919 15351
rect 10962 15348 10968 15360
rect 9907 15320 10968 15348
rect 9907 15317 9919 15320
rect 9861 15311 9919 15317
rect 10962 15308 10968 15320
rect 11020 15308 11026 15360
rect 11241 15351 11299 15357
rect 11241 15317 11253 15351
rect 11287 15348 11299 15351
rect 11974 15348 11980 15360
rect 11287 15320 11980 15348
rect 11287 15317 11299 15320
rect 11241 15311 11299 15317
rect 11974 15308 11980 15320
rect 12032 15308 12038 15360
rect 12710 15308 12716 15360
rect 12768 15348 12774 15360
rect 13354 15348 13360 15360
rect 12768 15320 12813 15348
rect 13315 15320 13360 15348
rect 12768 15308 12774 15320
rect 13354 15308 13360 15320
rect 13412 15308 13418 15360
rect 13722 15308 13728 15360
rect 13780 15348 13786 15360
rect 14553 15351 14611 15357
rect 14553 15348 14565 15351
rect 13780 15320 14565 15348
rect 13780 15308 13786 15320
rect 14553 15317 14565 15320
rect 14599 15348 14611 15351
rect 15010 15348 15016 15360
rect 14599 15320 15016 15348
rect 14599 15317 14611 15320
rect 14553 15311 14611 15317
rect 15010 15308 15016 15320
rect 15068 15308 15074 15360
rect 15562 15348 15568 15360
rect 15523 15320 15568 15348
rect 15562 15308 15568 15320
rect 15620 15308 15626 15360
rect 15654 15308 15660 15360
rect 15712 15348 15718 15360
rect 15712 15320 15757 15348
rect 15712 15308 15718 15320
rect 16390 15308 16396 15360
rect 16448 15348 16454 15360
rect 16868 15357 16896 15388
rect 17313 15385 17325 15388
rect 17359 15385 17371 15419
rect 20272 15416 20300 15447
rect 20530 15444 20536 15456
rect 20588 15444 20594 15496
rect 20640 15484 20668 15524
rect 20714 15512 20720 15564
rect 20772 15552 20778 15564
rect 21085 15555 21143 15561
rect 21085 15552 21097 15555
rect 20772 15524 21097 15552
rect 20772 15512 20778 15524
rect 21085 15521 21097 15524
rect 21131 15521 21143 15555
rect 21085 15515 21143 15521
rect 20809 15487 20867 15493
rect 20809 15484 20821 15487
rect 20640 15456 20821 15484
rect 20809 15453 20821 15456
rect 20855 15453 20867 15487
rect 20809 15447 20867 15453
rect 20990 15444 20996 15496
rect 21048 15484 21054 15496
rect 21269 15487 21327 15493
rect 21269 15484 21281 15487
rect 21048 15456 21281 15484
rect 21048 15444 21054 15456
rect 21269 15453 21281 15456
rect 21315 15453 21327 15487
rect 21269 15447 21327 15453
rect 17313 15379 17371 15385
rect 17696 15388 20300 15416
rect 17696 15357 17724 15388
rect 16485 15351 16543 15357
rect 16485 15348 16497 15351
rect 16448 15320 16497 15348
rect 16448 15308 16454 15320
rect 16485 15317 16497 15320
rect 16531 15317 16543 15351
rect 16485 15311 16543 15317
rect 16853 15351 16911 15357
rect 16853 15317 16865 15351
rect 16899 15317 16911 15351
rect 16853 15311 16911 15317
rect 17681 15351 17739 15357
rect 17681 15317 17693 15351
rect 17727 15317 17739 15351
rect 17681 15311 17739 15317
rect 17770 15308 17776 15360
rect 17828 15348 17834 15360
rect 18322 15348 18328 15360
rect 17828 15320 17873 15348
rect 18283 15320 18328 15348
rect 17828 15308 17834 15320
rect 18322 15308 18328 15320
rect 18380 15308 18386 15360
rect 18509 15351 18567 15357
rect 18509 15317 18521 15351
rect 18555 15348 18567 15351
rect 18690 15348 18696 15360
rect 18555 15320 18696 15348
rect 18555 15317 18567 15320
rect 18509 15311 18567 15317
rect 18690 15308 18696 15320
rect 18748 15308 18754 15360
rect 18874 15348 18880 15360
rect 18835 15320 18880 15348
rect 18874 15308 18880 15320
rect 18932 15308 18938 15360
rect 19337 15351 19395 15357
rect 19337 15317 19349 15351
rect 19383 15348 19395 15351
rect 19610 15348 19616 15360
rect 19383 15320 19616 15348
rect 19383 15317 19395 15320
rect 19337 15311 19395 15317
rect 19610 15308 19616 15320
rect 19668 15308 19674 15360
rect 20162 15348 20168 15360
rect 20123 15320 20168 15348
rect 20162 15308 20168 15320
rect 20220 15308 20226 15360
rect 20717 15351 20775 15357
rect 20717 15317 20729 15351
rect 20763 15348 20775 15351
rect 20806 15348 20812 15360
rect 20763 15320 20812 15348
rect 20763 15317 20775 15320
rect 20717 15311 20775 15317
rect 20806 15308 20812 15320
rect 20864 15308 20870 15360
rect 20990 15348 20996 15360
rect 20951 15320 20996 15348
rect 20990 15308 20996 15320
rect 21048 15308 21054 15360
rect 21450 15348 21456 15360
rect 21411 15320 21456 15348
rect 21450 15308 21456 15320
rect 21508 15308 21514 15360
rect 1104 15258 22056 15280
rect 1104 15206 6148 15258
rect 6200 15206 6212 15258
rect 6264 15206 6276 15258
rect 6328 15206 6340 15258
rect 6392 15206 6404 15258
rect 6456 15206 11346 15258
rect 11398 15206 11410 15258
rect 11462 15206 11474 15258
rect 11526 15206 11538 15258
rect 11590 15206 11602 15258
rect 11654 15206 16544 15258
rect 16596 15206 16608 15258
rect 16660 15206 16672 15258
rect 16724 15206 16736 15258
rect 16788 15206 16800 15258
rect 16852 15206 21742 15258
rect 21794 15206 21806 15258
rect 21858 15206 21870 15258
rect 21922 15206 21934 15258
rect 21986 15206 21998 15258
rect 22050 15206 22056 15258
rect 1104 15184 22056 15206
rect 2406 15104 2412 15156
rect 2464 15144 2470 15156
rect 3973 15147 4031 15153
rect 3973 15144 3985 15147
rect 2464 15116 3985 15144
rect 2464 15104 2470 15116
rect 3973 15113 3985 15116
rect 4019 15113 4031 15147
rect 5261 15147 5319 15153
rect 5261 15144 5273 15147
rect 3973 15107 4031 15113
rect 4080 15116 5273 15144
rect 2958 15036 2964 15088
rect 3016 15076 3022 15088
rect 4080 15076 4108 15116
rect 5261 15113 5273 15116
rect 5307 15113 5319 15147
rect 5261 15107 5319 15113
rect 5350 15104 5356 15156
rect 5408 15144 5414 15156
rect 6086 15144 6092 15156
rect 5408 15116 6092 15144
rect 5408 15104 5414 15116
rect 6086 15104 6092 15116
rect 6144 15104 6150 15156
rect 7558 15104 7564 15156
rect 7616 15144 7622 15156
rect 7837 15147 7895 15153
rect 7837 15144 7849 15147
rect 7616 15116 7849 15144
rect 7616 15104 7622 15116
rect 7837 15113 7849 15116
rect 7883 15113 7895 15147
rect 8386 15144 8392 15156
rect 8347 15116 8392 15144
rect 7837 15107 7895 15113
rect 8386 15104 8392 15116
rect 8444 15144 8450 15156
rect 8941 15147 8999 15153
rect 8444 15116 8892 15144
rect 8444 15104 8450 15116
rect 3016 15048 4108 15076
rect 4433 15079 4491 15085
rect 3016 15036 3022 15048
rect 4433 15045 4445 15079
rect 4479 15076 4491 15079
rect 4982 15076 4988 15088
rect 4479 15048 4988 15076
rect 4479 15045 4491 15048
rect 4433 15039 4491 15045
rect 4982 15036 4988 15048
rect 5040 15036 5046 15088
rect 8665 15079 8723 15085
rect 8665 15076 8677 15079
rect 5552 15048 8677 15076
rect 1670 15008 1676 15020
rect 1631 14980 1676 15008
rect 1670 14968 1676 14980
rect 1728 14968 1734 15020
rect 2041 15011 2099 15017
rect 2041 14977 2053 15011
rect 2087 15008 2099 15011
rect 2317 15011 2375 15017
rect 2087 14980 2176 15008
rect 2087 14977 2099 14980
rect 2041 14971 2099 14977
rect 1854 14872 1860 14884
rect 1815 14844 1860 14872
rect 1854 14832 1860 14844
rect 1912 14832 1918 14884
rect 2148 14881 2176 14980
rect 2317 14977 2329 15011
rect 2363 14977 2375 15011
rect 2498 15008 2504 15020
rect 2459 14980 2504 15008
rect 2317 14971 2375 14977
rect 2332 14940 2360 14971
rect 2498 14968 2504 14980
rect 2556 14968 2562 15020
rect 2768 15011 2826 15017
rect 2768 14977 2780 15011
rect 2814 15008 2826 15011
rect 3326 15008 3332 15020
rect 2814 14980 3332 15008
rect 2814 14977 2826 14980
rect 2768 14971 2826 14977
rect 3326 14968 3332 14980
rect 3384 15008 3390 15020
rect 4338 15008 4344 15020
rect 3384 14980 3740 15008
rect 4299 14980 4344 15008
rect 3384 14968 3390 14980
rect 2406 14940 2412 14952
rect 2332 14912 2412 14940
rect 2406 14900 2412 14912
rect 2464 14900 2470 14952
rect 2133 14875 2191 14881
rect 2133 14841 2145 14875
rect 2179 14841 2191 14875
rect 2133 14835 2191 14841
rect 1486 14804 1492 14816
rect 1447 14776 1492 14804
rect 1486 14764 1492 14776
rect 1544 14764 1550 14816
rect 2682 14764 2688 14816
rect 2740 14804 2746 14816
rect 3418 14804 3424 14816
rect 2740 14776 3424 14804
rect 2740 14764 2746 14776
rect 3418 14764 3424 14776
rect 3476 14764 3482 14816
rect 3712 14804 3740 14980
rect 4338 14968 4344 14980
rect 4396 14968 4402 15020
rect 4890 14968 4896 15020
rect 4948 15008 4954 15020
rect 5077 15011 5135 15017
rect 5077 15008 5089 15011
rect 4948 14980 5089 15008
rect 4948 14968 4954 14980
rect 5077 14977 5089 14980
rect 5123 14977 5135 15011
rect 5077 14971 5135 14977
rect 4525 14943 4583 14949
rect 4525 14909 4537 14943
rect 4571 14909 4583 14943
rect 4525 14903 4583 14909
rect 3878 14872 3884 14884
rect 3839 14844 3884 14872
rect 3878 14832 3884 14844
rect 3936 14872 3942 14884
rect 4540 14872 4568 14903
rect 4798 14900 4804 14952
rect 4856 14940 4862 14952
rect 5552 14940 5580 15048
rect 8665 15045 8677 15048
rect 8711 15045 8723 15079
rect 8864 15076 8892 15116
rect 8941 15113 8953 15147
rect 8987 15144 8999 15147
rect 9214 15144 9220 15156
rect 8987 15116 9220 15144
rect 8987 15113 8999 15116
rect 8941 15107 8999 15113
rect 9214 15104 9220 15116
rect 9272 15104 9278 15156
rect 9950 15104 9956 15156
rect 10008 15144 10014 15156
rect 10229 15147 10287 15153
rect 10229 15144 10241 15147
rect 10008 15116 10241 15144
rect 10008 15104 10014 15116
rect 10229 15113 10241 15116
rect 10275 15113 10287 15147
rect 10229 15107 10287 15113
rect 10778 15104 10784 15156
rect 10836 15144 10842 15156
rect 10836 15116 11100 15144
rect 10836 15104 10842 15116
rect 11072 15088 11100 15116
rect 12250 15104 12256 15156
rect 12308 15144 12314 15156
rect 12713 15147 12771 15153
rect 12713 15144 12725 15147
rect 12308 15116 12725 15144
rect 12308 15104 12314 15116
rect 12713 15113 12725 15116
rect 12759 15144 12771 15147
rect 13078 15144 13084 15156
rect 12759 15116 13084 15144
rect 12759 15113 12771 15116
rect 12713 15107 12771 15113
rect 13078 15104 13084 15116
rect 13136 15104 13142 15156
rect 13354 15104 13360 15156
rect 13412 15144 13418 15156
rect 13449 15147 13507 15153
rect 13449 15144 13461 15147
rect 13412 15116 13461 15144
rect 13412 15104 13418 15116
rect 13449 15113 13461 15116
rect 13495 15113 13507 15147
rect 13906 15144 13912 15156
rect 13867 15116 13912 15144
rect 13449 15107 13507 15113
rect 13906 15104 13912 15116
rect 13964 15104 13970 15156
rect 15746 15144 15752 15156
rect 14108 15116 15752 15144
rect 9861 15079 9919 15085
rect 8864 15048 9260 15076
rect 8665 15039 8723 15045
rect 9232 15020 9260 15048
rect 9861 15045 9873 15079
rect 9907 15076 9919 15079
rect 10870 15076 10876 15088
rect 9907 15048 10876 15076
rect 9907 15045 9919 15048
rect 9861 15039 9919 15045
rect 10870 15036 10876 15048
rect 10928 15036 10934 15088
rect 11054 15036 11060 15088
rect 11112 15036 11118 15088
rect 12069 15079 12127 15085
rect 12069 15045 12081 15079
rect 12115 15076 12127 15079
rect 13541 15079 13599 15085
rect 13541 15076 13553 15079
rect 12115 15048 13553 15076
rect 12115 15045 12127 15048
rect 12069 15039 12127 15045
rect 13541 15045 13553 15048
rect 13587 15076 13599 15079
rect 14108 15076 14136 15116
rect 15746 15104 15752 15116
rect 15804 15104 15810 15156
rect 16114 15144 16120 15156
rect 16075 15116 16120 15144
rect 16114 15104 16120 15116
rect 16172 15104 16178 15156
rect 20162 15104 20168 15156
rect 20220 15144 20226 15156
rect 20349 15147 20407 15153
rect 20349 15144 20361 15147
rect 20220 15116 20361 15144
rect 20220 15104 20226 15116
rect 20349 15113 20361 15116
rect 20395 15113 20407 15147
rect 20349 15107 20407 15113
rect 13587 15048 14136 15076
rect 13587 15045 13599 15048
rect 13541 15039 13599 15045
rect 14182 15036 14188 15088
rect 14240 15076 14246 15088
rect 14369 15079 14427 15085
rect 14369 15076 14381 15079
rect 14240 15048 14381 15076
rect 14240 15036 14246 15048
rect 14369 15045 14381 15048
rect 14415 15045 14427 15079
rect 18506 15076 18512 15088
rect 14369 15039 14427 15045
rect 17052 15048 18512 15076
rect 5629 15011 5687 15017
rect 5629 14977 5641 15011
rect 5675 15008 5687 15011
rect 5902 15008 5908 15020
rect 5675 14980 5908 15008
rect 5675 14977 5687 14980
rect 5629 14971 5687 14977
rect 5902 14968 5908 14980
rect 5960 14968 5966 15020
rect 5994 14968 6000 15020
rect 6052 15008 6058 15020
rect 6549 15011 6607 15017
rect 6549 15008 6561 15011
rect 6052 14980 6561 15008
rect 6052 14968 6058 14980
rect 6549 14977 6561 14980
rect 6595 14977 6607 15011
rect 6549 14971 6607 14977
rect 7377 15011 7435 15017
rect 7377 14977 7389 15011
rect 7423 14977 7435 15011
rect 7377 14971 7435 14977
rect 4856 14912 5580 14940
rect 5721 14943 5779 14949
rect 4856 14900 4862 14912
rect 5721 14909 5733 14943
rect 5767 14909 5779 14943
rect 5721 14903 5779 14909
rect 5813 14943 5871 14949
rect 5813 14909 5825 14943
rect 5859 14940 5871 14943
rect 7006 14940 7012 14952
rect 5859 14912 7012 14940
rect 5859 14909 5871 14912
rect 5813 14903 5871 14909
rect 3936 14844 4568 14872
rect 5736 14872 5764 14903
rect 7006 14900 7012 14912
rect 7064 14940 7070 14952
rect 7392 14940 7420 14971
rect 7650 14968 7656 15020
rect 7708 15008 7714 15020
rect 7745 15011 7803 15017
rect 7745 15008 7757 15011
rect 7708 14980 7757 15008
rect 7708 14968 7714 14980
rect 7745 14977 7757 14980
rect 7791 14977 7803 15011
rect 7745 14971 7803 14977
rect 8021 15011 8079 15017
rect 8021 14977 8033 15011
rect 8067 15008 8079 15011
rect 8294 15008 8300 15020
rect 8067 14980 8300 15008
rect 8067 14977 8079 14980
rect 8021 14971 8079 14977
rect 7064 14912 7420 14940
rect 7064 14900 7070 14912
rect 5994 14872 6000 14884
rect 5736 14844 6000 14872
rect 3936 14832 3942 14844
rect 5994 14832 6000 14844
rect 6052 14832 6058 14884
rect 6822 14872 6828 14884
rect 6380 14844 6828 14872
rect 6380 14816 6408 14844
rect 6822 14832 6828 14844
rect 6880 14832 6886 14884
rect 7760 14872 7788 14971
rect 8294 14968 8300 14980
rect 8352 14968 8358 15020
rect 9122 15008 9128 15020
rect 9083 14980 9128 15008
rect 9122 14968 9128 14980
rect 9180 14968 9186 15020
rect 9214 14968 9220 15020
rect 9272 14968 9278 15020
rect 9401 15011 9459 15017
rect 9401 14977 9413 15011
rect 9447 15008 9459 15011
rect 9447 14980 9812 15008
rect 9447 14977 9459 14980
rect 9401 14971 9459 14977
rect 9674 14940 9680 14952
rect 9635 14912 9680 14940
rect 9674 14900 9680 14912
rect 9732 14900 9738 14952
rect 9784 14949 9812 14980
rect 10594 14968 10600 15020
rect 10652 15008 10658 15020
rect 10689 15011 10747 15017
rect 10689 15008 10701 15011
rect 10652 14980 10701 15008
rect 10652 14968 10658 14980
rect 10689 14977 10701 14980
rect 10735 15008 10747 15011
rect 11149 15011 11207 15017
rect 11149 15008 11161 15011
rect 10735 14980 11161 15008
rect 10735 14977 10747 14980
rect 10689 14971 10747 14977
rect 11149 14977 11161 14980
rect 11195 14977 11207 15011
rect 11149 14971 11207 14977
rect 11977 15011 12035 15017
rect 11977 14977 11989 15011
rect 12023 15008 12035 15011
rect 12621 15011 12679 15017
rect 12621 15008 12633 15011
rect 12023 14980 12633 15008
rect 12023 14977 12035 14980
rect 11977 14971 12035 14977
rect 12621 14977 12633 14980
rect 12667 15008 12679 15011
rect 13354 15008 13360 15020
rect 12667 14980 13360 15008
rect 12667 14977 12679 14980
rect 12621 14971 12679 14977
rect 13354 14968 13360 14980
rect 13412 14968 13418 15020
rect 14274 15008 14280 15020
rect 13464 14980 13676 15008
rect 14235 14980 14280 15008
rect 9769 14943 9827 14949
rect 9769 14909 9781 14943
rect 9815 14940 9827 14943
rect 10410 14940 10416 14952
rect 9815 14912 10416 14940
rect 9815 14909 9827 14912
rect 9769 14903 9827 14909
rect 10410 14900 10416 14912
rect 10468 14900 10474 14952
rect 10781 14943 10839 14949
rect 10781 14940 10793 14943
rect 10520 14912 10793 14940
rect 8205 14875 8263 14881
rect 8205 14872 8217 14875
rect 6932 14844 7696 14872
rect 7760 14844 8217 14872
rect 4614 14804 4620 14816
rect 3712 14776 4620 14804
rect 4614 14764 4620 14776
rect 4672 14804 4678 14816
rect 4985 14807 5043 14813
rect 4985 14804 4997 14807
rect 4672 14776 4997 14804
rect 4672 14764 4678 14776
rect 4985 14773 4997 14776
rect 5031 14773 5043 14807
rect 6362 14804 6368 14816
rect 6323 14776 6368 14804
rect 4985 14767 5043 14773
rect 6362 14764 6368 14776
rect 6420 14764 6426 14816
rect 6638 14764 6644 14816
rect 6696 14804 6702 14816
rect 6932 14804 6960 14844
rect 7558 14804 7564 14816
rect 6696 14776 6960 14804
rect 7519 14776 7564 14804
rect 6696 14764 6702 14776
rect 7558 14764 7564 14776
rect 7616 14764 7622 14816
rect 7668 14804 7696 14844
rect 8205 14841 8217 14844
rect 8251 14841 8263 14875
rect 8205 14835 8263 14841
rect 8386 14832 8392 14884
rect 8444 14872 8450 14884
rect 8481 14875 8539 14881
rect 8481 14872 8493 14875
rect 8444 14844 8493 14872
rect 8444 14832 8450 14844
rect 8481 14841 8493 14844
rect 8527 14872 8539 14875
rect 9030 14872 9036 14884
rect 8527 14844 9036 14872
rect 8527 14841 8539 14844
rect 8481 14835 8539 14841
rect 9030 14832 9036 14844
rect 9088 14832 9094 14884
rect 9490 14832 9496 14884
rect 9548 14872 9554 14884
rect 10321 14875 10379 14881
rect 10321 14872 10333 14875
rect 9548 14844 10333 14872
rect 9548 14832 9554 14844
rect 10321 14841 10333 14844
rect 10367 14841 10379 14875
rect 10321 14835 10379 14841
rect 9122 14804 9128 14816
rect 7668 14776 9128 14804
rect 9122 14764 9128 14776
rect 9180 14764 9186 14816
rect 9398 14764 9404 14816
rect 9456 14804 9462 14816
rect 10520 14804 10548 14912
rect 10781 14909 10793 14912
rect 10827 14909 10839 14943
rect 10781 14903 10839 14909
rect 10965 14943 11023 14949
rect 10965 14909 10977 14943
rect 11011 14940 11023 14943
rect 11054 14940 11060 14952
rect 11011 14912 11060 14940
rect 11011 14909 11023 14912
rect 10965 14903 11023 14909
rect 10796 14872 10824 14903
rect 11054 14900 11060 14912
rect 11112 14900 11118 14952
rect 11793 14943 11851 14949
rect 11793 14909 11805 14943
rect 11839 14940 11851 14943
rect 12250 14940 12256 14952
rect 11839 14912 12256 14940
rect 11839 14909 11851 14912
rect 11793 14903 11851 14909
rect 12250 14900 12256 14912
rect 12308 14900 12314 14952
rect 12802 14900 12808 14952
rect 12860 14940 12866 14952
rect 13464 14940 13492 14980
rect 13648 14949 13676 14980
rect 14274 14968 14280 14980
rect 14332 14968 14338 15020
rect 14826 14968 14832 15020
rect 14884 15008 14890 15020
rect 17052 15017 17080 15048
rect 18506 15036 18512 15048
rect 18564 15036 18570 15088
rect 19518 15036 19524 15088
rect 19576 15076 19582 15088
rect 20257 15079 20315 15085
rect 20257 15076 20269 15079
rect 19576 15048 20269 15076
rect 19576 15036 19582 15048
rect 20257 15045 20269 15048
rect 20303 15045 20315 15079
rect 20257 15039 20315 15045
rect 14993 15011 15051 15017
rect 14993 15008 15005 15011
rect 14884 14980 15005 15008
rect 14884 14968 14890 14980
rect 14993 14977 15005 14980
rect 15039 14977 15051 15011
rect 14993 14971 15051 14977
rect 17037 15011 17095 15017
rect 17037 14977 17049 15011
rect 17083 14977 17095 15011
rect 17037 14971 17095 14977
rect 17126 14968 17132 15020
rect 17184 15008 17190 15020
rect 17293 15011 17351 15017
rect 17293 15008 17305 15011
rect 17184 14980 17305 15008
rect 17184 14968 17190 14980
rect 17293 14977 17305 14980
rect 17339 14977 17351 15011
rect 17293 14971 17351 14977
rect 18322 14968 18328 15020
rect 18380 15008 18386 15020
rect 18765 15011 18823 15017
rect 18765 15008 18777 15011
rect 18380 14980 18777 15008
rect 18380 14968 18386 14980
rect 18765 14977 18777 14980
rect 18811 14977 18823 15011
rect 18765 14971 18823 14977
rect 19058 14968 19064 15020
rect 19116 15008 19122 15020
rect 19116 14980 20208 15008
rect 19116 14968 19122 14980
rect 12860 14912 13492 14940
rect 13633 14943 13691 14949
rect 12860 14900 12866 14912
rect 13633 14909 13645 14943
rect 13679 14909 13691 14943
rect 14461 14943 14519 14949
rect 14461 14940 14473 14943
rect 13633 14903 13691 14909
rect 13731 14912 14473 14940
rect 11517 14875 11575 14881
rect 11517 14872 11529 14875
rect 10796 14844 11529 14872
rect 11517 14841 11529 14844
rect 11563 14841 11575 14875
rect 11517 14835 11575 14841
rect 12618 14832 12624 14884
rect 12676 14872 12682 14884
rect 13731 14872 13759 14912
rect 14461 14909 14473 14912
rect 14507 14909 14519 14943
rect 14461 14903 14519 14909
rect 14737 14943 14795 14949
rect 14737 14909 14749 14943
rect 14783 14909 14795 14943
rect 16850 14940 16856 14952
rect 16811 14912 16856 14940
rect 14737 14903 14795 14909
rect 12676 14844 13759 14872
rect 12676 14832 12682 14844
rect 9456 14776 10548 14804
rect 9456 14764 9462 14776
rect 12250 14764 12256 14816
rect 12308 14804 12314 14816
rect 12308 14776 12353 14804
rect 12308 14764 12314 14776
rect 12526 14764 12532 14816
rect 12584 14804 12590 14816
rect 13081 14807 13139 14813
rect 13081 14804 13093 14807
rect 12584 14776 13093 14804
rect 12584 14764 12590 14776
rect 13081 14773 13093 14776
rect 13127 14773 13139 14807
rect 13081 14767 13139 14773
rect 13814 14764 13820 14816
rect 13872 14804 13878 14816
rect 14458 14804 14464 14816
rect 13872 14776 14464 14804
rect 13872 14764 13878 14776
rect 14458 14764 14464 14776
rect 14516 14804 14522 14816
rect 14752 14804 14780 14903
rect 16850 14900 16856 14912
rect 16908 14900 16914 14952
rect 18506 14940 18512 14952
rect 18467 14912 18512 14940
rect 18506 14900 18512 14912
rect 18564 14900 18570 14952
rect 20073 14943 20131 14949
rect 20073 14940 20085 14943
rect 19904 14912 20085 14940
rect 15746 14804 15752 14816
rect 14516 14776 15752 14804
rect 14516 14764 14522 14776
rect 15746 14764 15752 14776
rect 15804 14804 15810 14816
rect 17770 14804 17776 14816
rect 15804 14776 17776 14804
rect 15804 14764 15810 14776
rect 17770 14764 17776 14776
rect 17828 14764 17834 14816
rect 18322 14764 18328 14816
rect 18380 14804 18386 14816
rect 18417 14807 18475 14813
rect 18417 14804 18429 14807
rect 18380 14776 18429 14804
rect 18380 14764 18386 14776
rect 18417 14773 18429 14776
rect 18463 14773 18475 14807
rect 18417 14767 18475 14773
rect 19518 14764 19524 14816
rect 19576 14804 19582 14816
rect 19904 14813 19932 14912
rect 20073 14909 20085 14912
rect 20119 14909 20131 14943
rect 20180 14940 20208 14980
rect 20806 14968 20812 15020
rect 20864 15008 20870 15020
rect 20901 15011 20959 15017
rect 20901 15008 20913 15011
rect 20864 14980 20913 15008
rect 20864 14968 20870 14980
rect 20901 14977 20913 14980
rect 20947 14977 20959 15011
rect 20901 14971 20959 14977
rect 20990 14968 20996 15020
rect 21048 15008 21054 15020
rect 21269 15011 21327 15017
rect 21269 15008 21281 15011
rect 21048 14980 21281 15008
rect 21048 14968 21054 14980
rect 21269 14977 21281 14980
rect 21315 14977 21327 15011
rect 21269 14971 21327 14977
rect 21358 14940 21364 14952
rect 20180 14912 21364 14940
rect 20073 14903 20131 14909
rect 21358 14900 21364 14912
rect 21416 14900 21422 14952
rect 21082 14872 21088 14884
rect 21043 14844 21088 14872
rect 21082 14832 21088 14844
rect 21140 14832 21146 14884
rect 19889 14807 19947 14813
rect 19889 14804 19901 14807
rect 19576 14776 19901 14804
rect 19576 14764 19582 14776
rect 19889 14773 19901 14776
rect 19935 14773 19947 14807
rect 19889 14767 19947 14773
rect 20438 14764 20444 14816
rect 20496 14804 20502 14816
rect 20717 14807 20775 14813
rect 20717 14804 20729 14807
rect 20496 14776 20729 14804
rect 20496 14764 20502 14776
rect 20717 14773 20729 14776
rect 20763 14773 20775 14807
rect 21450 14804 21456 14816
rect 21411 14776 21456 14804
rect 20717 14767 20775 14773
rect 21450 14764 21456 14776
rect 21508 14764 21514 14816
rect 1104 14714 21896 14736
rect 1104 14662 3549 14714
rect 3601 14662 3613 14714
rect 3665 14662 3677 14714
rect 3729 14662 3741 14714
rect 3793 14662 3805 14714
rect 3857 14662 8747 14714
rect 8799 14662 8811 14714
rect 8863 14662 8875 14714
rect 8927 14662 8939 14714
rect 8991 14662 9003 14714
rect 9055 14662 13945 14714
rect 13997 14662 14009 14714
rect 14061 14662 14073 14714
rect 14125 14662 14137 14714
rect 14189 14662 14201 14714
rect 14253 14662 19143 14714
rect 19195 14662 19207 14714
rect 19259 14662 19271 14714
rect 19323 14662 19335 14714
rect 19387 14662 19399 14714
rect 19451 14662 21896 14714
rect 1104 14640 21896 14662
rect 1762 14600 1768 14612
rect 1723 14572 1768 14600
rect 1762 14560 1768 14572
rect 1820 14560 1826 14612
rect 2133 14603 2191 14609
rect 2133 14569 2145 14603
rect 2179 14600 2191 14603
rect 2314 14600 2320 14612
rect 2179 14572 2320 14600
rect 2179 14569 2191 14572
rect 2133 14563 2191 14569
rect 2314 14560 2320 14572
rect 2372 14560 2378 14612
rect 3050 14600 3056 14612
rect 2700 14572 2943 14600
rect 3011 14572 3056 14600
rect 1670 14492 1676 14544
rect 1728 14532 1734 14544
rect 2501 14535 2559 14541
rect 2501 14532 2513 14535
rect 1728 14504 2513 14532
rect 1728 14492 1734 14504
rect 2501 14501 2513 14504
rect 2547 14501 2559 14535
rect 2501 14495 2559 14501
rect 1762 14424 1768 14476
rect 1820 14464 1826 14476
rect 2700 14464 2728 14572
rect 1820 14436 2728 14464
rect 2915 14464 2943 14572
rect 3050 14560 3056 14572
rect 3108 14560 3114 14612
rect 3329 14603 3387 14609
rect 3329 14569 3341 14603
rect 3375 14600 3387 14603
rect 5534 14600 5540 14612
rect 3375 14572 5540 14600
rect 3375 14569 3387 14572
rect 3329 14563 3387 14569
rect 5534 14560 5540 14572
rect 5592 14560 5598 14612
rect 7650 14600 7656 14612
rect 5644 14572 7656 14600
rect 3605 14535 3663 14541
rect 3605 14501 3617 14535
rect 3651 14532 3663 14535
rect 3970 14532 3976 14544
rect 3651 14504 3976 14532
rect 3651 14501 3663 14504
rect 3605 14495 3663 14501
rect 3970 14492 3976 14504
rect 4028 14492 4034 14544
rect 5644 14473 5672 14572
rect 7650 14560 7656 14572
rect 7708 14600 7714 14612
rect 7708 14572 8616 14600
rect 7708 14560 7714 14572
rect 8588 14473 8616 14572
rect 9122 14560 9128 14612
rect 9180 14600 9186 14612
rect 10502 14600 10508 14612
rect 9180 14572 10508 14600
rect 9180 14560 9186 14572
rect 10502 14560 10508 14572
rect 10560 14560 10566 14612
rect 11882 14600 11888 14612
rect 11795 14572 11888 14600
rect 11882 14560 11888 14572
rect 11940 14600 11946 14612
rect 12618 14600 12624 14612
rect 11940 14572 12624 14600
rect 11940 14560 11946 14572
rect 12618 14560 12624 14572
rect 12676 14560 12682 14612
rect 13262 14560 13268 14612
rect 13320 14600 13326 14612
rect 13357 14603 13415 14609
rect 13357 14600 13369 14603
rect 13320 14572 13369 14600
rect 13320 14560 13326 14572
rect 13357 14569 13369 14572
rect 13403 14569 13415 14603
rect 13357 14563 13415 14569
rect 9950 14532 9956 14544
rect 9232 14504 9956 14532
rect 9232 14476 9260 14504
rect 9950 14492 9956 14504
rect 10008 14532 10014 14544
rect 10318 14532 10324 14544
rect 10008 14504 10324 14532
rect 10008 14492 10014 14504
rect 10318 14492 10324 14504
rect 10376 14492 10382 14544
rect 5537 14467 5595 14473
rect 2915 14436 3464 14464
rect 1820 14424 1826 14436
rect 1673 14399 1731 14405
rect 1673 14365 1685 14399
rect 1719 14365 1731 14399
rect 1673 14359 1731 14365
rect 1949 14399 2007 14405
rect 1949 14365 1961 14399
rect 1995 14396 2007 14399
rect 2314 14396 2320 14408
rect 1995 14368 2320 14396
rect 1995 14365 2007 14368
rect 1949 14359 2007 14365
rect 1688 14328 1716 14359
rect 2314 14356 2320 14368
rect 2372 14356 2378 14408
rect 2409 14399 2467 14405
rect 2409 14365 2421 14399
rect 2455 14396 2467 14399
rect 2590 14396 2596 14408
rect 2455 14368 2596 14396
rect 2455 14365 2467 14368
rect 2409 14359 2467 14365
rect 2590 14356 2596 14368
rect 2648 14356 2654 14408
rect 2685 14399 2743 14405
rect 2685 14365 2697 14399
rect 2731 14365 2743 14399
rect 2685 14359 2743 14365
rect 2700 14328 2728 14359
rect 2774 14356 2780 14408
rect 2832 14392 2838 14408
rect 2869 14399 2927 14405
rect 2869 14392 2881 14399
rect 2832 14365 2881 14392
rect 2915 14365 2927 14399
rect 2832 14364 2927 14365
rect 2832 14356 2838 14364
rect 2869 14359 2927 14364
rect 2958 14356 2964 14408
rect 3016 14396 3022 14408
rect 3145 14399 3203 14405
rect 3145 14396 3157 14399
rect 3016 14368 3157 14396
rect 3016 14356 3022 14368
rect 3145 14365 3157 14368
rect 3191 14396 3203 14399
rect 3234 14396 3240 14408
rect 3191 14368 3240 14396
rect 3191 14365 3203 14368
rect 3145 14359 3203 14365
rect 3234 14356 3240 14368
rect 3292 14356 3298 14408
rect 3436 14405 3464 14436
rect 5537 14433 5549 14467
rect 5583 14464 5595 14467
rect 5629 14467 5687 14473
rect 5629 14464 5641 14467
rect 5583 14436 5641 14464
rect 5583 14433 5595 14436
rect 5537 14427 5595 14433
rect 5629 14433 5641 14436
rect 5675 14433 5687 14467
rect 5629 14427 5687 14433
rect 8573 14467 8631 14473
rect 8573 14433 8585 14467
rect 8619 14433 8631 14467
rect 8573 14427 8631 14433
rect 9214 14424 9220 14476
rect 9272 14424 9278 14476
rect 9493 14467 9551 14473
rect 9493 14433 9505 14467
rect 9539 14433 9551 14467
rect 10042 14464 10048 14476
rect 10003 14436 10048 14464
rect 9493 14427 9551 14433
rect 3421 14399 3479 14405
rect 3421 14365 3433 14399
rect 3467 14365 3479 14399
rect 3421 14359 3479 14365
rect 3789 14399 3847 14405
rect 3789 14365 3801 14399
rect 3835 14396 3847 14399
rect 4154 14396 4160 14408
rect 3835 14368 4160 14396
rect 3835 14365 3847 14368
rect 3789 14359 3847 14365
rect 4154 14356 4160 14368
rect 4212 14356 4218 14408
rect 6362 14396 6368 14408
rect 5184 14368 6368 14396
rect 1688 14300 2268 14328
rect 2700 14300 2912 14328
rect 1486 14260 1492 14272
rect 1447 14232 1492 14260
rect 1486 14220 1492 14232
rect 1544 14220 1550 14272
rect 2240 14269 2268 14300
rect 2884 14272 2912 14300
rect 4062 14288 4068 14340
rect 4120 14328 4126 14340
rect 5184 14328 5212 14368
rect 6362 14356 6368 14368
rect 6420 14356 6426 14408
rect 8294 14396 8300 14408
rect 8352 14405 8358 14408
rect 8352 14399 8375 14405
rect 8227 14368 8300 14396
rect 8294 14356 8300 14368
rect 8363 14396 8375 14399
rect 9508 14396 9536 14427
rect 10042 14424 10048 14436
rect 10100 14424 10106 14476
rect 11790 14424 11796 14476
rect 11848 14464 11854 14476
rect 11974 14464 11980 14476
rect 11848 14436 11980 14464
rect 11848 14424 11854 14436
rect 11974 14424 11980 14436
rect 12032 14424 12038 14476
rect 13372 14464 13400 14563
rect 16390 14560 16396 14612
rect 16448 14600 16454 14612
rect 17221 14603 17279 14609
rect 17221 14600 17233 14603
rect 16448 14572 17233 14600
rect 16448 14560 16454 14572
rect 17221 14569 17233 14572
rect 17267 14569 17279 14603
rect 18506 14600 18512 14612
rect 18467 14572 18512 14600
rect 17221 14563 17279 14569
rect 18506 14560 18512 14572
rect 18564 14560 18570 14612
rect 19886 14600 19892 14612
rect 18616 14572 19892 14600
rect 15473 14535 15531 14541
rect 15473 14501 15485 14535
rect 15519 14501 15531 14535
rect 17126 14532 17132 14544
rect 17087 14504 17132 14532
rect 15473 14495 15531 14501
rect 15488 14464 15516 14495
rect 17126 14492 17132 14504
rect 17184 14492 17190 14544
rect 18141 14535 18199 14541
rect 18141 14501 18153 14535
rect 18187 14532 18199 14535
rect 18616 14532 18644 14572
rect 19886 14560 19892 14572
rect 19944 14560 19950 14612
rect 18187 14504 18644 14532
rect 18187 14501 18199 14504
rect 18141 14495 18199 14501
rect 13372 14436 14228 14464
rect 15488 14436 15884 14464
rect 8363 14368 9536 14396
rect 8363 14365 8375 14368
rect 8352 14359 8375 14365
rect 8352 14356 8358 14359
rect 5350 14337 5356 14340
rect 4120 14300 5212 14328
rect 5292 14331 5356 14337
rect 4120 14288 4126 14300
rect 5292 14297 5304 14331
rect 5338 14297 5356 14331
rect 5292 14291 5356 14297
rect 5350 14288 5356 14291
rect 5408 14288 5414 14340
rect 5874 14331 5932 14337
rect 5874 14328 5886 14331
rect 5736 14300 5886 14328
rect 2225 14263 2283 14269
rect 2225 14229 2237 14263
rect 2271 14229 2283 14263
rect 2225 14223 2283 14229
rect 2866 14220 2872 14272
rect 2924 14220 2930 14272
rect 3418 14220 3424 14272
rect 3476 14260 3482 14272
rect 3973 14263 4031 14269
rect 3973 14260 3985 14263
rect 3476 14232 3985 14260
rect 3476 14220 3482 14232
rect 3973 14229 3985 14232
rect 4019 14229 4031 14263
rect 3973 14223 4031 14229
rect 4157 14263 4215 14269
rect 4157 14229 4169 14263
rect 4203 14260 4215 14263
rect 5166 14260 5172 14272
rect 4203 14232 5172 14260
rect 4203 14229 4215 14232
rect 4157 14223 4215 14229
rect 5166 14220 5172 14232
rect 5224 14260 5230 14272
rect 5736 14260 5764 14300
rect 5874 14297 5886 14300
rect 5920 14297 5932 14331
rect 5874 14291 5932 14297
rect 6546 14288 6552 14340
rect 6604 14328 6610 14340
rect 8570 14328 8576 14340
rect 6604 14300 8576 14328
rect 6604 14288 6610 14300
rect 8570 14288 8576 14300
rect 8628 14288 8634 14340
rect 9582 14328 9588 14340
rect 8680 14300 9588 14328
rect 7006 14260 7012 14272
rect 5224 14232 5764 14260
rect 6967 14232 7012 14260
rect 5224 14220 5230 14232
rect 7006 14220 7012 14232
rect 7064 14220 7070 14272
rect 7193 14263 7251 14269
rect 7193 14229 7205 14263
rect 7239 14260 7251 14263
rect 7742 14260 7748 14272
rect 7239 14232 7748 14260
rect 7239 14229 7251 14232
rect 7193 14223 7251 14229
rect 7742 14220 7748 14232
rect 7800 14220 7806 14272
rect 8018 14220 8024 14272
rect 8076 14260 8082 14272
rect 8680 14260 8708 14300
rect 9582 14288 9588 14300
rect 9640 14288 9646 14340
rect 10060 14328 10088 14424
rect 10318 14396 10324 14408
rect 10279 14368 10324 14396
rect 10318 14356 10324 14368
rect 10376 14356 10382 14408
rect 10505 14399 10563 14405
rect 10505 14365 10517 14399
rect 10551 14396 10563 14399
rect 11808 14396 11836 14424
rect 10551 14368 11836 14396
rect 12244 14399 12302 14405
rect 10551 14365 10563 14368
rect 10505 14359 10563 14365
rect 12244 14365 12256 14399
rect 12290 14396 12302 14399
rect 12618 14396 12624 14408
rect 12290 14368 12624 14396
rect 12290 14365 12302 14368
rect 12244 14359 12302 14365
rect 12618 14356 12624 14368
rect 12676 14356 12682 14408
rect 13814 14356 13820 14408
rect 13872 14396 13878 14408
rect 14093 14399 14151 14405
rect 14093 14396 14105 14399
rect 13872 14368 14105 14396
rect 13872 14356 13878 14368
rect 14093 14365 14105 14368
rect 14139 14365 14151 14399
rect 14200 14396 14228 14436
rect 14349 14399 14407 14405
rect 14349 14396 14361 14399
rect 14200 14368 14361 14396
rect 14093 14359 14151 14365
rect 14349 14365 14361 14368
rect 14395 14365 14407 14399
rect 15746 14396 15752 14408
rect 15707 14368 15752 14396
rect 14349 14359 14407 14365
rect 15746 14356 15752 14368
rect 15804 14356 15810 14408
rect 15856 14396 15884 14436
rect 17218 14424 17224 14476
rect 17276 14464 17282 14476
rect 17773 14467 17831 14473
rect 17773 14464 17785 14467
rect 17276 14436 17785 14464
rect 17276 14424 17282 14436
rect 17773 14433 17785 14436
rect 17819 14433 17831 14467
rect 17773 14427 17831 14433
rect 15856 14368 16804 14396
rect 10594 14328 10600 14340
rect 10060 14300 10600 14328
rect 10594 14288 10600 14300
rect 10652 14288 10658 14340
rect 10772 14331 10830 14337
rect 10772 14297 10784 14331
rect 10818 14328 10830 14331
rect 12802 14328 12808 14340
rect 10818 14300 12808 14328
rect 10818 14297 10830 14300
rect 10772 14291 10830 14297
rect 12802 14288 12808 14300
rect 12860 14288 12866 14340
rect 16016 14331 16074 14337
rect 16016 14297 16028 14331
rect 16062 14328 16074 14331
rect 16114 14328 16120 14340
rect 16062 14300 16120 14328
rect 16062 14297 16074 14300
rect 16016 14291 16074 14297
rect 16114 14288 16120 14300
rect 16172 14288 16178 14340
rect 16776 14328 16804 14368
rect 16850 14356 16856 14408
rect 16908 14396 16914 14408
rect 17589 14399 17647 14405
rect 17589 14396 17601 14399
rect 16908 14368 17601 14396
rect 16908 14356 16914 14368
rect 17589 14365 17601 14368
rect 17635 14365 17647 14399
rect 17589 14359 17647 14365
rect 17681 14399 17739 14405
rect 17681 14365 17693 14399
rect 17727 14396 17739 14399
rect 18156 14396 18184 14495
rect 18782 14492 18788 14544
rect 18840 14532 18846 14544
rect 18877 14535 18935 14541
rect 18877 14532 18889 14535
rect 18840 14504 18889 14532
rect 18840 14492 18846 14504
rect 18877 14501 18889 14504
rect 18923 14501 18935 14535
rect 18877 14495 18935 14501
rect 19794 14492 19800 14544
rect 19852 14532 19858 14544
rect 20346 14532 20352 14544
rect 19852 14504 20352 14532
rect 19852 14492 19858 14504
rect 20346 14492 20352 14504
rect 20404 14532 20410 14544
rect 20404 14504 20944 14532
rect 20404 14492 20410 14504
rect 19429 14467 19487 14473
rect 19429 14433 19441 14467
rect 19475 14464 19487 14467
rect 19518 14464 19524 14476
rect 19475 14436 19524 14464
rect 19475 14433 19487 14436
rect 19429 14427 19487 14433
rect 19518 14424 19524 14436
rect 19576 14424 19582 14476
rect 20622 14464 20628 14476
rect 20583 14436 20628 14464
rect 20622 14424 20628 14436
rect 20680 14424 20686 14476
rect 17727 14368 18184 14396
rect 18325 14399 18383 14405
rect 17727 14365 17739 14368
rect 17681 14359 17739 14365
rect 18325 14365 18337 14399
rect 18371 14396 18383 14399
rect 18414 14396 18420 14408
rect 18371 14368 18420 14396
rect 18371 14365 18383 14368
rect 18325 14359 18383 14365
rect 18414 14356 18420 14368
rect 18472 14356 18478 14408
rect 18785 14399 18843 14405
rect 18785 14365 18797 14399
rect 18831 14396 18843 14399
rect 19794 14396 19800 14408
rect 18831 14368 19800 14396
rect 18831 14365 18843 14368
rect 18785 14359 18843 14365
rect 19794 14356 19800 14368
rect 19852 14356 19858 14408
rect 20438 14396 20444 14408
rect 20399 14368 20444 14396
rect 20438 14356 20444 14368
rect 20496 14356 20502 14408
rect 20916 14405 20944 14504
rect 20901 14399 20959 14405
rect 20901 14365 20913 14399
rect 20947 14365 20959 14399
rect 21266 14396 21272 14408
rect 21227 14368 21272 14396
rect 20901 14359 20959 14365
rect 21266 14356 21272 14368
rect 21324 14356 21330 14408
rect 17402 14328 17408 14340
rect 16776 14300 17408 14328
rect 17402 14288 17408 14300
rect 17460 14288 17466 14340
rect 19610 14328 19616 14340
rect 19571 14300 19616 14328
rect 19610 14288 19616 14300
rect 19668 14288 19674 14340
rect 20533 14331 20591 14337
rect 20533 14328 20545 14331
rect 19996 14300 20545 14328
rect 8076 14232 8708 14260
rect 8076 14220 8082 14232
rect 8754 14220 8760 14272
rect 8812 14260 8818 14272
rect 8938 14260 8944 14272
rect 8812 14232 8857 14260
rect 8899 14232 8944 14260
rect 8812 14220 8818 14232
rect 8938 14220 8944 14232
rect 8996 14220 9002 14272
rect 9214 14220 9220 14272
rect 9272 14260 9278 14272
rect 9309 14263 9367 14269
rect 9309 14260 9321 14263
rect 9272 14232 9321 14260
rect 9272 14220 9278 14232
rect 9309 14229 9321 14232
rect 9355 14229 9367 14263
rect 9309 14223 9367 14229
rect 9401 14263 9459 14269
rect 9401 14229 9413 14263
rect 9447 14260 9459 14263
rect 9490 14260 9496 14272
rect 9447 14232 9496 14260
rect 9447 14229 9459 14232
rect 9401 14223 9459 14229
rect 9490 14220 9496 14232
rect 9548 14220 9554 14272
rect 9861 14263 9919 14269
rect 9861 14229 9873 14263
rect 9907 14260 9919 14263
rect 9950 14260 9956 14272
rect 9907 14232 9956 14260
rect 9907 14229 9919 14232
rect 9861 14223 9919 14229
rect 9950 14220 9956 14232
rect 10008 14220 10014 14272
rect 10134 14260 10140 14272
rect 10095 14232 10140 14260
rect 10134 14220 10140 14232
rect 10192 14220 10198 14272
rect 13446 14220 13452 14272
rect 13504 14260 13510 14272
rect 13504 14232 13549 14260
rect 13504 14220 13510 14232
rect 14090 14220 14096 14272
rect 14148 14260 14154 14272
rect 14550 14260 14556 14272
rect 14148 14232 14556 14260
rect 14148 14220 14154 14232
rect 14550 14220 14556 14232
rect 14608 14220 14614 14272
rect 18414 14220 18420 14272
rect 18472 14260 18478 14272
rect 18601 14263 18659 14269
rect 18601 14260 18613 14263
rect 18472 14232 18613 14260
rect 18472 14220 18478 14232
rect 18601 14229 18613 14232
rect 18647 14229 18659 14263
rect 18601 14223 18659 14229
rect 18782 14220 18788 14272
rect 18840 14260 18846 14272
rect 19996 14269 20024 14300
rect 20533 14297 20545 14300
rect 20579 14297 20591 14331
rect 20533 14291 20591 14297
rect 19521 14263 19579 14269
rect 19521 14260 19533 14263
rect 18840 14232 19533 14260
rect 18840 14220 18846 14232
rect 19521 14229 19533 14232
rect 19567 14229 19579 14263
rect 19521 14223 19579 14229
rect 19981 14263 20039 14269
rect 19981 14229 19993 14263
rect 20027 14229 20039 14263
rect 19981 14223 20039 14229
rect 20070 14220 20076 14272
rect 20128 14260 20134 14272
rect 20128 14232 20173 14260
rect 20128 14220 20134 14232
rect 20806 14220 20812 14272
rect 20864 14260 20870 14272
rect 21085 14263 21143 14269
rect 21085 14260 21097 14263
rect 20864 14232 21097 14260
rect 20864 14220 20870 14232
rect 21085 14229 21097 14232
rect 21131 14229 21143 14263
rect 21450 14260 21456 14272
rect 21411 14232 21456 14260
rect 21085 14223 21143 14229
rect 21450 14220 21456 14232
rect 21508 14220 21514 14272
rect 1104 14170 22056 14192
rect 1104 14118 6148 14170
rect 6200 14118 6212 14170
rect 6264 14118 6276 14170
rect 6328 14118 6340 14170
rect 6392 14118 6404 14170
rect 6456 14118 11346 14170
rect 11398 14118 11410 14170
rect 11462 14118 11474 14170
rect 11526 14118 11538 14170
rect 11590 14118 11602 14170
rect 11654 14118 16544 14170
rect 16596 14118 16608 14170
rect 16660 14118 16672 14170
rect 16724 14118 16736 14170
rect 16788 14118 16800 14170
rect 16852 14118 21742 14170
rect 21794 14118 21806 14170
rect 21858 14118 21870 14170
rect 21922 14118 21934 14170
rect 21986 14118 21998 14170
rect 22050 14118 22056 14170
rect 1104 14096 22056 14118
rect 2133 14059 2191 14065
rect 2133 14025 2145 14059
rect 2179 14025 2191 14059
rect 2133 14019 2191 14025
rect 2148 13988 2176 14019
rect 2314 14016 2320 14068
rect 2372 14056 2378 14068
rect 2593 14059 2651 14065
rect 2593 14056 2605 14059
rect 2372 14028 2605 14056
rect 2372 14016 2378 14028
rect 2593 14025 2605 14028
rect 2639 14025 2651 14059
rect 2593 14019 2651 14025
rect 3142 14016 3148 14068
rect 3200 14056 3206 14068
rect 4341 14059 4399 14065
rect 4341 14056 4353 14059
rect 3200 14028 4353 14056
rect 3200 14016 3206 14028
rect 4341 14025 4353 14028
rect 4387 14025 4399 14059
rect 4341 14019 4399 14025
rect 4522 14016 4528 14068
rect 4580 14056 4586 14068
rect 4709 14059 4767 14065
rect 4709 14056 4721 14059
rect 4580 14028 4721 14056
rect 4580 14016 4586 14028
rect 4709 14025 4721 14028
rect 4755 14056 4767 14059
rect 5902 14056 5908 14068
rect 4755 14028 5764 14056
rect 5863 14028 5908 14056
rect 4755 14025 4767 14028
rect 4709 14019 4767 14025
rect 1688 13960 2176 13988
rect 1688 13929 1716 13960
rect 2406 13948 2412 14000
rect 2464 13988 2470 14000
rect 3789 13991 3847 13997
rect 2464 13960 3740 13988
rect 2464 13948 2470 13960
rect 1673 13923 1731 13929
rect 1673 13889 1685 13923
rect 1719 13889 1731 13923
rect 1673 13883 1731 13889
rect 2041 13923 2099 13929
rect 2041 13889 2053 13923
rect 2087 13920 2099 13923
rect 2130 13920 2136 13932
rect 2087 13892 2136 13920
rect 2087 13889 2099 13892
rect 2041 13883 2099 13889
rect 2130 13880 2136 13892
rect 2188 13880 2194 13932
rect 2317 13923 2375 13929
rect 2317 13889 2329 13923
rect 2363 13889 2375 13923
rect 2958 13920 2964 13932
rect 2919 13892 2964 13920
rect 2317 13883 2375 13889
rect 1578 13812 1584 13864
rect 1636 13852 1642 13864
rect 2332 13852 2360 13883
rect 2958 13880 2964 13892
rect 3016 13880 3022 13932
rect 3712 13920 3740 13960
rect 3789 13957 3801 13991
rect 3835 13988 3847 13991
rect 3878 13988 3884 14000
rect 3835 13960 3884 13988
rect 3835 13957 3847 13960
rect 3789 13951 3847 13957
rect 3878 13948 3884 13960
rect 3936 13948 3942 14000
rect 5258 13948 5264 14000
rect 5316 13988 5322 14000
rect 5537 13991 5595 13997
rect 5537 13988 5549 13991
rect 5316 13960 5549 13988
rect 5316 13948 5322 13960
rect 5537 13957 5549 13960
rect 5583 13957 5595 13991
rect 5736 13988 5764 14028
rect 5902 14016 5908 14028
rect 5960 14016 5966 14068
rect 5994 14016 6000 14068
rect 6052 14056 6058 14068
rect 6365 14059 6423 14065
rect 6365 14056 6377 14059
rect 6052 14028 6377 14056
rect 6052 14016 6058 14028
rect 6365 14025 6377 14028
rect 6411 14025 6423 14059
rect 6365 14019 6423 14025
rect 6825 14059 6883 14065
rect 6825 14025 6837 14059
rect 6871 14056 6883 14059
rect 7193 14059 7251 14065
rect 7193 14056 7205 14059
rect 6871 14028 7205 14056
rect 6871 14025 6883 14028
rect 6825 14019 6883 14025
rect 7193 14025 7205 14028
rect 7239 14025 7251 14059
rect 7193 14019 7251 14025
rect 7561 14059 7619 14065
rect 7561 14025 7573 14059
rect 7607 14056 7619 14059
rect 8938 14056 8944 14068
rect 7607 14028 8944 14056
rect 7607 14025 7619 14028
rect 7561 14019 7619 14025
rect 8938 14016 8944 14028
rect 8996 14016 9002 14068
rect 9030 14016 9036 14068
rect 9088 14056 9094 14068
rect 9493 14059 9551 14065
rect 9493 14056 9505 14059
rect 9088 14028 9505 14056
rect 9088 14016 9094 14028
rect 9493 14025 9505 14028
rect 9539 14025 9551 14059
rect 9493 14019 9551 14025
rect 9582 14016 9588 14068
rect 9640 14056 9646 14068
rect 9640 14028 10732 14056
rect 9640 14016 9646 14028
rect 6546 13988 6552 14000
rect 5736 13960 6552 13988
rect 5537 13951 5595 13957
rect 6546 13948 6552 13960
rect 6604 13948 6610 14000
rect 6733 13991 6791 13997
rect 6733 13957 6745 13991
rect 6779 13988 6791 13991
rect 6914 13988 6920 14000
rect 6779 13960 6920 13988
rect 6779 13957 6791 13960
rect 6733 13951 6791 13957
rect 6914 13948 6920 13960
rect 6972 13948 6978 14000
rect 7006 13948 7012 14000
rect 7064 13988 7070 14000
rect 8266 13991 8324 13997
rect 8266 13988 8278 13991
rect 7064 13960 8278 13988
rect 7064 13948 7070 13960
rect 8266 13957 8278 13960
rect 8312 13957 8324 13991
rect 8266 13951 8324 13957
rect 8386 13948 8392 14000
rect 8444 13948 8450 14000
rect 8570 13948 8576 14000
rect 8628 13988 8634 14000
rect 10413 13991 10471 13997
rect 10413 13988 10425 13991
rect 8628 13960 10425 13988
rect 8628 13948 8634 13960
rect 10413 13957 10425 13960
rect 10459 13988 10471 13991
rect 10704 13988 10732 14028
rect 10778 14016 10784 14068
rect 10836 14056 10842 14068
rect 10873 14059 10931 14065
rect 10873 14056 10885 14059
rect 10836 14028 10885 14056
rect 10836 14016 10842 14028
rect 10873 14025 10885 14028
rect 10919 14025 10931 14059
rect 11054 14056 11060 14068
rect 11015 14028 11060 14056
rect 10873 14019 10931 14025
rect 11054 14016 11060 14028
rect 11112 14016 11118 14068
rect 11333 14059 11391 14065
rect 11333 14025 11345 14059
rect 11379 14056 11391 14059
rect 11422 14056 11428 14068
rect 11379 14028 11428 14056
rect 11379 14025 11391 14028
rect 11333 14019 11391 14025
rect 11422 14016 11428 14028
rect 11480 14016 11486 14068
rect 12345 14059 12403 14065
rect 12345 14025 12357 14059
rect 12391 14056 12403 14059
rect 12526 14056 12532 14068
rect 12391 14028 12532 14056
rect 12391 14025 12403 14028
rect 12345 14019 12403 14025
rect 12526 14016 12532 14028
rect 12584 14016 12590 14068
rect 12710 14056 12716 14068
rect 12671 14028 12716 14056
rect 12710 14016 12716 14028
rect 12768 14016 12774 14068
rect 13541 14059 13599 14065
rect 13541 14025 13553 14059
rect 13587 14056 13599 14059
rect 14274 14056 14280 14068
rect 13587 14028 14280 14056
rect 13587 14025 13599 14028
rect 13541 14019 13599 14025
rect 14274 14016 14280 14028
rect 14332 14016 14338 14068
rect 14550 14016 14556 14068
rect 14608 14056 14614 14068
rect 14918 14056 14924 14068
rect 14608 14028 14924 14056
rect 14608 14016 14614 14028
rect 14918 14016 14924 14028
rect 14976 14016 14982 14068
rect 15105 14059 15163 14065
rect 15105 14025 15117 14059
rect 15151 14056 15163 14059
rect 15933 14059 15991 14065
rect 15933 14056 15945 14059
rect 15151 14028 15945 14056
rect 15151 14025 15163 14028
rect 15105 14019 15163 14025
rect 15933 14025 15945 14028
rect 15979 14025 15991 14059
rect 15933 14019 15991 14025
rect 16669 14059 16727 14065
rect 16669 14025 16681 14059
rect 16715 14056 16727 14059
rect 16942 14056 16948 14068
rect 16715 14028 16948 14056
rect 16715 14025 16727 14028
rect 16669 14019 16727 14025
rect 16942 14016 16948 14028
rect 17000 14016 17006 14068
rect 17037 14059 17095 14065
rect 17037 14025 17049 14059
rect 17083 14056 17095 14059
rect 17954 14056 17960 14068
rect 17083 14028 17960 14056
rect 17083 14025 17095 14028
rect 17037 14019 17095 14025
rect 14645 13991 14703 13997
rect 14645 13988 14657 13991
rect 10459 13960 10640 13988
rect 10704 13960 14657 13988
rect 10459 13957 10471 13960
rect 10413 13951 10471 13957
rect 8021 13923 8079 13929
rect 3712 13892 5120 13920
rect 1636 13824 2360 13852
rect 1636 13812 1642 13824
rect 2406 13812 2412 13864
rect 2464 13852 2470 13864
rect 3050 13852 3056 13864
rect 2464 13824 2509 13852
rect 3011 13824 3056 13852
rect 2464 13812 2470 13824
rect 3050 13812 3056 13824
rect 3108 13812 3114 13864
rect 3145 13855 3203 13861
rect 3145 13821 3157 13855
rect 3191 13821 3203 13855
rect 3881 13855 3939 13861
rect 3881 13852 3893 13855
rect 3145 13815 3203 13821
rect 3252 13824 3893 13852
rect 2498 13744 2504 13796
rect 2556 13784 2562 13796
rect 3160 13784 3188 13815
rect 2556 13756 3188 13784
rect 2556 13744 2562 13756
rect 1486 13716 1492 13728
rect 1447 13688 1492 13716
rect 1486 13676 1492 13688
rect 1544 13676 1550 13728
rect 1854 13716 1860 13728
rect 1815 13688 1860 13716
rect 1854 13676 1860 13688
rect 1912 13676 1918 13728
rect 2406 13676 2412 13728
rect 2464 13716 2470 13728
rect 3252 13716 3280 13824
rect 3881 13821 3893 13824
rect 3927 13821 3939 13855
rect 3881 13815 3939 13821
rect 4065 13855 4123 13861
rect 4065 13821 4077 13855
rect 4111 13852 4123 13855
rect 4246 13852 4252 13864
rect 4111 13824 4252 13852
rect 4111 13821 4123 13824
rect 4065 13815 4123 13821
rect 4246 13812 4252 13824
rect 4304 13812 4310 13864
rect 4614 13812 4620 13864
rect 4672 13852 4678 13864
rect 4801 13855 4859 13861
rect 4801 13852 4813 13855
rect 4672 13824 4813 13852
rect 4672 13812 4678 13824
rect 4801 13821 4813 13824
rect 4847 13821 4859 13855
rect 4801 13815 4859 13821
rect 4890 13812 4896 13864
rect 4948 13852 4954 13864
rect 4948 13824 4993 13852
rect 4948 13812 4954 13824
rect 5092 13784 5120 13892
rect 5276 13892 6132 13920
rect 5166 13812 5172 13864
rect 5224 13852 5230 13864
rect 5276 13861 5304 13892
rect 5261 13855 5319 13861
rect 5261 13852 5273 13855
rect 5224 13824 5273 13852
rect 5224 13812 5230 13824
rect 5261 13821 5273 13824
rect 5307 13821 5319 13855
rect 5442 13852 5448 13864
rect 5403 13824 5448 13852
rect 5261 13815 5319 13821
rect 5442 13812 5448 13824
rect 5500 13812 5506 13864
rect 5994 13852 6000 13864
rect 5955 13824 6000 13852
rect 5994 13812 6000 13824
rect 6052 13812 6058 13864
rect 6104 13852 6132 13892
rect 8021 13889 8033 13923
rect 8067 13920 8079 13923
rect 8404 13920 8432 13948
rect 8067 13892 8432 13920
rect 9861 13923 9919 13929
rect 8067 13889 8079 13892
rect 8021 13883 8079 13889
rect 9861 13889 9873 13923
rect 9907 13920 9919 13923
rect 10502 13920 10508 13932
rect 9907 13892 10508 13920
rect 9907 13889 9919 13892
rect 9861 13883 9919 13889
rect 10502 13880 10508 13892
rect 10560 13880 10566 13932
rect 10612 13920 10640 13960
rect 14645 13957 14657 13960
rect 14691 13957 14703 13991
rect 14645 13951 14703 13957
rect 14737 13991 14795 13997
rect 14737 13957 14749 13991
rect 14783 13988 14795 13991
rect 16206 13988 16212 14000
rect 14783 13960 16212 13988
rect 14783 13957 14795 13960
rect 14737 13951 14795 13957
rect 12526 13920 12532 13932
rect 10612 13892 12532 13920
rect 12526 13880 12532 13892
rect 12584 13880 12590 13932
rect 13173 13923 13231 13929
rect 13173 13889 13185 13923
rect 13219 13920 13231 13923
rect 13538 13920 13544 13932
rect 13219 13892 13544 13920
rect 13219 13889 13231 13892
rect 13173 13883 13231 13889
rect 13538 13880 13544 13892
rect 13596 13880 13602 13932
rect 14090 13920 14096 13932
rect 14051 13892 14096 13920
rect 14090 13880 14096 13892
rect 14148 13880 14154 13932
rect 14277 13923 14335 13929
rect 14277 13889 14289 13923
rect 14323 13920 14335 13923
rect 14752 13920 14780 13951
rect 16206 13948 16212 13960
rect 16264 13948 16270 14000
rect 16298 13948 16304 14000
rect 16356 13988 16362 14000
rect 17052 13988 17080 14019
rect 17954 14016 17960 14028
rect 18012 14016 18018 14068
rect 18233 14059 18291 14065
rect 18233 14025 18245 14059
rect 18279 14056 18291 14059
rect 20162 14056 20168 14068
rect 18279 14028 20168 14056
rect 18279 14025 18291 14028
rect 18233 14019 18291 14025
rect 20162 14016 20168 14028
rect 20220 14016 20226 14068
rect 19518 13997 19524 14000
rect 16356 13960 17080 13988
rect 19460 13991 19524 13997
rect 16356 13948 16362 13960
rect 19460 13957 19472 13991
rect 19506 13957 19524 13991
rect 19460 13951 19524 13957
rect 19518 13948 19524 13951
rect 19576 13948 19582 14000
rect 20064 13991 20122 13997
rect 20064 13988 20076 13991
rect 19628 13960 20076 13988
rect 15838 13920 15844 13932
rect 14323 13892 14780 13920
rect 15799 13892 15844 13920
rect 14323 13889 14335 13892
rect 14277 13883 14335 13889
rect 15838 13880 15844 13892
rect 15896 13880 15902 13932
rect 17126 13880 17132 13932
rect 17184 13920 17190 13932
rect 17310 13920 17316 13932
rect 17184 13892 17316 13920
rect 17184 13880 17190 13892
rect 17310 13880 17316 13892
rect 17368 13880 17374 13932
rect 17865 13923 17923 13929
rect 17865 13889 17877 13923
rect 17911 13920 17923 13923
rect 18230 13920 18236 13932
rect 17911 13892 18236 13920
rect 17911 13889 17923 13892
rect 17865 13883 17923 13889
rect 18230 13880 18236 13892
rect 18288 13880 18294 13932
rect 19628 13920 19656 13960
rect 20064 13957 20076 13960
rect 20110 13988 20122 13991
rect 20622 13988 20628 14000
rect 20110 13960 20628 13988
rect 20110 13957 20122 13960
rect 20064 13951 20122 13957
rect 20622 13948 20628 13960
rect 20680 13948 20686 14000
rect 18708 13892 19656 13920
rect 19705 13923 19763 13929
rect 6917 13855 6975 13861
rect 6917 13852 6929 13855
rect 6104 13824 6929 13852
rect 6917 13821 6929 13824
rect 6963 13821 6975 13855
rect 7650 13852 7656 13864
rect 7611 13824 7656 13852
rect 6917 13815 6975 13821
rect 7650 13812 7656 13824
rect 7708 13812 7714 13864
rect 7742 13812 7748 13864
rect 7800 13852 7806 13864
rect 9398 13852 9404 13864
rect 7800 13824 7845 13852
rect 9048 13824 9404 13852
rect 7800 13812 7806 13824
rect 5902 13784 5908 13796
rect 5092 13756 5908 13784
rect 5902 13744 5908 13756
rect 5960 13744 5966 13796
rect 3418 13716 3424 13728
rect 2464 13688 3280 13716
rect 3379 13688 3424 13716
rect 2464 13676 2470 13688
rect 3418 13676 3424 13688
rect 3476 13676 3482 13728
rect 8202 13676 8208 13728
rect 8260 13716 8266 13728
rect 9048 13716 9076 13824
rect 9398 13812 9404 13824
rect 9456 13812 9462 13864
rect 9490 13812 9496 13864
rect 9548 13852 9554 13864
rect 9953 13855 10011 13861
rect 9953 13852 9965 13855
rect 9548 13824 9965 13852
rect 9548 13812 9554 13824
rect 9953 13821 9965 13824
rect 9999 13821 10011 13855
rect 9953 13815 10011 13821
rect 10045 13855 10103 13861
rect 10045 13821 10057 13855
rect 10091 13821 10103 13855
rect 10045 13815 10103 13821
rect 9582 13744 9588 13796
rect 9640 13784 9646 13796
rect 10060 13784 10088 13815
rect 10226 13812 10232 13864
rect 10284 13852 10290 13864
rect 10594 13852 10600 13864
rect 10284 13824 10456 13852
rect 10555 13824 10600 13852
rect 10284 13812 10290 13824
rect 9640 13756 10088 13784
rect 10428 13784 10456 13824
rect 10594 13812 10600 13824
rect 10652 13812 10658 13864
rect 10689 13855 10747 13861
rect 10689 13821 10701 13855
rect 10735 13821 10747 13855
rect 11514 13852 11520 13864
rect 11475 13824 11520 13852
rect 10689 13815 10747 13821
rect 10704 13784 10732 13815
rect 11514 13812 11520 13824
rect 11572 13812 11578 13864
rect 11698 13852 11704 13864
rect 11659 13824 11704 13852
rect 11698 13812 11704 13824
rect 11756 13812 11762 13864
rect 11882 13812 11888 13864
rect 11940 13852 11946 13864
rect 12069 13855 12127 13861
rect 12069 13852 12081 13855
rect 11940 13824 12081 13852
rect 11940 13812 11946 13824
rect 12069 13821 12081 13824
rect 12115 13821 12127 13855
rect 12250 13852 12256 13864
rect 12211 13824 12256 13852
rect 12069 13815 12127 13821
rect 12250 13812 12256 13824
rect 12308 13812 12314 13864
rect 12802 13812 12808 13864
rect 12860 13852 12866 13864
rect 12897 13855 12955 13861
rect 12897 13852 12909 13855
rect 12860 13824 12909 13852
rect 12860 13812 12866 13824
rect 12897 13821 12909 13824
rect 12943 13821 12955 13855
rect 12897 13815 12955 13821
rect 13081 13855 13139 13861
rect 13081 13821 13093 13855
rect 13127 13852 13139 13855
rect 13262 13852 13268 13864
rect 13127 13824 13268 13852
rect 13127 13821 13139 13824
rect 13081 13815 13139 13821
rect 13262 13812 13268 13824
rect 13320 13812 13326 13864
rect 13909 13855 13967 13861
rect 13909 13821 13921 13855
rect 13955 13852 13967 13855
rect 13998 13852 14004 13864
rect 13955 13824 14004 13852
rect 13955 13821 13967 13824
rect 13909 13815 13967 13821
rect 13998 13812 14004 13824
rect 14056 13812 14062 13864
rect 14553 13855 14611 13861
rect 14553 13821 14565 13855
rect 14599 13852 14611 13855
rect 14734 13852 14740 13864
rect 14599 13824 14740 13852
rect 14599 13821 14611 13824
rect 14553 13815 14611 13821
rect 14734 13812 14740 13824
rect 14792 13812 14798 13864
rect 15562 13852 15568 13864
rect 15488 13824 15568 13852
rect 10428 13756 10732 13784
rect 9640 13744 9646 13756
rect 10962 13744 10968 13796
rect 11020 13784 11026 13796
rect 15488 13793 15516 13824
rect 15562 13812 15568 13824
rect 15620 13812 15626 13864
rect 16025 13855 16083 13861
rect 16025 13821 16037 13855
rect 16071 13821 16083 13855
rect 17218 13852 17224 13864
rect 17131 13824 17224 13852
rect 16025 13815 16083 13821
rect 15473 13787 15531 13793
rect 11020 13756 14044 13784
rect 11020 13744 11026 13756
rect 8260 13688 9076 13716
rect 8260 13676 8266 13688
rect 9122 13676 9128 13728
rect 9180 13716 9186 13728
rect 9401 13719 9459 13725
rect 9401 13716 9413 13719
rect 9180 13688 9413 13716
rect 9180 13676 9186 13688
rect 9401 13685 9413 13688
rect 9447 13685 9459 13719
rect 9401 13679 9459 13685
rect 9766 13676 9772 13728
rect 9824 13716 9830 13728
rect 10594 13716 10600 13728
rect 9824 13688 10600 13716
rect 9824 13676 9830 13688
rect 10594 13676 10600 13688
rect 10652 13676 10658 13728
rect 11238 13676 11244 13728
rect 11296 13716 11302 13728
rect 11974 13716 11980 13728
rect 11296 13688 11980 13716
rect 11296 13676 11302 13688
rect 11974 13676 11980 13688
rect 12032 13676 12038 13728
rect 12710 13676 12716 13728
rect 12768 13716 12774 13728
rect 13354 13716 13360 13728
rect 12768 13688 13360 13716
rect 12768 13676 12774 13688
rect 13354 13676 13360 13688
rect 13412 13676 13418 13728
rect 13538 13676 13544 13728
rect 13596 13716 13602 13728
rect 13633 13719 13691 13725
rect 13633 13716 13645 13719
rect 13596 13688 13645 13716
rect 13596 13676 13602 13688
rect 13633 13685 13645 13688
rect 13679 13685 13691 13719
rect 14016 13716 14044 13756
rect 15473 13753 15485 13787
rect 15519 13753 15531 13787
rect 16040 13784 16068 13815
rect 17218 13812 17224 13824
rect 17276 13812 17282 13864
rect 17681 13855 17739 13861
rect 17681 13821 17693 13855
rect 17727 13821 17739 13855
rect 17681 13815 17739 13821
rect 17773 13855 17831 13861
rect 17773 13821 17785 13855
rect 17819 13852 17831 13855
rect 18046 13852 18052 13864
rect 17819 13824 18052 13852
rect 17819 13821 17831 13824
rect 17773 13815 17831 13821
rect 16114 13784 16120 13796
rect 16040 13756 16120 13784
rect 15473 13747 15531 13753
rect 16114 13744 16120 13756
rect 16172 13784 16178 13796
rect 17236 13784 17264 13812
rect 16172 13756 17264 13784
rect 17696 13784 17724 13815
rect 18046 13812 18052 13824
rect 18104 13812 18110 13864
rect 18708 13852 18736 13892
rect 19705 13889 19717 13923
rect 19751 13920 19763 13923
rect 19794 13920 19800 13932
rect 19751 13892 19800 13920
rect 19751 13889 19763 13892
rect 19705 13883 19763 13889
rect 19794 13880 19800 13892
rect 19852 13880 19858 13932
rect 20346 13880 20352 13932
rect 20404 13920 20410 13932
rect 21269 13923 21327 13929
rect 21269 13920 21281 13923
rect 20404 13892 21281 13920
rect 20404 13880 20410 13892
rect 21269 13889 21281 13892
rect 21315 13889 21327 13923
rect 21269 13883 21327 13889
rect 21542 13880 21548 13932
rect 21600 13920 21606 13932
rect 22646 13920 22652 13932
rect 21600 13892 22652 13920
rect 21600 13880 21606 13892
rect 22646 13880 22652 13892
rect 22704 13880 22710 13932
rect 18340 13824 18736 13852
rect 18340 13793 18368 13824
rect 18325 13787 18383 13793
rect 18325 13784 18337 13787
rect 17696 13756 18337 13784
rect 16172 13744 16178 13756
rect 18325 13753 18337 13756
rect 18371 13753 18383 13787
rect 18325 13747 18383 13753
rect 16301 13719 16359 13725
rect 16301 13716 16313 13719
rect 14016 13688 16313 13716
rect 13633 13679 13691 13685
rect 16301 13685 16313 13688
rect 16347 13716 16359 13719
rect 17126 13716 17132 13728
rect 16347 13688 17132 13716
rect 16347 13685 16359 13688
rect 16301 13679 16359 13685
rect 17126 13676 17132 13688
rect 17184 13676 17190 13728
rect 21174 13716 21180 13728
rect 21135 13688 21180 13716
rect 21174 13676 21180 13688
rect 21232 13676 21238 13728
rect 21450 13716 21456 13728
rect 21411 13688 21456 13716
rect 21450 13676 21456 13688
rect 21508 13676 21514 13728
rect 1104 13626 21896 13648
rect 1104 13574 3549 13626
rect 3601 13574 3613 13626
rect 3665 13574 3677 13626
rect 3729 13574 3741 13626
rect 3793 13574 3805 13626
rect 3857 13574 8747 13626
rect 8799 13574 8811 13626
rect 8863 13574 8875 13626
rect 8927 13574 8939 13626
rect 8991 13574 9003 13626
rect 9055 13574 13945 13626
rect 13997 13574 14009 13626
rect 14061 13574 14073 13626
rect 14125 13574 14137 13626
rect 14189 13574 14201 13626
rect 14253 13574 19143 13626
rect 19195 13574 19207 13626
rect 19259 13574 19271 13626
rect 19323 13574 19335 13626
rect 19387 13574 19399 13626
rect 19451 13574 21896 13626
rect 1104 13552 21896 13574
rect 1765 13515 1823 13521
rect 1765 13481 1777 13515
rect 1811 13512 1823 13515
rect 2498 13512 2504 13524
rect 1811 13484 2504 13512
rect 1811 13481 1823 13484
rect 1765 13475 1823 13481
rect 2498 13472 2504 13484
rect 2556 13472 2562 13524
rect 4154 13512 4160 13524
rect 4115 13484 4160 13512
rect 4154 13472 4160 13484
rect 4212 13472 4218 13524
rect 5258 13512 5264 13524
rect 5219 13484 5264 13512
rect 5258 13472 5264 13484
rect 5316 13472 5322 13524
rect 5353 13515 5411 13521
rect 5353 13481 5365 13515
rect 5399 13512 5411 13515
rect 5442 13512 5448 13524
rect 5399 13484 5448 13512
rect 5399 13481 5411 13484
rect 5353 13475 5411 13481
rect 5442 13472 5448 13484
rect 5500 13472 5506 13524
rect 6457 13515 6515 13521
rect 6457 13481 6469 13515
rect 6503 13512 6515 13515
rect 6546 13512 6552 13524
rect 6503 13484 6552 13512
rect 6503 13481 6515 13484
rect 6457 13475 6515 13481
rect 6546 13472 6552 13484
rect 6604 13472 6610 13524
rect 6914 13512 6920 13524
rect 6875 13484 6920 13512
rect 6914 13472 6920 13484
rect 6972 13472 6978 13524
rect 7650 13472 7656 13524
rect 7708 13512 7714 13524
rect 7745 13515 7803 13521
rect 7745 13512 7757 13515
rect 7708 13484 7757 13512
rect 7708 13472 7714 13484
rect 7745 13481 7757 13484
rect 7791 13481 7803 13515
rect 7745 13475 7803 13481
rect 8386 13472 8392 13524
rect 8444 13472 8450 13524
rect 8570 13472 8576 13524
rect 8628 13512 8634 13524
rect 10502 13512 10508 13524
rect 8628 13484 10180 13512
rect 10463 13484 10508 13512
rect 8628 13472 8634 13484
rect 3605 13447 3663 13453
rect 3605 13444 3617 13447
rect 3252 13416 3617 13444
rect 1673 13311 1731 13317
rect 1673 13277 1685 13311
rect 1719 13308 1731 13311
rect 1719 13280 2452 13308
rect 1719 13277 1731 13280
rect 1673 13271 1731 13277
rect 198 13200 204 13252
rect 256 13240 262 13252
rect 1762 13240 1768 13252
rect 256 13212 1768 13240
rect 256 13200 262 13212
rect 1762 13200 1768 13212
rect 1820 13200 1826 13252
rect 1486 13172 1492 13184
rect 1447 13144 1492 13172
rect 1486 13132 1492 13144
rect 1544 13132 1550 13184
rect 2424 13172 2452 13280
rect 2590 13268 2596 13320
rect 2648 13308 2654 13320
rect 3145 13311 3203 13317
rect 3145 13308 3157 13311
rect 2648 13280 3157 13308
rect 2648 13268 2654 13280
rect 3145 13277 3157 13280
rect 3191 13277 3203 13311
rect 3252 13308 3280 13416
rect 3605 13413 3617 13416
rect 3651 13444 3663 13447
rect 4522 13444 4528 13456
rect 3651 13416 4528 13444
rect 3651 13413 3663 13416
rect 3605 13407 3663 13413
rect 4522 13404 4528 13416
rect 4580 13404 4586 13456
rect 5626 13404 5632 13456
rect 5684 13444 5690 13456
rect 6733 13447 6791 13453
rect 6733 13444 6745 13447
rect 5684 13416 6745 13444
rect 5684 13404 5690 13416
rect 6733 13413 6745 13416
rect 6779 13444 6791 13447
rect 7282 13444 7288 13456
rect 6779 13416 7288 13444
rect 6779 13413 6791 13416
rect 6733 13407 6791 13413
rect 7282 13404 7288 13416
rect 7340 13444 7346 13456
rect 7340 13416 8156 13444
rect 7340 13404 7346 13416
rect 3326 13336 3332 13388
rect 3384 13376 3390 13388
rect 3789 13379 3847 13385
rect 3384 13348 3556 13376
rect 3384 13336 3390 13348
rect 3421 13311 3479 13317
rect 3421 13308 3433 13311
rect 3252 13280 3433 13308
rect 3145 13271 3203 13277
rect 3421 13277 3433 13280
rect 3467 13277 3479 13311
rect 3528 13308 3556 13348
rect 3789 13345 3801 13379
rect 3835 13376 3847 13379
rect 3878 13376 3884 13388
rect 3835 13348 3884 13376
rect 3835 13345 3847 13348
rect 3789 13339 3847 13345
rect 3878 13336 3884 13348
rect 3936 13336 3942 13388
rect 4433 13379 4491 13385
rect 4433 13345 4445 13379
rect 4479 13376 4491 13379
rect 4614 13376 4620 13388
rect 4479 13348 4620 13376
rect 4479 13345 4491 13348
rect 4433 13339 4491 13345
rect 4614 13336 4620 13348
rect 4672 13336 4678 13388
rect 4709 13379 4767 13385
rect 4709 13345 4721 13379
rect 4755 13376 4767 13379
rect 5350 13376 5356 13388
rect 4755 13348 5356 13376
rect 4755 13345 4767 13348
rect 4709 13339 4767 13345
rect 5350 13336 5356 13348
rect 5408 13376 5414 13388
rect 5905 13379 5963 13385
rect 5905 13376 5917 13379
rect 5408 13348 5917 13376
rect 5408 13336 5414 13348
rect 5905 13345 5917 13348
rect 5951 13376 5963 13379
rect 7469 13379 7527 13385
rect 7469 13376 7481 13379
rect 5951 13348 7481 13376
rect 5951 13345 5963 13348
rect 5905 13339 5963 13345
rect 7469 13345 7481 13348
rect 7515 13376 7527 13379
rect 7742 13376 7748 13388
rect 7515 13348 7748 13376
rect 7515 13345 7527 13348
rect 7469 13339 7527 13345
rect 7742 13336 7748 13348
rect 7800 13336 7806 13388
rect 4893 13311 4951 13317
rect 3528 13280 4476 13308
rect 3421 13271 3479 13277
rect 2900 13243 2958 13249
rect 2900 13209 2912 13243
rect 2946 13240 2958 13243
rect 3970 13240 3976 13252
rect 2946 13212 3976 13240
rect 2946 13209 2958 13212
rect 2900 13203 2958 13209
rect 3970 13200 3976 13212
rect 4028 13200 4034 13252
rect 3237 13175 3295 13181
rect 3237 13172 3249 13175
rect 2424 13144 3249 13172
rect 3237 13141 3249 13144
rect 3283 13141 3295 13175
rect 4448 13172 4476 13280
rect 4893 13277 4905 13311
rect 4939 13308 4951 13311
rect 5994 13308 6000 13320
rect 4939 13280 6000 13308
rect 4939 13277 4951 13280
rect 4893 13271 4951 13277
rect 5994 13268 6000 13280
rect 6052 13268 6058 13320
rect 6273 13311 6331 13317
rect 6273 13277 6285 13311
rect 6319 13308 6331 13311
rect 6546 13308 6552 13320
rect 6319 13280 6552 13308
rect 6319 13277 6331 13280
rect 6273 13271 6331 13277
rect 4801 13243 4859 13249
rect 4801 13209 4813 13243
rect 4847 13240 4859 13243
rect 5258 13240 5264 13252
rect 4847 13212 5264 13240
rect 4847 13209 4859 13212
rect 4801 13203 4859 13209
rect 5258 13200 5264 13212
rect 5316 13200 5322 13252
rect 5721 13175 5779 13181
rect 5721 13172 5733 13175
rect 4448 13144 5733 13172
rect 3237 13135 3295 13141
rect 5721 13141 5733 13144
rect 5767 13141 5779 13175
rect 5721 13135 5779 13141
rect 5813 13175 5871 13181
rect 5813 13141 5825 13175
rect 5859 13172 5871 13175
rect 6288 13172 6316 13271
rect 6546 13268 6552 13280
rect 6604 13268 6610 13320
rect 8128 13317 8156 13416
rect 8294 13376 8300 13388
rect 8255 13348 8300 13376
rect 8294 13336 8300 13348
rect 8352 13336 8358 13388
rect 8404 13376 8432 13472
rect 10152 13444 10180 13484
rect 10502 13472 10508 13484
rect 10560 13472 10566 13524
rect 11330 13512 11336 13524
rect 11291 13484 11336 13512
rect 11330 13472 11336 13484
rect 11388 13472 11394 13524
rect 11606 13512 11612 13524
rect 11567 13484 11612 13512
rect 11606 13472 11612 13484
rect 11664 13472 11670 13524
rect 11974 13512 11980 13524
rect 11935 13484 11980 13512
rect 11974 13472 11980 13484
rect 12032 13472 12038 13524
rect 13081 13515 13139 13521
rect 13081 13481 13093 13515
rect 13127 13512 13139 13515
rect 13722 13512 13728 13524
rect 13127 13484 13728 13512
rect 13127 13481 13139 13484
rect 13081 13475 13139 13481
rect 13722 13472 13728 13484
rect 13780 13472 13786 13524
rect 13817 13515 13875 13521
rect 13817 13481 13829 13515
rect 13863 13512 13875 13515
rect 14366 13512 14372 13524
rect 13863 13484 14372 13512
rect 13863 13481 13875 13484
rect 13817 13475 13875 13481
rect 14366 13472 14372 13484
rect 14424 13472 14430 13524
rect 14476 13484 15792 13512
rect 12069 13447 12127 13453
rect 12069 13444 12081 13447
rect 10152 13416 12081 13444
rect 12069 13413 12081 13416
rect 12115 13413 12127 13447
rect 14476 13444 14504 13484
rect 12069 13407 12127 13413
rect 12360 13416 14504 13444
rect 15764 13444 15792 13484
rect 15838 13472 15844 13524
rect 15896 13512 15902 13524
rect 16485 13515 16543 13521
rect 16485 13512 16497 13515
rect 15896 13484 16497 13512
rect 15896 13472 15902 13484
rect 16485 13481 16497 13484
rect 16531 13481 16543 13515
rect 18230 13512 18236 13524
rect 18191 13484 18236 13512
rect 16485 13475 16543 13481
rect 18230 13472 18236 13484
rect 18288 13472 18294 13524
rect 19702 13512 19708 13524
rect 19663 13484 19708 13512
rect 19702 13472 19708 13484
rect 19760 13472 19766 13524
rect 20809 13515 20867 13521
rect 20809 13481 20821 13515
rect 20855 13512 20867 13515
rect 21266 13512 21272 13524
rect 20855 13484 21272 13512
rect 20855 13481 20867 13484
rect 20809 13475 20867 13481
rect 21266 13472 21272 13484
rect 21324 13472 21330 13524
rect 16298 13444 16304 13456
rect 15764 13416 16059 13444
rect 16259 13416 16304 13444
rect 9033 13379 9091 13385
rect 9033 13376 9045 13379
rect 8404 13348 9045 13376
rect 9033 13345 9045 13348
rect 9079 13345 9091 13379
rect 10502 13376 10508 13388
rect 9033 13339 9091 13345
rect 10060 13348 10508 13376
rect 8113 13311 8171 13317
rect 8113 13277 8125 13311
rect 8159 13277 8171 13311
rect 8113 13271 8171 13277
rect 8938 13268 8944 13320
rect 8996 13308 9002 13320
rect 9122 13308 9128 13320
rect 8996 13280 9128 13308
rect 8996 13268 9002 13280
rect 9122 13268 9128 13280
rect 9180 13308 9186 13320
rect 9289 13311 9347 13317
rect 9289 13308 9301 13311
rect 9180 13280 9301 13308
rect 9180 13268 9186 13280
rect 9289 13277 9301 13280
rect 9335 13308 9347 13311
rect 10060 13308 10088 13348
rect 10502 13336 10508 13348
rect 10560 13376 10566 13388
rect 11057 13379 11115 13385
rect 11057 13376 11069 13379
rect 10560 13348 11069 13376
rect 10560 13336 10566 13348
rect 11057 13345 11069 13348
rect 11103 13345 11115 13379
rect 11057 13339 11115 13345
rect 9335 13280 10088 13308
rect 10965 13311 11023 13317
rect 9335 13277 9347 13280
rect 9289 13271 9347 13277
rect 10965 13277 10977 13311
rect 11011 13308 11023 13311
rect 11606 13308 11612 13320
rect 11011 13280 11612 13308
rect 11011 13277 11023 13280
rect 10965 13271 11023 13277
rect 11606 13268 11612 13280
rect 11664 13268 11670 13320
rect 11793 13311 11851 13317
rect 11793 13277 11805 13311
rect 11839 13308 11851 13311
rect 11882 13308 11888 13320
rect 11839 13280 11888 13308
rect 11839 13277 11851 13280
rect 11793 13271 11851 13277
rect 11882 13268 11888 13280
rect 11940 13268 11946 13320
rect 7300 13212 8524 13240
rect 5859 13144 6316 13172
rect 6641 13175 6699 13181
rect 5859 13141 5871 13144
rect 5813 13135 5871 13141
rect 6641 13141 6653 13175
rect 6687 13172 6699 13175
rect 6822 13172 6828 13184
rect 6687 13144 6828 13172
rect 6687 13141 6699 13144
rect 6641 13135 6699 13141
rect 6822 13132 6828 13144
rect 6880 13172 6886 13184
rect 7300 13181 7328 13212
rect 7285 13175 7343 13181
rect 7285 13172 7297 13175
rect 6880 13144 7297 13172
rect 6880 13132 6886 13144
rect 7285 13141 7297 13144
rect 7331 13141 7343 13175
rect 7285 13135 7343 13141
rect 7377 13175 7435 13181
rect 7377 13141 7389 13175
rect 7423 13172 7435 13175
rect 7834 13172 7840 13184
rect 7423 13144 7840 13172
rect 7423 13141 7435 13144
rect 7377 13135 7435 13141
rect 7834 13132 7840 13144
rect 7892 13132 7898 13184
rect 8018 13132 8024 13184
rect 8076 13172 8082 13184
rect 8205 13175 8263 13181
rect 8205 13172 8217 13175
rect 8076 13144 8217 13172
rect 8076 13132 8082 13144
rect 8205 13141 8217 13144
rect 8251 13141 8263 13175
rect 8496 13172 8524 13212
rect 8570 13200 8576 13252
rect 8628 13240 8634 13252
rect 12360 13240 12388 13416
rect 12618 13376 12624 13388
rect 12579 13348 12624 13376
rect 12618 13336 12624 13348
rect 12676 13336 12682 13388
rect 14458 13376 14464 13388
rect 14419 13348 14464 13376
rect 14458 13336 14464 13348
rect 14516 13336 14522 13388
rect 13078 13268 13084 13320
rect 13136 13308 13142 13320
rect 14734 13317 14740 13320
rect 14728 13308 14740 13317
rect 13136 13280 14320 13308
rect 14647 13280 14740 13308
rect 13136 13268 13142 13280
rect 8628 13212 12388 13240
rect 8628 13200 8634 13212
rect 12434 13200 12440 13252
rect 12492 13240 12498 13252
rect 12618 13240 12624 13252
rect 12492 13212 12624 13240
rect 12492 13200 12498 13212
rect 12618 13200 12624 13212
rect 12676 13200 12682 13252
rect 13265 13243 13323 13249
rect 13265 13209 13277 13243
rect 13311 13240 13323 13243
rect 13630 13240 13636 13252
rect 13311 13212 13636 13240
rect 13311 13209 13323 13212
rect 13265 13203 13323 13209
rect 13630 13200 13636 13212
rect 13688 13200 13694 13252
rect 8846 13172 8852 13184
rect 8496 13144 8852 13172
rect 8205 13135 8263 13141
rect 8846 13132 8852 13144
rect 8904 13132 8910 13184
rect 9030 13132 9036 13184
rect 9088 13172 9094 13184
rect 9582 13172 9588 13184
rect 9088 13144 9588 13172
rect 9088 13132 9094 13144
rect 9582 13132 9588 13144
rect 9640 13172 9646 13184
rect 10413 13175 10471 13181
rect 10413 13172 10425 13175
rect 9640 13144 10425 13172
rect 9640 13132 9646 13144
rect 10413 13141 10425 13144
rect 10459 13141 10471 13175
rect 10413 13135 10471 13141
rect 10873 13175 10931 13181
rect 10873 13141 10885 13175
rect 10919 13172 10931 13175
rect 11330 13172 11336 13184
rect 10919 13144 11336 13172
rect 10919 13141 10931 13144
rect 10873 13135 10931 13141
rect 11330 13132 11336 13144
rect 11388 13172 11394 13184
rect 12066 13172 12072 13184
rect 11388 13144 12072 13172
rect 11388 13132 11394 13144
rect 12066 13132 12072 13144
rect 12124 13132 12130 13184
rect 12250 13132 12256 13184
rect 12308 13172 12314 13184
rect 12345 13175 12403 13181
rect 12345 13172 12357 13175
rect 12308 13144 12357 13172
rect 12308 13132 12314 13144
rect 12345 13141 12357 13144
rect 12391 13141 12403 13175
rect 12802 13172 12808 13184
rect 12763 13144 12808 13172
rect 12345 13135 12403 13141
rect 12802 13132 12808 13144
rect 12860 13132 12866 13184
rect 13354 13172 13360 13184
rect 13315 13144 13360 13172
rect 13354 13132 13360 13144
rect 13412 13132 13418 13184
rect 13538 13172 13544 13184
rect 13499 13144 13544 13172
rect 13538 13132 13544 13144
rect 13596 13132 13602 13184
rect 14182 13172 14188 13184
rect 14143 13144 14188 13172
rect 14182 13132 14188 13144
rect 14240 13132 14246 13184
rect 14292 13172 14320 13280
rect 14728 13271 14740 13280
rect 14792 13308 14798 13320
rect 15286 13308 15292 13320
rect 14792 13280 15292 13308
rect 14734 13268 14740 13271
rect 14792 13268 14798 13280
rect 15286 13268 15292 13280
rect 15344 13268 15350 13320
rect 15930 13308 15936 13320
rect 15891 13280 15936 13308
rect 15930 13268 15936 13280
rect 15988 13268 15994 13320
rect 16031 13308 16059 13416
rect 16298 13404 16304 13416
rect 16356 13404 16362 13456
rect 19613 13447 19671 13453
rect 19613 13413 19625 13447
rect 19659 13444 19671 13447
rect 20346 13444 20352 13456
rect 19659 13416 20352 13444
rect 19659 13413 19671 13416
rect 19613 13407 19671 13413
rect 20346 13404 20352 13416
rect 20404 13404 20410 13456
rect 16942 13336 16948 13388
rect 17000 13376 17006 13388
rect 17037 13379 17095 13385
rect 17037 13376 17049 13379
rect 17000 13348 17049 13376
rect 17000 13336 17006 13348
rect 17037 13345 17049 13348
rect 17083 13345 17095 13379
rect 17037 13339 17095 13345
rect 17589 13379 17647 13385
rect 17589 13345 17601 13379
rect 17635 13376 17647 13379
rect 18230 13376 18236 13388
rect 17635 13348 18236 13376
rect 17635 13345 17647 13348
rect 17589 13339 17647 13345
rect 18230 13336 18236 13348
rect 18288 13336 18294 13388
rect 18782 13376 18788 13388
rect 18743 13348 18788 13376
rect 18782 13336 18788 13348
rect 18840 13376 18846 13388
rect 19518 13376 19524 13388
rect 18840 13348 19524 13376
rect 18840 13336 18846 13348
rect 19518 13336 19524 13348
rect 19576 13336 19582 13388
rect 20162 13376 20168 13388
rect 20123 13348 20168 13376
rect 20162 13336 20168 13348
rect 20220 13336 20226 13388
rect 20257 13379 20315 13385
rect 20257 13345 20269 13379
rect 20303 13376 20315 13379
rect 21174 13376 21180 13388
rect 20303 13348 21180 13376
rect 20303 13345 20315 13348
rect 20257 13339 20315 13345
rect 21174 13336 21180 13348
rect 21232 13336 21238 13388
rect 17494 13308 17500 13320
rect 16031 13280 17500 13308
rect 17494 13268 17500 13280
rect 17552 13308 17558 13320
rect 18601 13311 18659 13317
rect 18601 13308 18613 13311
rect 17552 13280 18613 13308
rect 17552 13268 17558 13280
rect 18601 13277 18613 13280
rect 18647 13308 18659 13311
rect 19245 13311 19303 13317
rect 19245 13308 19257 13311
rect 18647 13280 19257 13308
rect 18647 13277 18659 13280
rect 18601 13271 18659 13277
rect 19245 13277 19257 13280
rect 19291 13277 19303 13311
rect 19245 13271 19303 13277
rect 19429 13311 19487 13317
rect 19429 13277 19441 13311
rect 19475 13308 19487 13311
rect 19886 13308 19892 13320
rect 19475 13280 19892 13308
rect 19475 13277 19487 13280
rect 19429 13271 19487 13277
rect 19886 13268 19892 13280
rect 19944 13268 19950 13320
rect 20070 13308 20076 13320
rect 20031 13280 20076 13308
rect 20070 13268 20076 13280
rect 20128 13268 20134 13320
rect 20530 13268 20536 13320
rect 20588 13308 20594 13320
rect 20625 13311 20683 13317
rect 20625 13308 20637 13311
rect 20588 13280 20637 13308
rect 20588 13268 20594 13280
rect 20625 13277 20637 13280
rect 20671 13308 20683 13311
rect 20714 13308 20720 13320
rect 20671 13280 20720 13308
rect 20671 13277 20683 13280
rect 20625 13271 20683 13277
rect 20714 13268 20720 13280
rect 20772 13268 20778 13320
rect 20901 13311 20959 13317
rect 20901 13277 20913 13311
rect 20947 13277 20959 13311
rect 21266 13308 21272 13320
rect 21227 13280 21272 13308
rect 20901 13271 20959 13277
rect 14369 13243 14427 13249
rect 14369 13209 14381 13243
rect 14415 13240 14427 13243
rect 14642 13240 14648 13252
rect 14415 13212 14648 13240
rect 14415 13209 14427 13212
rect 14369 13203 14427 13209
rect 14642 13200 14648 13212
rect 14700 13200 14706 13252
rect 15470 13200 15476 13252
rect 15528 13240 15534 13252
rect 16853 13243 16911 13249
rect 15528 13212 16252 13240
rect 15528 13200 15534 13212
rect 14550 13172 14556 13184
rect 14292 13144 14556 13172
rect 14550 13132 14556 13144
rect 14608 13132 14614 13184
rect 14826 13132 14832 13184
rect 14884 13172 14890 13184
rect 15194 13172 15200 13184
rect 14884 13144 15200 13172
rect 14884 13132 14890 13144
rect 15194 13132 15200 13144
rect 15252 13172 15258 13184
rect 15841 13175 15899 13181
rect 15841 13172 15853 13175
rect 15252 13144 15853 13172
rect 15252 13132 15258 13144
rect 15841 13141 15853 13144
rect 15887 13172 15899 13175
rect 16114 13172 16120 13184
rect 15887 13144 16120 13172
rect 15887 13141 15899 13144
rect 15841 13135 15899 13141
rect 16114 13132 16120 13144
rect 16172 13132 16178 13184
rect 16224 13181 16252 13212
rect 16853 13209 16865 13243
rect 16899 13240 16911 13243
rect 17218 13240 17224 13252
rect 16899 13212 17224 13240
rect 16899 13209 16911 13212
rect 16853 13203 16911 13209
rect 17218 13200 17224 13212
rect 17276 13200 17282 13252
rect 17310 13200 17316 13252
rect 17368 13240 17374 13252
rect 17773 13243 17831 13249
rect 17773 13240 17785 13243
rect 17368 13212 17785 13240
rect 17368 13200 17374 13212
rect 17773 13209 17785 13212
rect 17819 13209 17831 13243
rect 17773 13203 17831 13209
rect 19058 13200 19064 13252
rect 19116 13240 19122 13252
rect 20916 13240 20944 13271
rect 21266 13268 21272 13280
rect 21324 13268 21330 13320
rect 19116 13212 20944 13240
rect 19116 13200 19122 13212
rect 16209 13175 16267 13181
rect 16209 13141 16221 13175
rect 16255 13172 16267 13175
rect 16945 13175 17003 13181
rect 16945 13172 16957 13175
rect 16255 13144 16957 13172
rect 16255 13141 16267 13144
rect 16209 13135 16267 13141
rect 16945 13141 16957 13144
rect 16991 13172 17003 13175
rect 17034 13172 17040 13184
rect 16991 13144 17040 13172
rect 16991 13141 17003 13144
rect 16945 13135 17003 13141
rect 17034 13132 17040 13144
rect 17092 13132 17098 13184
rect 17586 13132 17592 13184
rect 17644 13172 17650 13184
rect 17681 13175 17739 13181
rect 17681 13172 17693 13175
rect 17644 13144 17693 13172
rect 17644 13132 17650 13144
rect 17681 13141 17693 13144
rect 17727 13141 17739 13175
rect 17681 13135 17739 13141
rect 18141 13175 18199 13181
rect 18141 13141 18153 13175
rect 18187 13172 18199 13175
rect 18322 13172 18328 13184
rect 18187 13144 18328 13172
rect 18187 13141 18199 13144
rect 18141 13135 18199 13141
rect 18322 13132 18328 13144
rect 18380 13132 18386 13184
rect 18690 13132 18696 13184
rect 18748 13172 18754 13184
rect 21082 13172 21088 13184
rect 18748 13144 18793 13172
rect 21043 13144 21088 13172
rect 18748 13132 18754 13144
rect 21082 13132 21088 13144
rect 21140 13132 21146 13184
rect 21450 13172 21456 13184
rect 21411 13144 21456 13172
rect 21450 13132 21456 13144
rect 21508 13132 21514 13184
rect 22002 13132 22008 13184
rect 22060 13172 22066 13184
rect 22830 13172 22836 13184
rect 22060 13144 22836 13172
rect 22060 13132 22066 13144
rect 22830 13132 22836 13144
rect 22888 13132 22894 13184
rect 1104 13082 22056 13104
rect 1104 13030 6148 13082
rect 6200 13030 6212 13082
rect 6264 13030 6276 13082
rect 6328 13030 6340 13082
rect 6392 13030 6404 13082
rect 6456 13030 11346 13082
rect 11398 13030 11410 13082
rect 11462 13030 11474 13082
rect 11526 13030 11538 13082
rect 11590 13030 11602 13082
rect 11654 13030 16544 13082
rect 16596 13030 16608 13082
rect 16660 13030 16672 13082
rect 16724 13030 16736 13082
rect 16788 13030 16800 13082
rect 16852 13030 21742 13082
rect 21794 13030 21806 13082
rect 21858 13030 21870 13082
rect 21922 13030 21934 13082
rect 21986 13030 21998 13082
rect 22050 13030 22056 13082
rect 1104 13008 22056 13030
rect 1486 12968 1492 12980
rect 1447 12940 1492 12968
rect 1486 12928 1492 12940
rect 1544 12928 1550 12980
rect 3050 12928 3056 12980
rect 3108 12968 3114 12980
rect 4249 12971 4307 12977
rect 4249 12968 4261 12971
rect 3108 12940 4261 12968
rect 3108 12928 3114 12940
rect 4249 12937 4261 12940
rect 4295 12937 4307 12971
rect 6914 12968 6920 12980
rect 4249 12931 4307 12937
rect 4356 12940 6920 12968
rect 2498 12900 2504 12912
rect 1964 12872 2504 12900
rect 1964 12844 1992 12872
rect 2498 12860 2504 12872
rect 2556 12860 2562 12912
rect 4062 12860 4068 12912
rect 4120 12900 4126 12912
rect 4356 12900 4384 12940
rect 6914 12928 6920 12940
rect 6972 12928 6978 12980
rect 7834 12968 7840 12980
rect 7795 12940 7840 12968
rect 7834 12928 7840 12940
rect 7892 12928 7898 12980
rect 8202 12968 8208 12980
rect 8163 12940 8208 12968
rect 8202 12928 8208 12940
rect 8260 12928 8266 12980
rect 9048 12940 9343 12968
rect 4120 12872 4384 12900
rect 4709 12903 4767 12909
rect 4120 12860 4126 12872
rect 4709 12869 4721 12903
rect 4755 12900 4767 12903
rect 8754 12900 8760 12912
rect 4755 12872 8760 12900
rect 4755 12869 4767 12872
rect 4709 12863 4767 12869
rect 8754 12860 8760 12872
rect 8812 12860 8818 12912
rect 8846 12860 8852 12912
rect 8904 12900 8910 12912
rect 9048 12900 9076 12940
rect 8904 12872 9076 12900
rect 9125 12903 9183 12909
rect 8904 12860 8910 12872
rect 9125 12869 9137 12903
rect 9171 12869 9183 12903
rect 9315 12900 9343 12940
rect 9398 12928 9404 12980
rect 9456 12968 9462 12980
rect 9585 12971 9643 12977
rect 9585 12968 9597 12971
rect 9456 12940 9597 12968
rect 9456 12928 9462 12940
rect 9585 12937 9597 12940
rect 9631 12937 9643 12971
rect 9585 12931 9643 12937
rect 10045 12971 10103 12977
rect 10045 12937 10057 12971
rect 10091 12968 10103 12971
rect 10594 12968 10600 12980
rect 10091 12940 10600 12968
rect 10091 12937 10103 12940
rect 10045 12931 10103 12937
rect 10594 12928 10600 12940
rect 10652 12928 10658 12980
rect 10778 12968 10784 12980
rect 10739 12940 10784 12968
rect 10778 12928 10784 12940
rect 10836 12928 10842 12980
rect 11054 12968 11060 12980
rect 11015 12940 11060 12968
rect 11054 12928 11060 12940
rect 11112 12928 11118 12980
rect 12066 12928 12072 12980
rect 12124 12968 12130 12980
rect 13357 12971 13415 12977
rect 13357 12968 13369 12971
rect 12124 12940 13369 12968
rect 12124 12928 12130 12940
rect 13357 12937 13369 12940
rect 13403 12968 13415 12971
rect 13817 12971 13875 12977
rect 13817 12968 13829 12971
rect 13403 12940 13829 12968
rect 13403 12937 13415 12940
rect 13357 12931 13415 12937
rect 13817 12937 13829 12940
rect 13863 12937 13875 12971
rect 14090 12968 14096 12980
rect 14051 12940 14096 12968
rect 13817 12931 13875 12937
rect 14090 12928 14096 12940
rect 14148 12928 14154 12980
rect 15381 12971 15439 12977
rect 15381 12937 15393 12971
rect 15427 12968 15439 12971
rect 15654 12968 15660 12980
rect 15427 12940 15660 12968
rect 15427 12937 15439 12940
rect 15381 12931 15439 12937
rect 15654 12928 15660 12940
rect 15712 12928 15718 12980
rect 16669 12971 16727 12977
rect 16669 12968 16681 12971
rect 15755 12940 16681 12968
rect 9766 12900 9772 12912
rect 9315 12872 9772 12900
rect 9125 12863 9183 12869
rect 1670 12832 1676 12844
rect 1631 12804 1676 12832
rect 1670 12792 1676 12804
rect 1728 12792 1734 12844
rect 1946 12832 1952 12844
rect 1859 12804 1952 12832
rect 1946 12792 1952 12804
rect 2004 12792 2010 12844
rect 2590 12792 2596 12844
rect 2648 12832 2654 12844
rect 2777 12835 2835 12841
rect 2777 12832 2789 12835
rect 2648 12804 2789 12832
rect 2648 12792 2654 12804
rect 2777 12801 2789 12804
rect 2823 12801 2835 12835
rect 2777 12795 2835 12801
rect 3044 12835 3102 12841
rect 3044 12801 3056 12835
rect 3090 12832 3102 12835
rect 4246 12832 4252 12844
rect 3090 12804 4252 12832
rect 3090 12801 3102 12804
rect 3044 12795 3102 12801
rect 4246 12792 4252 12804
rect 4304 12792 4310 12844
rect 4617 12835 4675 12841
rect 4617 12801 4629 12835
rect 4663 12832 4675 12835
rect 5721 12835 5779 12841
rect 4663 12804 5120 12832
rect 4663 12801 4675 12804
rect 4617 12795 4675 12801
rect 1762 12724 1768 12776
rect 1820 12764 1826 12776
rect 2608 12764 2636 12792
rect 1820 12736 2636 12764
rect 4801 12767 4859 12773
rect 1820 12724 1826 12736
rect 4801 12733 4813 12767
rect 4847 12733 4859 12767
rect 4801 12727 4859 12733
rect 382 12656 388 12708
rect 440 12696 446 12708
rect 1486 12696 1492 12708
rect 440 12668 1492 12696
rect 440 12656 446 12668
rect 1486 12656 1492 12668
rect 1544 12656 1550 12708
rect 3970 12656 3976 12708
rect 4028 12696 4034 12708
rect 4157 12699 4215 12705
rect 4157 12696 4169 12699
rect 4028 12668 4169 12696
rect 4028 12656 4034 12668
rect 4157 12665 4169 12668
rect 4203 12696 4215 12699
rect 4816 12696 4844 12727
rect 4203 12668 4844 12696
rect 5092 12696 5120 12804
rect 5721 12801 5733 12835
rect 5767 12832 5779 12835
rect 6454 12832 6460 12844
rect 5767 12804 6460 12832
rect 5767 12801 5779 12804
rect 5721 12795 5779 12801
rect 5166 12724 5172 12776
rect 5224 12764 5230 12776
rect 5736 12764 5764 12795
rect 6454 12792 6460 12804
rect 6512 12832 6518 12844
rect 6632 12836 6690 12841
rect 6564 12835 6690 12836
rect 6564 12832 6644 12835
rect 6512 12808 6644 12832
rect 6512 12804 6592 12808
rect 6512 12792 6518 12804
rect 6632 12801 6644 12808
rect 6678 12801 6690 12835
rect 6632 12795 6690 12801
rect 6914 12792 6920 12844
rect 6972 12832 6978 12844
rect 6972 12804 7420 12832
rect 6972 12792 6978 12804
rect 5902 12764 5908 12776
rect 5224 12736 5764 12764
rect 5863 12736 5908 12764
rect 5224 12724 5230 12736
rect 5902 12724 5908 12736
rect 5960 12724 5966 12776
rect 6365 12767 6423 12773
rect 6365 12733 6377 12767
rect 6411 12733 6423 12767
rect 6365 12727 6423 12733
rect 6178 12696 6184 12708
rect 5092 12668 6184 12696
rect 4203 12665 4215 12668
rect 4157 12659 4215 12665
rect 6178 12656 6184 12668
rect 6236 12656 6242 12708
rect 6380 12640 6408 12727
rect 7392 12696 7420 12804
rect 7466 12792 7472 12844
rect 7524 12832 7530 12844
rect 8297 12835 8355 12841
rect 8297 12832 8309 12835
rect 7524 12804 8309 12832
rect 7524 12792 7530 12804
rect 8297 12801 8309 12804
rect 8343 12832 8355 12835
rect 8662 12832 8668 12844
rect 8343 12804 8668 12832
rect 8343 12801 8355 12804
rect 8297 12795 8355 12801
rect 8662 12792 8668 12804
rect 8720 12792 8726 12844
rect 9140 12832 9168 12863
rect 9766 12860 9772 12872
rect 9824 12860 9830 12912
rect 10226 12860 10232 12912
rect 10284 12860 10290 12912
rect 10612 12900 10640 12928
rect 13262 12900 13268 12912
rect 10612 12872 12020 12900
rect 13223 12872 13268 12900
rect 8772 12804 9168 12832
rect 9953 12835 10011 12841
rect 8386 12724 8392 12776
rect 8444 12764 8450 12776
rect 8444 12736 8489 12764
rect 8444 12724 8450 12736
rect 8570 12724 8576 12776
rect 8628 12764 8634 12776
rect 8772 12764 8800 12804
rect 9953 12801 9965 12835
rect 9999 12832 10011 12835
rect 10042 12832 10048 12844
rect 9999 12804 10048 12832
rect 9999 12801 10011 12804
rect 9953 12795 10011 12801
rect 10042 12792 10048 12804
rect 10100 12792 10106 12844
rect 10244 12832 10272 12860
rect 10244 12804 11192 12832
rect 8938 12764 8944 12776
rect 8628 12736 8800 12764
rect 8899 12736 8944 12764
rect 8628 12724 8634 12736
rect 8938 12724 8944 12736
rect 8996 12724 9002 12776
rect 9033 12767 9091 12773
rect 9033 12733 9045 12767
rect 9079 12764 9091 12767
rect 10229 12767 10287 12773
rect 9079 12736 10189 12764
rect 9079 12733 9091 12736
rect 9033 12727 9091 12733
rect 7745 12699 7803 12705
rect 7392 12668 7696 12696
rect 2498 12588 2504 12640
rect 2556 12628 2562 12640
rect 6089 12631 6147 12637
rect 6089 12628 6101 12631
rect 2556 12600 6101 12628
rect 2556 12588 2562 12600
rect 6089 12597 6101 12600
rect 6135 12597 6147 12631
rect 6362 12628 6368 12640
rect 6275 12600 6368 12628
rect 6089 12591 6147 12597
rect 6362 12588 6368 12600
rect 6420 12628 6426 12640
rect 7558 12628 7564 12640
rect 6420 12600 7564 12628
rect 6420 12588 6426 12600
rect 7558 12588 7564 12600
rect 7616 12588 7622 12640
rect 7668 12628 7696 12668
rect 7745 12665 7757 12699
rect 7791 12696 7803 12699
rect 8404 12696 8432 12724
rect 7791 12668 8432 12696
rect 7791 12665 7803 12668
rect 7745 12659 7803 12665
rect 8478 12656 8484 12708
rect 8536 12696 8542 12708
rect 9048 12696 9076 12727
rect 9766 12696 9772 12708
rect 8536 12668 9076 12696
rect 9232 12668 9772 12696
rect 8536 12656 8542 12668
rect 9232 12628 9260 12668
rect 9766 12656 9772 12668
rect 9824 12656 9830 12708
rect 7668 12600 9260 12628
rect 9398 12588 9404 12640
rect 9456 12628 9462 12640
rect 9493 12631 9551 12637
rect 9493 12628 9505 12631
rect 9456 12600 9505 12628
rect 9456 12588 9462 12600
rect 9493 12597 9505 12600
rect 9539 12597 9551 12631
rect 10161 12628 10189 12736
rect 10229 12733 10241 12767
rect 10275 12764 10287 12767
rect 10502 12764 10508 12776
rect 10275 12736 10508 12764
rect 10275 12733 10287 12736
rect 10229 12727 10287 12733
rect 10502 12724 10508 12736
rect 10560 12724 10566 12776
rect 10594 12696 10600 12708
rect 10555 12668 10600 12696
rect 10594 12656 10600 12668
rect 10652 12656 10658 12708
rect 11164 12696 11192 12804
rect 11238 12792 11244 12844
rect 11296 12832 11302 12844
rect 11790 12841 11796 12844
rect 11333 12835 11391 12841
rect 11333 12832 11345 12835
rect 11296 12804 11345 12832
rect 11296 12792 11302 12804
rect 11333 12801 11345 12804
rect 11379 12832 11391 12835
rect 11517 12835 11575 12841
rect 11517 12832 11529 12835
rect 11379 12804 11529 12832
rect 11379 12801 11391 12804
rect 11333 12795 11391 12801
rect 11517 12801 11529 12804
rect 11563 12801 11575 12835
rect 11517 12795 11575 12801
rect 11784 12795 11796 12841
rect 11848 12832 11854 12844
rect 11992 12832 12020 12872
rect 13262 12860 13268 12872
rect 13320 12900 13326 12912
rect 13446 12900 13452 12912
rect 13320 12872 13452 12900
rect 13320 12860 13326 12872
rect 13446 12860 13452 12872
rect 13504 12860 13510 12912
rect 15013 12903 15071 12909
rect 15013 12900 15025 12903
rect 14200 12872 15025 12900
rect 13170 12832 13176 12844
rect 11848 12804 11884 12832
rect 11992 12804 13176 12832
rect 11790 12792 11796 12795
rect 11848 12792 11854 12804
rect 13170 12792 13176 12804
rect 13228 12792 13234 12844
rect 13078 12764 13084 12776
rect 13039 12736 13084 12764
rect 13078 12724 13084 12736
rect 13136 12724 13142 12776
rect 13722 12724 13728 12776
rect 13780 12724 13786 12776
rect 13740 12696 13768 12724
rect 14200 12696 14228 12872
rect 15013 12869 15025 12872
rect 15059 12869 15071 12903
rect 15013 12863 15071 12869
rect 15286 12860 15292 12912
rect 15344 12900 15350 12912
rect 15755 12900 15783 12940
rect 16669 12937 16681 12940
rect 16715 12968 16727 12971
rect 16942 12968 16948 12980
rect 16715 12940 16948 12968
rect 16715 12937 16727 12940
rect 16669 12931 16727 12937
rect 16942 12928 16948 12940
rect 17000 12928 17006 12980
rect 18046 12928 18052 12980
rect 18104 12968 18110 12980
rect 18141 12971 18199 12977
rect 18141 12968 18153 12971
rect 18104 12940 18153 12968
rect 18104 12928 18110 12940
rect 18141 12937 18153 12940
rect 18187 12937 18199 12971
rect 18141 12931 18199 12937
rect 18509 12971 18567 12977
rect 18509 12937 18521 12971
rect 18555 12968 18567 12971
rect 18969 12971 19027 12977
rect 18969 12968 18981 12971
rect 18555 12940 18981 12968
rect 18555 12937 18567 12940
rect 18509 12931 18567 12937
rect 18969 12937 18981 12940
rect 19015 12937 19027 12971
rect 19886 12968 19892 12980
rect 19847 12940 19892 12968
rect 18969 12931 19027 12937
rect 19886 12928 19892 12940
rect 19944 12928 19950 12980
rect 20349 12971 20407 12977
rect 20349 12937 20361 12971
rect 20395 12968 20407 12971
rect 21266 12968 21272 12980
rect 20395 12940 21272 12968
rect 20395 12937 20407 12940
rect 20349 12931 20407 12937
rect 21266 12928 21272 12940
rect 21324 12928 21330 12980
rect 15344 12872 15783 12900
rect 15344 12860 15350 12872
rect 16482 12860 16488 12912
rect 16540 12900 16546 12912
rect 16540 12872 17908 12900
rect 16540 12860 16546 12872
rect 14366 12832 14372 12844
rect 14327 12804 14372 12832
rect 14366 12792 14372 12804
rect 14424 12792 14430 12844
rect 15194 12832 15200 12844
rect 14752 12804 15200 12832
rect 14274 12724 14280 12776
rect 14332 12764 14338 12776
rect 14752 12773 14780 12804
rect 15194 12792 15200 12804
rect 15252 12792 15258 12844
rect 15470 12792 15476 12844
rect 15528 12832 15534 12844
rect 15654 12832 15660 12844
rect 15528 12804 15660 12832
rect 15528 12792 15534 12804
rect 15654 12792 15660 12804
rect 15712 12792 15718 12844
rect 15841 12835 15899 12841
rect 15841 12801 15853 12835
rect 15887 12832 15899 12835
rect 16393 12835 16451 12841
rect 16393 12832 16405 12835
rect 15887 12804 16405 12832
rect 15887 12801 15899 12804
rect 15841 12795 15899 12801
rect 16393 12801 16405 12804
rect 16439 12832 16451 12835
rect 16850 12832 16856 12844
rect 16439 12804 16856 12832
rect 16439 12801 16451 12804
rect 16393 12795 16451 12801
rect 14737 12767 14795 12773
rect 14332 12736 14688 12764
rect 14332 12724 14338 12736
rect 14461 12699 14519 12705
rect 14461 12696 14473 12699
rect 11164 12668 11560 12696
rect 10502 12628 10508 12640
rect 10161 12600 10508 12628
rect 9493 12591 9551 12597
rect 10502 12588 10508 12600
rect 10560 12588 10566 12640
rect 11054 12588 11060 12640
rect 11112 12628 11118 12640
rect 11149 12631 11207 12637
rect 11149 12628 11161 12631
rect 11112 12600 11161 12628
rect 11112 12588 11118 12600
rect 11149 12597 11161 12600
rect 11195 12597 11207 12631
rect 11532 12628 11560 12668
rect 12820 12668 14473 12696
rect 12820 12628 12848 12668
rect 14461 12665 14473 12668
rect 14507 12665 14519 12699
rect 14660 12696 14688 12736
rect 14737 12733 14749 12767
rect 14783 12733 14795 12767
rect 14918 12764 14924 12776
rect 14879 12736 14924 12764
rect 14737 12727 14795 12733
rect 14918 12724 14924 12736
rect 14976 12724 14982 12776
rect 15562 12724 15568 12776
rect 15620 12764 15626 12776
rect 15856 12764 15884 12795
rect 16850 12792 16856 12804
rect 16908 12832 16914 12844
rect 17782 12835 17840 12841
rect 17782 12832 17794 12835
rect 16908 12804 17794 12832
rect 16908 12792 16914 12804
rect 17782 12801 17794 12804
rect 17828 12801 17840 12835
rect 17880 12832 17908 12872
rect 18322 12860 18328 12912
rect 18380 12900 18386 12912
rect 18601 12903 18659 12909
rect 18601 12900 18613 12903
rect 18380 12872 18613 12900
rect 18380 12860 18386 12872
rect 18601 12869 18613 12872
rect 18647 12869 18659 12903
rect 18601 12863 18659 12869
rect 19337 12903 19395 12909
rect 19337 12869 19349 12903
rect 19383 12900 19395 12903
rect 20254 12900 20260 12912
rect 19383 12872 20260 12900
rect 19383 12869 19395 12872
rect 19337 12863 19395 12869
rect 20254 12860 20260 12872
rect 20312 12860 20318 12912
rect 21085 12903 21143 12909
rect 21085 12900 21097 12903
rect 20548 12872 21097 12900
rect 20548 12841 20576 12872
rect 21085 12869 21097 12872
rect 21131 12900 21143 12903
rect 21174 12900 21180 12912
rect 21131 12872 21180 12900
rect 21131 12869 21143 12872
rect 21085 12863 21143 12869
rect 21174 12860 21180 12872
rect 21232 12860 21238 12912
rect 20073 12835 20131 12841
rect 20073 12832 20085 12835
rect 17880 12804 20085 12832
rect 17782 12795 17840 12801
rect 20073 12801 20085 12804
rect 20119 12801 20131 12835
rect 20073 12795 20131 12801
rect 20165 12835 20223 12841
rect 20165 12801 20177 12835
rect 20211 12801 20223 12835
rect 20165 12795 20223 12801
rect 20533 12835 20591 12841
rect 20533 12801 20545 12835
rect 20579 12801 20591 12835
rect 21266 12832 21272 12844
rect 21227 12804 21272 12832
rect 20533 12795 20591 12801
rect 18049 12767 18107 12773
rect 15620 12736 15884 12764
rect 16500 12736 17080 12764
rect 15620 12724 15626 12736
rect 15473 12699 15531 12705
rect 15473 12696 15485 12699
rect 14660 12668 15485 12696
rect 14461 12659 14519 12665
rect 15473 12665 15485 12668
rect 15519 12665 15531 12699
rect 15473 12659 15531 12665
rect 15654 12656 15660 12708
rect 15712 12696 15718 12708
rect 16500 12696 16528 12736
rect 15712 12668 16528 12696
rect 15712 12656 15718 12668
rect 11532 12600 12848 12628
rect 12897 12631 12955 12637
rect 11149 12591 11207 12597
rect 12897 12597 12909 12631
rect 12943 12628 12955 12631
rect 13538 12628 13544 12640
rect 12943 12600 13544 12628
rect 12943 12597 12955 12600
rect 12897 12591 12955 12597
rect 13538 12588 13544 12600
rect 13596 12588 13602 12640
rect 13722 12628 13728 12640
rect 13683 12600 13728 12628
rect 13722 12588 13728 12600
rect 13780 12588 13786 12640
rect 13814 12588 13820 12640
rect 13872 12628 13878 12640
rect 13998 12628 14004 12640
rect 13872 12600 14004 12628
rect 13872 12588 13878 12600
rect 13998 12588 14004 12600
rect 14056 12588 14062 12640
rect 14826 12588 14832 12640
rect 14884 12628 14890 12640
rect 15930 12628 15936 12640
rect 14884 12600 15936 12628
rect 14884 12588 14890 12600
rect 15930 12588 15936 12600
rect 15988 12628 15994 12640
rect 16942 12628 16948 12640
rect 15988 12600 16948 12628
rect 15988 12588 15994 12600
rect 16942 12588 16948 12600
rect 17000 12588 17006 12640
rect 17052 12628 17080 12736
rect 18049 12733 18061 12767
rect 18095 12764 18107 12767
rect 18414 12764 18420 12776
rect 18095 12736 18420 12764
rect 18095 12733 18107 12736
rect 18049 12727 18107 12733
rect 18064 12628 18092 12727
rect 18414 12724 18420 12736
rect 18472 12724 18478 12776
rect 18782 12764 18788 12776
rect 18743 12736 18788 12764
rect 18782 12724 18788 12736
rect 18840 12724 18846 12776
rect 19426 12764 19432 12776
rect 19387 12736 19432 12764
rect 19426 12724 19432 12736
rect 19484 12724 19490 12776
rect 19521 12767 19579 12773
rect 19521 12733 19533 12767
rect 19567 12733 19579 12767
rect 19521 12727 19579 12733
rect 18230 12656 18236 12708
rect 18288 12696 18294 12708
rect 19536 12696 19564 12727
rect 19610 12724 19616 12776
rect 19668 12764 19674 12776
rect 20180 12764 20208 12795
rect 21266 12792 21272 12804
rect 21324 12792 21330 12844
rect 19668 12736 20208 12764
rect 19668 12724 19674 12736
rect 18288 12668 19564 12696
rect 18288 12656 18294 12668
rect 17052 12600 18092 12628
rect 18322 12588 18328 12640
rect 18380 12628 18386 12640
rect 19426 12628 19432 12640
rect 18380 12600 19432 12628
rect 18380 12588 18386 12600
rect 19426 12588 19432 12600
rect 19484 12628 19490 12640
rect 20346 12628 20352 12640
rect 19484 12600 20352 12628
rect 19484 12588 19490 12600
rect 20346 12588 20352 12600
rect 20404 12588 20410 12640
rect 20714 12588 20720 12640
rect 20772 12628 20778 12640
rect 20898 12628 20904 12640
rect 20772 12600 20904 12628
rect 20772 12588 20778 12600
rect 20898 12588 20904 12600
rect 20956 12588 20962 12640
rect 21450 12628 21456 12640
rect 21411 12600 21456 12628
rect 21450 12588 21456 12600
rect 21508 12588 21514 12640
rect 1104 12538 21896 12560
rect 1104 12486 3549 12538
rect 3601 12486 3613 12538
rect 3665 12486 3677 12538
rect 3729 12486 3741 12538
rect 3793 12486 3805 12538
rect 3857 12486 8747 12538
rect 8799 12486 8811 12538
rect 8863 12486 8875 12538
rect 8927 12486 8939 12538
rect 8991 12486 9003 12538
rect 9055 12486 13945 12538
rect 13997 12486 14009 12538
rect 14061 12486 14073 12538
rect 14125 12486 14137 12538
rect 14189 12486 14201 12538
rect 14253 12486 19143 12538
rect 19195 12486 19207 12538
rect 19259 12486 19271 12538
rect 19323 12486 19335 12538
rect 19387 12486 19399 12538
rect 19451 12486 21896 12538
rect 1104 12464 21896 12486
rect 1578 12424 1584 12436
rect 1539 12396 1584 12424
rect 1578 12384 1584 12396
rect 1636 12384 1642 12436
rect 1670 12384 1676 12436
rect 1728 12424 1734 12436
rect 3145 12427 3203 12433
rect 3145 12424 3157 12427
rect 1728 12396 3157 12424
rect 1728 12384 1734 12396
rect 3145 12393 3157 12396
rect 3191 12393 3203 12427
rect 3145 12387 3203 12393
rect 3234 12384 3240 12436
rect 3292 12424 3298 12436
rect 3421 12427 3479 12433
rect 3421 12424 3433 12427
rect 3292 12396 3433 12424
rect 3292 12384 3298 12396
rect 3421 12393 3433 12396
rect 3467 12393 3479 12427
rect 3421 12387 3479 12393
rect 4801 12427 4859 12433
rect 4801 12393 4813 12427
rect 4847 12424 4859 12427
rect 5166 12424 5172 12436
rect 4847 12396 5172 12424
rect 4847 12393 4859 12396
rect 4801 12387 4859 12393
rect 5166 12384 5172 12396
rect 5224 12384 5230 12436
rect 9214 12424 9220 12436
rect 5276 12396 9220 12424
rect 2866 12316 2872 12368
rect 2924 12356 2930 12368
rect 3881 12359 3939 12365
rect 3881 12356 3893 12359
rect 2924 12328 3893 12356
rect 2924 12316 2930 12328
rect 3881 12325 3893 12328
rect 3927 12356 3939 12359
rect 3970 12356 3976 12368
rect 3927 12328 3976 12356
rect 3927 12325 3939 12328
rect 3881 12319 3939 12325
rect 3970 12316 3976 12328
rect 4028 12316 4034 12368
rect 5276 12356 5304 12396
rect 9214 12384 9220 12396
rect 9272 12424 9278 12436
rect 9490 12424 9496 12436
rect 9272 12396 9496 12424
rect 9272 12384 9278 12396
rect 9490 12384 9496 12396
rect 9548 12384 9554 12436
rect 10042 12424 10048 12436
rect 10003 12396 10048 12424
rect 10042 12384 10048 12396
rect 10100 12424 10106 12436
rect 12802 12424 12808 12436
rect 10100 12396 12808 12424
rect 10100 12384 10106 12396
rect 12802 12384 12808 12396
rect 12860 12424 12866 12436
rect 13633 12427 13691 12433
rect 13633 12424 13645 12427
rect 12860 12396 13645 12424
rect 12860 12384 12866 12396
rect 13633 12393 13645 12396
rect 13679 12393 13691 12427
rect 13633 12387 13691 12393
rect 4540 12328 5304 12356
rect 4246 12248 4252 12300
rect 4304 12288 4310 12300
rect 4540 12297 4568 12328
rect 7190 12316 7196 12368
rect 7248 12356 7254 12368
rect 7469 12359 7527 12365
rect 7469 12356 7481 12359
rect 7248 12328 7481 12356
rect 7248 12316 7254 12328
rect 7469 12325 7481 12328
rect 7515 12356 7527 12359
rect 7558 12356 7564 12368
rect 7515 12328 7564 12356
rect 7515 12325 7527 12328
rect 7469 12319 7527 12325
rect 7558 12316 7564 12328
rect 7616 12316 7622 12368
rect 7834 12316 7840 12368
rect 7892 12356 7898 12368
rect 10321 12359 10379 12365
rect 10321 12356 10333 12359
rect 7892 12328 10333 12356
rect 7892 12316 7898 12328
rect 10321 12325 10333 12328
rect 10367 12325 10379 12359
rect 13648 12356 13676 12387
rect 13814 12384 13820 12436
rect 13872 12424 13878 12436
rect 14461 12427 14519 12433
rect 14461 12424 14473 12427
rect 13872 12396 14473 12424
rect 13872 12384 13878 12396
rect 14461 12393 14473 12396
rect 14507 12393 14519 12427
rect 14826 12424 14832 12436
rect 14461 12387 14519 12393
rect 14568 12396 14832 12424
rect 14568 12356 14596 12396
rect 14826 12384 14832 12396
rect 14884 12384 14890 12436
rect 14918 12384 14924 12436
rect 14976 12424 14982 12436
rect 15381 12427 15439 12433
rect 15381 12424 15393 12427
rect 14976 12396 15393 12424
rect 14976 12384 14982 12396
rect 15381 12393 15393 12396
rect 15427 12393 15439 12427
rect 16850 12424 16856 12436
rect 15381 12387 15439 12393
rect 15488 12396 16712 12424
rect 16811 12396 16856 12424
rect 15488 12356 15516 12396
rect 13648 12328 14596 12356
rect 14660 12328 15516 12356
rect 16684 12356 16712 12396
rect 16850 12384 16856 12396
rect 16908 12384 16914 12436
rect 16942 12384 16948 12436
rect 17000 12424 17006 12436
rect 17037 12427 17095 12433
rect 17037 12424 17049 12427
rect 17000 12396 17049 12424
rect 17000 12384 17006 12396
rect 17037 12393 17049 12396
rect 17083 12424 17095 12427
rect 17586 12424 17592 12436
rect 17083 12396 17592 12424
rect 17083 12393 17095 12396
rect 17037 12387 17095 12393
rect 17586 12384 17592 12396
rect 17644 12384 17650 12436
rect 18322 12424 18328 12436
rect 17788 12396 18328 12424
rect 17788 12368 17816 12396
rect 18322 12384 18328 12396
rect 18380 12384 18386 12436
rect 18690 12424 18696 12436
rect 18651 12396 18696 12424
rect 18690 12384 18696 12396
rect 18748 12384 18754 12436
rect 17770 12356 17776 12368
rect 16684 12328 17776 12356
rect 10321 12319 10379 12325
rect 4525 12291 4583 12297
rect 4525 12288 4537 12291
rect 4304 12260 4537 12288
rect 4304 12248 4310 12260
rect 4525 12257 4537 12260
rect 4571 12257 4583 12291
rect 4525 12251 4583 12257
rect 6181 12291 6239 12297
rect 6181 12257 6193 12291
rect 6227 12288 6239 12291
rect 6362 12288 6368 12300
rect 6227 12260 6368 12288
rect 6227 12257 6239 12260
rect 6181 12251 6239 12257
rect 1397 12223 1455 12229
rect 1397 12189 1409 12223
rect 1443 12189 1455 12223
rect 1397 12183 1455 12189
rect 1673 12223 1731 12229
rect 1673 12189 1685 12223
rect 1719 12220 1731 12223
rect 1762 12220 1768 12232
rect 1719 12192 1768 12220
rect 1719 12189 1731 12192
rect 1673 12183 1731 12189
rect 1412 12152 1440 12183
rect 1762 12180 1768 12192
rect 1820 12180 1826 12232
rect 1946 12229 1952 12232
rect 1940 12220 1952 12229
rect 1907 12192 1952 12220
rect 1940 12183 1952 12192
rect 1946 12180 1952 12183
rect 2004 12180 2010 12232
rect 3326 12220 3332 12232
rect 3287 12192 3332 12220
rect 3326 12180 3332 12192
rect 3384 12180 3390 12232
rect 3786 12180 3792 12232
rect 3844 12220 3850 12232
rect 4341 12223 4399 12229
rect 4341 12220 4353 12223
rect 3844 12192 4353 12220
rect 3844 12180 3850 12192
rect 4341 12189 4353 12192
rect 4387 12189 4399 12223
rect 4341 12183 4399 12189
rect 4433 12223 4491 12229
rect 4433 12189 4445 12223
rect 4479 12220 4491 12223
rect 4798 12220 4804 12232
rect 4479 12192 4804 12220
rect 4479 12189 4491 12192
rect 4433 12183 4491 12189
rect 4798 12180 4804 12192
rect 4856 12180 4862 12232
rect 5534 12180 5540 12232
rect 5592 12220 5598 12232
rect 6196 12220 6224 12251
rect 6362 12248 6368 12260
rect 6420 12248 6426 12300
rect 6454 12248 6460 12300
rect 6512 12288 6518 12300
rect 6825 12291 6883 12297
rect 6825 12288 6837 12291
rect 6512 12260 6837 12288
rect 6512 12248 6518 12260
rect 6825 12257 6837 12260
rect 6871 12257 6883 12291
rect 6825 12251 6883 12257
rect 7282 12248 7288 12300
rect 7340 12288 7346 12300
rect 7742 12288 7748 12300
rect 7340 12260 7748 12288
rect 7340 12248 7346 12260
rect 7742 12248 7748 12260
rect 7800 12248 7806 12300
rect 7926 12248 7932 12300
rect 7984 12288 7990 12300
rect 8386 12288 8392 12300
rect 7984 12260 8392 12288
rect 7984 12248 7990 12260
rect 8386 12248 8392 12260
rect 8444 12248 8450 12300
rect 9398 12288 9404 12300
rect 9359 12260 9404 12288
rect 9398 12248 9404 12260
rect 9456 12248 9462 12300
rect 9490 12248 9496 12300
rect 9548 12288 9554 12300
rect 12897 12291 12955 12297
rect 12897 12288 12909 12291
rect 9548 12260 9593 12288
rect 12406 12260 12909 12288
rect 9548 12248 9554 12260
rect 5592 12192 6224 12220
rect 5592 12180 5598 12192
rect 6546 12180 6552 12232
rect 6604 12220 6610 12232
rect 7653 12223 7711 12229
rect 7653 12220 7665 12223
rect 6604 12192 7665 12220
rect 6604 12180 6610 12192
rect 7653 12189 7665 12192
rect 7699 12189 7711 12223
rect 8662 12220 8668 12232
rect 7653 12183 7711 12189
rect 7760 12192 7972 12220
rect 8623 12192 8668 12220
rect 1412 12124 4568 12152
rect 3050 12084 3056 12096
rect 3011 12056 3056 12084
rect 3050 12044 3056 12056
rect 3108 12044 3114 12096
rect 3970 12084 3976 12096
rect 3931 12056 3976 12084
rect 3970 12044 3976 12056
rect 4028 12044 4034 12096
rect 4540 12084 4568 12124
rect 5626 12112 5632 12164
rect 5684 12152 5690 12164
rect 5914 12155 5972 12161
rect 5914 12152 5926 12155
rect 5684 12124 5926 12152
rect 5684 12112 5690 12124
rect 5914 12121 5926 12124
rect 5960 12121 5972 12155
rect 5914 12115 5972 12121
rect 6178 12112 6184 12164
rect 6236 12152 6242 12164
rect 7760 12152 7788 12192
rect 6236 12124 7788 12152
rect 7944 12152 7972 12192
rect 8662 12180 8668 12192
rect 8720 12180 8726 12232
rect 9950 12220 9956 12232
rect 9863 12192 9956 12220
rect 9950 12180 9956 12192
rect 10008 12220 10014 12232
rect 11054 12220 11060 12232
rect 10008 12192 11060 12220
rect 10008 12180 10014 12192
rect 11054 12180 11060 12192
rect 11112 12180 11118 12232
rect 11324 12223 11382 12229
rect 11324 12189 11336 12223
rect 11370 12220 11382 12223
rect 11790 12220 11796 12232
rect 11370 12192 11796 12220
rect 11370 12189 11382 12192
rect 11324 12183 11382 12189
rect 11790 12180 11796 12192
rect 11848 12220 11854 12232
rect 12406 12220 12434 12260
rect 12897 12257 12909 12260
rect 12943 12288 12955 12291
rect 13078 12288 13084 12300
rect 12943 12260 13084 12288
rect 12943 12257 12955 12260
rect 12897 12251 12955 12257
rect 13078 12248 13084 12260
rect 13136 12248 13142 12300
rect 14660 12288 14688 12328
rect 17770 12316 17776 12328
rect 17828 12316 17834 12368
rect 17865 12359 17923 12365
rect 17865 12325 17877 12359
rect 17911 12356 17923 12359
rect 21266 12356 21272 12368
rect 17911 12328 21272 12356
rect 17911 12325 17923 12328
rect 17865 12319 17923 12325
rect 21266 12316 21272 12328
rect 21324 12316 21330 12368
rect 13740 12260 14688 12288
rect 11848 12192 12434 12220
rect 11848 12180 11854 12192
rect 12802 12180 12808 12232
rect 12860 12220 12866 12232
rect 12989 12223 13047 12229
rect 12989 12220 13001 12223
rect 12860 12192 13001 12220
rect 12860 12180 12866 12192
rect 12989 12189 13001 12192
rect 13035 12189 13047 12223
rect 12989 12183 13047 12189
rect 13354 12180 13360 12232
rect 13412 12220 13418 12232
rect 13630 12220 13636 12232
rect 13412 12192 13636 12220
rect 13412 12180 13418 12192
rect 13630 12180 13636 12192
rect 13688 12180 13694 12232
rect 7944 12124 8984 12152
rect 6236 12112 6242 12124
rect 6273 12087 6331 12093
rect 6273 12084 6285 12087
rect 4540 12056 6285 12084
rect 6273 12053 6285 12056
rect 6319 12053 6331 12087
rect 6638 12084 6644 12096
rect 6599 12056 6644 12084
rect 6273 12047 6331 12053
rect 6638 12044 6644 12056
rect 6696 12044 6702 12096
rect 6730 12044 6736 12096
rect 6788 12084 6794 12096
rect 6788 12056 6833 12084
rect 6788 12044 6794 12056
rect 7006 12044 7012 12096
rect 7064 12084 7070 12096
rect 7101 12087 7159 12093
rect 7101 12084 7113 12087
rect 7064 12056 7113 12084
rect 7064 12044 7070 12056
rect 7101 12053 7113 12056
rect 7147 12053 7159 12087
rect 7374 12084 7380 12096
rect 7335 12056 7380 12084
rect 7101 12047 7159 12053
rect 7374 12044 7380 12056
rect 7432 12044 7438 12096
rect 7466 12044 7472 12096
rect 7524 12084 7530 12096
rect 7834 12084 7840 12096
rect 7524 12056 7840 12084
rect 7524 12044 7530 12056
rect 7834 12044 7840 12056
rect 7892 12044 7898 12096
rect 7929 12087 7987 12093
rect 7929 12053 7941 12087
rect 7975 12084 7987 12087
rect 8018 12084 8024 12096
rect 7975 12056 8024 12084
rect 7975 12053 7987 12056
rect 7929 12047 7987 12053
rect 8018 12044 8024 12056
rect 8076 12044 8082 12096
rect 8113 12087 8171 12093
rect 8113 12053 8125 12087
rect 8159 12084 8171 12087
rect 8202 12084 8208 12096
rect 8159 12056 8208 12084
rect 8159 12053 8171 12056
rect 8113 12047 8171 12053
rect 8202 12044 8208 12056
rect 8260 12044 8266 12096
rect 8386 12044 8392 12096
rect 8444 12084 8450 12096
rect 8956 12093 8984 12124
rect 10594 12112 10600 12164
rect 10652 12152 10658 12164
rect 10781 12155 10839 12161
rect 10781 12152 10793 12155
rect 10652 12124 10793 12152
rect 10652 12112 10658 12124
rect 10781 12121 10793 12124
rect 10827 12121 10839 12155
rect 10781 12115 10839 12121
rect 11606 12112 11612 12164
rect 11664 12152 11670 12164
rect 12529 12155 12587 12161
rect 12529 12152 12541 12155
rect 11664 12124 12541 12152
rect 11664 12112 11670 12124
rect 12529 12121 12541 12124
rect 12575 12152 12587 12155
rect 13081 12155 13139 12161
rect 13081 12152 13093 12155
rect 12575 12124 13093 12152
rect 12575 12121 12587 12124
rect 12529 12115 12587 12121
rect 13081 12121 13093 12124
rect 13127 12152 13139 12155
rect 13740 12152 13768 12260
rect 14734 12248 14740 12300
rect 14792 12288 14798 12300
rect 14921 12291 14979 12297
rect 14792 12260 14837 12288
rect 14792 12248 14798 12260
rect 14921 12257 14933 12291
rect 14967 12288 14979 12291
rect 15194 12288 15200 12300
rect 14967 12260 15200 12288
rect 14967 12257 14979 12260
rect 14921 12251 14979 12257
rect 15194 12248 15200 12260
rect 15252 12248 15258 12300
rect 15470 12288 15476 12300
rect 15431 12260 15476 12288
rect 15470 12248 15476 12260
rect 15528 12248 15534 12300
rect 18141 12291 18199 12297
rect 18141 12257 18153 12291
rect 18187 12288 18199 12291
rect 18230 12288 18236 12300
rect 18187 12260 18236 12288
rect 18187 12257 18199 12260
rect 18141 12251 18199 12257
rect 18230 12248 18236 12260
rect 18288 12248 18294 12300
rect 20898 12288 20904 12300
rect 19444 12260 20904 12288
rect 13814 12180 13820 12232
rect 13872 12220 13878 12232
rect 17497 12223 17555 12229
rect 17497 12220 17509 12223
rect 13872 12192 17509 12220
rect 13872 12180 13878 12192
rect 17497 12189 17509 12192
rect 17543 12189 17555 12223
rect 17497 12183 17555 12189
rect 14093 12155 14151 12161
rect 14093 12152 14105 12155
rect 13127 12124 14105 12152
rect 13127 12121 13139 12124
rect 13081 12115 13139 12121
rect 14093 12121 14105 12124
rect 14139 12121 14151 12155
rect 14093 12115 14151 12121
rect 15740 12155 15798 12161
rect 15740 12121 15752 12155
rect 15786 12121 15798 12155
rect 15740 12115 15798 12121
rect 8481 12087 8539 12093
rect 8481 12084 8493 12087
rect 8444 12056 8493 12084
rect 8444 12044 8450 12056
rect 8481 12053 8493 12056
rect 8527 12053 8539 12087
rect 8481 12047 8539 12053
rect 8941 12087 8999 12093
rect 8941 12053 8953 12087
rect 8987 12053 8999 12087
rect 9306 12084 9312 12096
rect 9267 12056 9312 12084
rect 8941 12047 8999 12053
rect 9306 12044 9312 12056
rect 9364 12044 9370 12096
rect 9398 12044 9404 12096
rect 9456 12084 9462 12096
rect 9769 12087 9827 12093
rect 9769 12084 9781 12087
rect 9456 12056 9781 12084
rect 9456 12044 9462 12056
rect 9769 12053 9781 12056
rect 9815 12053 9827 12087
rect 9769 12047 9827 12053
rect 10134 12044 10140 12096
rect 10192 12084 10198 12096
rect 10413 12087 10471 12093
rect 10413 12084 10425 12087
rect 10192 12056 10425 12084
rect 10192 12044 10198 12056
rect 10413 12053 10425 12056
rect 10459 12053 10471 12087
rect 10686 12084 10692 12096
rect 10647 12056 10692 12084
rect 10413 12047 10471 12053
rect 10686 12044 10692 12056
rect 10744 12044 10750 12096
rect 12342 12044 12348 12096
rect 12400 12084 12406 12096
rect 12437 12087 12495 12093
rect 12437 12084 12449 12087
rect 12400 12056 12449 12084
rect 12400 12044 12406 12056
rect 12437 12053 12449 12056
rect 12483 12053 12495 12087
rect 13446 12084 13452 12096
rect 13407 12056 13452 12084
rect 12437 12047 12495 12053
rect 13446 12044 13452 12056
rect 13504 12044 13510 12096
rect 13906 12084 13912 12096
rect 13867 12056 13912 12084
rect 13906 12044 13912 12056
rect 13964 12044 13970 12096
rect 14369 12087 14427 12093
rect 14369 12053 14381 12087
rect 14415 12084 14427 12087
rect 14550 12084 14556 12096
rect 14415 12056 14556 12084
rect 14415 12053 14427 12056
rect 14369 12047 14427 12053
rect 14550 12044 14556 12056
rect 14608 12044 14614 12096
rect 15010 12044 15016 12096
rect 15068 12084 15074 12096
rect 15755 12084 15783 12115
rect 16206 12112 16212 12164
rect 16264 12152 16270 12164
rect 17221 12155 17279 12161
rect 17221 12152 17233 12155
rect 16264 12124 17233 12152
rect 16264 12112 16270 12124
rect 17221 12121 17233 12124
rect 17267 12152 17279 12155
rect 17310 12152 17316 12164
rect 17267 12124 17316 12152
rect 17267 12121 17279 12124
rect 17221 12115 17279 12121
rect 17310 12112 17316 12124
rect 17368 12112 17374 12164
rect 17512 12152 17540 12183
rect 17586 12180 17592 12232
rect 17644 12220 17650 12232
rect 17681 12223 17739 12229
rect 17681 12220 17693 12223
rect 17644 12192 17693 12220
rect 17644 12180 17650 12192
rect 17681 12189 17693 12192
rect 17727 12189 17739 12223
rect 18325 12223 18383 12229
rect 18325 12220 18337 12223
rect 17681 12183 17739 12189
rect 17788 12192 18337 12220
rect 17788 12152 17816 12192
rect 18325 12189 18337 12192
rect 18371 12189 18383 12223
rect 18325 12183 18383 12189
rect 18598 12180 18604 12232
rect 18656 12220 18662 12232
rect 19444 12229 19472 12260
rect 20898 12248 20904 12260
rect 20956 12248 20962 12300
rect 18877 12223 18935 12229
rect 18877 12220 18889 12223
rect 18656 12192 18889 12220
rect 18656 12180 18662 12192
rect 18877 12189 18889 12192
rect 18923 12220 18935 12223
rect 19245 12223 19303 12229
rect 19245 12220 19257 12223
rect 18923 12192 19257 12220
rect 18923 12189 18935 12192
rect 18877 12183 18935 12189
rect 19245 12189 19257 12192
rect 19291 12189 19303 12223
rect 19245 12183 19303 12189
rect 19429 12223 19487 12229
rect 19429 12189 19441 12223
rect 19475 12189 19487 12223
rect 19429 12183 19487 12189
rect 19794 12180 19800 12232
rect 19852 12220 19858 12232
rect 20165 12223 20223 12229
rect 20165 12220 20177 12223
rect 19852 12192 20177 12220
rect 19852 12180 19858 12192
rect 20165 12189 20177 12192
rect 20211 12220 20223 12223
rect 20533 12223 20591 12229
rect 20533 12220 20545 12223
rect 20211 12192 20545 12220
rect 20211 12189 20223 12192
rect 20165 12183 20223 12189
rect 20533 12189 20545 12192
rect 20579 12189 20591 12223
rect 20533 12183 20591 12189
rect 20990 12180 20996 12232
rect 21048 12220 21054 12232
rect 21269 12223 21327 12229
rect 21269 12220 21281 12223
rect 21048 12192 21281 12220
rect 21048 12180 21054 12192
rect 21269 12189 21281 12192
rect 21315 12189 21327 12223
rect 21269 12183 21327 12189
rect 17512 12124 17816 12152
rect 18046 12112 18052 12164
rect 18104 12152 18110 12164
rect 18966 12152 18972 12164
rect 18104 12124 18972 12152
rect 18104 12112 18110 12124
rect 18966 12112 18972 12124
rect 19024 12152 19030 12164
rect 19889 12155 19947 12161
rect 19889 12152 19901 12155
rect 19024 12124 19901 12152
rect 19024 12112 19030 12124
rect 19889 12121 19901 12124
rect 19935 12121 19947 12155
rect 19889 12115 19947 12121
rect 20714 12112 20720 12164
rect 20772 12152 20778 12164
rect 20901 12155 20959 12161
rect 20901 12152 20913 12155
rect 20772 12124 20913 12152
rect 20772 12112 20778 12124
rect 20901 12121 20913 12124
rect 20947 12121 20959 12155
rect 21082 12152 21088 12164
rect 21043 12124 21088 12152
rect 20901 12115 20959 12121
rect 21082 12112 21088 12124
rect 21140 12112 21146 12164
rect 15838 12084 15844 12096
rect 15068 12056 15113 12084
rect 15755 12056 15844 12084
rect 15068 12044 15074 12056
rect 15838 12044 15844 12056
rect 15896 12044 15902 12096
rect 18138 12044 18144 12096
rect 18196 12084 18202 12096
rect 18233 12087 18291 12093
rect 18233 12084 18245 12087
rect 18196 12056 18245 12084
rect 18196 12044 18202 12056
rect 18233 12053 18245 12056
rect 18279 12053 18291 12087
rect 18233 12047 18291 12053
rect 18874 12044 18880 12096
rect 18932 12084 18938 12096
rect 19061 12087 19119 12093
rect 19061 12084 19073 12087
rect 18932 12056 19073 12084
rect 18932 12044 18938 12056
rect 19061 12053 19073 12056
rect 19107 12053 19119 12087
rect 19061 12047 19119 12053
rect 19334 12044 19340 12096
rect 19392 12084 19398 12096
rect 19797 12087 19855 12093
rect 19797 12084 19809 12087
rect 19392 12056 19809 12084
rect 19392 12044 19398 12056
rect 19797 12053 19809 12056
rect 19843 12053 19855 12087
rect 21450 12084 21456 12096
rect 21411 12056 21456 12084
rect 19797 12047 19855 12053
rect 21450 12044 21456 12056
rect 21508 12044 21514 12096
rect 21726 12044 21732 12096
rect 21784 12084 21790 12096
rect 22738 12084 22744 12096
rect 21784 12056 22744 12084
rect 21784 12044 21790 12056
rect 22738 12044 22744 12056
rect 22796 12044 22802 12096
rect 1104 11994 22056 12016
rect 1104 11942 6148 11994
rect 6200 11942 6212 11994
rect 6264 11942 6276 11994
rect 6328 11942 6340 11994
rect 6392 11942 6404 11994
rect 6456 11942 11346 11994
rect 11398 11942 11410 11994
rect 11462 11942 11474 11994
rect 11526 11942 11538 11994
rect 11590 11942 11602 11994
rect 11654 11942 16544 11994
rect 16596 11942 16608 11994
rect 16660 11942 16672 11994
rect 16724 11942 16736 11994
rect 16788 11942 16800 11994
rect 16852 11942 21742 11994
rect 21794 11942 21806 11994
rect 21858 11942 21870 11994
rect 21922 11942 21934 11994
rect 21986 11942 21998 11994
rect 22050 11942 22056 11994
rect 1104 11920 22056 11942
rect 1854 11840 1860 11892
rect 1912 11880 1918 11892
rect 2498 11880 2504 11892
rect 1912 11852 2504 11880
rect 1912 11840 1918 11852
rect 2498 11840 2504 11852
rect 2556 11840 2562 11892
rect 2958 11840 2964 11892
rect 3016 11880 3022 11892
rect 3237 11883 3295 11889
rect 3237 11880 3249 11883
rect 3016 11852 3249 11880
rect 3016 11840 3022 11852
rect 3237 11849 3249 11852
rect 3283 11849 3295 11883
rect 3237 11843 3295 11849
rect 3418 11840 3424 11892
rect 3476 11880 3482 11892
rect 3605 11883 3663 11889
rect 3605 11880 3617 11883
rect 3476 11852 3617 11880
rect 3476 11840 3482 11852
rect 3605 11849 3617 11852
rect 3651 11849 3663 11883
rect 3605 11843 3663 11849
rect 3697 11883 3755 11889
rect 3697 11849 3709 11883
rect 3743 11880 3755 11883
rect 3970 11880 3976 11892
rect 3743 11852 3976 11880
rect 3743 11849 3755 11852
rect 3697 11843 3755 11849
rect 3970 11840 3976 11852
rect 4028 11840 4034 11892
rect 4338 11880 4344 11892
rect 4299 11852 4344 11880
rect 4338 11840 4344 11852
rect 4396 11840 4402 11892
rect 5721 11883 5779 11889
rect 5721 11849 5733 11883
rect 5767 11880 5779 11883
rect 6457 11883 6515 11889
rect 6457 11880 6469 11883
rect 5767 11852 6469 11880
rect 5767 11849 5779 11852
rect 5721 11843 5779 11849
rect 6457 11849 6469 11852
rect 6503 11849 6515 11883
rect 6457 11843 6515 11849
rect 6917 11883 6975 11889
rect 6917 11849 6929 11883
rect 6963 11880 6975 11883
rect 7285 11883 7343 11889
rect 7285 11880 7297 11883
rect 6963 11852 7297 11880
rect 6963 11849 6975 11852
rect 6917 11843 6975 11849
rect 7285 11849 7297 11852
rect 7331 11849 7343 11883
rect 7285 11843 7343 11849
rect 7374 11840 7380 11892
rect 7432 11880 7438 11892
rect 7745 11883 7803 11889
rect 7745 11880 7757 11883
rect 7432 11852 7757 11880
rect 7432 11840 7438 11852
rect 7745 11849 7757 11852
rect 7791 11849 7803 11883
rect 7745 11843 7803 11849
rect 7834 11840 7840 11892
rect 7892 11880 7898 11892
rect 8018 11880 8024 11892
rect 7892 11852 8024 11880
rect 7892 11840 7898 11852
rect 8018 11840 8024 11852
rect 8076 11840 8082 11892
rect 8113 11883 8171 11889
rect 8113 11849 8125 11883
rect 8159 11849 8171 11883
rect 8113 11843 8171 11849
rect 5169 11815 5227 11821
rect 5169 11812 5181 11815
rect 2240 11784 5181 11812
rect 2240 11756 2268 11784
rect 5169 11781 5181 11784
rect 5215 11781 5227 11815
rect 6546 11812 6552 11824
rect 5169 11775 5227 11781
rect 5276 11784 6552 11812
rect 1946 11744 1952 11756
rect 1907 11716 1952 11744
rect 1946 11704 1952 11716
rect 2004 11704 2010 11756
rect 2222 11744 2228 11756
rect 2135 11716 2228 11744
rect 2222 11704 2228 11716
rect 2280 11704 2286 11756
rect 2682 11744 2688 11756
rect 2643 11716 2688 11744
rect 2682 11704 2688 11716
rect 2740 11704 2746 11756
rect 2774 11704 2780 11756
rect 2832 11744 2838 11756
rect 4065 11747 4123 11753
rect 4065 11744 4077 11747
rect 2832 11716 4077 11744
rect 2832 11704 2838 11716
rect 4065 11713 4077 11716
rect 4111 11713 4123 11747
rect 4065 11707 4123 11713
rect 2498 11676 2504 11688
rect 2459 11648 2504 11676
rect 2498 11636 2504 11648
rect 2556 11636 2562 11688
rect 2590 11636 2596 11688
rect 2648 11676 2654 11688
rect 3878 11676 3884 11688
rect 2648 11648 2693 11676
rect 3839 11648 3884 11676
rect 2648 11636 2654 11648
rect 3878 11636 3884 11648
rect 3936 11636 3942 11688
rect 3970 11636 3976 11688
rect 4028 11676 4034 11688
rect 5276 11676 5304 11784
rect 6546 11772 6552 11784
rect 6604 11772 6610 11824
rect 6825 11815 6883 11821
rect 6825 11781 6837 11815
rect 6871 11812 6883 11815
rect 8128 11812 8156 11843
rect 8294 11840 8300 11892
rect 8352 11880 8358 11892
rect 8481 11883 8539 11889
rect 8481 11880 8493 11883
rect 8352 11852 8493 11880
rect 8352 11840 8358 11852
rect 8481 11849 8493 11852
rect 8527 11880 8539 11883
rect 8662 11880 8668 11892
rect 8527 11852 8668 11880
rect 8527 11849 8539 11852
rect 8481 11843 8539 11849
rect 8662 11840 8668 11852
rect 8720 11840 8726 11892
rect 11333 11883 11391 11889
rect 11333 11849 11345 11883
rect 11379 11880 11391 11883
rect 11606 11880 11612 11892
rect 11379 11852 11612 11880
rect 11379 11849 11391 11852
rect 11333 11843 11391 11849
rect 11606 11840 11612 11852
rect 11664 11880 11670 11892
rect 11790 11880 11796 11892
rect 11664 11852 11796 11880
rect 11664 11840 11670 11852
rect 11790 11840 11796 11852
rect 11848 11840 11854 11892
rect 11885 11883 11943 11889
rect 11885 11849 11897 11883
rect 11931 11880 11943 11883
rect 12250 11880 12256 11892
rect 11931 11852 12256 11880
rect 11931 11849 11943 11852
rect 11885 11843 11943 11849
rect 12250 11840 12256 11852
rect 12308 11840 12314 11892
rect 12710 11880 12716 11892
rect 12671 11852 12716 11880
rect 12710 11840 12716 11852
rect 12768 11880 12774 11892
rect 13262 11880 13268 11892
rect 12768 11852 13268 11880
rect 12768 11840 12774 11852
rect 13262 11840 13268 11852
rect 13320 11840 13326 11892
rect 13446 11840 13452 11892
rect 13504 11880 13510 11892
rect 13633 11883 13691 11889
rect 13633 11880 13645 11883
rect 13504 11852 13645 11880
rect 13504 11840 13510 11852
rect 13633 11849 13645 11852
rect 13679 11849 13691 11883
rect 13633 11843 13691 11849
rect 14090 11840 14096 11892
rect 14148 11880 14154 11892
rect 15102 11880 15108 11892
rect 14148 11852 15108 11880
rect 14148 11840 14154 11852
rect 15102 11840 15108 11852
rect 15160 11840 15166 11892
rect 15194 11840 15200 11892
rect 15252 11880 15258 11892
rect 15930 11880 15936 11892
rect 15252 11852 15936 11880
rect 15252 11840 15258 11852
rect 15930 11840 15936 11852
rect 15988 11840 15994 11892
rect 16209 11883 16267 11889
rect 16209 11849 16221 11883
rect 16255 11880 16267 11883
rect 16390 11880 16396 11892
rect 16255 11852 16396 11880
rect 16255 11849 16267 11852
rect 16209 11843 16267 11849
rect 16390 11840 16396 11852
rect 16448 11840 16454 11892
rect 16942 11880 16948 11892
rect 16903 11852 16948 11880
rect 16942 11840 16948 11852
rect 17000 11840 17006 11892
rect 18046 11880 18052 11892
rect 18007 11852 18052 11880
rect 18046 11840 18052 11852
rect 18104 11840 18110 11892
rect 18322 11840 18328 11892
rect 18380 11880 18386 11892
rect 18601 11883 18659 11889
rect 18601 11880 18613 11883
rect 18380 11852 18613 11880
rect 18380 11840 18386 11852
rect 18601 11849 18613 11852
rect 18647 11849 18659 11883
rect 18601 11843 18659 11849
rect 18690 11840 18696 11892
rect 18748 11880 18754 11892
rect 21266 11880 21272 11892
rect 18748 11852 21272 11880
rect 18748 11840 18754 11852
rect 21266 11840 21272 11852
rect 21324 11840 21330 11892
rect 6871 11784 8156 11812
rect 8496 11784 11652 11812
rect 6871 11781 6883 11784
rect 6825 11775 6883 11781
rect 5810 11744 5816 11756
rect 5771 11716 5816 11744
rect 5810 11704 5816 11716
rect 5868 11704 5874 11756
rect 7006 11704 7012 11756
rect 7064 11744 7070 11756
rect 7653 11747 7711 11753
rect 7653 11744 7665 11747
rect 7064 11716 7665 11744
rect 7064 11704 7070 11716
rect 7653 11713 7665 11716
rect 7699 11744 7711 11747
rect 8496 11744 8524 11784
rect 7699 11716 8524 11744
rect 8573 11747 8631 11753
rect 7699 11713 7711 11716
rect 7653 11707 7711 11713
rect 8573 11713 8585 11747
rect 8619 11744 8631 11747
rect 8846 11744 8852 11756
rect 8619 11716 8852 11744
rect 8619 11713 8631 11716
rect 8573 11707 8631 11713
rect 8846 11704 8852 11716
rect 8904 11704 8910 11756
rect 9122 11704 9128 11756
rect 9180 11744 9186 11756
rect 9401 11747 9459 11753
rect 9401 11744 9413 11747
rect 9180 11716 9413 11744
rect 9180 11704 9186 11716
rect 9401 11713 9413 11716
rect 9447 11744 9459 11747
rect 9769 11747 9827 11753
rect 9769 11744 9781 11747
rect 9447 11716 9781 11744
rect 9447 11713 9459 11716
rect 9401 11707 9459 11713
rect 9769 11713 9781 11716
rect 9815 11744 9827 11747
rect 10209 11747 10267 11753
rect 10209 11744 10221 11747
rect 9815 11716 10221 11744
rect 9815 11713 9827 11716
rect 9769 11707 9827 11713
rect 10209 11713 10221 11716
rect 10255 11713 10267 11747
rect 11624 11744 11652 11784
rect 11698 11772 11704 11824
rect 11756 11812 11762 11824
rect 12342 11812 12348 11824
rect 11756 11784 12348 11812
rect 11756 11772 11762 11784
rect 12342 11772 12348 11784
rect 12400 11812 12406 11824
rect 13541 11815 13599 11821
rect 12400 11784 13032 11812
rect 12400 11772 12406 11784
rect 12710 11744 12716 11756
rect 11624 11716 12716 11744
rect 10209 11707 10267 11713
rect 12710 11704 12716 11716
rect 12768 11704 12774 11756
rect 5626 11676 5632 11688
rect 4028 11648 5304 11676
rect 5587 11648 5632 11676
rect 4028 11636 4034 11648
rect 5626 11636 5632 11648
rect 5684 11636 5690 11688
rect 5718 11636 5724 11688
rect 5776 11676 5782 11688
rect 7101 11679 7159 11685
rect 5776 11648 6868 11676
rect 5776 11636 5782 11648
rect 3418 11568 3424 11620
rect 3476 11608 3482 11620
rect 4433 11611 4491 11617
rect 4433 11608 4445 11611
rect 3476 11580 4445 11608
rect 3476 11568 3482 11580
rect 4433 11577 4445 11580
rect 4479 11577 4491 11611
rect 4433 11571 4491 11577
rect 6181 11611 6239 11617
rect 6181 11577 6193 11611
rect 6227 11608 6239 11611
rect 6730 11608 6736 11620
rect 6227 11580 6736 11608
rect 6227 11577 6239 11580
rect 6181 11571 6239 11577
rect 6730 11568 6736 11580
rect 6788 11568 6794 11620
rect 6840 11608 6868 11648
rect 7101 11645 7113 11679
rect 7147 11676 7159 11679
rect 7190 11676 7196 11688
rect 7147 11648 7196 11676
rect 7147 11645 7159 11648
rect 7101 11639 7159 11645
rect 7190 11636 7196 11648
rect 7248 11636 7254 11688
rect 7929 11679 7987 11685
rect 7929 11645 7941 11679
rect 7975 11676 7987 11679
rect 8018 11676 8024 11688
rect 7975 11648 8024 11676
rect 7975 11645 7987 11648
rect 7929 11639 7987 11645
rect 8018 11636 8024 11648
rect 8076 11636 8082 11688
rect 8665 11679 8723 11685
rect 8665 11645 8677 11679
rect 8711 11645 8723 11679
rect 9950 11676 9956 11688
rect 9911 11648 9956 11676
rect 8665 11639 8723 11645
rect 7834 11608 7840 11620
rect 6840 11580 7840 11608
rect 7834 11568 7840 11580
rect 7892 11568 7898 11620
rect 8036 11608 8064 11636
rect 8680 11608 8708 11639
rect 9950 11636 9956 11648
rect 10008 11636 10014 11688
rect 11698 11676 11704 11688
rect 11659 11648 11704 11676
rect 11698 11636 11704 11648
rect 11756 11636 11762 11688
rect 11790 11636 11796 11688
rect 11848 11676 11854 11688
rect 11848 11648 11893 11676
rect 11848 11636 11854 11648
rect 12066 11636 12072 11688
rect 12124 11676 12130 11688
rect 13004 11685 13032 11784
rect 13541 11781 13553 11815
rect 13587 11812 13599 11815
rect 13722 11812 13728 11824
rect 13587 11784 13728 11812
rect 13587 11781 13599 11784
rect 13541 11775 13599 11781
rect 13722 11772 13728 11784
rect 13780 11772 13786 11824
rect 13906 11772 13912 11824
rect 13964 11812 13970 11824
rect 14369 11815 14427 11821
rect 14369 11812 14381 11815
rect 13964 11784 14381 11812
rect 13964 11772 13970 11784
rect 14369 11781 14381 11784
rect 14415 11812 14427 11815
rect 16669 11815 16727 11821
rect 16669 11812 16681 11815
rect 14415 11784 16681 11812
rect 14415 11781 14427 11784
rect 14369 11775 14427 11781
rect 16669 11781 16681 11784
rect 16715 11781 16727 11815
rect 16669 11775 16727 11781
rect 17770 11772 17776 11824
rect 17828 11812 17834 11824
rect 18141 11815 18199 11821
rect 18141 11812 18153 11815
rect 17828 11784 18153 11812
rect 17828 11772 17834 11784
rect 18141 11781 18153 11784
rect 18187 11781 18199 11815
rect 18141 11775 18199 11781
rect 18248 11784 18920 11812
rect 13170 11704 13176 11756
rect 13228 11744 13234 11756
rect 14277 11747 14335 11753
rect 14277 11744 14289 11747
rect 13228 11716 14289 11744
rect 13228 11704 13234 11716
rect 14277 11713 14289 11716
rect 14323 11713 14335 11747
rect 14277 11707 14335 11713
rect 15562 11704 15568 11756
rect 15620 11748 15626 11756
rect 15749 11748 15807 11753
rect 15620 11747 15807 11748
rect 15620 11720 15761 11747
rect 15620 11704 15626 11720
rect 15744 11716 15761 11720
rect 15749 11713 15761 11716
rect 15795 11713 15807 11747
rect 15749 11707 15807 11713
rect 15841 11747 15899 11753
rect 15841 11713 15853 11747
rect 15887 11744 15899 11747
rect 16114 11744 16120 11756
rect 15887 11716 16120 11744
rect 15887 11713 15899 11716
rect 15841 11707 15899 11713
rect 16114 11704 16120 11716
rect 16172 11704 16178 11756
rect 17218 11704 17224 11756
rect 17276 11744 17282 11756
rect 17494 11744 17500 11756
rect 17276 11716 17500 11744
rect 17276 11704 17282 11716
rect 17494 11704 17500 11716
rect 17552 11704 17558 11756
rect 17865 11747 17923 11753
rect 17865 11713 17877 11747
rect 17911 11744 17923 11747
rect 18248 11744 18276 11784
rect 17911 11716 18276 11744
rect 17911 11713 17923 11716
rect 17865 11707 17923 11713
rect 18322 11704 18328 11756
rect 18380 11744 18386 11756
rect 18782 11744 18788 11756
rect 18380 11716 18425 11744
rect 18743 11716 18788 11744
rect 18380 11704 18386 11716
rect 18782 11704 18788 11716
rect 18840 11704 18846 11756
rect 18892 11744 18920 11784
rect 19242 11772 19248 11824
rect 19300 11812 19306 11824
rect 19518 11812 19524 11824
rect 19300 11784 19524 11812
rect 19300 11772 19306 11784
rect 19518 11772 19524 11784
rect 19576 11772 19582 11824
rect 19794 11772 19800 11824
rect 19852 11812 19858 11824
rect 19990 11815 20048 11821
rect 19990 11812 20002 11815
rect 19852 11784 20002 11812
rect 19852 11772 19858 11784
rect 19990 11781 20002 11784
rect 20036 11781 20048 11815
rect 21082 11812 21088 11824
rect 19990 11775 20048 11781
rect 20364 11784 21088 11812
rect 20364 11744 20392 11784
rect 21082 11772 21088 11784
rect 21140 11772 21146 11824
rect 18892 11716 20392 11744
rect 20438 11704 20444 11756
rect 20496 11744 20502 11756
rect 20533 11747 20591 11753
rect 20533 11744 20545 11747
rect 20496 11716 20545 11744
rect 20496 11704 20502 11716
rect 20533 11713 20545 11716
rect 20579 11713 20591 11747
rect 20714 11744 20720 11756
rect 20675 11716 20720 11744
rect 20533 11707 20591 11713
rect 20714 11704 20720 11716
rect 20772 11704 20778 11756
rect 20806 11704 20812 11756
rect 20864 11744 20870 11756
rect 20993 11747 21051 11753
rect 20993 11744 21005 11747
rect 20864 11716 21005 11744
rect 20864 11704 20870 11716
rect 20993 11713 21005 11716
rect 21039 11744 21051 11747
rect 22462 11744 22468 11756
rect 21039 11716 22468 11744
rect 21039 11713 21051 11716
rect 20993 11707 21051 11713
rect 22462 11704 22468 11716
rect 22520 11704 22526 11756
rect 12805 11679 12863 11685
rect 12805 11676 12817 11679
rect 12124 11648 12817 11676
rect 12124 11636 12130 11648
rect 12805 11645 12817 11648
rect 12851 11645 12863 11679
rect 12805 11639 12863 11645
rect 12989 11679 13047 11685
rect 12989 11645 13001 11679
rect 13035 11676 13047 11679
rect 13725 11679 13783 11685
rect 13725 11676 13737 11679
rect 13035 11648 13737 11676
rect 13035 11645 13047 11648
rect 12989 11639 13047 11645
rect 13725 11645 13737 11648
rect 13771 11645 13783 11679
rect 13725 11639 13783 11645
rect 14185 11679 14243 11685
rect 14185 11645 14197 11679
rect 14231 11676 14243 11679
rect 14550 11676 14556 11688
rect 14231 11648 14556 11676
rect 14231 11645 14243 11648
rect 14185 11639 14243 11645
rect 12253 11611 12311 11617
rect 8036 11580 8708 11608
rect 8772 11580 9352 11608
rect 3053 11543 3111 11549
rect 3053 11509 3065 11543
rect 3099 11540 3111 11543
rect 3142 11540 3148 11552
rect 3099 11512 3148 11540
rect 3099 11509 3111 11512
rect 3053 11503 3111 11509
rect 3142 11500 3148 11512
rect 3200 11500 3206 11552
rect 3786 11500 3792 11552
rect 3844 11540 3850 11552
rect 3878 11540 3884 11552
rect 3844 11512 3884 11540
rect 3844 11500 3850 11512
rect 3878 11500 3884 11512
rect 3936 11500 3942 11552
rect 4522 11500 4528 11552
rect 4580 11540 4586 11552
rect 4617 11543 4675 11549
rect 4617 11540 4629 11543
rect 4580 11512 4629 11540
rect 4580 11500 4586 11512
rect 4617 11509 4629 11512
rect 4663 11509 4675 11543
rect 4798 11540 4804 11552
rect 4759 11512 4804 11540
rect 4617 11503 4675 11509
rect 4798 11500 4804 11512
rect 4856 11500 4862 11552
rect 5074 11540 5080 11552
rect 5035 11512 5080 11540
rect 5074 11500 5080 11512
rect 5132 11500 5138 11552
rect 7006 11500 7012 11552
rect 7064 11540 7070 11552
rect 8202 11540 8208 11552
rect 7064 11512 8208 11540
rect 7064 11500 7070 11512
rect 8202 11500 8208 11512
rect 8260 11540 8266 11552
rect 8772 11540 8800 11580
rect 8260 11512 8800 11540
rect 8260 11500 8266 11512
rect 8846 11500 8852 11552
rect 8904 11540 8910 11552
rect 9033 11543 9091 11549
rect 9033 11540 9045 11543
rect 8904 11512 9045 11540
rect 8904 11500 8910 11512
rect 9033 11509 9045 11512
rect 9079 11540 9091 11543
rect 9214 11540 9220 11552
rect 9079 11512 9220 11540
rect 9079 11509 9091 11512
rect 9033 11503 9091 11509
rect 9214 11500 9220 11512
rect 9272 11500 9278 11552
rect 9324 11540 9352 11580
rect 12253 11577 12265 11611
rect 12299 11608 12311 11611
rect 12820 11608 12848 11639
rect 14550 11636 14556 11648
rect 14608 11636 14614 11688
rect 15654 11636 15660 11688
rect 15712 11676 15718 11688
rect 19150 11676 19156 11688
rect 15712 11648 15757 11676
rect 18524 11648 19156 11676
rect 15712 11636 15718 11648
rect 14366 11608 14372 11620
rect 12299 11580 12664 11608
rect 12820 11580 14372 11608
rect 12299 11577 12311 11580
rect 12253 11571 12311 11577
rect 11790 11540 11796 11552
rect 9324 11512 11796 11540
rect 11790 11500 11796 11512
rect 11848 11500 11854 11552
rect 12342 11540 12348 11552
rect 12303 11512 12348 11540
rect 12342 11500 12348 11512
rect 12400 11500 12406 11552
rect 12636 11540 12664 11580
rect 14366 11568 14372 11580
rect 14424 11568 14430 11620
rect 14737 11611 14795 11617
rect 14737 11577 14749 11611
rect 14783 11608 14795 11611
rect 16942 11608 16948 11620
rect 14783 11580 15608 11608
rect 14783 11577 14795 11580
rect 14737 11571 14795 11577
rect 12802 11540 12808 11552
rect 12636 11512 12808 11540
rect 12802 11500 12808 11512
rect 12860 11500 12866 11552
rect 13173 11543 13231 11549
rect 13173 11509 13185 11543
rect 13219 11540 13231 11543
rect 13354 11540 13360 11552
rect 13219 11512 13360 11540
rect 13219 11509 13231 11512
rect 13173 11503 13231 11509
rect 13354 11500 13360 11512
rect 13412 11500 13418 11552
rect 13722 11500 13728 11552
rect 13780 11540 13786 11552
rect 14826 11540 14832 11552
rect 13780 11512 14832 11540
rect 13780 11500 13786 11512
rect 14826 11500 14832 11512
rect 14884 11540 14890 11552
rect 14921 11543 14979 11549
rect 14921 11540 14933 11543
rect 14884 11512 14933 11540
rect 14884 11500 14890 11512
rect 14921 11509 14933 11512
rect 14967 11509 14979 11543
rect 15194 11540 15200 11552
rect 15155 11512 15200 11540
rect 14921 11503 14979 11509
rect 15194 11500 15200 11512
rect 15252 11500 15258 11552
rect 15381 11543 15439 11549
rect 15381 11509 15393 11543
rect 15427 11540 15439 11543
rect 15470 11540 15476 11552
rect 15427 11512 15476 11540
rect 15427 11509 15439 11512
rect 15381 11503 15439 11509
rect 15470 11500 15476 11512
rect 15528 11500 15534 11552
rect 15580 11540 15608 11580
rect 16233 11580 16948 11608
rect 16233 11540 16261 11580
rect 16942 11568 16948 11580
rect 17000 11568 17006 11620
rect 17681 11611 17739 11617
rect 17681 11577 17693 11611
rect 17727 11608 17739 11611
rect 18046 11608 18052 11620
rect 17727 11580 18052 11608
rect 17727 11577 17739 11580
rect 17681 11571 17739 11577
rect 18046 11568 18052 11580
rect 18104 11568 18110 11620
rect 18524 11617 18552 11648
rect 19150 11636 19156 11648
rect 19208 11636 19214 11688
rect 20257 11679 20315 11685
rect 20257 11645 20269 11679
rect 20303 11645 20315 11679
rect 20257 11639 20315 11645
rect 18509 11611 18567 11617
rect 18509 11577 18521 11611
rect 18555 11577 18567 11611
rect 20272 11608 20300 11639
rect 20898 11608 20904 11620
rect 20272 11580 20904 11608
rect 18509 11571 18567 11577
rect 20898 11568 20904 11580
rect 20956 11568 20962 11620
rect 16390 11540 16396 11552
rect 15580 11512 16261 11540
rect 16351 11512 16396 11540
rect 16390 11500 16396 11512
rect 16448 11500 16454 11552
rect 17034 11540 17040 11552
rect 16995 11512 17040 11540
rect 17034 11500 17040 11512
rect 17092 11500 17098 11552
rect 17310 11540 17316 11552
rect 17271 11512 17316 11540
rect 17310 11500 17316 11512
rect 17368 11500 17374 11552
rect 17497 11543 17555 11549
rect 17497 11509 17509 11543
rect 17543 11540 17555 11543
rect 17770 11540 17776 11552
rect 17543 11512 17776 11540
rect 17543 11509 17555 11512
rect 17497 11503 17555 11509
rect 17770 11500 17776 11512
rect 17828 11500 17834 11552
rect 18230 11500 18236 11552
rect 18288 11540 18294 11552
rect 18877 11543 18935 11549
rect 18877 11540 18889 11543
rect 18288 11512 18889 11540
rect 18288 11500 18294 11512
rect 18877 11509 18889 11512
rect 18923 11509 18935 11543
rect 18877 11503 18935 11509
rect 19518 11500 19524 11552
rect 19576 11540 19582 11552
rect 20070 11540 20076 11552
rect 19576 11512 20076 11540
rect 19576 11500 19582 11512
rect 20070 11500 20076 11512
rect 20128 11500 20134 11552
rect 20441 11543 20499 11549
rect 20441 11509 20453 11543
rect 20487 11540 20499 11543
rect 20530 11540 20536 11552
rect 20487 11512 20536 11540
rect 20487 11509 20499 11512
rect 20441 11503 20499 11509
rect 20530 11500 20536 11512
rect 20588 11500 20594 11552
rect 1104 11450 21896 11472
rect 1104 11398 3549 11450
rect 3601 11398 3613 11450
rect 3665 11398 3677 11450
rect 3729 11398 3741 11450
rect 3793 11398 3805 11450
rect 3857 11398 8747 11450
rect 8799 11398 8811 11450
rect 8863 11398 8875 11450
rect 8927 11398 8939 11450
rect 8991 11398 9003 11450
rect 9055 11398 13945 11450
rect 13997 11398 14009 11450
rect 14061 11398 14073 11450
rect 14125 11398 14137 11450
rect 14189 11398 14201 11450
rect 14253 11398 19143 11450
rect 19195 11398 19207 11450
rect 19259 11398 19271 11450
rect 19323 11398 19335 11450
rect 19387 11398 19399 11450
rect 19451 11398 21896 11450
rect 1104 11376 21896 11398
rect 1486 11336 1492 11348
rect 1447 11308 1492 11336
rect 1486 11296 1492 11308
rect 1544 11296 1550 11348
rect 2225 11339 2283 11345
rect 2225 11305 2237 11339
rect 2271 11336 2283 11339
rect 2314 11336 2320 11348
rect 2271 11308 2320 11336
rect 2271 11305 2283 11308
rect 2225 11299 2283 11305
rect 2314 11296 2320 11308
rect 2372 11296 2378 11348
rect 5626 11336 5632 11348
rect 2746 11308 3556 11336
rect 5587 11308 5632 11336
rect 2038 11268 2044 11280
rect 1999 11240 2044 11268
rect 2038 11228 2044 11240
rect 2096 11228 2102 11280
rect 2332 11268 2360 11296
rect 2746 11268 2774 11308
rect 2332 11240 2774 11268
rect 3142 11228 3148 11280
rect 3200 11268 3206 11280
rect 3200 11240 3280 11268
rect 3200 11228 3206 11240
rect 2498 11200 2504 11212
rect 2459 11172 2504 11200
rect 2498 11160 2504 11172
rect 2556 11200 2562 11212
rect 2556 11172 3004 11200
rect 2556 11160 2562 11172
rect 2976 11144 3004 11172
rect 1670 11132 1676 11144
rect 1631 11104 1676 11132
rect 1670 11092 1676 11104
rect 1728 11092 1734 11144
rect 1854 11132 1860 11144
rect 1815 11104 1860 11132
rect 1854 11092 1860 11104
rect 1912 11092 1918 11144
rect 2958 11092 2964 11144
rect 3016 11132 3022 11144
rect 3153 11135 3211 11141
rect 3016 11104 3109 11132
rect 3016 11092 3022 11104
rect 3153 11101 3165 11135
rect 3199 11132 3211 11135
rect 3252 11132 3280 11240
rect 3326 11228 3332 11280
rect 3384 11268 3390 11280
rect 3528 11268 3556 11308
rect 5626 11296 5632 11308
rect 5684 11296 5690 11348
rect 6457 11339 6515 11345
rect 6457 11305 6469 11339
rect 6503 11336 6515 11339
rect 6638 11336 6644 11348
rect 6503 11308 6644 11336
rect 6503 11305 6515 11308
rect 6457 11299 6515 11305
rect 6638 11296 6644 11308
rect 6696 11296 6702 11348
rect 6730 11296 6736 11348
rect 6788 11336 6794 11348
rect 10594 11336 10600 11348
rect 6788 11308 10600 11336
rect 6788 11296 6794 11308
rect 10594 11296 10600 11308
rect 10652 11296 10658 11348
rect 11149 11339 11207 11345
rect 11149 11305 11161 11339
rect 11195 11336 11207 11339
rect 12066 11336 12072 11348
rect 11195 11308 12072 11336
rect 11195 11305 11207 11308
rect 11149 11299 11207 11305
rect 12066 11296 12072 11308
rect 12124 11296 12130 11348
rect 12452 11308 12664 11336
rect 4246 11268 4252 11280
rect 3384 11240 3429 11268
rect 3528 11240 4252 11268
rect 3384 11228 3390 11240
rect 4246 11228 4252 11240
rect 4304 11228 4310 11280
rect 5534 11200 5540 11212
rect 5276 11172 5540 11200
rect 3199 11104 3280 11132
rect 3605 11135 3663 11141
rect 3199 11101 3211 11104
rect 3153 11095 3211 11101
rect 3605 11101 3617 11135
rect 3651 11101 3663 11135
rect 3605 11095 3663 11101
rect 4157 11135 4215 11141
rect 4157 11101 4169 11135
rect 4203 11132 4215 11135
rect 4249 11135 4307 11141
rect 4249 11132 4261 11135
rect 4203 11104 4261 11132
rect 4203 11101 4215 11104
rect 4157 11095 4215 11101
rect 4249 11101 4261 11104
rect 4295 11132 4307 11135
rect 5276 11132 5304 11172
rect 5534 11160 5540 11172
rect 5592 11160 5598 11212
rect 5644 11200 5672 11296
rect 7469 11271 7527 11277
rect 7469 11268 7481 11271
rect 7116 11240 7481 11268
rect 7116 11209 7144 11240
rect 7469 11237 7481 11240
rect 7515 11237 7527 11271
rect 7469 11231 7527 11237
rect 8386 11228 8392 11280
rect 8444 11268 8450 11280
rect 8481 11271 8539 11277
rect 8481 11268 8493 11271
rect 8444 11240 8493 11268
rect 8444 11228 8450 11240
rect 8481 11237 8493 11240
rect 8527 11237 8539 11271
rect 8662 11268 8668 11280
rect 8623 11240 8668 11268
rect 8481 11231 8539 11237
rect 8662 11228 8668 11240
rect 8720 11268 8726 11280
rect 8938 11268 8944 11280
rect 8720 11240 8944 11268
rect 8720 11228 8726 11240
rect 8938 11228 8944 11240
rect 8996 11228 9002 11280
rect 9033 11271 9091 11277
rect 9033 11237 9045 11271
rect 9079 11268 9091 11271
rect 9122 11268 9128 11280
rect 9079 11240 9128 11268
rect 9079 11237 9091 11240
rect 9033 11231 9091 11237
rect 9122 11228 9128 11240
rect 9180 11228 9186 11280
rect 10870 11228 10876 11280
rect 10928 11268 10934 11280
rect 11974 11268 11980 11280
rect 10928 11240 11980 11268
rect 10928 11228 10934 11240
rect 11974 11228 11980 11240
rect 12032 11228 12038 11280
rect 5813 11203 5871 11209
rect 5813 11200 5825 11203
rect 5644 11172 5825 11200
rect 5813 11169 5825 11172
rect 5859 11169 5871 11203
rect 5813 11163 5871 11169
rect 7101 11203 7159 11209
rect 7101 11169 7113 11203
rect 7147 11169 7159 11203
rect 7101 11163 7159 11169
rect 7190 11160 7196 11212
rect 7248 11200 7254 11212
rect 8018 11200 8024 11212
rect 7248 11172 7293 11200
rect 7979 11172 8024 11200
rect 7248 11160 7254 11172
rect 8018 11160 8024 11172
rect 8076 11160 8082 11212
rect 9398 11160 9404 11212
rect 9456 11160 9462 11212
rect 10413 11203 10471 11209
rect 10413 11169 10425 11203
rect 10459 11200 10471 11203
rect 11054 11200 11060 11212
rect 10459 11172 11060 11200
rect 10459 11169 10471 11172
rect 10413 11163 10471 11169
rect 11054 11160 11060 11172
rect 11112 11160 11118 11212
rect 11425 11203 11483 11209
rect 11425 11169 11437 11203
rect 11471 11200 11483 11203
rect 11606 11200 11612 11212
rect 11471 11172 11612 11200
rect 11471 11169 11483 11172
rect 11425 11163 11483 11169
rect 11606 11160 11612 11172
rect 11664 11160 11670 11212
rect 12253 11203 12311 11209
rect 12253 11169 12265 11203
rect 12299 11200 12311 11203
rect 12452 11200 12480 11308
rect 12636 11268 12664 11308
rect 13262 11296 13268 11348
rect 13320 11336 13326 11348
rect 13725 11339 13783 11345
rect 13725 11336 13737 11339
rect 13320 11308 13737 11336
rect 13320 11296 13326 11308
rect 13725 11305 13737 11308
rect 13771 11305 13783 11339
rect 13725 11299 13783 11305
rect 15562 11296 15568 11348
rect 15620 11336 15626 11348
rect 15749 11339 15807 11345
rect 15749 11336 15761 11339
rect 15620 11308 15761 11336
rect 15620 11296 15626 11308
rect 15749 11305 15761 11308
rect 15795 11305 15807 11339
rect 19061 11339 19119 11345
rect 15749 11299 15807 11305
rect 15856 11308 18644 11336
rect 12636 11240 13584 11268
rect 13556 11212 13584 11240
rect 13354 11200 13360 11212
rect 12299 11172 12480 11200
rect 13315 11172 13360 11200
rect 12299 11169 12311 11172
rect 12253 11163 12311 11169
rect 13354 11160 13360 11172
rect 13412 11160 13418 11212
rect 13538 11200 13544 11212
rect 13499 11172 13544 11200
rect 13538 11160 13544 11172
rect 13596 11160 13602 11212
rect 14274 11200 14280 11212
rect 14235 11172 14280 11200
rect 14274 11160 14280 11172
rect 14332 11160 14338 11212
rect 15856 11200 15884 11308
rect 16577 11271 16635 11277
rect 16577 11268 16589 11271
rect 16224 11240 16589 11268
rect 16224 11209 16252 11240
rect 16577 11237 16589 11240
rect 16623 11237 16635 11271
rect 16577 11231 16635 11237
rect 16850 11228 16856 11280
rect 16908 11268 16914 11280
rect 17405 11271 17463 11277
rect 17405 11268 17417 11271
rect 16908 11240 17417 11268
rect 16908 11228 16914 11240
rect 17405 11237 17417 11240
rect 17451 11237 17463 11271
rect 18616 11268 18644 11308
rect 19061 11305 19073 11339
rect 19107 11336 19119 11339
rect 19886 11336 19892 11348
rect 19107 11308 19892 11336
rect 19107 11305 19119 11308
rect 19061 11299 19119 11305
rect 19886 11296 19892 11308
rect 19944 11296 19950 11348
rect 19242 11268 19248 11280
rect 18616 11240 19248 11268
rect 17405 11231 17463 11237
rect 19242 11228 19248 11240
rect 19300 11228 19306 11280
rect 15304 11172 15884 11200
rect 16209 11203 16267 11209
rect 4295 11104 5304 11132
rect 4295 11101 4307 11104
rect 4249 11095 4307 11101
rect 2866 11024 2872 11076
rect 2924 11064 2930 11076
rect 3620 11064 3648 11095
rect 5350 11092 5356 11144
rect 5408 11132 5414 11144
rect 6089 11135 6147 11141
rect 6089 11132 6101 11135
rect 5408 11104 6101 11132
rect 5408 11092 5414 11104
rect 6089 11101 6101 11104
rect 6135 11101 6147 11135
rect 6089 11095 6147 11101
rect 6546 11092 6552 11144
rect 6604 11132 6610 11144
rect 7208 11132 7236 11160
rect 7926 11132 7932 11144
rect 6604 11104 7236 11132
rect 7887 11104 7932 11132
rect 6604 11092 6610 11104
rect 7926 11092 7932 11104
rect 7984 11092 7990 11144
rect 8297 11135 8355 11141
rect 8297 11132 8309 11135
rect 8036 11104 8309 11132
rect 3789 11067 3847 11073
rect 3789 11064 3801 11067
rect 2924 11036 3801 11064
rect 2924 11024 2930 11036
rect 3789 11033 3801 11036
rect 3835 11033 3847 11067
rect 3789 11027 3847 11033
rect 4516 11067 4574 11073
rect 4516 11033 4528 11067
rect 4562 11064 4574 11067
rect 5534 11064 5540 11076
rect 4562 11036 5540 11064
rect 4562 11033 4574 11036
rect 4516 11027 4574 11033
rect 5534 11024 5540 11036
rect 5592 11024 5598 11076
rect 5810 11024 5816 11076
rect 5868 11064 5874 11076
rect 7834 11064 7840 11076
rect 5868 11036 6684 11064
rect 7795 11036 7840 11064
rect 5868 11024 5874 11036
rect 3326 10956 3332 11008
rect 3384 10996 3390 11008
rect 3421 10999 3479 11005
rect 3421 10996 3433 10999
rect 3384 10968 3433 10996
rect 3384 10956 3390 10968
rect 3421 10965 3433 10968
rect 3467 10996 3479 10999
rect 3694 10996 3700 11008
rect 3467 10968 3700 10996
rect 3467 10965 3479 10968
rect 3421 10959 3479 10965
rect 3694 10956 3700 10968
rect 3752 10956 3758 11008
rect 3970 10996 3976 11008
rect 3931 10968 3976 10996
rect 3970 10956 3976 10968
rect 4028 10956 4034 11008
rect 5994 10996 6000 11008
rect 5955 10968 6000 10996
rect 5994 10956 6000 10968
rect 6052 10956 6058 11008
rect 6656 11005 6684 11036
rect 7834 11024 7840 11036
rect 7892 11024 7898 11076
rect 8036 11064 8064 11104
rect 8297 11101 8309 11104
rect 8343 11132 8355 11135
rect 9416 11132 9444 11160
rect 8343 11104 9444 11132
rect 8343 11101 8355 11104
rect 8297 11095 8355 11101
rect 10134 11092 10140 11144
rect 10192 11141 10198 11144
rect 10192 11132 10204 11141
rect 10192 11104 10237 11132
rect 10192 11095 10204 11104
rect 10192 11092 10198 11095
rect 10502 11092 10508 11144
rect 10560 11132 10566 11144
rect 11514 11132 11520 11144
rect 10560 11104 11520 11132
rect 10560 11092 10566 11104
rect 11514 11092 11520 11104
rect 11572 11092 11578 11144
rect 11790 11092 11796 11144
rect 11848 11132 11854 11144
rect 12437 11135 12495 11141
rect 11848 11104 12296 11132
rect 11848 11092 11854 11104
rect 7944 11036 8064 11064
rect 7944 11008 7972 11036
rect 8202 11024 8208 11076
rect 8260 11064 8266 11076
rect 8260 11036 8800 11064
rect 8260 11024 8266 11036
rect 6641 10999 6699 11005
rect 6641 10965 6653 10999
rect 6687 10965 6699 10999
rect 6641 10959 6699 10965
rect 6914 10956 6920 11008
rect 6972 10996 6978 11008
rect 7009 10999 7067 11005
rect 7009 10996 7021 10999
rect 6972 10968 7021 10996
rect 6972 10956 6978 10968
rect 7009 10965 7021 10968
rect 7055 10965 7067 10999
rect 7009 10959 7067 10965
rect 7926 10956 7932 11008
rect 7984 10956 7990 11008
rect 8294 10956 8300 11008
rect 8352 10996 8358 11008
rect 8662 10996 8668 11008
rect 8352 10968 8668 10996
rect 8352 10956 8358 10968
rect 8662 10956 8668 10968
rect 8720 10956 8726 11008
rect 8772 10996 8800 11036
rect 9582 11024 9588 11076
rect 9640 11024 9646 11076
rect 10686 11024 10692 11076
rect 10744 11064 10750 11076
rect 10965 11067 11023 11073
rect 10965 11064 10977 11067
rect 10744 11036 10977 11064
rect 10744 11024 10750 11036
rect 10965 11033 10977 11036
rect 11011 11064 11023 11067
rect 11609 11067 11667 11073
rect 11609 11064 11621 11067
rect 11011 11036 11621 11064
rect 11011 11033 11023 11036
rect 10965 11027 11023 11033
rect 11609 11033 11621 11036
rect 11655 11064 11667 11067
rect 12158 11064 12164 11076
rect 11655 11036 12164 11064
rect 11655 11033 11667 11036
rect 11609 11027 11667 11033
rect 12158 11024 12164 11036
rect 12216 11024 12222 11076
rect 12268 11064 12296 11104
rect 12437 11101 12449 11135
rect 12483 11132 12495 11135
rect 12802 11132 12808 11144
rect 12483 11104 12808 11132
rect 12483 11101 12495 11104
rect 12437 11095 12495 11101
rect 12802 11092 12808 11104
rect 12860 11092 12866 11144
rect 13446 11092 13452 11144
rect 13504 11132 13510 11144
rect 14093 11135 14151 11141
rect 14093 11132 14105 11135
rect 13504 11104 14105 11132
rect 13504 11092 13510 11104
rect 14093 11101 14105 11104
rect 14139 11101 14151 11135
rect 15304 11132 15332 11172
rect 16209 11169 16221 11203
rect 16255 11169 16267 11203
rect 16209 11163 16267 11169
rect 16301 11203 16359 11209
rect 16301 11169 16313 11203
rect 16347 11169 16359 11203
rect 16301 11163 16359 11169
rect 14093 11095 14151 11101
rect 14200 11104 15332 11132
rect 13814 11064 13820 11076
rect 12268 11036 13820 11064
rect 13814 11024 13820 11036
rect 13872 11024 13878 11076
rect 14200 11064 14228 11104
rect 15838 11092 15844 11144
rect 15896 11132 15902 11144
rect 16316 11132 16344 11163
rect 16942 11160 16948 11212
rect 17000 11200 17006 11212
rect 17037 11203 17095 11209
rect 17037 11200 17049 11203
rect 17000 11172 17049 11200
rect 17000 11160 17006 11172
rect 17037 11169 17049 11172
rect 17083 11169 17095 11203
rect 17218 11200 17224 11212
rect 17179 11172 17224 11200
rect 17037 11163 17095 11169
rect 17218 11160 17224 11172
rect 17276 11160 17282 11212
rect 21266 11200 21272 11212
rect 17604 11172 17825 11200
rect 21227 11172 21272 11200
rect 17604 11132 17632 11172
rect 15896 11104 16344 11132
rect 16776 11104 17632 11132
rect 17681 11135 17739 11141
rect 15896 11092 15902 11104
rect 13924 11036 14228 11064
rect 14544 11067 14602 11073
rect 9600 10996 9628 11024
rect 8772 10968 9628 10996
rect 9674 10956 9680 11008
rect 9732 10996 9738 11008
rect 10505 10999 10563 11005
rect 10505 10996 10517 10999
rect 9732 10968 10517 10996
rect 9732 10956 9738 10968
rect 10505 10965 10517 10968
rect 10551 10965 10563 10999
rect 11974 10996 11980 11008
rect 11935 10968 11980 10996
rect 10505 10959 10563 10965
rect 11974 10956 11980 10968
rect 12032 10956 12038 11008
rect 12342 10996 12348 11008
rect 12303 10968 12348 10996
rect 12342 10956 12348 10968
rect 12400 10956 12406 11008
rect 12802 10996 12808 11008
rect 12763 10968 12808 10996
rect 12802 10956 12808 10968
rect 12860 10956 12866 11008
rect 12894 10956 12900 11008
rect 12952 10996 12958 11008
rect 13262 10996 13268 11008
rect 12952 10968 12997 10996
rect 13223 10968 13268 10996
rect 12952 10956 12958 10968
rect 13262 10956 13268 10968
rect 13320 10956 13326 11008
rect 13354 10956 13360 11008
rect 13412 10996 13418 11008
rect 13924 10996 13952 11036
rect 14544 11033 14556 11067
rect 14590 11064 14602 11067
rect 14642 11064 14648 11076
rect 14590 11036 14648 11064
rect 14590 11033 14602 11036
rect 14544 11027 14602 11033
rect 14642 11024 14648 11036
rect 14700 11024 14706 11076
rect 15286 11024 15292 11076
rect 15344 11064 15350 11076
rect 16117 11067 16175 11073
rect 16117 11064 16129 11067
rect 15344 11036 16129 11064
rect 15344 11024 15350 11036
rect 16117 11033 16129 11036
rect 16163 11033 16175 11067
rect 16117 11027 16175 11033
rect 16206 11024 16212 11076
rect 16264 11064 16270 11076
rect 16776 11064 16804 11104
rect 17681 11101 17693 11135
rect 17727 11101 17739 11135
rect 17797 11132 17825 11172
rect 21266 11160 21272 11172
rect 21324 11160 21330 11212
rect 19150 11132 19156 11144
rect 17797 11104 19156 11132
rect 17681 11095 17739 11101
rect 16264 11036 16804 11064
rect 16264 11024 16270 11036
rect 13412 10968 13952 10996
rect 15657 10999 15715 11005
rect 13412 10956 13418 10968
rect 15657 10965 15669 10999
rect 15703 10996 15715 10999
rect 15838 10996 15844 11008
rect 15703 10968 15844 10996
rect 15703 10965 15715 10968
rect 15657 10959 15715 10965
rect 15838 10956 15844 10968
rect 15896 10956 15902 11008
rect 16942 10996 16948 11008
rect 16903 10968 16948 10996
rect 16942 10956 16948 10968
rect 17000 10956 17006 11008
rect 17696 10996 17724 11095
rect 19150 11092 19156 11104
rect 19208 11092 19214 11144
rect 19245 11135 19303 11141
rect 19245 11101 19257 11135
rect 19291 11132 19303 11135
rect 20898 11132 20904 11144
rect 19291 11104 20904 11132
rect 19291 11101 19303 11104
rect 19245 11095 19303 11101
rect 20898 11092 20904 11104
rect 20956 11092 20962 11144
rect 17948 11067 18006 11073
rect 17948 11033 17960 11067
rect 17994 11064 18006 11067
rect 18690 11064 18696 11076
rect 17994 11036 18696 11064
rect 17994 11033 18006 11036
rect 17948 11027 18006 11033
rect 18690 11024 18696 11036
rect 18748 11024 18754 11076
rect 19512 11067 19570 11073
rect 19512 11033 19524 11067
rect 19558 11064 19570 11067
rect 19886 11064 19892 11076
rect 19558 11036 19892 11064
rect 19558 11033 19570 11036
rect 19512 11027 19570 11033
rect 19886 11024 19892 11036
rect 19944 11024 19950 11076
rect 21082 11064 21088 11076
rect 21043 11036 21088 11064
rect 21082 11024 21088 11036
rect 21140 11024 21146 11076
rect 21177 11067 21235 11073
rect 21177 11033 21189 11067
rect 21223 11064 21235 11067
rect 21358 11064 21364 11076
rect 21223 11036 21364 11064
rect 21223 11033 21235 11036
rect 21177 11027 21235 11033
rect 21358 11024 21364 11036
rect 21416 11024 21422 11076
rect 18046 10996 18052 11008
rect 17696 10968 18052 10996
rect 18046 10956 18052 10968
rect 18104 10996 18110 11008
rect 18598 10996 18604 11008
rect 18104 10968 18604 10996
rect 18104 10956 18110 10968
rect 18598 10956 18604 10968
rect 18656 10956 18662 11008
rect 19794 10956 19800 11008
rect 19852 10996 19858 11008
rect 20625 10999 20683 11005
rect 20625 10996 20637 10999
rect 19852 10968 20637 10996
rect 19852 10956 19858 10968
rect 20625 10965 20637 10968
rect 20671 10965 20683 10999
rect 20625 10959 20683 10965
rect 20717 10999 20775 11005
rect 20717 10965 20729 10999
rect 20763 10996 20775 10999
rect 20806 10996 20812 11008
rect 20763 10968 20812 10996
rect 20763 10965 20775 10968
rect 20717 10959 20775 10965
rect 20806 10956 20812 10968
rect 20864 10956 20870 11008
rect 1104 10906 22056 10928
rect 1104 10854 6148 10906
rect 6200 10854 6212 10906
rect 6264 10854 6276 10906
rect 6328 10854 6340 10906
rect 6392 10854 6404 10906
rect 6456 10854 11346 10906
rect 11398 10854 11410 10906
rect 11462 10854 11474 10906
rect 11526 10854 11538 10906
rect 11590 10854 11602 10906
rect 11654 10854 16544 10906
rect 16596 10854 16608 10906
rect 16660 10854 16672 10906
rect 16724 10854 16736 10906
rect 16788 10854 16800 10906
rect 16852 10854 21742 10906
rect 21794 10854 21806 10906
rect 21858 10854 21870 10906
rect 21922 10854 21934 10906
rect 21986 10854 21998 10906
rect 22050 10854 22056 10906
rect 1104 10832 22056 10854
rect 2958 10752 2964 10804
rect 3016 10792 3022 10804
rect 3145 10795 3203 10801
rect 3145 10792 3157 10795
rect 3016 10764 3157 10792
rect 3016 10752 3022 10764
rect 3145 10761 3157 10764
rect 3191 10761 3203 10795
rect 3145 10755 3203 10761
rect 5368 10764 5957 10792
rect 3160 10724 3188 10755
rect 3482 10727 3540 10733
rect 3482 10724 3494 10727
rect 1596 10696 2176 10724
rect 3160 10696 3494 10724
rect 1486 10656 1492 10668
rect 1399 10628 1492 10656
rect 1486 10616 1492 10628
rect 1544 10616 1550 10668
rect 1504 10520 1532 10616
rect 1596 10588 1624 10696
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10656 1731 10659
rect 1854 10656 1860 10668
rect 1719 10628 1860 10656
rect 1719 10625 1731 10628
rect 1673 10619 1731 10625
rect 1854 10616 1860 10628
rect 1912 10616 1918 10668
rect 2038 10665 2044 10668
rect 2032 10656 2044 10665
rect 1999 10628 2044 10656
rect 2032 10619 2044 10628
rect 2038 10616 2044 10619
rect 2096 10616 2102 10668
rect 2148 10656 2176 10696
rect 3482 10693 3494 10696
rect 3528 10693 3540 10727
rect 3482 10687 3540 10693
rect 3237 10659 3295 10665
rect 3237 10656 3249 10659
rect 2148 10628 3249 10656
rect 3237 10625 3249 10628
rect 3283 10656 3295 10659
rect 3970 10656 3976 10668
rect 3283 10628 3976 10656
rect 3283 10625 3295 10628
rect 3237 10619 3295 10625
rect 3970 10616 3976 10628
rect 4028 10616 4034 10668
rect 5368 10665 5396 10764
rect 5718 10724 5724 10736
rect 5460 10696 5724 10724
rect 5353 10659 5411 10665
rect 4540 10628 4936 10656
rect 1762 10588 1768 10600
rect 1596 10560 1768 10588
rect 1762 10548 1768 10560
rect 1820 10548 1826 10600
rect 1504 10492 1624 10520
rect 1596 10452 1624 10492
rect 4540 10452 4568 10628
rect 4798 10588 4804 10600
rect 4759 10560 4804 10588
rect 4798 10548 4804 10560
rect 4856 10548 4862 10600
rect 4908 10588 4936 10628
rect 5353 10625 5365 10659
rect 5399 10625 5411 10659
rect 5353 10619 5411 10625
rect 5460 10588 5488 10696
rect 5718 10684 5724 10696
rect 5776 10684 5782 10736
rect 5929 10724 5957 10764
rect 5994 10752 6000 10804
rect 6052 10792 6058 10804
rect 6181 10795 6239 10801
rect 6181 10792 6193 10795
rect 6052 10764 6193 10792
rect 6052 10752 6058 10764
rect 6181 10761 6193 10764
rect 6227 10761 6239 10795
rect 6181 10755 6239 10761
rect 6365 10795 6423 10801
rect 6365 10761 6377 10795
rect 6411 10792 6423 10795
rect 6546 10792 6552 10804
rect 6411 10764 6552 10792
rect 6411 10761 6423 10764
rect 6365 10755 6423 10761
rect 6546 10752 6552 10764
rect 6604 10752 6610 10804
rect 7098 10752 7104 10804
rect 7156 10792 7162 10804
rect 9674 10792 9680 10804
rect 7156 10764 9536 10792
rect 9635 10764 9680 10792
rect 7156 10752 7162 10764
rect 7834 10724 7840 10736
rect 5929 10696 7840 10724
rect 7834 10684 7840 10696
rect 7892 10724 7898 10736
rect 7892 10696 8156 10724
rect 7892 10684 7898 10696
rect 5810 10656 5816 10668
rect 5771 10628 5816 10656
rect 5810 10616 5816 10628
rect 5868 10616 5874 10668
rect 7478 10659 7536 10665
rect 7478 10656 7490 10659
rect 6748 10628 7490 10656
rect 4908 10560 5488 10588
rect 5534 10548 5540 10600
rect 5592 10588 5598 10600
rect 5721 10591 5779 10597
rect 5592 10560 5637 10588
rect 5592 10548 5598 10560
rect 5721 10557 5733 10591
rect 5767 10588 5779 10591
rect 6362 10588 6368 10600
rect 5767 10560 6368 10588
rect 5767 10557 5779 10560
rect 5721 10551 5779 10557
rect 6362 10548 6368 10560
rect 6420 10548 6426 10600
rect 4617 10523 4675 10529
rect 4617 10489 4629 10523
rect 4663 10520 4675 10523
rect 6748 10520 6776 10628
rect 7478 10625 7490 10628
rect 7524 10656 7536 10659
rect 8018 10656 8024 10668
rect 7524 10628 8024 10656
rect 7524 10625 7536 10628
rect 7478 10619 7536 10625
rect 8018 10616 8024 10628
rect 8076 10616 8082 10668
rect 8128 10656 8156 10696
rect 8294 10684 8300 10736
rect 8352 10724 8358 10736
rect 8950 10727 9008 10733
rect 8950 10724 8962 10727
rect 8352 10696 8962 10724
rect 8352 10684 8358 10696
rect 8950 10693 8962 10696
rect 8996 10724 9008 10727
rect 9508 10724 9536 10764
rect 9674 10752 9680 10764
rect 9732 10752 9738 10804
rect 10045 10795 10103 10801
rect 10045 10761 10057 10795
rect 10091 10792 10103 10795
rect 10505 10795 10563 10801
rect 10505 10792 10517 10795
rect 10091 10764 10517 10792
rect 10091 10761 10103 10764
rect 10045 10755 10103 10761
rect 10505 10761 10517 10764
rect 10551 10761 10563 10795
rect 10505 10755 10563 10761
rect 10686 10752 10692 10804
rect 10744 10792 10750 10804
rect 10965 10795 11023 10801
rect 10965 10792 10977 10795
rect 10744 10764 10977 10792
rect 10744 10752 10750 10764
rect 10965 10761 10977 10764
rect 11011 10761 11023 10795
rect 10965 10755 11023 10761
rect 11885 10795 11943 10801
rect 11885 10761 11897 10795
rect 11931 10792 11943 10795
rect 11974 10792 11980 10804
rect 11931 10764 11980 10792
rect 11931 10761 11943 10764
rect 11885 10755 11943 10761
rect 11974 10752 11980 10764
rect 12032 10752 12038 10804
rect 12345 10795 12403 10801
rect 12345 10761 12357 10795
rect 12391 10792 12403 10795
rect 13262 10792 13268 10804
rect 12391 10764 13268 10792
rect 12391 10761 12403 10764
rect 12345 10755 12403 10761
rect 13262 10752 13268 10764
rect 13320 10752 13326 10804
rect 13722 10792 13728 10804
rect 13464 10764 13728 10792
rect 13464 10724 13492 10764
rect 13722 10752 13728 10764
rect 13780 10752 13786 10804
rect 14093 10795 14151 10801
rect 14093 10761 14105 10795
rect 14139 10792 14151 10795
rect 14458 10792 14464 10804
rect 14139 10764 14464 10792
rect 14139 10761 14151 10764
rect 14093 10755 14151 10761
rect 14458 10752 14464 10764
rect 14516 10752 14522 10804
rect 14921 10795 14979 10801
rect 14921 10792 14933 10795
rect 14559 10764 14933 10792
rect 8996 10696 9444 10724
rect 9508 10696 13492 10724
rect 8996 10693 9008 10696
rect 8950 10687 9008 10693
rect 9217 10659 9275 10665
rect 9217 10656 9229 10659
rect 8128 10628 9229 10656
rect 9217 10625 9229 10628
rect 9263 10625 9275 10659
rect 9217 10619 9275 10625
rect 7745 10591 7803 10597
rect 7745 10557 7757 10591
rect 7791 10588 7803 10591
rect 7834 10588 7840 10600
rect 7791 10560 7840 10588
rect 7791 10557 7803 10560
rect 7745 10551 7803 10557
rect 7834 10548 7840 10560
rect 7892 10548 7898 10600
rect 9416 10597 9444 10696
rect 13538 10684 13544 10736
rect 13596 10733 13602 10736
rect 13596 10724 13608 10733
rect 14274 10724 14280 10736
rect 13596 10696 13641 10724
rect 13924 10696 14280 10724
rect 13596 10687 13608 10696
rect 13596 10684 13602 10687
rect 10870 10656 10876 10668
rect 9968 10628 10876 10656
rect 9968 10600 9996 10628
rect 10870 10616 10876 10628
rect 10928 10616 10934 10668
rect 11238 10656 11244 10668
rect 11199 10628 11244 10656
rect 11238 10616 11244 10628
rect 11296 10616 11302 10668
rect 11974 10656 11980 10668
rect 11935 10628 11980 10656
rect 11974 10616 11980 10628
rect 12032 10616 12038 10668
rect 13924 10665 13952 10696
rect 14274 10684 14280 10696
rect 14332 10684 14338 10736
rect 14559 10724 14587 10764
rect 14921 10761 14933 10764
rect 14967 10761 14979 10795
rect 15286 10792 15292 10804
rect 15247 10764 15292 10792
rect 14921 10755 14979 10761
rect 15286 10752 15292 10764
rect 15344 10752 15350 10804
rect 16114 10792 16120 10804
rect 16075 10764 16120 10792
rect 16114 10752 16120 10764
rect 16172 10752 16178 10804
rect 16669 10795 16727 10801
rect 16669 10761 16681 10795
rect 16715 10761 16727 10795
rect 16669 10755 16727 10761
rect 14384 10696 14587 10724
rect 13817 10659 13875 10665
rect 13817 10625 13829 10659
rect 13863 10656 13875 10659
rect 13909 10659 13967 10665
rect 13909 10656 13921 10659
rect 13863 10628 13921 10656
rect 13863 10625 13875 10628
rect 13817 10619 13875 10625
rect 13909 10625 13921 10628
rect 13955 10625 13967 10659
rect 13909 10619 13967 10625
rect 14182 10616 14188 10668
rect 14240 10656 14246 10668
rect 14384 10665 14412 10696
rect 14642 10684 14648 10736
rect 14700 10724 14706 10736
rect 15102 10724 15108 10736
rect 14700 10696 15108 10724
rect 14700 10684 14706 10696
rect 15102 10684 15108 10696
rect 15160 10684 15166 10736
rect 15749 10727 15807 10733
rect 15749 10693 15761 10727
rect 15795 10724 15807 10727
rect 16684 10724 16712 10755
rect 16942 10752 16948 10804
rect 17000 10792 17006 10804
rect 17497 10795 17555 10801
rect 17497 10792 17509 10795
rect 17000 10764 17509 10792
rect 17000 10752 17006 10764
rect 17497 10761 17509 10764
rect 17543 10761 17555 10795
rect 17862 10792 17868 10804
rect 17497 10755 17555 10761
rect 17696 10764 17868 10792
rect 15795 10696 16712 10724
rect 15795 10693 15807 10696
rect 15749 10687 15807 10693
rect 16758 10684 16764 10736
rect 16816 10724 16822 10736
rect 17126 10724 17132 10736
rect 16816 10696 17132 10724
rect 16816 10684 16822 10696
rect 17126 10684 17132 10696
rect 17184 10684 17190 10736
rect 14369 10659 14427 10665
rect 14369 10656 14381 10659
rect 14240 10628 14381 10656
rect 14240 10616 14246 10628
rect 14369 10625 14381 10628
rect 14415 10625 14427 10659
rect 15838 10656 15844 10668
rect 14369 10619 14427 10625
rect 15488 10628 15844 10656
rect 9401 10591 9459 10597
rect 9401 10557 9413 10591
rect 9447 10557 9459 10591
rect 9401 10551 9459 10557
rect 9585 10591 9643 10597
rect 9585 10557 9597 10591
rect 9631 10588 9643 10591
rect 9674 10588 9680 10600
rect 9631 10560 9680 10588
rect 9631 10557 9643 10560
rect 9585 10551 9643 10557
rect 9674 10548 9680 10560
rect 9732 10588 9738 10600
rect 9950 10588 9956 10600
rect 9732 10560 9956 10588
rect 9732 10548 9738 10560
rect 9950 10548 9956 10560
rect 10008 10548 10014 10600
rect 10134 10548 10140 10600
rect 10192 10548 10198 10600
rect 10594 10588 10600 10600
rect 10555 10560 10600 10588
rect 10594 10548 10600 10560
rect 10652 10548 10658 10600
rect 10689 10591 10747 10597
rect 10689 10557 10701 10591
rect 10735 10557 10747 10591
rect 11698 10588 11704 10600
rect 11659 10560 11704 10588
rect 10689 10551 10747 10557
rect 10152 10520 10180 10548
rect 10704 10520 10732 10551
rect 11698 10548 11704 10560
rect 11756 10548 11762 10600
rect 14642 10588 14648 10600
rect 14603 10560 14648 10588
rect 14642 10548 14648 10560
rect 14700 10548 14706 10600
rect 14826 10588 14832 10600
rect 14787 10560 14832 10588
rect 14826 10548 14832 10560
rect 14884 10548 14890 10600
rect 15488 10597 15516 10628
rect 15838 10616 15844 10628
rect 15896 10616 15902 10668
rect 16393 10659 16451 10665
rect 16393 10625 16405 10659
rect 16439 10656 16451 10659
rect 17037 10659 17095 10665
rect 17037 10656 17049 10659
rect 16439 10628 17049 10656
rect 16439 10625 16451 10628
rect 16393 10619 16451 10625
rect 17037 10625 17049 10628
rect 17083 10625 17095 10659
rect 17037 10619 17095 10625
rect 15473 10591 15531 10597
rect 15473 10557 15485 10591
rect 15519 10557 15531 10591
rect 15654 10588 15660 10600
rect 15615 10560 15660 10588
rect 15473 10551 15531 10557
rect 15654 10548 15660 10560
rect 15712 10548 15718 10600
rect 17218 10588 17224 10600
rect 17179 10560 17224 10588
rect 17218 10548 17224 10560
rect 17276 10548 17282 10600
rect 17696 10588 17724 10764
rect 17862 10752 17868 10764
rect 17920 10792 17926 10804
rect 17957 10795 18015 10801
rect 17957 10792 17969 10795
rect 17920 10764 17969 10792
rect 17920 10752 17926 10764
rect 17957 10761 17969 10764
rect 18003 10761 18015 10795
rect 17957 10755 18015 10761
rect 18782 10752 18788 10804
rect 18840 10792 18846 10804
rect 19153 10795 19211 10801
rect 19153 10792 19165 10795
rect 18840 10764 19165 10792
rect 18840 10752 18846 10764
rect 19153 10761 19165 10764
rect 19199 10761 19211 10795
rect 19153 10755 19211 10761
rect 19610 10752 19616 10804
rect 19668 10792 19674 10804
rect 19981 10795 20039 10801
rect 19981 10792 19993 10795
rect 19668 10764 19993 10792
rect 19668 10752 19674 10764
rect 19981 10761 19993 10764
rect 20027 10761 20039 10795
rect 19981 10755 20039 10761
rect 17770 10684 17776 10736
rect 17828 10724 17834 10736
rect 20714 10724 20720 10736
rect 17828 10696 20720 10724
rect 17828 10684 17834 10696
rect 20714 10684 20720 10696
rect 20772 10684 20778 10736
rect 21174 10684 21180 10736
rect 21232 10724 21238 10736
rect 21278 10727 21336 10733
rect 21278 10724 21290 10727
rect 21232 10696 21290 10724
rect 21232 10684 21238 10696
rect 21278 10693 21290 10696
rect 21324 10693 21336 10727
rect 21278 10687 21336 10693
rect 17865 10659 17923 10665
rect 17865 10625 17877 10659
rect 17911 10656 17923 10659
rect 18322 10656 18328 10668
rect 17911 10628 18328 10656
rect 17911 10625 17923 10628
rect 17865 10619 17923 10625
rect 18322 10616 18328 10628
rect 18380 10616 18386 10668
rect 18693 10659 18751 10665
rect 18693 10625 18705 10659
rect 18739 10656 18751 10659
rect 18782 10656 18788 10668
rect 18739 10628 18788 10656
rect 18739 10625 18751 10628
rect 18693 10619 18751 10625
rect 18782 10616 18788 10628
rect 18840 10616 18846 10668
rect 19518 10656 19524 10668
rect 19479 10628 19524 10656
rect 19518 10616 19524 10628
rect 19576 10616 19582 10668
rect 20898 10616 20904 10668
rect 20956 10656 20962 10668
rect 21545 10659 21603 10665
rect 21545 10656 21557 10659
rect 20956 10628 21557 10656
rect 20956 10616 20962 10628
rect 21545 10625 21557 10628
rect 21591 10625 21603 10659
rect 21545 10619 21603 10625
rect 17770 10588 17776 10600
rect 17696 10560 17776 10588
rect 17770 10548 17776 10560
rect 17828 10548 17834 10600
rect 18141 10591 18199 10597
rect 18141 10557 18153 10591
rect 18187 10588 18199 10591
rect 18230 10588 18236 10600
rect 18187 10560 18236 10588
rect 18187 10557 18199 10560
rect 18141 10551 18199 10557
rect 18230 10548 18236 10560
rect 18288 10548 18294 10600
rect 18506 10588 18512 10600
rect 18467 10560 18512 10588
rect 18506 10548 18512 10560
rect 18564 10548 18570 10600
rect 18601 10591 18659 10597
rect 18601 10557 18613 10591
rect 18647 10557 18659 10591
rect 19610 10588 19616 10600
rect 19571 10560 19616 10588
rect 18601 10551 18659 10557
rect 4663 10492 6776 10520
rect 9416 10492 10732 10520
rect 4663 10489 4675 10492
rect 4617 10483 4675 10489
rect 5166 10452 5172 10464
rect 1596 10424 4568 10452
rect 5127 10424 5172 10452
rect 5166 10412 5172 10424
rect 5224 10412 5230 10464
rect 5534 10412 5540 10464
rect 5592 10452 5598 10464
rect 6546 10452 6552 10464
rect 5592 10424 6552 10452
rect 5592 10412 5598 10424
rect 6546 10412 6552 10424
rect 6604 10412 6610 10464
rect 7834 10452 7840 10464
rect 7795 10424 7840 10452
rect 7834 10412 7840 10424
rect 7892 10452 7898 10464
rect 9416 10452 9444 10492
rect 13814 10480 13820 10532
rect 13872 10520 13878 10532
rect 18616 10520 18644 10551
rect 19610 10548 19616 10560
rect 19668 10548 19674 10600
rect 19794 10588 19800 10600
rect 19755 10560 19800 10588
rect 19794 10548 19800 10560
rect 19852 10548 19858 10600
rect 20165 10523 20223 10529
rect 20165 10520 20177 10523
rect 13872 10492 18644 10520
rect 18708 10492 20177 10520
rect 13872 10480 13878 10492
rect 7892 10424 9444 10452
rect 7892 10412 7898 10424
rect 9490 10412 9496 10464
rect 9548 10452 9554 10464
rect 10137 10455 10195 10461
rect 10137 10452 10149 10455
rect 9548 10424 10149 10452
rect 9548 10412 9554 10424
rect 10137 10421 10149 10424
rect 10183 10421 10195 10455
rect 10137 10415 10195 10421
rect 12434 10412 12440 10464
rect 12492 10452 12498 10464
rect 14277 10455 14335 10461
rect 12492 10424 12537 10452
rect 12492 10412 12498 10424
rect 14277 10421 14289 10455
rect 14323 10452 14335 10455
rect 18138 10452 18144 10464
rect 14323 10424 18144 10452
rect 14323 10421 14335 10424
rect 14277 10415 14335 10421
rect 18138 10412 18144 10424
rect 18196 10412 18202 10464
rect 18598 10412 18604 10464
rect 18656 10452 18662 10464
rect 18708 10452 18736 10492
rect 20165 10489 20177 10492
rect 20211 10489 20223 10523
rect 20165 10483 20223 10489
rect 18656 10424 18736 10452
rect 19061 10455 19119 10461
rect 18656 10412 18662 10424
rect 19061 10421 19073 10455
rect 19107 10452 19119 10455
rect 19702 10452 19708 10464
rect 19107 10424 19708 10452
rect 19107 10421 19119 10424
rect 19061 10415 19119 10421
rect 19702 10412 19708 10424
rect 19760 10412 19766 10464
rect 1104 10362 21896 10384
rect 1104 10310 3549 10362
rect 3601 10310 3613 10362
rect 3665 10310 3677 10362
rect 3729 10310 3741 10362
rect 3793 10310 3805 10362
rect 3857 10310 8747 10362
rect 8799 10310 8811 10362
rect 8863 10310 8875 10362
rect 8927 10310 8939 10362
rect 8991 10310 9003 10362
rect 9055 10310 13945 10362
rect 13997 10310 14009 10362
rect 14061 10310 14073 10362
rect 14125 10310 14137 10362
rect 14189 10310 14201 10362
rect 14253 10310 19143 10362
rect 19195 10310 19207 10362
rect 19259 10310 19271 10362
rect 19323 10310 19335 10362
rect 19387 10310 19399 10362
rect 19451 10310 21896 10362
rect 1104 10288 21896 10310
rect 750 10208 756 10260
rect 808 10248 814 10260
rect 934 10248 940 10260
rect 808 10220 940 10248
rect 808 10208 814 10220
rect 934 10208 940 10220
rect 992 10208 998 10260
rect 2130 10208 2136 10260
rect 2188 10248 2194 10260
rect 3421 10251 3479 10257
rect 3421 10248 3433 10251
rect 2188 10220 3433 10248
rect 2188 10208 2194 10220
rect 3421 10217 3433 10220
rect 3467 10217 3479 10251
rect 3421 10211 3479 10217
rect 3602 10208 3608 10260
rect 3660 10248 3666 10260
rect 4614 10248 4620 10260
rect 3660 10220 4620 10248
rect 3660 10208 3666 10220
rect 4614 10208 4620 10220
rect 4672 10208 4678 10260
rect 5169 10251 5227 10257
rect 5169 10217 5181 10251
rect 5215 10248 5227 10251
rect 5350 10248 5356 10260
rect 5215 10220 5356 10248
rect 5215 10217 5227 10220
rect 5169 10211 5227 10217
rect 5350 10208 5356 10220
rect 5408 10208 5414 10260
rect 6362 10248 6368 10260
rect 6275 10220 6368 10248
rect 6362 10208 6368 10220
rect 6420 10248 6426 10260
rect 8202 10248 8208 10260
rect 6420 10220 8208 10248
rect 6420 10208 6426 10220
rect 8202 10208 8208 10220
rect 8260 10208 8266 10260
rect 8757 10251 8815 10257
rect 8757 10217 8769 10251
rect 8803 10248 8815 10251
rect 10594 10248 10600 10260
rect 8803 10220 10600 10248
rect 8803 10217 8815 10220
rect 8757 10211 8815 10217
rect 10594 10208 10600 10220
rect 10652 10208 10658 10260
rect 11885 10251 11943 10257
rect 11885 10217 11897 10251
rect 11931 10248 11943 10251
rect 13814 10248 13820 10260
rect 11931 10220 13820 10248
rect 11931 10217 11943 10220
rect 11885 10211 11943 10217
rect 13814 10208 13820 10220
rect 13872 10208 13878 10260
rect 14274 10248 14280 10260
rect 14108 10220 14280 10248
rect 1673 10183 1731 10189
rect 1673 10149 1685 10183
rect 1719 10180 1731 10183
rect 1854 10180 1860 10192
rect 1719 10152 1860 10180
rect 1719 10149 1731 10152
rect 1673 10143 1731 10149
rect 1854 10140 1860 10152
rect 1912 10140 1918 10192
rect 3329 10183 3387 10189
rect 3329 10149 3341 10183
rect 3375 10180 3387 10183
rect 4338 10180 4344 10192
rect 3375 10152 4344 10180
rect 3375 10149 3387 10152
rect 3329 10143 3387 10149
rect 1762 10072 1768 10124
rect 1820 10112 1826 10124
rect 1949 10115 2007 10121
rect 1949 10112 1961 10115
rect 1820 10084 1961 10112
rect 1820 10072 1826 10084
rect 1949 10081 1961 10084
rect 1995 10081 2007 10115
rect 1949 10075 2007 10081
rect 566 10004 572 10056
rect 624 10044 630 10056
rect 1026 10044 1032 10056
rect 624 10016 1032 10044
rect 624 10004 630 10016
rect 1026 10004 1032 10016
rect 1084 10004 1090 10056
rect 1486 10044 1492 10056
rect 1399 10016 1492 10044
rect 1486 10004 1492 10016
rect 1544 10044 1550 10056
rect 3234 10044 3240 10056
rect 1544 10016 3240 10044
rect 1544 10004 1550 10016
rect 3234 10004 3240 10016
rect 3292 10004 3298 10056
rect 2222 9985 2228 9988
rect 2216 9939 2228 9985
rect 2280 9976 2286 9988
rect 2280 9948 2316 9976
rect 2222 9936 2228 9939
rect 2280 9936 2286 9948
rect 2774 9936 2780 9988
rect 2832 9976 2838 9988
rect 3050 9976 3056 9988
rect 2832 9948 3056 9976
rect 2832 9936 2838 9948
rect 3050 9936 3056 9948
rect 3108 9936 3114 9988
rect 1854 9908 1860 9920
rect 1815 9880 1860 9908
rect 1854 9868 1860 9880
rect 1912 9868 1918 9920
rect 1946 9868 1952 9920
rect 2004 9908 2010 9920
rect 3344 9908 3372 10143
rect 4338 10140 4344 10152
rect 4396 10140 4402 10192
rect 5261 10183 5319 10189
rect 5261 10180 5273 10183
rect 4448 10152 5273 10180
rect 3510 10072 3516 10124
rect 3568 10112 3574 10124
rect 3568 10084 3832 10112
rect 3568 10072 3574 10084
rect 3602 10044 3608 10056
rect 3563 10016 3608 10044
rect 3602 10004 3608 10016
rect 3660 10004 3666 10056
rect 3804 10053 3832 10084
rect 3878 10072 3884 10124
rect 3936 10112 3942 10124
rect 4448 10112 4476 10152
rect 5261 10149 5273 10152
rect 5307 10149 5319 10183
rect 5261 10143 5319 10149
rect 5718 10140 5724 10192
rect 5776 10180 5782 10192
rect 6181 10183 6239 10189
rect 6181 10180 6193 10183
rect 5776 10152 6193 10180
rect 5776 10140 5782 10152
rect 6181 10149 6193 10152
rect 6227 10180 6239 10183
rect 7098 10180 7104 10192
rect 6227 10152 7104 10180
rect 6227 10149 6239 10152
rect 6181 10143 6239 10149
rect 7098 10140 7104 10152
rect 7156 10140 7162 10192
rect 7282 10140 7288 10192
rect 7340 10180 7346 10192
rect 9950 10180 9956 10192
rect 7340 10152 9812 10180
rect 9911 10152 9956 10180
rect 7340 10140 7346 10152
rect 3936 10084 4476 10112
rect 4617 10115 4675 10121
rect 3936 10072 3942 10084
rect 4617 10081 4629 10115
rect 4663 10112 4675 10115
rect 5626 10112 5632 10124
rect 4663 10084 5632 10112
rect 4663 10081 4675 10084
rect 4617 10075 4675 10081
rect 5626 10072 5632 10084
rect 5684 10072 5690 10124
rect 5813 10115 5871 10121
rect 5813 10081 5825 10115
rect 5859 10081 5871 10115
rect 5813 10075 5871 10081
rect 3789 10047 3847 10053
rect 3789 10013 3801 10047
rect 3835 10013 3847 10047
rect 3789 10007 3847 10013
rect 4065 10047 4123 10053
rect 4065 10013 4077 10047
rect 4111 10013 4123 10047
rect 4798 10044 4804 10056
rect 4759 10016 4804 10044
rect 4065 10007 4123 10013
rect 4080 9976 4108 10007
rect 4798 10004 4804 10016
rect 4856 10004 4862 10056
rect 5350 10004 5356 10056
rect 5408 10044 5414 10056
rect 5828 10044 5856 10075
rect 5902 10072 5908 10124
rect 5960 10072 5966 10124
rect 6546 10112 6552 10124
rect 6507 10084 6552 10112
rect 6546 10072 6552 10084
rect 6604 10112 6610 10124
rect 6914 10112 6920 10124
rect 6604 10084 6920 10112
rect 6604 10072 6610 10084
rect 6914 10072 6920 10084
rect 6972 10072 6978 10124
rect 7377 10115 7435 10121
rect 7377 10081 7389 10115
rect 7423 10112 7435 10115
rect 7834 10112 7840 10124
rect 7423 10084 7840 10112
rect 7423 10081 7435 10084
rect 7377 10075 7435 10081
rect 7834 10072 7840 10084
rect 7892 10072 7898 10124
rect 8205 10115 8263 10121
rect 8205 10081 8217 10115
rect 8251 10112 8263 10115
rect 8294 10112 8300 10124
rect 8251 10084 8300 10112
rect 8251 10081 8263 10084
rect 8205 10075 8263 10081
rect 8294 10072 8300 10084
rect 8352 10072 8358 10124
rect 8846 10072 8852 10124
rect 8904 10112 8910 10124
rect 8904 10084 9343 10112
rect 8904 10072 8910 10084
rect 5408 10016 5856 10044
rect 5408 10004 5414 10016
rect 5534 9976 5540 9988
rect 3620 9948 4108 9976
rect 4264 9948 5540 9976
rect 3620 9920 3648 9948
rect 2004 9880 3372 9908
rect 2004 9868 2010 9880
rect 3602 9868 3608 9920
rect 3660 9868 3666 9920
rect 3973 9911 4031 9917
rect 3973 9877 3985 9911
rect 4019 9908 4031 9911
rect 4154 9908 4160 9920
rect 4019 9880 4160 9908
rect 4019 9877 4031 9880
rect 3973 9871 4031 9877
rect 4154 9868 4160 9880
rect 4212 9868 4218 9920
rect 4264 9917 4292 9948
rect 5534 9936 5540 9948
rect 5592 9976 5598 9988
rect 5810 9976 5816 9988
rect 5592 9948 5816 9976
rect 5592 9936 5598 9948
rect 5810 9936 5816 9948
rect 5868 9936 5874 9988
rect 4249 9911 4307 9917
rect 4249 9877 4261 9911
rect 4295 9877 4307 9911
rect 4249 9871 4307 9877
rect 4706 9868 4712 9920
rect 4764 9908 4770 9920
rect 5626 9908 5632 9920
rect 4764 9880 4809 9908
rect 5587 9880 5632 9908
rect 4764 9868 4770 9880
rect 5626 9868 5632 9880
rect 5684 9868 5690 9920
rect 5721 9911 5779 9917
rect 5721 9877 5733 9911
rect 5767 9908 5779 9911
rect 5920 9908 5948 10072
rect 6454 10004 6460 10056
rect 6512 10044 6518 10056
rect 6512 10016 9260 10044
rect 6512 10004 6518 10016
rect 5994 9936 6000 9988
rect 6052 9976 6058 9988
rect 7101 9979 7159 9985
rect 7101 9976 7113 9979
rect 6052 9948 7113 9976
rect 6052 9936 6058 9948
rect 7101 9945 7113 9948
rect 7147 9976 7159 9979
rect 7834 9976 7840 9988
rect 7147 9948 7840 9976
rect 7147 9945 7159 9948
rect 7101 9939 7159 9945
rect 7834 9936 7840 9948
rect 7892 9936 7898 9988
rect 8846 9976 8852 9988
rect 7944 9948 8852 9976
rect 6454 9908 6460 9920
rect 5767 9880 6460 9908
rect 5767 9877 5779 9880
rect 5721 9871 5779 9877
rect 6454 9868 6460 9880
rect 6512 9868 6518 9920
rect 6638 9908 6644 9920
rect 6599 9880 6644 9908
rect 6638 9868 6644 9880
rect 6696 9868 6702 9920
rect 6914 9908 6920 9920
rect 6875 9880 6920 9908
rect 6914 9868 6920 9880
rect 6972 9868 6978 9920
rect 7466 9908 7472 9920
rect 7427 9880 7472 9908
rect 7466 9868 7472 9880
rect 7524 9868 7530 9920
rect 7558 9868 7564 9920
rect 7616 9908 7622 9920
rect 7944 9917 7972 9948
rect 8846 9936 8852 9948
rect 8904 9936 8910 9988
rect 7929 9911 7987 9917
rect 7616 9880 7661 9908
rect 7616 9868 7622 9880
rect 7929 9877 7941 9911
rect 7975 9877 7987 9911
rect 7929 9871 7987 9877
rect 8202 9868 8208 9920
rect 8260 9908 8266 9920
rect 8297 9911 8355 9917
rect 8297 9908 8309 9911
rect 8260 9880 8309 9908
rect 8260 9868 8266 9880
rect 8297 9877 8309 9880
rect 8343 9877 8355 9911
rect 8297 9871 8355 9877
rect 8389 9911 8447 9917
rect 8389 9877 8401 9911
rect 8435 9908 8447 9911
rect 8662 9908 8668 9920
rect 8435 9880 8668 9908
rect 8435 9877 8447 9880
rect 8389 9871 8447 9877
rect 8662 9868 8668 9880
rect 8720 9868 8726 9920
rect 8938 9908 8944 9920
rect 8899 9880 8944 9908
rect 8938 9868 8944 9880
rect 8996 9868 9002 9920
rect 9122 9908 9128 9920
rect 9083 9880 9128 9908
rect 9122 9868 9128 9880
rect 9180 9868 9186 9920
rect 9232 9908 9260 10016
rect 9315 9976 9343 10084
rect 9582 10072 9588 10124
rect 9640 10112 9646 10124
rect 9677 10115 9735 10121
rect 9677 10112 9689 10115
rect 9640 10084 9689 10112
rect 9640 10072 9646 10084
rect 9677 10081 9689 10084
rect 9723 10081 9735 10115
rect 9677 10075 9735 10081
rect 9490 10044 9496 10056
rect 9451 10016 9496 10044
rect 9490 10004 9496 10016
rect 9548 10004 9554 10056
rect 9784 10044 9812 10152
rect 9950 10140 9956 10152
rect 10008 10140 10014 10192
rect 13998 10180 14004 10192
rect 10520 10152 14004 10180
rect 10520 10121 10548 10152
rect 13998 10140 14004 10152
rect 14056 10140 14062 10192
rect 10505 10115 10563 10121
rect 10505 10081 10517 10115
rect 10551 10081 10563 10115
rect 10505 10075 10563 10081
rect 11333 10115 11391 10121
rect 11333 10081 11345 10115
rect 11379 10112 11391 10115
rect 11698 10112 11704 10124
rect 11379 10084 11704 10112
rect 11379 10081 11391 10084
rect 11333 10075 11391 10081
rect 11698 10072 11704 10084
rect 11756 10072 11762 10124
rect 12066 10112 12072 10124
rect 12027 10084 12072 10112
rect 12066 10072 12072 10084
rect 12124 10072 12130 10124
rect 12434 10072 12440 10124
rect 12492 10112 12498 10124
rect 12529 10115 12587 10121
rect 12529 10112 12541 10115
rect 12492 10084 12541 10112
rect 12492 10072 12498 10084
rect 12529 10081 12541 10084
rect 12575 10081 12587 10115
rect 12529 10075 12587 10081
rect 12713 10115 12771 10121
rect 12713 10081 12725 10115
rect 12759 10112 12771 10115
rect 12894 10112 12900 10124
rect 12759 10084 12900 10112
rect 12759 10081 12771 10084
rect 12713 10075 12771 10081
rect 12894 10072 12900 10084
rect 12952 10072 12958 10124
rect 13262 10112 13268 10124
rect 13223 10084 13268 10112
rect 13262 10072 13268 10084
rect 13320 10072 13326 10124
rect 14108 10121 14136 10220
rect 14274 10208 14280 10220
rect 14332 10208 14338 10260
rect 15654 10248 15660 10260
rect 15615 10220 15660 10248
rect 15654 10208 15660 10220
rect 15712 10208 15718 10260
rect 17218 10248 17224 10260
rect 16408 10220 17224 10248
rect 15102 10140 15108 10192
rect 15160 10180 15166 10192
rect 15473 10183 15531 10189
rect 15473 10180 15485 10183
rect 15160 10152 15485 10180
rect 15160 10140 15166 10152
rect 15473 10149 15485 10152
rect 15519 10180 15531 10183
rect 16408 10180 16436 10220
rect 17218 10208 17224 10220
rect 17276 10208 17282 10260
rect 18233 10251 18291 10257
rect 18233 10217 18245 10251
rect 18279 10248 18291 10251
rect 18506 10248 18512 10260
rect 18279 10220 18512 10248
rect 18279 10217 18291 10220
rect 18233 10211 18291 10217
rect 18506 10208 18512 10220
rect 18564 10208 18570 10260
rect 19245 10251 19303 10257
rect 19245 10217 19257 10251
rect 19291 10248 19303 10251
rect 19610 10248 19616 10260
rect 19291 10220 19616 10248
rect 19291 10217 19303 10220
rect 19245 10211 19303 10217
rect 19610 10208 19616 10220
rect 19668 10208 19674 10260
rect 16758 10180 16764 10192
rect 15519 10152 16436 10180
rect 16719 10152 16764 10180
rect 15519 10149 15531 10152
rect 15473 10143 15531 10149
rect 14093 10115 14151 10121
rect 14093 10081 14105 10115
rect 14139 10081 14151 10115
rect 14093 10075 14151 10081
rect 15654 10072 15660 10124
rect 15712 10112 15718 10124
rect 16022 10112 16028 10124
rect 15712 10084 16028 10112
rect 15712 10072 15718 10084
rect 16022 10072 16028 10084
rect 16080 10072 16086 10124
rect 16301 10115 16359 10121
rect 16301 10081 16313 10115
rect 16347 10112 16359 10115
rect 16408 10112 16436 10152
rect 16758 10140 16764 10152
rect 16816 10140 16822 10192
rect 19061 10183 19119 10189
rect 19061 10149 19073 10183
rect 19107 10180 19119 10183
rect 20898 10180 20904 10192
rect 19107 10152 20904 10180
rect 19107 10149 19119 10152
rect 19061 10143 19119 10149
rect 20898 10140 20904 10152
rect 20956 10140 20962 10192
rect 18417 10115 18475 10121
rect 18417 10112 18429 10115
rect 16347 10084 16436 10112
rect 17880 10084 18429 10112
rect 16347 10081 16359 10084
rect 16301 10075 16359 10081
rect 12253 10047 12311 10053
rect 12253 10044 12265 10047
rect 9784 10016 12265 10044
rect 12253 10013 12265 10016
rect 12299 10013 12311 10047
rect 12802 10044 12808 10056
rect 12763 10016 12808 10044
rect 12253 10007 12311 10013
rect 12802 10004 12808 10016
rect 12860 10004 12866 10056
rect 16853 10047 16911 10053
rect 12912 10016 16804 10044
rect 9585 9979 9643 9985
rect 9585 9976 9597 9979
rect 9315 9948 9597 9976
rect 9585 9945 9597 9948
rect 9631 9945 9643 9979
rect 10597 9979 10655 9985
rect 10597 9976 10609 9979
rect 9585 9939 9643 9945
rect 9692 9948 10609 9976
rect 9692 9908 9720 9948
rect 10597 9945 10609 9948
rect 10643 9945 10655 9979
rect 10597 9939 10655 9945
rect 10689 9979 10747 9985
rect 10689 9945 10701 9979
rect 10735 9976 10747 9979
rect 10778 9976 10784 9988
rect 10735 9948 10784 9976
rect 10735 9945 10747 9948
rect 10689 9939 10747 9945
rect 10778 9936 10784 9948
rect 10836 9936 10842 9988
rect 11238 9936 11244 9988
rect 11296 9976 11302 9988
rect 11514 9976 11520 9988
rect 11296 9948 11520 9976
rect 11296 9936 11302 9948
rect 11514 9936 11520 9948
rect 11572 9936 11578 9988
rect 11698 9936 11704 9988
rect 11756 9976 11762 9988
rect 12912 9976 12940 10016
rect 13541 9979 13599 9985
rect 13541 9976 13553 9979
rect 11756 9948 12940 9976
rect 13004 9948 13553 9976
rect 11756 9936 11762 9948
rect 9232 9880 9720 9908
rect 9766 9868 9772 9920
rect 9824 9908 9830 9920
rect 9950 9908 9956 9920
rect 9824 9880 9956 9908
rect 9824 9868 9830 9880
rect 9950 9868 9956 9880
rect 10008 9908 10014 9920
rect 10137 9911 10195 9917
rect 10137 9908 10149 9911
rect 10008 9880 10149 9908
rect 10008 9868 10014 9880
rect 10137 9877 10149 9880
rect 10183 9877 10195 9911
rect 10137 9871 10195 9877
rect 11057 9911 11115 9917
rect 11057 9877 11069 9911
rect 11103 9908 11115 9911
rect 11425 9911 11483 9917
rect 11425 9908 11437 9911
rect 11103 9880 11437 9908
rect 11103 9877 11115 9880
rect 11057 9871 11115 9877
rect 11425 9877 11437 9880
rect 11471 9877 11483 9911
rect 11425 9871 11483 9877
rect 12066 9868 12072 9920
rect 12124 9908 12130 9920
rect 13004 9908 13032 9948
rect 13541 9945 13553 9948
rect 13587 9945 13599 9979
rect 13541 9939 13599 9945
rect 13630 9936 13636 9988
rect 13688 9976 13694 9988
rect 13817 9979 13875 9985
rect 13817 9976 13829 9979
rect 13688 9948 13829 9976
rect 13688 9936 13694 9948
rect 13817 9945 13829 9948
rect 13863 9945 13875 9979
rect 13817 9939 13875 9945
rect 14360 9979 14418 9985
rect 14360 9945 14372 9979
rect 14406 9976 14418 9979
rect 14550 9976 14556 9988
rect 14406 9948 14556 9976
rect 14406 9945 14418 9948
rect 14360 9939 14418 9945
rect 14550 9936 14556 9948
rect 14608 9976 14614 9988
rect 16298 9976 16304 9988
rect 14608 9948 16304 9976
rect 14608 9936 14614 9948
rect 16298 9936 16304 9948
rect 16356 9936 16362 9988
rect 16776 9976 16804 10016
rect 16853 10013 16865 10047
rect 16899 10044 16911 10047
rect 16942 10044 16948 10056
rect 16899 10016 16948 10044
rect 16899 10013 16911 10016
rect 16853 10007 16911 10013
rect 16942 10004 16948 10016
rect 17000 10004 17006 10056
rect 17098 9979 17156 9985
rect 17098 9976 17110 9979
rect 16776 9948 17110 9976
rect 17098 9945 17110 9948
rect 17144 9976 17156 9979
rect 17880 9976 17908 10084
rect 18417 10081 18429 10084
rect 18463 10081 18475 10115
rect 19702 10112 19708 10124
rect 19663 10084 19708 10112
rect 18417 10075 18475 10081
rect 17144 9948 17908 9976
rect 18432 9976 18460 10075
rect 19702 10072 19708 10084
rect 19760 10072 19766 10124
rect 19794 10072 19800 10124
rect 19852 10112 19858 10124
rect 20806 10112 20812 10124
rect 19852 10084 19897 10112
rect 20180 10084 20812 10112
rect 19852 10072 19858 10084
rect 18690 10044 18696 10056
rect 18651 10016 18696 10044
rect 18690 10004 18696 10016
rect 18748 10004 18754 10056
rect 19613 10047 19671 10053
rect 19613 10013 19625 10047
rect 19659 10044 19671 10047
rect 20180 10044 20208 10084
rect 20806 10072 20812 10084
rect 20864 10072 20870 10124
rect 20993 10115 21051 10121
rect 20993 10081 21005 10115
rect 21039 10112 21051 10115
rect 21542 10112 21548 10124
rect 21039 10084 21548 10112
rect 21039 10081 21051 10084
rect 20993 10075 21051 10081
rect 21542 10072 21548 10084
rect 21600 10072 21606 10124
rect 19659 10016 20208 10044
rect 20441 10047 20499 10053
rect 19659 10013 19671 10016
rect 19613 10007 19671 10013
rect 20441 10013 20453 10047
rect 20487 10044 20499 10047
rect 20714 10044 20720 10056
rect 20487 10016 20521 10044
rect 20675 10016 20720 10044
rect 20487 10013 20499 10016
rect 20441 10007 20499 10013
rect 20073 9979 20131 9985
rect 20073 9976 20085 9979
rect 18432 9948 20085 9976
rect 17144 9945 17156 9948
rect 17098 9939 17156 9945
rect 20073 9945 20085 9948
rect 20119 9945 20131 9979
rect 20073 9939 20131 9945
rect 20257 9979 20315 9985
rect 20257 9945 20269 9979
rect 20303 9976 20315 9979
rect 20456 9976 20484 10007
rect 20714 10004 20720 10016
rect 20772 10004 20778 10056
rect 20530 9976 20536 9988
rect 20303 9948 20536 9976
rect 20303 9945 20315 9948
rect 20257 9939 20315 9945
rect 20530 9936 20536 9948
rect 20588 9936 20594 9988
rect 12124 9880 13032 9908
rect 13173 9911 13231 9917
rect 12124 9868 12130 9880
rect 13173 9877 13185 9911
rect 13219 9908 13231 9911
rect 13722 9908 13728 9920
rect 13219 9880 13728 9908
rect 13219 9877 13231 9880
rect 13173 9871 13231 9877
rect 13722 9868 13728 9880
rect 13780 9868 13786 9920
rect 16022 9908 16028 9920
rect 15983 9880 16028 9908
rect 16022 9868 16028 9880
rect 16080 9868 16086 9920
rect 16114 9868 16120 9920
rect 16172 9908 16178 9920
rect 16485 9911 16543 9917
rect 16485 9908 16497 9911
rect 16172 9880 16497 9908
rect 16172 9868 16178 9880
rect 16485 9877 16497 9880
rect 16531 9877 16543 9911
rect 16485 9871 16543 9877
rect 16942 9868 16948 9920
rect 17000 9908 17006 9920
rect 18046 9908 18052 9920
rect 17000 9880 18052 9908
rect 17000 9868 17006 9880
rect 18046 9868 18052 9880
rect 18104 9908 18110 9920
rect 18506 9908 18512 9920
rect 18104 9880 18512 9908
rect 18104 9868 18110 9880
rect 18506 9868 18512 9880
rect 18564 9868 18570 9920
rect 18601 9911 18659 9917
rect 18601 9877 18613 9911
rect 18647 9908 18659 9911
rect 18690 9908 18696 9920
rect 18647 9880 18696 9908
rect 18647 9877 18659 9880
rect 18601 9871 18659 9877
rect 18690 9868 18696 9880
rect 18748 9868 18754 9920
rect 18782 9868 18788 9920
rect 18840 9908 18846 9920
rect 19886 9908 19892 9920
rect 18840 9880 19892 9908
rect 18840 9868 18846 9880
rect 19886 9868 19892 9880
rect 19944 9868 19950 9920
rect 20625 9911 20683 9917
rect 20625 9877 20637 9911
rect 20671 9908 20683 9911
rect 20806 9908 20812 9920
rect 20671 9880 20812 9908
rect 20671 9877 20683 9880
rect 20625 9871 20683 9877
rect 20806 9868 20812 9880
rect 20864 9868 20870 9920
rect 1104 9818 22056 9840
rect 1104 9766 6148 9818
rect 6200 9766 6212 9818
rect 6264 9766 6276 9818
rect 6328 9766 6340 9818
rect 6392 9766 6404 9818
rect 6456 9766 11346 9818
rect 11398 9766 11410 9818
rect 11462 9766 11474 9818
rect 11526 9766 11538 9818
rect 11590 9766 11602 9818
rect 11654 9766 16544 9818
rect 16596 9766 16608 9818
rect 16660 9766 16672 9818
rect 16724 9766 16736 9818
rect 16788 9766 16800 9818
rect 16852 9766 21742 9818
rect 21794 9766 21806 9818
rect 21858 9766 21870 9818
rect 21922 9766 21934 9818
rect 21986 9766 21998 9818
rect 22050 9766 22056 9818
rect 1104 9744 22056 9766
rect 1854 9664 1860 9716
rect 1912 9704 1918 9716
rect 3050 9704 3056 9716
rect 1912 9676 3056 9704
rect 1912 9664 1918 9676
rect 3050 9664 3056 9676
rect 3108 9664 3114 9716
rect 3234 9664 3240 9716
rect 3292 9704 3298 9716
rect 7282 9704 7288 9716
rect 3292 9676 7288 9704
rect 3292 9664 3298 9676
rect 7282 9664 7288 9676
rect 7340 9664 7346 9716
rect 7466 9664 7472 9716
rect 7524 9704 7530 9716
rect 7561 9707 7619 9713
rect 7561 9704 7573 9707
rect 7524 9676 7573 9704
rect 7524 9664 7530 9676
rect 7561 9673 7573 9676
rect 7607 9673 7619 9707
rect 7561 9667 7619 9673
rect 8294 9664 8300 9716
rect 8352 9704 8358 9716
rect 9769 9707 9827 9713
rect 9769 9704 9781 9707
rect 8352 9676 9781 9704
rect 8352 9664 8358 9676
rect 9769 9673 9781 9676
rect 9815 9673 9827 9707
rect 9769 9667 9827 9673
rect 9861 9707 9919 9713
rect 9861 9673 9873 9707
rect 9907 9673 9919 9707
rect 9861 9667 9919 9673
rect 1486 9636 1492 9648
rect 1399 9608 1492 9636
rect 1486 9596 1492 9608
rect 1544 9636 1550 9648
rect 3418 9636 3424 9648
rect 1544 9608 3424 9636
rect 1544 9596 1550 9608
rect 3418 9596 3424 9608
rect 3476 9596 3482 9648
rect 7101 9639 7159 9645
rect 3804 9608 6500 9636
rect 2225 9571 2283 9577
rect 2225 9537 2237 9571
rect 2271 9568 2283 9571
rect 2314 9568 2320 9580
rect 2271 9540 2320 9568
rect 2271 9537 2283 9540
rect 2225 9531 2283 9537
rect 2314 9528 2320 9540
rect 2372 9528 2378 9580
rect 2498 9528 2504 9580
rect 2556 9568 2562 9580
rect 2685 9571 2743 9577
rect 2685 9568 2697 9571
rect 2556 9540 2697 9568
rect 2556 9528 2562 9540
rect 2685 9537 2697 9540
rect 2731 9537 2743 9571
rect 3602 9568 3608 9580
rect 2685 9531 2743 9537
rect 2792 9540 3608 9568
rect 1946 9500 1952 9512
rect 1907 9472 1952 9500
rect 1946 9460 1952 9472
rect 2004 9460 2010 9512
rect 2130 9500 2136 9512
rect 2091 9472 2136 9500
rect 2130 9460 2136 9472
rect 2188 9460 2194 9512
rect 2792 9500 2820 9540
rect 3602 9528 3608 9540
rect 3660 9528 3666 9580
rect 3694 9528 3700 9580
rect 3752 9568 3758 9580
rect 3804 9577 3832 9608
rect 3789 9571 3847 9577
rect 3789 9568 3801 9571
rect 3752 9540 3801 9568
rect 3752 9528 3758 9540
rect 3789 9537 3801 9540
rect 3835 9537 3847 9571
rect 3789 9531 3847 9537
rect 3881 9571 3939 9577
rect 3881 9537 3893 9571
rect 3927 9568 3939 9571
rect 4154 9568 4160 9580
rect 3927 9540 4160 9568
rect 3927 9537 3939 9540
rect 3881 9531 3939 9537
rect 4154 9528 4160 9540
rect 4212 9568 4218 9580
rect 4522 9568 4528 9580
rect 4212 9540 4528 9568
rect 4212 9528 4218 9540
rect 4522 9528 4528 9540
rect 4580 9528 4586 9580
rect 4706 9568 4712 9580
rect 4667 9540 4712 9568
rect 4706 9528 4712 9540
rect 4764 9528 4770 9580
rect 5258 9528 5264 9580
rect 5316 9568 5322 9580
rect 5537 9571 5595 9577
rect 5537 9568 5549 9571
rect 5316 9540 5549 9568
rect 5316 9528 5322 9540
rect 5537 9537 5549 9540
rect 5583 9537 5595 9571
rect 6178 9568 6184 9580
rect 6139 9540 6184 9568
rect 5537 9531 5595 9537
rect 6178 9528 6184 9540
rect 6236 9528 6242 9580
rect 2231 9472 2820 9500
rect 1673 9435 1731 9441
rect 1673 9401 1685 9435
rect 1719 9432 1731 9435
rect 1854 9432 1860 9444
rect 1719 9404 1860 9432
rect 1719 9401 1731 9404
rect 1673 9395 1731 9401
rect 1854 9392 1860 9404
rect 1912 9392 1918 9444
rect 2231 9432 2259 9472
rect 3050 9460 3056 9512
rect 3108 9500 3114 9512
rect 3513 9503 3571 9509
rect 3513 9500 3525 9503
rect 3108 9472 3525 9500
rect 3108 9460 3114 9472
rect 3513 9469 3525 9472
rect 3559 9469 3571 9503
rect 4798 9500 4804 9512
rect 3513 9463 3571 9469
rect 3896 9472 4568 9500
rect 4759 9472 4804 9500
rect 1964 9404 2259 9432
rect 2593 9435 2651 9441
rect 1486 9324 1492 9376
rect 1544 9364 1550 9376
rect 1964 9364 1992 9404
rect 2593 9401 2605 9435
rect 2639 9432 2651 9435
rect 2682 9432 2688 9444
rect 2639 9404 2688 9432
rect 2639 9401 2651 9404
rect 2593 9395 2651 9401
rect 2682 9392 2688 9404
rect 2740 9392 2746 9444
rect 3896 9432 3924 9472
rect 4062 9432 4068 9444
rect 2792 9404 3924 9432
rect 4023 9404 4068 9432
rect 1544 9336 1992 9364
rect 1544 9324 1550 9336
rect 2222 9324 2228 9376
rect 2280 9364 2286 9376
rect 2792 9364 2820 9404
rect 4062 9392 4068 9404
rect 4120 9392 4126 9444
rect 4540 9432 4568 9472
rect 4798 9460 4804 9472
rect 4856 9460 4862 9512
rect 4893 9503 4951 9509
rect 4893 9469 4905 9503
rect 4939 9469 4951 9503
rect 5626 9500 5632 9512
rect 5587 9472 5632 9500
rect 4893 9463 4951 9469
rect 4908 9432 4936 9463
rect 5626 9460 5632 9472
rect 5684 9460 5690 9512
rect 5721 9503 5779 9509
rect 5721 9469 5733 9503
rect 5767 9469 5779 9503
rect 5721 9463 5779 9469
rect 5736 9432 5764 9463
rect 4540 9404 5764 9432
rect 6472 9376 6500 9608
rect 7101 9605 7113 9639
rect 7147 9636 7159 9639
rect 7834 9636 7840 9648
rect 7147 9608 7840 9636
rect 7147 9605 7159 9608
rect 7101 9599 7159 9605
rect 7834 9596 7840 9608
rect 7892 9596 7898 9648
rect 7929 9639 7987 9645
rect 7929 9605 7941 9639
rect 7975 9636 7987 9639
rect 8202 9636 8208 9648
rect 7975 9608 8208 9636
rect 7975 9605 7987 9608
rect 7929 9599 7987 9605
rect 8202 9596 8208 9608
rect 8260 9596 8266 9648
rect 8590 9608 8892 9636
rect 6638 9568 6644 9580
rect 6599 9540 6644 9568
rect 6638 9528 6644 9540
rect 6696 9528 6702 9580
rect 8386 9568 8392 9580
rect 7392 9540 8156 9568
rect 8347 9540 8392 9568
rect 6825 9503 6883 9509
rect 6825 9469 6837 9503
rect 6871 9469 6883 9503
rect 7006 9500 7012 9512
rect 6967 9472 7012 9500
rect 6825 9463 6883 9469
rect 6840 9432 6868 9463
rect 7006 9460 7012 9472
rect 7064 9460 7070 9512
rect 7392 9432 7420 9540
rect 8018 9500 8024 9512
rect 7979 9472 8024 9500
rect 8018 9460 8024 9472
rect 8076 9460 8082 9512
rect 8128 9509 8156 9540
rect 8386 9528 8392 9540
rect 8444 9528 8450 9580
rect 8590 9568 8618 9608
rect 8496 9540 8618 9568
rect 8113 9503 8171 9509
rect 8113 9469 8125 9503
rect 8159 9500 8171 9503
rect 8294 9500 8300 9512
rect 8159 9472 8300 9500
rect 8159 9469 8171 9472
rect 8113 9463 8171 9469
rect 8294 9460 8300 9472
rect 8352 9460 8358 9512
rect 8496 9500 8524 9540
rect 8653 9528 8659 9580
rect 8711 9568 8717 9580
rect 8864 9568 8892 9608
rect 9122 9596 9128 9648
rect 9180 9636 9186 9648
rect 9876 9636 9904 9667
rect 10686 9664 10692 9716
rect 10744 9704 10750 9716
rect 12526 9704 12532 9716
rect 10744 9676 12532 9704
rect 10744 9664 10750 9676
rect 12526 9664 12532 9676
rect 12584 9664 12590 9716
rect 12897 9707 12955 9713
rect 12897 9673 12909 9707
rect 12943 9704 12955 9707
rect 13262 9704 13268 9716
rect 12943 9676 13268 9704
rect 12943 9673 12955 9676
rect 12897 9667 12955 9673
rect 13262 9664 13268 9676
rect 13320 9664 13326 9716
rect 15378 9704 15384 9716
rect 15212 9676 15384 9704
rect 10226 9636 10232 9648
rect 9180 9608 9904 9636
rect 10187 9608 10232 9636
rect 9180 9596 9186 9608
rect 10226 9596 10232 9608
rect 10284 9636 10290 9648
rect 10870 9636 10876 9648
rect 10284 9608 10876 9636
rect 10284 9596 10290 9608
rect 10870 9596 10876 9608
rect 10928 9596 10934 9648
rect 12345 9639 12403 9645
rect 12345 9605 12357 9639
rect 12391 9636 12403 9639
rect 12805 9639 12863 9645
rect 12805 9636 12817 9639
rect 12391 9608 12817 9636
rect 12391 9605 12403 9608
rect 12345 9599 12403 9605
rect 12805 9605 12817 9608
rect 12851 9636 12863 9639
rect 12986 9636 12992 9648
rect 12851 9608 12992 9636
rect 12851 9605 12863 9608
rect 12805 9599 12863 9605
rect 12986 9596 12992 9608
rect 13044 9596 13050 9648
rect 13630 9596 13636 9648
rect 13688 9636 13694 9648
rect 14384 9646 14964 9674
rect 14384 9636 14412 9646
rect 13688 9608 14412 9636
rect 14936 9636 14964 9646
rect 15212 9636 15240 9676
rect 15378 9664 15384 9676
rect 15436 9704 15442 9716
rect 15436 9676 15792 9704
rect 15436 9664 15442 9676
rect 14936 9608 15240 9636
rect 13688 9596 13694 9608
rect 15562 9596 15568 9648
rect 15620 9636 15626 9648
rect 15657 9639 15715 9645
rect 15657 9636 15669 9639
rect 15620 9608 15669 9636
rect 15620 9596 15626 9608
rect 15657 9605 15669 9608
rect 15703 9605 15715 9639
rect 15764 9636 15792 9676
rect 16298 9664 16304 9716
rect 16356 9704 16362 9716
rect 18230 9704 18236 9716
rect 16356 9676 18236 9704
rect 16356 9664 16362 9676
rect 18230 9664 18236 9676
rect 18288 9664 18294 9716
rect 18322 9664 18328 9716
rect 18380 9704 18386 9716
rect 18380 9676 19012 9704
rect 18380 9664 18386 9676
rect 16022 9636 16028 9648
rect 15764 9608 16028 9636
rect 15657 9599 15715 9605
rect 16022 9596 16028 9608
rect 16080 9636 16086 9648
rect 16117 9639 16175 9645
rect 16117 9636 16129 9639
rect 16080 9608 16129 9636
rect 16080 9596 16086 9608
rect 16117 9605 16129 9608
rect 16163 9605 16175 9639
rect 16117 9599 16175 9605
rect 16206 9596 16212 9648
rect 16264 9636 16270 9648
rect 16393 9639 16451 9645
rect 16393 9636 16405 9639
rect 16264 9608 16405 9636
rect 16264 9596 16270 9608
rect 16393 9605 16405 9608
rect 16439 9605 16451 9639
rect 16393 9599 16451 9605
rect 8711 9540 8756 9568
rect 8864 9540 9674 9568
rect 8711 9528 8717 9540
rect 8404 9472 8524 9500
rect 6840 9404 7420 9432
rect 7469 9435 7527 9441
rect 7469 9401 7481 9435
rect 7515 9432 7527 9435
rect 7558 9432 7564 9444
rect 7515 9404 7564 9432
rect 7515 9401 7527 9404
rect 7469 9395 7527 9401
rect 7558 9392 7564 9404
rect 7616 9392 7622 9444
rect 7650 9392 7656 9444
rect 7708 9432 7714 9444
rect 8404 9432 8432 9472
rect 7708 9404 8432 9432
rect 9646 9432 9674 9540
rect 10134 9528 10140 9580
rect 10192 9568 10198 9580
rect 10321 9571 10379 9577
rect 10321 9568 10333 9571
rect 10192 9540 10333 9568
rect 10192 9528 10198 9540
rect 10321 9537 10333 9540
rect 10367 9568 10379 9571
rect 10686 9568 10692 9580
rect 10367 9540 10692 9568
rect 10367 9537 10379 9540
rect 10321 9531 10379 9537
rect 10686 9528 10692 9540
rect 10744 9528 10750 9580
rect 11330 9568 11336 9580
rect 10796 9540 11336 9568
rect 10410 9500 10416 9512
rect 10371 9472 10416 9500
rect 10410 9460 10416 9472
rect 10468 9460 10474 9512
rect 10502 9460 10508 9512
rect 10560 9500 10566 9512
rect 10796 9500 10824 9540
rect 11330 9528 11336 9540
rect 11388 9528 11394 9580
rect 11606 9528 11612 9580
rect 11664 9568 11670 9580
rect 11885 9571 11943 9577
rect 11885 9568 11897 9571
rect 11664 9540 11897 9568
rect 11664 9528 11670 9540
rect 11885 9537 11897 9540
rect 11931 9537 11943 9571
rect 11885 9531 11943 9537
rect 12434 9528 12440 9580
rect 12492 9568 12498 9580
rect 13449 9571 13507 9577
rect 13449 9568 13461 9571
rect 12492 9540 13461 9568
rect 12492 9528 12498 9540
rect 13449 9537 13461 9540
rect 13495 9568 13507 9571
rect 13722 9568 13728 9580
rect 13495 9540 13728 9568
rect 13495 9537 13507 9540
rect 13449 9531 13507 9537
rect 13722 9528 13728 9540
rect 13780 9568 13786 9580
rect 13817 9571 13875 9577
rect 13817 9568 13829 9571
rect 13780 9540 13829 9568
rect 13780 9528 13786 9540
rect 13817 9537 13829 9540
rect 13863 9537 13875 9571
rect 13817 9531 13875 9537
rect 14461 9571 14519 9577
rect 14461 9537 14473 9571
rect 14507 9568 14519 9571
rect 15013 9571 15071 9577
rect 14507 9540 14872 9568
rect 14507 9537 14519 9540
rect 14461 9531 14519 9537
rect 10560 9472 10824 9500
rect 10560 9460 10566 9472
rect 11054 9460 11060 9512
rect 11112 9500 11118 9512
rect 11149 9503 11207 9509
rect 11149 9500 11161 9503
rect 11112 9472 11161 9500
rect 11112 9460 11118 9472
rect 11149 9469 11161 9472
rect 11195 9500 11207 9503
rect 11514 9500 11520 9512
rect 11195 9472 11520 9500
rect 11195 9469 11207 9472
rect 11149 9463 11207 9469
rect 11514 9460 11520 9472
rect 11572 9460 11578 9512
rect 11698 9500 11704 9512
rect 11659 9472 11704 9500
rect 11698 9460 11704 9472
rect 11756 9460 11762 9512
rect 11793 9503 11851 9509
rect 11793 9469 11805 9503
rect 11839 9469 11851 9503
rect 12618 9500 12624 9512
rect 12579 9472 12624 9500
rect 11793 9463 11851 9469
rect 11241 9435 11299 9441
rect 11241 9432 11253 9435
rect 9646 9404 11253 9432
rect 7708 9392 7714 9404
rect 11241 9401 11253 9404
rect 11287 9432 11299 9435
rect 11808 9432 11836 9463
rect 12618 9460 12624 9472
rect 12676 9460 12682 9512
rect 14844 9500 14872 9540
rect 15013 9537 15025 9571
rect 15059 9568 15071 9571
rect 15470 9568 15476 9580
rect 15059 9540 15476 9568
rect 15059 9537 15071 9540
rect 15013 9531 15071 9537
rect 15470 9528 15476 9540
rect 15528 9528 15534 9580
rect 15746 9568 15752 9580
rect 15707 9540 15752 9568
rect 15746 9528 15752 9540
rect 15804 9528 15810 9580
rect 16298 9568 16304 9580
rect 15948 9540 16304 9568
rect 14918 9500 14924 9512
rect 14844 9472 14924 9500
rect 14918 9460 14924 9472
rect 14976 9460 14982 9512
rect 15948 9509 15976 9540
rect 16298 9528 16304 9540
rect 16356 9528 16362 9580
rect 17126 9568 17132 9580
rect 17087 9540 17132 9568
rect 17126 9528 17132 9540
rect 17184 9528 17190 9580
rect 17954 9568 17960 9580
rect 17915 9540 17960 9568
rect 17954 9528 17960 9540
rect 18012 9528 18018 9580
rect 18782 9568 18788 9580
rect 18743 9540 18788 9568
rect 18782 9528 18788 9540
rect 18840 9528 18846 9580
rect 18984 9568 19012 9676
rect 19518 9664 19524 9716
rect 19576 9704 19582 9716
rect 19705 9707 19763 9713
rect 19705 9704 19717 9707
rect 19576 9676 19717 9704
rect 19576 9664 19582 9676
rect 19705 9673 19717 9676
rect 19751 9673 19763 9707
rect 19705 9667 19763 9673
rect 19794 9664 19800 9716
rect 19852 9704 19858 9716
rect 20622 9704 20628 9716
rect 19852 9676 20628 9704
rect 19852 9664 19858 9676
rect 20622 9664 20628 9676
rect 20680 9664 20686 9716
rect 20990 9664 20996 9716
rect 21048 9704 21054 9716
rect 21174 9704 21180 9716
rect 21048 9676 21180 9704
rect 21048 9664 21054 9676
rect 21174 9664 21180 9676
rect 21232 9664 21238 9716
rect 19245 9639 19303 9645
rect 19245 9605 19257 9639
rect 19291 9636 19303 9639
rect 20714 9636 20720 9648
rect 19291 9608 20720 9636
rect 19291 9605 19303 9608
rect 19245 9599 19303 9605
rect 20714 9596 20720 9608
rect 20772 9596 20778 9648
rect 20898 9596 20904 9648
rect 20956 9636 20962 9648
rect 21085 9639 21143 9645
rect 21085 9636 21097 9639
rect 20956 9608 21097 9636
rect 20956 9596 20962 9608
rect 21085 9605 21097 9608
rect 21131 9605 21143 9639
rect 21085 9599 21143 9605
rect 19337 9571 19395 9577
rect 18984 9540 19288 9568
rect 15933 9503 15991 9509
rect 15120 9472 15792 9500
rect 11287 9404 11836 9432
rect 12253 9435 12311 9441
rect 11287 9401 11299 9404
rect 11241 9395 11299 9401
rect 12253 9401 12265 9435
rect 12299 9432 12311 9435
rect 15120 9432 15148 9472
rect 15286 9432 15292 9444
rect 12299 9404 15148 9432
rect 15247 9404 15292 9432
rect 12299 9401 12311 9404
rect 12253 9395 12311 9401
rect 15286 9392 15292 9404
rect 15344 9392 15350 9444
rect 15764 9432 15792 9472
rect 15933 9469 15945 9503
rect 15979 9469 15991 9503
rect 16942 9500 16948 9512
rect 16903 9472 16948 9500
rect 15933 9463 15991 9469
rect 16942 9460 16948 9472
rect 17000 9460 17006 9512
rect 17037 9503 17095 9509
rect 17037 9469 17049 9503
rect 17083 9500 17095 9503
rect 17083 9472 17632 9500
rect 17083 9469 17095 9472
rect 17037 9463 17095 9469
rect 17402 9432 17408 9444
rect 15764 9404 17408 9432
rect 17402 9392 17408 9404
rect 17460 9392 17466 9444
rect 17604 9441 17632 9472
rect 17770 9460 17776 9512
rect 17828 9460 17834 9512
rect 18046 9500 18052 9512
rect 18007 9472 18052 9500
rect 18046 9460 18052 9472
rect 18104 9460 18110 9512
rect 18138 9460 18144 9512
rect 18196 9500 18202 9512
rect 19153 9503 19211 9509
rect 18196 9472 18241 9500
rect 18196 9460 18202 9472
rect 19153 9469 19165 9503
rect 19199 9469 19211 9503
rect 19260 9500 19288 9540
rect 19337 9537 19349 9571
rect 19383 9568 19395 9571
rect 19610 9568 19616 9580
rect 19383 9540 19616 9568
rect 19383 9537 19395 9540
rect 19337 9531 19395 9537
rect 19610 9528 19616 9540
rect 19668 9528 19674 9580
rect 20165 9571 20223 9577
rect 20165 9537 20177 9571
rect 20211 9568 20223 9571
rect 20990 9568 20996 9580
rect 20211 9540 20760 9568
rect 20951 9540 20996 9568
rect 20211 9537 20223 9540
rect 20165 9531 20223 9537
rect 20257 9503 20315 9509
rect 20257 9500 20269 9503
rect 19260 9472 19334 9500
rect 19153 9463 19211 9469
rect 17589 9435 17647 9441
rect 17589 9401 17601 9435
rect 17635 9401 17647 9435
rect 17788 9432 17816 9460
rect 18601 9435 18659 9441
rect 18601 9432 18613 9435
rect 17788 9404 18613 9432
rect 17589 9395 17647 9401
rect 18601 9401 18613 9404
rect 18647 9401 18659 9435
rect 18601 9395 18659 9401
rect 2280 9336 2820 9364
rect 2869 9367 2927 9373
rect 2280 9324 2286 9336
rect 2869 9333 2881 9367
rect 2915 9364 2927 9367
rect 3786 9364 3792 9376
rect 2915 9336 3792 9364
rect 2915 9333 2927 9336
rect 2869 9327 2927 9333
rect 3786 9324 3792 9336
rect 3844 9324 3850 9376
rect 4246 9324 4252 9376
rect 4304 9364 4310 9376
rect 4341 9367 4399 9373
rect 4341 9364 4353 9367
rect 4304 9336 4353 9364
rect 4304 9324 4310 9336
rect 4341 9333 4353 9336
rect 4387 9333 4399 9367
rect 4341 9327 4399 9333
rect 4430 9324 4436 9376
rect 4488 9364 4494 9376
rect 5169 9367 5227 9373
rect 5169 9364 5181 9367
rect 4488 9336 5181 9364
rect 4488 9324 4494 9336
rect 5169 9333 5181 9336
rect 5215 9333 5227 9367
rect 5169 9327 5227 9333
rect 5442 9324 5448 9376
rect 5500 9364 5506 9376
rect 5997 9367 6055 9373
rect 5997 9364 6009 9367
rect 5500 9336 6009 9364
rect 5500 9324 5506 9336
rect 5997 9333 6009 9336
rect 6043 9333 6055 9367
rect 6454 9364 6460 9376
rect 6415 9336 6460 9364
rect 5997 9327 6055 9333
rect 6454 9324 6460 9336
rect 6512 9324 6518 9376
rect 6546 9324 6552 9376
rect 6604 9364 6610 9376
rect 12802 9364 12808 9376
rect 6604 9336 12808 9364
rect 6604 9324 6610 9336
rect 12802 9324 12808 9336
rect 12860 9324 12866 9376
rect 12894 9324 12900 9376
rect 12952 9364 12958 9376
rect 13265 9367 13323 9373
rect 13265 9364 13277 9367
rect 12952 9336 13277 9364
rect 12952 9324 12958 9336
rect 13265 9333 13277 9336
rect 13311 9333 13323 9367
rect 14274 9364 14280 9376
rect 14235 9336 14280 9364
rect 13265 9327 13323 9333
rect 14274 9324 14280 9336
rect 14332 9324 14338 9376
rect 14642 9324 14648 9376
rect 14700 9364 14706 9376
rect 14829 9367 14887 9373
rect 14700 9336 14745 9364
rect 14700 9324 14706 9336
rect 14829 9333 14841 9367
rect 14875 9364 14887 9367
rect 15102 9364 15108 9376
rect 14875 9336 15108 9364
rect 14875 9333 14887 9336
rect 14829 9327 14887 9333
rect 15102 9324 15108 9336
rect 15160 9324 15166 9376
rect 15197 9367 15255 9373
rect 15197 9333 15209 9367
rect 15243 9364 15255 9367
rect 15562 9364 15568 9376
rect 15243 9336 15568 9364
rect 15243 9333 15255 9336
rect 15197 9327 15255 9333
rect 15562 9324 15568 9336
rect 15620 9324 15626 9376
rect 17497 9367 17555 9373
rect 17497 9333 17509 9367
rect 17543 9364 17555 9367
rect 17678 9364 17684 9376
rect 17543 9336 17684 9364
rect 17543 9333 17555 9336
rect 17497 9327 17555 9333
rect 17678 9324 17684 9336
rect 17736 9324 17742 9376
rect 17770 9324 17776 9376
rect 17828 9364 17834 9376
rect 18322 9364 18328 9376
rect 17828 9336 18328 9364
rect 17828 9324 17834 9336
rect 18322 9324 18328 9336
rect 18380 9324 18386 9376
rect 18509 9367 18567 9373
rect 18509 9333 18521 9367
rect 18555 9364 18567 9367
rect 18690 9364 18696 9376
rect 18555 9336 18696 9364
rect 18555 9333 18567 9336
rect 18509 9327 18567 9333
rect 18690 9324 18696 9336
rect 18748 9324 18754 9376
rect 19168 9364 19196 9463
rect 19306 9432 19334 9472
rect 19444 9472 20269 9500
rect 19444 9432 19472 9472
rect 20257 9469 20269 9472
rect 20303 9469 20315 9503
rect 20257 9463 20315 9469
rect 20441 9503 20499 9509
rect 20441 9469 20453 9503
rect 20487 9500 20499 9503
rect 20530 9500 20536 9512
rect 20487 9472 20536 9500
rect 20487 9469 20499 9472
rect 20441 9463 20499 9469
rect 20530 9460 20536 9472
rect 20588 9460 20594 9512
rect 19306 9404 19472 9432
rect 19610 9392 19616 9444
rect 19668 9432 19674 9444
rect 20625 9435 20683 9441
rect 20625 9432 20637 9435
rect 19668 9404 20637 9432
rect 19668 9392 19674 9404
rect 20625 9401 20637 9404
rect 20671 9401 20683 9435
rect 20732 9432 20760 9540
rect 20990 9528 20996 9540
rect 21048 9528 21054 9580
rect 21542 9528 21548 9580
rect 21600 9568 21606 9580
rect 22922 9568 22928 9580
rect 21600 9540 22928 9568
rect 21600 9528 21606 9540
rect 22922 9528 22928 9540
rect 22980 9528 22986 9580
rect 21266 9500 21272 9512
rect 21227 9472 21272 9500
rect 21266 9460 21272 9472
rect 21324 9460 21330 9512
rect 22922 9432 22928 9444
rect 20732 9404 22928 9432
rect 20625 9395 20683 9401
rect 22922 9392 22928 9404
rect 22980 9392 22986 9444
rect 19702 9364 19708 9376
rect 19168 9336 19708 9364
rect 19702 9324 19708 9336
rect 19760 9324 19766 9376
rect 19797 9367 19855 9373
rect 19797 9333 19809 9367
rect 19843 9364 19855 9367
rect 19886 9364 19892 9376
rect 19843 9336 19892 9364
rect 19843 9333 19855 9336
rect 19797 9327 19855 9333
rect 19886 9324 19892 9336
rect 19944 9324 19950 9376
rect 20438 9324 20444 9376
rect 20496 9364 20502 9376
rect 21453 9367 21511 9373
rect 21453 9364 21465 9367
rect 20496 9336 21465 9364
rect 20496 9324 20502 9336
rect 21453 9333 21465 9336
rect 21499 9333 21511 9367
rect 21453 9327 21511 9333
rect 1104 9274 21896 9296
rect 1104 9222 3549 9274
rect 3601 9222 3613 9274
rect 3665 9222 3677 9274
rect 3729 9222 3741 9274
rect 3793 9222 3805 9274
rect 3857 9222 8747 9274
rect 8799 9222 8811 9274
rect 8863 9222 8875 9274
rect 8927 9222 8939 9274
rect 8991 9222 9003 9274
rect 9055 9222 13945 9274
rect 13997 9222 14009 9274
rect 14061 9222 14073 9274
rect 14125 9222 14137 9274
rect 14189 9222 14201 9274
rect 14253 9222 19143 9274
rect 19195 9222 19207 9274
rect 19259 9222 19271 9274
rect 19323 9222 19335 9274
rect 19387 9222 19399 9274
rect 19451 9222 21896 9274
rect 1104 9200 21896 9222
rect 2130 9160 2136 9172
rect 2091 9132 2136 9160
rect 2130 9120 2136 9132
rect 2188 9120 2194 9172
rect 2222 9120 2228 9172
rect 2280 9160 2286 9172
rect 2280 9132 2325 9160
rect 2280 9120 2286 9132
rect 2590 9120 2596 9172
rect 2648 9160 2654 9172
rect 3789 9163 3847 9169
rect 3789 9160 3801 9163
rect 2648 9132 3801 9160
rect 2648 9120 2654 9132
rect 3789 9129 3801 9132
rect 3835 9129 3847 9163
rect 4614 9160 4620 9172
rect 4575 9132 4620 9160
rect 3789 9123 3847 9129
rect 4614 9120 4620 9132
rect 4672 9120 4678 9172
rect 5258 9160 5264 9172
rect 5219 9132 5264 9160
rect 5258 9120 5264 9132
rect 5316 9120 5322 9172
rect 5626 9120 5632 9172
rect 5684 9160 5690 9172
rect 6089 9163 6147 9169
rect 6089 9160 6101 9163
rect 5684 9132 6101 9160
rect 5684 9120 5690 9132
rect 6089 9129 6101 9132
rect 6135 9129 6147 9163
rect 6089 9123 6147 9129
rect 7006 9120 7012 9172
rect 7064 9160 7070 9172
rect 8021 9163 8079 9169
rect 8021 9160 8033 9163
rect 7064 9132 8033 9160
rect 7064 9120 7070 9132
rect 8021 9129 8033 9132
rect 8067 9129 8079 9163
rect 8021 9123 8079 9129
rect 8662 9120 8668 9172
rect 8720 9160 8726 9172
rect 10321 9163 10379 9169
rect 10321 9160 10333 9163
rect 8720 9132 10333 9160
rect 8720 9120 8726 9132
rect 10321 9129 10333 9132
rect 10367 9160 10379 9163
rect 10410 9160 10416 9172
rect 10367 9132 10416 9160
rect 10367 9129 10379 9132
rect 10321 9123 10379 9129
rect 10410 9120 10416 9132
rect 10468 9120 10474 9172
rect 10505 9163 10563 9169
rect 10505 9129 10517 9163
rect 10551 9160 10563 9163
rect 10962 9160 10968 9172
rect 10551 9132 10968 9160
rect 10551 9129 10563 9132
rect 10505 9123 10563 9129
rect 1578 9024 1584 9036
rect 1491 8996 1584 9024
rect 1578 8984 1584 8996
rect 1636 9024 1642 9036
rect 2240 9024 2268 9120
rect 3694 9052 3700 9104
rect 3752 9092 3758 9104
rect 4154 9092 4160 9104
rect 3752 9064 4160 9092
rect 3752 9052 3758 9064
rect 4154 9052 4160 9064
rect 4212 9052 4218 9104
rect 4798 9052 4804 9104
rect 4856 9092 4862 9104
rect 6917 9095 6975 9101
rect 6917 9092 6929 9095
rect 4856 9064 6929 9092
rect 4856 9052 4862 9064
rect 6917 9061 6929 9064
rect 6963 9061 6975 9095
rect 7834 9092 7840 9104
rect 7795 9064 7840 9092
rect 6917 9055 6975 9061
rect 7834 9052 7840 9064
rect 7892 9052 7898 9104
rect 8570 9092 8576 9104
rect 8483 9064 8576 9092
rect 1636 8996 2268 9024
rect 3605 9027 3663 9033
rect 1636 8984 1642 8996
rect 3605 8993 3617 9027
rect 3651 9024 3663 9027
rect 3970 9024 3976 9036
rect 3651 8996 3976 9024
rect 3651 8993 3663 8996
rect 3605 8987 3663 8993
rect 3970 8984 3976 8996
rect 4028 8984 4034 9036
rect 4246 9024 4252 9036
rect 4207 8996 4252 9024
rect 4246 8984 4252 8996
rect 4304 8984 4310 9036
rect 4338 8984 4344 9036
rect 4396 9024 4402 9036
rect 4396 8996 4441 9024
rect 4396 8984 4402 8996
rect 5902 8984 5908 9036
rect 5960 9024 5966 9036
rect 6454 9024 6460 9036
rect 5960 8996 6460 9024
rect 5960 8984 5966 8996
rect 6454 8984 6460 8996
rect 6512 8984 6518 9036
rect 6638 8984 6644 9036
rect 6696 9024 6702 9036
rect 6733 9027 6791 9033
rect 6733 9024 6745 9027
rect 6696 8996 6745 9024
rect 6696 8984 6702 8996
rect 6733 8993 6745 8996
rect 6779 9024 6791 9027
rect 7558 9024 7564 9036
rect 6779 8996 7564 9024
rect 6779 8993 6791 8996
rect 6733 8987 6791 8993
rect 7558 8984 7564 8996
rect 7616 8984 7622 9036
rect 1394 8916 1400 8968
rect 1452 8956 1458 8968
rect 2958 8956 2964 8968
rect 1452 8928 2964 8956
rect 1452 8916 1458 8928
rect 2958 8916 2964 8928
rect 3016 8916 3022 8968
rect 3326 8916 3332 8968
rect 3384 8965 3390 8968
rect 3384 8956 3396 8965
rect 4157 8959 4215 8965
rect 3384 8928 3429 8956
rect 3384 8919 3396 8928
rect 4157 8925 4169 8959
rect 4203 8956 4215 8959
rect 4430 8956 4436 8968
rect 4203 8928 4436 8956
rect 4203 8925 4215 8928
rect 4157 8919 4215 8925
rect 3384 8916 3390 8919
rect 4430 8916 4436 8928
rect 4488 8916 4494 8968
rect 4801 8959 4859 8965
rect 4801 8925 4813 8959
rect 4847 8925 4859 8959
rect 4801 8919 4859 8925
rect 4893 8959 4951 8965
rect 4893 8925 4905 8959
rect 4939 8956 4951 8959
rect 5074 8956 5080 8968
rect 4939 8928 5080 8956
rect 4939 8925 4951 8928
rect 4893 8919 4951 8925
rect 1673 8891 1731 8897
rect 1673 8857 1685 8891
rect 1719 8888 1731 8891
rect 2406 8888 2412 8900
rect 1719 8860 2412 8888
rect 1719 8857 1731 8860
rect 1673 8851 1731 8857
rect 2406 8848 2412 8860
rect 2464 8848 2470 8900
rect 1762 8780 1768 8832
rect 1820 8820 1826 8832
rect 1820 8792 1865 8820
rect 1820 8780 1826 8792
rect 4154 8780 4160 8832
rect 4212 8820 4218 8832
rect 4816 8820 4844 8919
rect 5074 8916 5080 8928
rect 5132 8916 5138 8968
rect 7006 8956 7012 8968
rect 6472 8928 7012 8956
rect 5810 8888 5816 8900
rect 5644 8860 5816 8888
rect 4212 8792 4844 8820
rect 5077 8823 5135 8829
rect 4212 8780 4218 8792
rect 5077 8789 5089 8823
rect 5123 8820 5135 8823
rect 5258 8820 5264 8832
rect 5123 8792 5264 8820
rect 5123 8789 5135 8792
rect 5077 8783 5135 8789
rect 5258 8780 5264 8792
rect 5316 8780 5322 8832
rect 5534 8780 5540 8832
rect 5592 8820 5598 8832
rect 5644 8829 5672 8860
rect 5810 8848 5816 8860
rect 5868 8848 5874 8900
rect 6472 8888 6500 8928
rect 7006 8916 7012 8928
rect 7064 8916 7070 8968
rect 7285 8959 7343 8965
rect 7285 8925 7297 8959
rect 7331 8956 7343 8959
rect 7852 8956 7880 9052
rect 8496 9033 8524 9064
rect 8570 9052 8576 9064
rect 8628 9092 8634 9104
rect 8628 9064 8800 9092
rect 8628 9052 8634 9064
rect 8481 9027 8539 9033
rect 8481 8993 8493 9027
rect 8527 8993 8539 9027
rect 8662 9024 8668 9036
rect 8623 8996 8668 9024
rect 8481 8987 8539 8993
rect 8662 8984 8668 8996
rect 8720 8984 8726 9036
rect 8772 9024 8800 9064
rect 8772 8996 9076 9024
rect 7331 8928 7880 8956
rect 7331 8925 7343 8928
rect 7285 8919 7343 8925
rect 8386 8916 8392 8968
rect 8444 8956 8450 8968
rect 8941 8959 8999 8965
rect 8941 8956 8953 8959
rect 8444 8928 8953 8956
rect 8444 8916 8450 8928
rect 8941 8925 8953 8928
rect 8987 8925 8999 8959
rect 9048 8956 9076 8996
rect 10520 8956 10548 9123
rect 10962 9120 10968 9132
rect 11020 9120 11026 9172
rect 11330 9120 11336 9172
rect 11388 9160 11394 9172
rect 13630 9160 13636 9172
rect 11388 9132 13636 9160
rect 11388 9120 11394 9132
rect 13630 9120 13636 9132
rect 13688 9120 13694 9172
rect 14090 9120 14096 9172
rect 14148 9160 14154 9172
rect 14458 9160 14464 9172
rect 14148 9132 14464 9160
rect 14148 9120 14154 9132
rect 14458 9120 14464 9132
rect 14516 9120 14522 9172
rect 16850 9160 16856 9172
rect 15672 9132 16856 9160
rect 13081 9027 13139 9033
rect 13081 9024 13093 9027
rect 12360 8996 13093 9024
rect 9048 8928 10548 8956
rect 10965 8959 11023 8965
rect 8941 8919 8999 8925
rect 10965 8925 10977 8959
rect 11011 8956 11023 8959
rect 12360 8956 12388 8996
rect 13081 8993 13093 8996
rect 13127 8993 13139 9027
rect 13081 8987 13139 8993
rect 13354 8984 13360 9036
rect 13412 9024 13418 9036
rect 13814 9024 13820 9036
rect 13412 8996 13820 9024
rect 13412 8984 13418 8996
rect 13814 8984 13820 8996
rect 13872 8984 13878 9036
rect 15672 9033 15700 9132
rect 16850 9120 16856 9132
rect 16908 9120 16914 9172
rect 17126 9160 17132 9172
rect 17087 9132 17132 9160
rect 17126 9120 17132 9132
rect 17184 9120 17190 9172
rect 17310 9120 17316 9172
rect 17368 9160 17374 9172
rect 18690 9160 18696 9172
rect 17368 9132 18696 9160
rect 17368 9120 17374 9132
rect 18690 9120 18696 9132
rect 18748 9120 18754 9172
rect 18782 9120 18788 9172
rect 18840 9160 18846 9172
rect 20254 9160 20260 9172
rect 18840 9132 20260 9160
rect 18840 9120 18846 9132
rect 20254 9120 20260 9132
rect 20312 9120 20318 9172
rect 20714 9160 20720 9172
rect 20675 9132 20720 9160
rect 20714 9120 20720 9132
rect 20772 9120 20778 9172
rect 17037 9095 17095 9101
rect 17037 9061 17049 9095
rect 17083 9061 17095 9095
rect 17037 9055 17095 9061
rect 15657 9027 15715 9033
rect 15657 8993 15669 9027
rect 15703 8993 15715 9027
rect 17052 9024 17080 9055
rect 17402 9052 17408 9104
rect 17460 9092 17466 9104
rect 17460 9064 18920 9092
rect 17460 9052 17466 9064
rect 17126 9024 17132 9036
rect 17039 8996 17132 9024
rect 15657 8987 15715 8993
rect 17126 8984 17132 8996
rect 17184 9024 17190 9036
rect 17773 9027 17831 9033
rect 17773 9024 17785 9027
rect 17184 8996 17785 9024
rect 17184 8984 17190 8996
rect 17773 8993 17785 8996
rect 17819 9024 17831 9027
rect 18138 9024 18144 9036
rect 17819 8996 18144 9024
rect 17819 8993 17831 8996
rect 17773 8987 17831 8993
rect 18138 8984 18144 8996
rect 18196 8984 18202 9036
rect 18509 9027 18567 9033
rect 18509 8993 18521 9027
rect 18555 8993 18567 9027
rect 18782 9024 18788 9036
rect 18743 8996 18788 9024
rect 18509 8987 18567 8993
rect 11011 8928 11652 8956
rect 11011 8925 11023 8928
rect 10965 8919 11023 8925
rect 6380 8860 6500 8888
rect 6549 8891 6607 8897
rect 5629 8823 5687 8829
rect 5629 8820 5641 8823
rect 5592 8792 5641 8820
rect 5592 8780 5598 8792
rect 5629 8789 5641 8792
rect 5675 8789 5687 8823
rect 5629 8783 5687 8789
rect 5721 8823 5779 8829
rect 5721 8789 5733 8823
rect 5767 8820 5779 8823
rect 6380 8820 6408 8860
rect 6549 8857 6561 8891
rect 6595 8888 6607 8891
rect 6638 8888 6644 8900
rect 6595 8860 6644 8888
rect 6595 8857 6607 8860
rect 6549 8851 6607 8857
rect 6638 8848 6644 8860
rect 6696 8848 6702 8900
rect 9030 8848 9036 8900
rect 9088 8888 9094 8900
rect 9208 8891 9266 8897
rect 9208 8888 9220 8891
rect 9088 8860 9220 8888
rect 9088 8848 9094 8860
rect 9208 8857 9220 8860
rect 9254 8888 9266 8891
rect 9254 8860 11100 8888
rect 9254 8857 9266 8860
rect 9208 8851 9266 8857
rect 11072 8832 11100 8860
rect 5767 8792 6408 8820
rect 6457 8823 6515 8829
rect 5767 8789 5779 8792
rect 5721 8783 5779 8789
rect 6457 8789 6469 8823
rect 6503 8820 6515 8823
rect 6914 8820 6920 8832
rect 6503 8792 6920 8820
rect 6503 8789 6515 8792
rect 6457 8783 6515 8789
rect 6914 8780 6920 8792
rect 6972 8780 6978 8832
rect 7374 8780 7380 8832
rect 7432 8820 7438 8832
rect 7432 8792 7477 8820
rect 7432 8780 7438 8792
rect 7650 8780 7656 8832
rect 7708 8820 7714 8832
rect 8389 8823 8447 8829
rect 8389 8820 8401 8823
rect 7708 8792 8401 8820
rect 7708 8780 7714 8792
rect 8389 8789 8401 8792
rect 8435 8789 8447 8823
rect 8389 8783 8447 8789
rect 8570 8780 8576 8832
rect 8628 8820 8634 8832
rect 10597 8823 10655 8829
rect 10597 8820 10609 8823
rect 8628 8792 10609 8820
rect 8628 8780 8634 8792
rect 10597 8789 10609 8792
rect 10643 8789 10655 8823
rect 10778 8820 10784 8832
rect 10739 8792 10784 8820
rect 10597 8783 10655 8789
rect 10778 8780 10784 8792
rect 10836 8780 10842 8832
rect 11054 8820 11060 8832
rect 11015 8792 11060 8820
rect 11054 8780 11060 8792
rect 11112 8780 11118 8832
rect 11624 8820 11652 8928
rect 12268 8928 12388 8956
rect 12437 8959 12495 8965
rect 11698 8848 11704 8900
rect 11756 8888 11762 8900
rect 12170 8891 12228 8897
rect 12170 8888 12182 8891
rect 11756 8860 12182 8888
rect 11756 8848 11762 8860
rect 12170 8857 12182 8860
rect 12216 8888 12228 8891
rect 12268 8888 12296 8928
rect 12437 8925 12449 8959
rect 12483 8925 12495 8959
rect 12894 8956 12900 8968
rect 12855 8928 12900 8956
rect 12437 8919 12495 8925
rect 12452 8888 12480 8919
rect 12894 8916 12900 8928
rect 12952 8916 12958 8968
rect 14090 8956 14096 8968
rect 13004 8928 14096 8956
rect 12802 8888 12808 8900
rect 12216 8860 12296 8888
rect 12348 8860 12808 8888
rect 12216 8857 12228 8860
rect 12170 8851 12228 8857
rect 12348 8820 12376 8860
rect 12802 8848 12808 8860
rect 12860 8888 12866 8900
rect 13004 8888 13032 8928
rect 14090 8916 14096 8928
rect 14148 8916 14154 8968
rect 15470 8956 15476 8968
rect 15120 8928 15476 8956
rect 12860 8860 13032 8888
rect 12860 8848 12866 8860
rect 13354 8848 13360 8900
rect 13412 8888 13418 8900
rect 13633 8891 13691 8897
rect 13633 8888 13645 8891
rect 13412 8860 13645 8888
rect 13412 8848 13418 8860
rect 13633 8857 13645 8860
rect 13679 8857 13691 8891
rect 13633 8851 13691 8857
rect 13722 8848 13728 8900
rect 13780 8888 13786 8900
rect 14338 8891 14396 8897
rect 14338 8888 14350 8891
rect 13780 8860 14350 8888
rect 13780 8848 13786 8860
rect 14338 8857 14350 8860
rect 14384 8857 14396 8891
rect 14338 8851 14396 8857
rect 12526 8820 12532 8832
rect 11624 8792 12376 8820
rect 12487 8792 12532 8820
rect 12526 8780 12532 8792
rect 12584 8780 12590 8832
rect 12894 8780 12900 8832
rect 12952 8820 12958 8832
rect 12989 8823 13047 8829
rect 12989 8820 13001 8823
rect 12952 8792 13001 8820
rect 12952 8780 12958 8792
rect 12989 8789 13001 8792
rect 13035 8789 13047 8823
rect 13538 8820 13544 8832
rect 13499 8792 13544 8820
rect 12989 8783 13047 8789
rect 13538 8780 13544 8792
rect 13596 8780 13602 8832
rect 13909 8823 13967 8829
rect 13909 8789 13921 8823
rect 13955 8820 13967 8823
rect 15120 8820 15148 8928
rect 15470 8916 15476 8928
rect 15528 8916 15534 8968
rect 15924 8959 15982 8965
rect 15924 8956 15936 8959
rect 15672 8928 15936 8956
rect 15194 8848 15200 8900
rect 15252 8888 15258 8900
rect 15672 8888 15700 8928
rect 15924 8925 15936 8928
rect 15970 8956 15982 8959
rect 18524 8956 18552 8987
rect 18782 8984 18788 8996
rect 18840 8984 18846 9036
rect 18892 9024 18920 9064
rect 21266 9024 21272 9036
rect 18892 8996 19380 9024
rect 21227 8996 21272 9024
rect 18598 8956 18604 8968
rect 15970 8928 18604 8956
rect 15970 8925 15982 8928
rect 15924 8919 15982 8925
rect 18598 8916 18604 8928
rect 18656 8916 18662 8968
rect 19058 8916 19064 8968
rect 19116 8956 19122 8968
rect 19245 8959 19303 8965
rect 19245 8956 19257 8959
rect 19116 8928 19257 8956
rect 19116 8916 19122 8928
rect 19245 8925 19257 8928
rect 19291 8925 19303 8959
rect 19352 8956 19380 8996
rect 21266 8984 21272 8996
rect 21324 8984 21330 9036
rect 21085 8959 21143 8965
rect 21085 8956 21097 8959
rect 19352 8928 21097 8956
rect 19245 8919 19303 8925
rect 21085 8925 21097 8928
rect 21131 8925 21143 8959
rect 21085 8919 21143 8925
rect 15252 8860 15700 8888
rect 15252 8848 15258 8860
rect 16022 8848 16028 8900
rect 16080 8888 16086 8900
rect 17589 8891 17647 8897
rect 17589 8888 17601 8891
rect 16080 8860 17601 8888
rect 16080 8848 16086 8860
rect 17589 8857 17601 8860
rect 17635 8857 17647 8891
rect 17589 8851 17647 8857
rect 18138 8848 18144 8900
rect 18196 8888 18202 8900
rect 18417 8891 18475 8897
rect 18417 8888 18429 8891
rect 18196 8860 18429 8888
rect 18196 8848 18202 8860
rect 18417 8857 18429 8860
rect 18463 8857 18475 8891
rect 18966 8888 18972 8900
rect 18927 8860 18972 8888
rect 18417 8851 18475 8857
rect 18966 8848 18972 8860
rect 19024 8848 19030 8900
rect 19490 8891 19548 8897
rect 19490 8888 19502 8891
rect 19076 8860 19502 8888
rect 13955 8792 15148 8820
rect 13955 8789 13967 8792
rect 13909 8783 13967 8789
rect 15286 8780 15292 8832
rect 15344 8820 15350 8832
rect 15473 8823 15531 8829
rect 15473 8820 15485 8823
rect 15344 8792 15485 8820
rect 15344 8780 15350 8792
rect 15473 8789 15485 8792
rect 15519 8789 15531 8823
rect 15473 8783 15531 8789
rect 15746 8780 15752 8832
rect 15804 8820 15810 8832
rect 16114 8820 16120 8832
rect 15804 8792 16120 8820
rect 15804 8780 15810 8792
rect 16114 8780 16120 8792
rect 16172 8780 16178 8832
rect 17497 8823 17555 8829
rect 17497 8789 17509 8823
rect 17543 8820 17555 8823
rect 17957 8823 18015 8829
rect 17957 8820 17969 8823
rect 17543 8792 17969 8820
rect 17543 8789 17555 8792
rect 17497 8783 17555 8789
rect 17957 8789 17969 8792
rect 18003 8789 18015 8823
rect 18322 8820 18328 8832
rect 18283 8792 18328 8820
rect 17957 8783 18015 8789
rect 18322 8780 18328 8792
rect 18380 8780 18386 8832
rect 18782 8780 18788 8832
rect 18840 8820 18846 8832
rect 19076 8820 19104 8860
rect 19490 8857 19502 8860
rect 19536 8857 19548 8891
rect 19490 8851 19548 8857
rect 19886 8848 19892 8900
rect 19944 8888 19950 8900
rect 21542 8888 21548 8900
rect 19944 8860 21548 8888
rect 19944 8848 19950 8860
rect 21542 8848 21548 8860
rect 21600 8848 21606 8900
rect 18840 8792 19104 8820
rect 18840 8780 18846 8792
rect 19242 8780 19248 8832
rect 19300 8820 19306 8832
rect 19794 8820 19800 8832
rect 19300 8792 19800 8820
rect 19300 8780 19306 8792
rect 19794 8780 19800 8792
rect 19852 8780 19858 8832
rect 20622 8820 20628 8832
rect 20583 8792 20628 8820
rect 20622 8780 20628 8792
rect 20680 8780 20686 8832
rect 21174 8780 21180 8832
rect 21232 8820 21238 8832
rect 21232 8792 21277 8820
rect 21232 8780 21238 8792
rect 1104 8730 22056 8752
rect 1104 8678 6148 8730
rect 6200 8678 6212 8730
rect 6264 8678 6276 8730
rect 6328 8678 6340 8730
rect 6392 8678 6404 8730
rect 6456 8678 11346 8730
rect 11398 8678 11410 8730
rect 11462 8678 11474 8730
rect 11526 8678 11538 8730
rect 11590 8678 11602 8730
rect 11654 8678 16544 8730
rect 16596 8678 16608 8730
rect 16660 8678 16672 8730
rect 16724 8678 16736 8730
rect 16788 8678 16800 8730
rect 16852 8678 21742 8730
rect 21794 8678 21806 8730
rect 21858 8678 21870 8730
rect 21922 8678 21934 8730
rect 21986 8678 21998 8730
rect 22050 8678 22056 8730
rect 1104 8656 22056 8678
rect 1489 8619 1547 8625
rect 1489 8585 1501 8619
rect 1535 8616 1547 8619
rect 2130 8616 2136 8628
rect 1535 8588 2136 8616
rect 1535 8585 1547 8588
rect 1489 8579 1547 8585
rect 2130 8576 2136 8588
rect 2188 8576 2194 8628
rect 2314 8616 2320 8628
rect 2275 8588 2320 8616
rect 2314 8576 2320 8588
rect 2372 8576 2378 8628
rect 2406 8576 2412 8628
rect 2464 8616 2470 8628
rect 2869 8619 2927 8625
rect 2464 8588 2509 8616
rect 2464 8576 2470 8588
rect 2869 8585 2881 8619
rect 2915 8616 2927 8619
rect 3142 8616 3148 8628
rect 2915 8588 3148 8616
rect 2915 8585 2927 8588
rect 2869 8579 2927 8585
rect 3142 8576 3148 8588
rect 3200 8616 3206 8628
rect 3326 8616 3332 8628
rect 3200 8588 3332 8616
rect 3200 8576 3206 8588
rect 3326 8576 3332 8588
rect 3384 8576 3390 8628
rect 3878 8616 3884 8628
rect 3839 8588 3884 8616
rect 3878 8576 3884 8588
rect 3936 8576 3942 8628
rect 3973 8619 4031 8625
rect 3973 8585 3985 8619
rect 4019 8616 4031 8619
rect 4433 8619 4491 8625
rect 4433 8616 4445 8619
rect 4019 8588 4445 8616
rect 4019 8585 4031 8588
rect 3973 8579 4031 8585
rect 4433 8585 4445 8588
rect 4479 8585 4491 8619
rect 4433 8579 4491 8585
rect 4706 8576 4712 8628
rect 4764 8616 4770 8628
rect 5261 8619 5319 8625
rect 5261 8616 5273 8619
rect 4764 8588 5273 8616
rect 4764 8576 4770 8588
rect 5261 8585 5273 8588
rect 5307 8585 5319 8619
rect 5626 8616 5632 8628
rect 5587 8588 5632 8616
rect 5261 8579 5319 8585
rect 5626 8576 5632 8588
rect 5684 8576 5690 8628
rect 6086 8576 6092 8628
rect 6144 8576 6150 8628
rect 6181 8619 6239 8625
rect 6181 8585 6193 8619
rect 6227 8616 6239 8619
rect 7006 8616 7012 8628
rect 6227 8588 7012 8616
rect 6227 8585 6239 8588
rect 6181 8579 6239 8585
rect 7006 8576 7012 8588
rect 7064 8576 7070 8628
rect 7558 8576 7564 8628
rect 7616 8616 7622 8628
rect 7745 8619 7803 8625
rect 7745 8616 7757 8619
rect 7616 8588 7757 8616
rect 7616 8576 7622 8588
rect 7745 8585 7757 8588
rect 7791 8585 7803 8619
rect 7745 8579 7803 8585
rect 8018 8576 8024 8628
rect 8076 8616 8082 8628
rect 9217 8619 9275 8625
rect 9217 8616 9229 8619
rect 8076 8588 9229 8616
rect 8076 8576 8082 8588
rect 9217 8585 9229 8588
rect 9263 8585 9275 8619
rect 9582 8616 9588 8628
rect 9543 8588 9588 8616
rect 9217 8579 9275 8585
rect 9582 8576 9588 8588
rect 9640 8576 9646 8628
rect 10134 8616 10140 8628
rect 10095 8588 10140 8616
rect 10134 8576 10140 8588
rect 10192 8576 10198 8628
rect 10502 8616 10508 8628
rect 10463 8588 10508 8616
rect 10502 8576 10508 8588
rect 10560 8576 10566 8628
rect 10594 8576 10600 8628
rect 10652 8616 10658 8628
rect 10965 8619 11023 8625
rect 10965 8616 10977 8619
rect 10652 8588 10977 8616
rect 10652 8576 10658 8588
rect 10965 8585 10977 8588
rect 11011 8585 11023 8619
rect 10965 8579 11023 8585
rect 11333 8619 11391 8625
rect 11333 8585 11345 8619
rect 11379 8616 11391 8619
rect 12894 8616 12900 8628
rect 11379 8588 12900 8616
rect 11379 8585 11391 8588
rect 11333 8579 11391 8585
rect 12894 8576 12900 8588
rect 12952 8576 12958 8628
rect 12989 8619 13047 8625
rect 12989 8585 13001 8619
rect 13035 8616 13047 8619
rect 13262 8616 13268 8628
rect 13035 8588 13268 8616
rect 13035 8585 13047 8588
rect 12989 8579 13047 8585
rect 13262 8576 13268 8588
rect 13320 8576 13326 8628
rect 13814 8576 13820 8628
rect 13872 8616 13878 8628
rect 14645 8619 14703 8625
rect 14645 8616 14657 8619
rect 13872 8588 14657 8616
rect 13872 8576 13878 8588
rect 14645 8585 14657 8588
rect 14691 8616 14703 8619
rect 15381 8619 15439 8625
rect 15381 8616 15393 8619
rect 14691 8588 15393 8616
rect 14691 8585 14703 8588
rect 14645 8579 14703 8585
rect 15381 8585 15393 8588
rect 15427 8585 15439 8619
rect 15381 8579 15439 8585
rect 15749 8619 15807 8625
rect 15749 8585 15761 8619
rect 15795 8616 15807 8619
rect 18046 8616 18052 8628
rect 15795 8588 18052 8616
rect 15795 8585 15807 8588
rect 15749 8579 15807 8585
rect 18046 8576 18052 8588
rect 18104 8576 18110 8628
rect 18322 8616 18328 8628
rect 18283 8588 18328 8616
rect 18322 8576 18328 8588
rect 18380 8576 18386 8628
rect 18414 8576 18420 8628
rect 18472 8616 18478 8628
rect 18693 8619 18751 8625
rect 18693 8616 18705 8619
rect 18472 8588 18705 8616
rect 18472 8576 18478 8588
rect 18693 8585 18705 8588
rect 18739 8616 18751 8619
rect 18782 8616 18788 8628
rect 18739 8588 18788 8616
rect 18739 8585 18751 8588
rect 18693 8579 18751 8585
rect 18782 8576 18788 8588
rect 18840 8576 18846 8628
rect 18874 8576 18880 8628
rect 18932 8616 18938 8628
rect 18932 8588 19104 8616
rect 18932 8576 18938 8588
rect 3513 8551 3571 8557
rect 3513 8517 3525 8551
rect 3559 8548 3571 8551
rect 6104 8548 6132 8576
rect 3559 8520 6132 8548
rect 6632 8551 6690 8557
rect 3559 8517 3571 8520
rect 3513 8511 3571 8517
rect 6632 8517 6644 8551
rect 6678 8548 6690 8551
rect 6822 8548 6828 8560
rect 6678 8520 6828 8548
rect 6678 8517 6690 8520
rect 6632 8511 6690 8517
rect 6822 8508 6828 8520
rect 6880 8508 6886 8560
rect 7466 8508 7472 8560
rect 7524 8548 7530 8560
rect 7837 8551 7895 8557
rect 7837 8548 7849 8551
rect 7524 8520 7849 8548
rect 7524 8508 7530 8520
rect 1946 8480 1952 8492
rect 1907 8452 1952 8480
rect 1946 8440 1952 8452
rect 2004 8440 2010 8492
rect 2777 8483 2835 8489
rect 2777 8449 2789 8483
rect 2823 8480 2835 8483
rect 3142 8480 3148 8492
rect 2823 8452 3148 8480
rect 2823 8449 2835 8452
rect 2777 8443 2835 8449
rect 3142 8440 3148 8452
rect 3200 8440 3206 8492
rect 3329 8483 3387 8489
rect 3329 8449 3341 8483
rect 3375 8480 3387 8483
rect 3878 8480 3884 8492
rect 3375 8452 3884 8480
rect 3375 8449 3387 8452
rect 3329 8443 3387 8449
rect 3878 8440 3884 8452
rect 3936 8480 3942 8492
rect 4522 8480 4528 8492
rect 3936 8452 4528 8480
rect 3936 8440 3942 8452
rect 4522 8440 4528 8452
rect 4580 8440 4586 8492
rect 4798 8480 4804 8492
rect 4759 8452 4804 8480
rect 4798 8440 4804 8452
rect 4856 8440 4862 8492
rect 5721 8483 5779 8489
rect 5721 8449 5733 8483
rect 5767 8480 5779 8483
rect 6086 8480 6092 8492
rect 5767 8452 6092 8480
rect 5767 8449 5779 8452
rect 5721 8443 5779 8449
rect 6086 8440 6092 8452
rect 6144 8480 6150 8492
rect 7558 8480 7564 8492
rect 6144 8452 7564 8480
rect 6144 8440 6150 8452
rect 7558 8440 7564 8452
rect 7616 8440 7622 8492
rect 1578 8372 1584 8424
rect 1636 8412 1642 8424
rect 1673 8415 1731 8421
rect 1673 8412 1685 8415
rect 1636 8384 1685 8412
rect 1636 8372 1642 8384
rect 1673 8381 1685 8384
rect 1719 8381 1731 8415
rect 1854 8412 1860 8424
rect 1815 8384 1860 8412
rect 1673 8375 1731 8381
rect 1854 8372 1860 8384
rect 1912 8372 1918 8424
rect 3050 8412 3056 8424
rect 3011 8384 3056 8412
rect 3050 8372 3056 8384
rect 3108 8372 3114 8424
rect 3510 8372 3516 8424
rect 3568 8412 3574 8424
rect 3697 8415 3755 8421
rect 3697 8412 3709 8415
rect 3568 8384 3709 8412
rect 3568 8372 3574 8384
rect 3697 8381 3709 8384
rect 3743 8381 3755 8415
rect 3697 8375 3755 8381
rect 4614 8372 4620 8424
rect 4672 8412 4678 8424
rect 4893 8415 4951 8421
rect 4893 8412 4905 8415
rect 4672 8384 4905 8412
rect 4672 8372 4678 8384
rect 4893 8381 4905 8384
rect 4939 8381 4951 8415
rect 4893 8375 4951 8381
rect 4985 8415 5043 8421
rect 4985 8381 4997 8415
rect 5031 8412 5043 8415
rect 5258 8412 5264 8424
rect 5031 8384 5264 8412
rect 5031 8381 5043 8384
rect 4985 8375 5043 8381
rect 5258 8372 5264 8384
rect 5316 8372 5322 8424
rect 5902 8412 5908 8424
rect 5863 8384 5908 8412
rect 5902 8372 5908 8384
rect 5960 8372 5966 8424
rect 6365 8415 6423 8421
rect 6365 8381 6377 8415
rect 6411 8381 6423 8415
rect 6365 8375 6423 8381
rect 2314 8304 2320 8356
rect 2372 8344 2378 8356
rect 5074 8344 5080 8356
rect 2372 8316 5080 8344
rect 2372 8304 2378 8316
rect 5074 8304 5080 8316
rect 5132 8304 5138 8356
rect 5626 8304 5632 8356
rect 5684 8344 5690 8356
rect 6178 8344 6184 8356
rect 5684 8316 6184 8344
rect 5684 8304 5690 8316
rect 6178 8304 6184 8316
rect 6236 8304 6242 8356
rect 4246 8236 4252 8288
rect 4304 8276 4310 8288
rect 4341 8279 4399 8285
rect 4341 8276 4353 8279
rect 4304 8248 4353 8276
rect 4304 8236 4310 8248
rect 4341 8245 4353 8248
rect 4387 8245 4399 8279
rect 4341 8239 4399 8245
rect 4798 8236 4804 8288
rect 4856 8276 4862 8288
rect 5166 8276 5172 8288
rect 4856 8248 5172 8276
rect 4856 8236 4862 8248
rect 5166 8236 5172 8248
rect 5224 8276 5230 8288
rect 6380 8276 6408 8375
rect 7668 8344 7696 8520
rect 7837 8517 7849 8520
rect 7883 8517 7895 8551
rect 7837 8511 7895 8517
rect 8297 8551 8355 8557
rect 8297 8517 8309 8551
rect 8343 8548 8355 8551
rect 9600 8548 9628 8576
rect 13449 8551 13507 8557
rect 8343 8520 9628 8548
rect 9692 8520 13400 8548
rect 8343 8517 8355 8520
rect 8297 8511 8355 8517
rect 7742 8440 7748 8492
rect 7800 8480 7806 8492
rect 8021 8483 8079 8489
rect 8021 8480 8033 8483
rect 7800 8452 8033 8480
rect 7800 8440 7806 8452
rect 8021 8449 8033 8452
rect 8067 8449 8079 8483
rect 8021 8443 8079 8449
rect 8665 8483 8723 8489
rect 8665 8449 8677 8483
rect 8711 8480 8723 8483
rect 9030 8480 9036 8492
rect 8711 8452 9036 8480
rect 8711 8449 8723 8452
rect 8665 8443 8723 8449
rect 8036 8412 8064 8443
rect 9030 8440 9036 8452
rect 9088 8440 9094 8492
rect 9214 8440 9220 8492
rect 9272 8480 9278 8492
rect 9692 8480 9720 8520
rect 9272 8452 9720 8480
rect 9272 8440 9278 8452
rect 10502 8440 10508 8492
rect 10560 8480 10566 8492
rect 10873 8483 10931 8489
rect 10873 8480 10885 8483
rect 10560 8452 10885 8480
rect 10560 8440 10566 8452
rect 10873 8449 10885 8452
rect 10919 8449 10931 8483
rect 12618 8480 12624 8492
rect 12676 8489 12682 8492
rect 10873 8443 10931 8449
rect 11532 8452 12624 8480
rect 9674 8412 9680 8424
rect 8036 8384 9680 8412
rect 9674 8372 9680 8384
rect 9732 8412 9738 8424
rect 9861 8415 9919 8421
rect 9732 8384 9777 8412
rect 9732 8372 9738 8384
rect 9861 8381 9873 8415
rect 9907 8412 9919 8415
rect 10410 8412 10416 8424
rect 9907 8384 10416 8412
rect 9907 8381 9919 8384
rect 9861 8375 9919 8381
rect 10410 8372 10416 8384
rect 10468 8372 10474 8424
rect 10781 8415 10839 8421
rect 10781 8381 10793 8415
rect 10827 8412 10839 8415
rect 11532 8412 11560 8452
rect 12618 8440 12624 8452
rect 12676 8480 12688 8489
rect 12676 8452 12769 8480
rect 12676 8443 12688 8452
rect 12676 8440 12682 8443
rect 12802 8440 12808 8492
rect 12860 8480 12866 8492
rect 13372 8489 13400 8520
rect 13449 8517 13461 8551
rect 13495 8548 13507 8551
rect 13630 8548 13636 8560
rect 13495 8520 13636 8548
rect 13495 8517 13507 8520
rect 13449 8511 13507 8517
rect 13630 8508 13636 8520
rect 13688 8508 13694 8560
rect 13998 8508 14004 8560
rect 14056 8548 14062 8560
rect 15838 8548 15844 8560
rect 14056 8520 15844 8548
rect 14056 8508 14062 8520
rect 15838 8508 15844 8520
rect 15896 8548 15902 8560
rect 16206 8548 16212 8560
rect 15896 8520 16212 8548
rect 15896 8508 15902 8520
rect 16206 8508 16212 8520
rect 16264 8508 16270 8560
rect 17126 8508 17132 8560
rect 17184 8548 17190 8560
rect 17782 8551 17840 8557
rect 17782 8548 17794 8551
rect 17184 8520 17794 8548
rect 17184 8508 17190 8520
rect 17782 8517 17794 8520
rect 17828 8517 17840 8551
rect 18966 8548 18972 8560
rect 17782 8511 17840 8517
rect 18340 8520 18972 8548
rect 12897 8483 12955 8489
rect 12897 8480 12909 8483
rect 12860 8452 12909 8480
rect 12860 8440 12866 8452
rect 12897 8449 12909 8452
rect 12943 8449 12955 8483
rect 12897 8443 12955 8449
rect 13357 8483 13415 8489
rect 13357 8449 13369 8483
rect 13403 8480 13415 8483
rect 14090 8480 14096 8492
rect 13403 8452 14096 8480
rect 13403 8449 13415 8452
rect 13357 8443 13415 8449
rect 14090 8440 14096 8452
rect 14148 8440 14154 8492
rect 14918 8440 14924 8492
rect 14976 8480 14982 8492
rect 16485 8483 16543 8489
rect 14976 8452 16436 8480
rect 14976 8440 14982 8452
rect 10827 8384 11560 8412
rect 10827 8381 10839 8384
rect 10781 8375 10839 8381
rect 11606 8372 11612 8424
rect 11664 8412 11670 8424
rect 11790 8412 11796 8424
rect 11664 8384 11796 8412
rect 11664 8372 11670 8384
rect 11790 8372 11796 8384
rect 11848 8372 11854 8424
rect 12986 8372 12992 8424
rect 13044 8412 13050 8424
rect 13541 8415 13599 8421
rect 13541 8412 13553 8415
rect 13044 8384 13553 8412
rect 13044 8372 13050 8384
rect 13541 8381 13553 8384
rect 13587 8381 13599 8415
rect 13541 8375 13599 8381
rect 13630 8372 13636 8424
rect 13688 8412 13694 8424
rect 13817 8415 13875 8421
rect 13817 8412 13829 8415
rect 13688 8384 13829 8412
rect 13688 8372 13694 8384
rect 13817 8381 13829 8384
rect 13863 8412 13875 8415
rect 14734 8412 14740 8424
rect 13863 8384 14740 8412
rect 13863 8381 13875 8384
rect 13817 8375 13875 8381
rect 14734 8372 14740 8384
rect 14792 8372 14798 8424
rect 15194 8412 15200 8424
rect 15155 8384 15200 8412
rect 15194 8372 15200 8384
rect 15252 8372 15258 8424
rect 15289 8415 15347 8421
rect 15289 8381 15301 8415
rect 15335 8381 15347 8415
rect 15289 8375 15347 8381
rect 8018 8344 8024 8356
rect 7668 8316 8024 8344
rect 8018 8304 8024 8316
rect 8076 8304 8082 8356
rect 8294 8304 8300 8356
rect 8352 8344 8358 8356
rect 9122 8344 9128 8356
rect 8352 8316 9128 8344
rect 8352 8304 8358 8316
rect 9122 8304 9128 8316
rect 9180 8304 9186 8356
rect 10226 8304 10232 8356
rect 10284 8344 10290 8356
rect 10321 8347 10379 8353
rect 10321 8344 10333 8347
rect 10284 8316 10333 8344
rect 10284 8304 10290 8316
rect 10321 8313 10333 8316
rect 10367 8344 10379 8347
rect 10367 8316 12020 8344
rect 10367 8313 10379 8316
rect 10321 8307 10379 8313
rect 5224 8248 6408 8276
rect 5224 8236 5230 8248
rect 7006 8236 7012 8288
rect 7064 8276 7070 8288
rect 9766 8276 9772 8288
rect 7064 8248 9772 8276
rect 7064 8236 7070 8248
rect 9766 8236 9772 8248
rect 9824 8236 9830 8288
rect 11054 8236 11060 8288
rect 11112 8276 11118 8288
rect 11330 8276 11336 8288
rect 11112 8248 11336 8276
rect 11112 8236 11118 8248
rect 11330 8236 11336 8248
rect 11388 8236 11394 8288
rect 11517 8279 11575 8285
rect 11517 8245 11529 8279
rect 11563 8276 11575 8279
rect 11698 8276 11704 8288
rect 11563 8248 11704 8276
rect 11563 8245 11575 8248
rect 11517 8239 11575 8245
rect 11698 8236 11704 8248
rect 11756 8236 11762 8288
rect 11992 8276 12020 8316
rect 12894 8304 12900 8356
rect 12952 8344 12958 8356
rect 13998 8344 14004 8356
rect 12952 8316 14004 8344
rect 12952 8304 12958 8316
rect 13998 8304 14004 8316
rect 14056 8304 14062 8356
rect 14182 8304 14188 8356
rect 14240 8344 14246 8356
rect 14277 8347 14335 8353
rect 14277 8344 14289 8347
rect 14240 8316 14289 8344
rect 14240 8304 14246 8316
rect 14277 8313 14289 8316
rect 14323 8313 14335 8347
rect 14277 8307 14335 8313
rect 14553 8347 14611 8353
rect 14553 8313 14565 8347
rect 14599 8344 14611 8347
rect 15010 8344 15016 8356
rect 14599 8316 15016 8344
rect 14599 8313 14611 8316
rect 14553 8307 14611 8313
rect 15010 8304 15016 8316
rect 15068 8304 15074 8356
rect 13814 8276 13820 8288
rect 11992 8248 13820 8276
rect 13814 8236 13820 8248
rect 13872 8236 13878 8288
rect 14826 8236 14832 8288
rect 14884 8276 14890 8288
rect 14921 8279 14979 8285
rect 14921 8276 14933 8279
rect 14884 8248 14933 8276
rect 14884 8236 14890 8248
rect 14921 8245 14933 8248
rect 14967 8276 14979 8279
rect 15304 8276 15332 8375
rect 15562 8372 15568 8424
rect 15620 8412 15626 8424
rect 15746 8412 15752 8424
rect 15620 8384 15752 8412
rect 15620 8372 15626 8384
rect 15746 8372 15752 8384
rect 15804 8372 15810 8424
rect 16408 8412 16436 8452
rect 16485 8449 16497 8483
rect 16531 8480 16543 8483
rect 18340 8480 18368 8520
rect 18966 8508 18972 8520
rect 19024 8508 19030 8560
rect 19076 8548 19104 8588
rect 19334 8576 19340 8628
rect 19392 8616 19398 8628
rect 19886 8616 19892 8628
rect 19392 8588 19892 8616
rect 19392 8576 19398 8588
rect 19886 8576 19892 8588
rect 19944 8576 19950 8628
rect 20254 8616 20260 8628
rect 20215 8588 20260 8616
rect 20254 8576 20260 8588
rect 20312 8576 20318 8628
rect 20438 8616 20444 8628
rect 20399 8588 20444 8616
rect 20438 8576 20444 8588
rect 20496 8576 20502 8628
rect 20533 8551 20591 8557
rect 20533 8548 20545 8551
rect 19076 8520 20545 8548
rect 20533 8517 20545 8520
rect 20579 8517 20591 8551
rect 20533 8511 20591 8517
rect 16531 8452 18368 8480
rect 16531 8449 16543 8452
rect 16485 8443 16543 8449
rect 18414 8440 18420 8492
rect 18472 8480 18478 8492
rect 18472 8452 18517 8480
rect 18472 8440 18478 8452
rect 18874 8440 18880 8492
rect 18932 8480 18938 8492
rect 19242 8480 19248 8492
rect 18932 8452 19248 8480
rect 18932 8440 18938 8452
rect 19242 8440 19248 8452
rect 19300 8440 19306 8492
rect 19794 8480 19800 8492
rect 19852 8489 19858 8492
rect 19764 8452 19800 8480
rect 19794 8440 19800 8452
rect 19852 8443 19864 8489
rect 20714 8480 20720 8492
rect 20675 8452 20720 8480
rect 19852 8440 19858 8443
rect 20714 8440 20720 8452
rect 20772 8440 20778 8492
rect 16574 8412 16580 8424
rect 16408 8384 16580 8412
rect 16574 8372 16580 8384
rect 16632 8372 16638 8424
rect 18049 8415 18107 8421
rect 18049 8381 18061 8415
rect 18095 8412 18107 8415
rect 18506 8412 18512 8424
rect 18095 8384 18512 8412
rect 18095 8381 18107 8384
rect 18049 8375 18107 8381
rect 18506 8372 18512 8384
rect 18564 8372 18570 8424
rect 20073 8415 20131 8421
rect 20073 8381 20085 8415
rect 20119 8381 20131 8415
rect 20073 8375 20131 8381
rect 20993 8415 21051 8421
rect 20993 8381 21005 8415
rect 21039 8381 21051 8415
rect 20993 8375 21051 8381
rect 15654 8304 15660 8356
rect 15712 8344 15718 8356
rect 16025 8347 16083 8353
rect 16025 8344 16037 8347
rect 15712 8316 16037 8344
rect 15712 8304 15718 8316
rect 16025 8313 16037 8316
rect 16071 8313 16083 8347
rect 16298 8344 16304 8356
rect 16259 8316 16304 8344
rect 16025 8307 16083 8313
rect 16298 8304 16304 8316
rect 16356 8304 16362 8356
rect 16669 8347 16727 8353
rect 16669 8313 16681 8347
rect 16715 8344 16727 8347
rect 16942 8344 16948 8356
rect 16715 8316 16948 8344
rect 16715 8313 16727 8316
rect 16669 8307 16727 8313
rect 16942 8304 16948 8316
rect 17000 8304 17006 8356
rect 18230 8304 18236 8356
rect 18288 8344 18294 8356
rect 18601 8347 18659 8353
rect 18601 8344 18613 8347
rect 18288 8316 18613 8344
rect 18288 8304 18294 8316
rect 18601 8313 18613 8316
rect 18647 8313 18659 8347
rect 18601 8307 18659 8313
rect 15838 8276 15844 8288
rect 14967 8248 15844 8276
rect 14967 8245 14979 8248
rect 14921 8239 14979 8245
rect 15838 8236 15844 8248
rect 15896 8236 15902 8288
rect 16206 8236 16212 8288
rect 16264 8276 16270 8288
rect 18138 8276 18144 8288
rect 16264 8248 18144 8276
rect 16264 8236 16270 8248
rect 18138 8236 18144 8248
rect 18196 8236 18202 8288
rect 18690 8236 18696 8288
rect 18748 8276 18754 8288
rect 19058 8276 19064 8288
rect 18748 8248 19064 8276
rect 18748 8236 18754 8248
rect 19058 8236 19064 8248
rect 19116 8276 19122 8288
rect 20088 8276 20116 8375
rect 20714 8304 20720 8356
rect 20772 8344 20778 8356
rect 21008 8344 21036 8375
rect 20772 8316 21036 8344
rect 20772 8304 20778 8316
rect 21726 8304 21732 8356
rect 21784 8344 21790 8356
rect 22922 8344 22928 8356
rect 21784 8316 22928 8344
rect 21784 8304 21790 8316
rect 22922 8304 22928 8316
rect 22980 8304 22986 8356
rect 19116 8248 20116 8276
rect 19116 8236 19122 8248
rect 1104 8186 21896 8208
rect 1104 8134 3549 8186
rect 3601 8134 3613 8186
rect 3665 8134 3677 8186
rect 3729 8134 3741 8186
rect 3793 8134 3805 8186
rect 3857 8134 8747 8186
rect 8799 8134 8811 8186
rect 8863 8134 8875 8186
rect 8927 8134 8939 8186
rect 8991 8134 9003 8186
rect 9055 8134 13945 8186
rect 13997 8134 14009 8186
rect 14061 8134 14073 8186
rect 14125 8134 14137 8186
rect 14189 8134 14201 8186
rect 14253 8134 19143 8186
rect 19195 8134 19207 8186
rect 19259 8134 19271 8186
rect 19323 8134 19335 8186
rect 19387 8134 19399 8186
rect 19451 8134 21896 8186
rect 1104 8112 21896 8134
rect 1489 8075 1547 8081
rect 1489 8041 1501 8075
rect 1535 8072 1547 8075
rect 1762 8072 1768 8084
rect 1535 8044 1768 8072
rect 1535 8041 1547 8044
rect 1489 8035 1547 8041
rect 1762 8032 1768 8044
rect 1820 8032 1826 8084
rect 1854 8032 1860 8084
rect 1912 8072 1918 8084
rect 2317 8075 2375 8081
rect 2317 8072 2329 8075
rect 1912 8044 2329 8072
rect 1912 8032 1918 8044
rect 2317 8041 2329 8044
rect 2363 8041 2375 8075
rect 2317 8035 2375 8041
rect 2958 8032 2964 8084
rect 3016 8072 3022 8084
rect 3789 8075 3847 8081
rect 3789 8072 3801 8075
rect 3016 8044 3801 8072
rect 3016 8032 3022 8044
rect 3789 8041 3801 8044
rect 3835 8041 3847 8075
rect 3789 8035 3847 8041
rect 4982 8032 4988 8084
rect 5040 8072 5046 8084
rect 5169 8075 5227 8081
rect 5169 8072 5181 8075
rect 5040 8044 5181 8072
rect 5040 8032 5046 8044
rect 5169 8041 5181 8044
rect 5215 8041 5227 8075
rect 5169 8035 5227 8041
rect 5350 8032 5356 8084
rect 5408 8072 5414 8084
rect 5718 8072 5724 8084
rect 5408 8044 5724 8072
rect 5408 8032 5414 8044
rect 5718 8032 5724 8044
rect 5776 8072 5782 8084
rect 6549 8075 6607 8081
rect 6549 8072 6561 8075
rect 5776 8044 6561 8072
rect 5776 8032 5782 8044
rect 6549 8041 6561 8044
rect 6595 8041 6607 8075
rect 6549 8035 6607 8041
rect 7374 8032 7380 8084
rect 7432 8072 7438 8084
rect 7561 8075 7619 8081
rect 7561 8072 7573 8075
rect 7432 8044 7573 8072
rect 7432 8032 7438 8044
rect 7561 8041 7573 8044
rect 7607 8041 7619 8075
rect 7561 8035 7619 8041
rect 7742 8032 7748 8084
rect 7800 8072 7806 8084
rect 9306 8072 9312 8084
rect 7800 8044 9312 8072
rect 7800 8032 7806 8044
rect 9306 8032 9312 8044
rect 9364 8032 9370 8084
rect 9766 8032 9772 8084
rect 9824 8072 9830 8084
rect 10137 8075 10195 8081
rect 10137 8072 10149 8075
rect 9824 8044 10149 8072
rect 9824 8032 9830 8044
rect 10137 8041 10149 8044
rect 10183 8041 10195 8075
rect 10137 8035 10195 8041
rect 10597 8075 10655 8081
rect 10597 8041 10609 8075
rect 10643 8072 10655 8075
rect 11790 8072 11796 8084
rect 10643 8044 11796 8072
rect 10643 8041 10655 8044
rect 10597 8035 10655 8041
rect 11790 8032 11796 8044
rect 11848 8032 11854 8084
rect 12434 8032 12440 8084
rect 12492 8072 12498 8084
rect 13262 8072 13268 8084
rect 12492 8044 13268 8072
rect 12492 8032 12498 8044
rect 13262 8032 13268 8044
rect 13320 8032 13326 8084
rect 13906 8032 13912 8084
rect 13964 8072 13970 8084
rect 15102 8072 15108 8084
rect 13964 8044 15108 8072
rect 13964 8032 13970 8044
rect 15102 8032 15108 8044
rect 15160 8032 15166 8084
rect 15565 8075 15623 8081
rect 15565 8041 15577 8075
rect 15611 8072 15623 8075
rect 16022 8072 16028 8084
rect 15611 8044 16028 8072
rect 15611 8041 15623 8044
rect 15565 8035 15623 8041
rect 16022 8032 16028 8044
rect 16080 8032 16086 8084
rect 16114 8032 16120 8084
rect 16172 8072 16178 8084
rect 17221 8075 17279 8081
rect 17221 8072 17233 8075
rect 16172 8044 17233 8072
rect 16172 8032 16178 8044
rect 17221 8041 17233 8044
rect 17267 8072 17279 8075
rect 17310 8072 17316 8084
rect 17267 8044 17316 8072
rect 17267 8041 17279 8044
rect 17221 8035 17279 8041
rect 17310 8032 17316 8044
rect 17368 8032 17374 8084
rect 17954 8032 17960 8084
rect 18012 8072 18018 8084
rect 18325 8075 18383 8081
rect 18325 8072 18337 8075
rect 18012 8044 18337 8072
rect 18012 8032 18018 8044
rect 18325 8041 18337 8044
rect 18371 8041 18383 8075
rect 18325 8035 18383 8041
rect 18414 8032 18420 8084
rect 18472 8072 18478 8084
rect 19245 8075 19303 8081
rect 19245 8072 19257 8075
rect 18472 8044 19257 8072
rect 18472 8032 18478 8044
rect 19245 8041 19257 8044
rect 19291 8041 19303 8075
rect 19245 8035 19303 8041
rect 20349 8075 20407 8081
rect 20349 8041 20361 8075
rect 20395 8072 20407 8075
rect 20990 8072 20996 8084
rect 20395 8044 20996 8072
rect 20395 8041 20407 8044
rect 20349 8035 20407 8041
rect 20990 8032 20996 8044
rect 21048 8032 21054 8084
rect 21082 8032 21088 8084
rect 21140 8072 21146 8084
rect 21269 8075 21327 8081
rect 21269 8072 21281 8075
rect 21140 8044 21281 8072
rect 21140 8032 21146 8044
rect 21269 8041 21281 8044
rect 21315 8041 21327 8075
rect 21269 8035 21327 8041
rect 3234 8004 3240 8016
rect 1964 7976 3240 8004
rect 1964 7945 1992 7976
rect 3234 7964 3240 7976
rect 3292 8004 3298 8016
rect 5442 8004 5448 8016
rect 3292 7976 5448 8004
rect 3292 7964 3298 7976
rect 5442 7964 5448 7976
rect 5500 7964 5506 8016
rect 6270 8004 6276 8016
rect 5644 7976 6276 8004
rect 1949 7939 2007 7945
rect 1949 7905 1961 7939
rect 1995 7905 2007 7939
rect 1949 7899 2007 7905
rect 2133 7939 2191 7945
rect 2133 7905 2145 7939
rect 2179 7936 2191 7939
rect 2682 7936 2688 7948
rect 2179 7908 2688 7936
rect 2179 7905 2191 7908
rect 2133 7899 2191 7905
rect 2682 7896 2688 7908
rect 2740 7936 2746 7948
rect 2961 7939 3019 7945
rect 2961 7936 2973 7939
rect 2740 7908 2973 7936
rect 2740 7896 2746 7908
rect 2961 7905 2973 7908
rect 3007 7936 3019 7939
rect 3050 7936 3056 7948
rect 3007 7908 3056 7936
rect 3007 7905 3019 7908
rect 2961 7899 3019 7905
rect 3050 7896 3056 7908
rect 3108 7896 3114 7948
rect 3510 7896 3516 7948
rect 3568 7936 3574 7948
rect 3970 7936 3976 7948
rect 3568 7908 3976 7936
rect 3568 7896 3574 7908
rect 3970 7896 3976 7908
rect 4028 7896 4034 7948
rect 4246 7936 4252 7948
rect 4207 7908 4252 7936
rect 4246 7896 4252 7908
rect 4304 7896 4310 7948
rect 4338 7896 4344 7948
rect 4396 7936 4402 7948
rect 4396 7908 4441 7936
rect 4396 7896 4402 7908
rect 4890 7896 4896 7948
rect 4948 7936 4954 7948
rect 5166 7936 5172 7948
rect 4948 7908 5172 7936
rect 4948 7896 4954 7908
rect 5166 7896 5172 7908
rect 5224 7896 5230 7948
rect 1857 7871 1915 7877
rect 1857 7837 1869 7871
rect 1903 7868 1915 7871
rect 2038 7868 2044 7880
rect 1903 7840 2044 7868
rect 1903 7837 1915 7840
rect 1857 7831 1915 7837
rect 2038 7828 2044 7840
rect 2096 7828 2102 7880
rect 2222 7828 2228 7880
rect 2280 7868 2286 7880
rect 4617 7871 4675 7877
rect 4617 7868 4629 7871
rect 2280 7840 4629 7868
rect 2280 7828 2286 7840
rect 4617 7837 4629 7840
rect 4663 7837 4675 7871
rect 4617 7831 4675 7837
rect 4798 7828 4804 7880
rect 4856 7868 4862 7880
rect 5077 7871 5135 7877
rect 5077 7868 5089 7871
rect 4856 7840 5089 7868
rect 4856 7828 4862 7840
rect 5077 7837 5089 7840
rect 5123 7837 5135 7871
rect 5077 7831 5135 7837
rect 5442 7828 5448 7880
rect 5500 7868 5506 7880
rect 5644 7868 5672 7976
rect 6270 7964 6276 7976
rect 6328 7964 6334 8016
rect 9953 8007 10011 8013
rect 9953 8004 9965 8007
rect 6748 7976 9965 8004
rect 5721 7939 5779 7945
rect 5721 7905 5733 7939
rect 5767 7936 5779 7939
rect 5994 7936 6000 7948
rect 5767 7908 6000 7936
rect 5767 7905 5779 7908
rect 5721 7899 5779 7905
rect 5994 7896 6000 7908
rect 6052 7896 6058 7948
rect 6748 7936 6776 7976
rect 9953 7973 9965 7976
rect 9999 7973 10011 8007
rect 11238 8004 11244 8016
rect 9953 7967 10011 7973
rect 10244 7976 11244 8004
rect 6104 7908 6776 7936
rect 5500 7840 5672 7868
rect 5500 7828 5506 7840
rect 5810 7828 5816 7880
rect 5868 7868 5874 7880
rect 6104 7868 6132 7908
rect 5868 7840 6132 7868
rect 5868 7828 5874 7840
rect 6178 7828 6184 7880
rect 6236 7868 6242 7880
rect 6748 7877 6776 7908
rect 6822 7896 6828 7948
rect 6880 7936 6886 7948
rect 6917 7939 6975 7945
rect 6917 7936 6929 7939
rect 6880 7908 6929 7936
rect 6880 7896 6886 7908
rect 6917 7905 6929 7908
rect 6963 7905 6975 7939
rect 6917 7899 6975 7905
rect 7101 7939 7159 7945
rect 7101 7905 7113 7939
rect 7147 7936 7159 7939
rect 7834 7936 7840 7948
rect 7147 7908 7840 7936
rect 7147 7905 7159 7908
rect 7101 7899 7159 7905
rect 7834 7896 7840 7908
rect 7892 7896 7898 7948
rect 8110 7896 8116 7948
rect 8168 7936 8174 7948
rect 8205 7939 8263 7945
rect 8205 7936 8217 7939
rect 8168 7908 8217 7936
rect 8168 7896 8174 7908
rect 8205 7905 8217 7908
rect 8251 7905 8263 7939
rect 8205 7899 8263 7905
rect 8389 7939 8447 7945
rect 8389 7905 8401 7939
rect 8435 7936 8447 7939
rect 8754 7936 8760 7948
rect 8435 7908 8760 7936
rect 8435 7905 8447 7908
rect 8389 7899 8447 7905
rect 8754 7896 8760 7908
rect 8812 7896 8818 7948
rect 8846 7896 8852 7948
rect 8904 7936 8910 7948
rect 9493 7939 9551 7945
rect 9493 7936 9505 7939
rect 8904 7908 9505 7936
rect 8904 7896 8910 7908
rect 9493 7905 9505 7908
rect 9539 7905 9551 7939
rect 9493 7899 9551 7905
rect 6457 7871 6515 7877
rect 6236 7840 6281 7868
rect 6236 7828 6242 7840
rect 6457 7837 6469 7871
rect 6503 7868 6515 7871
rect 6733 7871 6791 7877
rect 6503 7840 6675 7868
rect 6503 7837 6515 7840
rect 6457 7831 6515 7837
rect 2590 7760 2596 7812
rect 2648 7800 2654 7812
rect 2777 7803 2835 7809
rect 2777 7800 2789 7803
rect 2648 7772 2789 7800
rect 2648 7760 2654 7772
rect 2777 7769 2789 7772
rect 2823 7769 2835 7803
rect 2777 7763 2835 7769
rect 3237 7803 3295 7809
rect 3237 7769 3249 7803
rect 3283 7769 3295 7803
rect 3237 7763 3295 7769
rect 3421 7803 3479 7809
rect 3421 7769 3433 7803
rect 3467 7800 3479 7803
rect 3786 7800 3792 7812
rect 3467 7772 3792 7800
rect 3467 7769 3479 7772
rect 3421 7763 3479 7769
rect 2498 7692 2504 7744
rect 2556 7732 2562 7744
rect 2685 7735 2743 7741
rect 2685 7732 2697 7735
rect 2556 7704 2697 7732
rect 2556 7692 2562 7704
rect 2685 7701 2697 7704
rect 2731 7701 2743 7735
rect 3252 7732 3280 7763
rect 3786 7760 3792 7772
rect 3844 7760 3850 7812
rect 3896 7772 4384 7800
rect 3510 7732 3516 7744
rect 3252 7704 3516 7732
rect 2685 7695 2743 7701
rect 3510 7692 3516 7704
rect 3568 7692 3574 7744
rect 3605 7735 3663 7741
rect 3605 7701 3617 7735
rect 3651 7732 3663 7735
rect 3896 7732 3924 7772
rect 3651 7704 3924 7732
rect 3651 7701 3663 7704
rect 3605 7695 3663 7701
rect 3970 7692 3976 7744
rect 4028 7732 4034 7744
rect 4157 7735 4215 7741
rect 4157 7732 4169 7735
rect 4028 7704 4169 7732
rect 4028 7692 4034 7704
rect 4157 7701 4169 7704
rect 4203 7701 4215 7735
rect 4356 7732 4384 7772
rect 4522 7760 4528 7812
rect 4580 7800 4586 7812
rect 5350 7800 5356 7812
rect 4580 7772 5356 7800
rect 4580 7760 4586 7772
rect 5350 7760 5356 7772
rect 5408 7760 5414 7812
rect 5537 7803 5595 7809
rect 5537 7769 5549 7803
rect 5583 7800 5595 7803
rect 6546 7800 6552 7812
rect 5583 7772 6552 7800
rect 5583 7769 5595 7772
rect 5537 7763 5595 7769
rect 6546 7760 6552 7772
rect 6604 7760 6610 7812
rect 6647 7800 6675 7840
rect 6733 7837 6745 7871
rect 6779 7837 6791 7871
rect 6733 7831 6791 7837
rect 7193 7871 7251 7877
rect 7193 7837 7205 7871
rect 7239 7868 7251 7871
rect 7742 7868 7748 7880
rect 7239 7840 7748 7868
rect 7239 7837 7251 7840
rect 7193 7831 7251 7837
rect 7742 7828 7748 7840
rect 7800 7828 7806 7880
rect 9306 7868 9312 7880
rect 9267 7840 9312 7868
rect 9306 7828 9312 7840
rect 9364 7868 9370 7880
rect 10244 7868 10272 7976
rect 11238 7964 11244 7976
rect 11296 7964 11302 8016
rect 12618 7964 12624 8016
rect 12676 8004 12682 8016
rect 12897 8007 12955 8013
rect 12897 8004 12909 8007
rect 12676 7976 12909 8004
rect 12676 7964 12682 7976
rect 12897 7973 12909 7976
rect 12943 7973 12955 8007
rect 15120 8004 15148 8032
rect 16574 8004 16580 8016
rect 15120 7976 16344 8004
rect 16535 7976 16580 8004
rect 12897 7967 12955 7973
rect 10873 7939 10931 7945
rect 10873 7905 10885 7939
rect 10919 7936 10931 7939
rect 11330 7936 11336 7948
rect 10919 7908 11336 7936
rect 10919 7905 10931 7908
rect 10873 7899 10931 7905
rect 11330 7896 11336 7908
rect 11388 7896 11394 7948
rect 12912 7936 12940 7967
rect 13633 7939 13691 7945
rect 13633 7936 13645 7939
rect 12912 7908 13645 7936
rect 13633 7905 13645 7908
rect 13679 7936 13691 7939
rect 13722 7936 13728 7948
rect 13679 7908 13728 7936
rect 13679 7905 13691 7908
rect 13633 7899 13691 7905
rect 13722 7896 13728 7908
rect 13780 7896 13786 7948
rect 13909 7939 13967 7945
rect 13909 7905 13921 7939
rect 13955 7936 13967 7939
rect 14734 7936 14740 7948
rect 13955 7908 14740 7936
rect 13955 7905 13967 7908
rect 13909 7899 13967 7905
rect 14734 7896 14740 7908
rect 14792 7896 14798 7948
rect 15013 7939 15071 7945
rect 15013 7905 15025 7939
rect 15059 7936 15071 7939
rect 15194 7936 15200 7948
rect 15059 7908 15200 7936
rect 15059 7905 15071 7908
rect 15013 7899 15071 7905
rect 15194 7896 15200 7908
rect 15252 7896 15258 7948
rect 15286 7896 15292 7948
rect 15344 7936 15350 7948
rect 16209 7939 16267 7945
rect 16209 7936 16221 7939
rect 15344 7908 16221 7936
rect 15344 7896 15350 7908
rect 16209 7905 16221 7908
rect 16255 7905 16267 7939
rect 16316 7936 16344 7976
rect 16574 7964 16580 7976
rect 16632 7964 16638 8016
rect 18233 8007 18291 8013
rect 18233 7973 18245 8007
rect 18279 8004 18291 8007
rect 20438 8004 20444 8016
rect 18279 7976 20444 8004
rect 18279 7973 18291 7976
rect 18233 7967 18291 7973
rect 20438 7964 20444 7976
rect 20496 7964 20502 8016
rect 20530 7964 20536 8016
rect 20588 8004 20594 8016
rect 21450 8004 21456 8016
rect 20588 7976 21456 8004
rect 20588 7964 20594 7976
rect 21450 7964 21456 7976
rect 21508 7964 21514 8016
rect 16669 7939 16727 7945
rect 16669 7936 16681 7939
rect 16316 7908 16681 7936
rect 16209 7899 16267 7905
rect 16669 7905 16681 7908
rect 16715 7936 16727 7939
rect 17218 7936 17224 7948
rect 16715 7908 17224 7936
rect 16715 7905 16727 7908
rect 16669 7899 16727 7905
rect 17218 7896 17224 7908
rect 17276 7896 17282 7948
rect 17681 7939 17739 7945
rect 17681 7905 17693 7939
rect 17727 7905 17739 7939
rect 17681 7899 17739 7905
rect 9364 7840 10272 7868
rect 9364 7828 9370 7840
rect 10594 7828 10600 7880
rect 10652 7868 10658 7880
rect 10778 7868 10784 7880
rect 10652 7840 10784 7868
rect 10652 7828 10658 7840
rect 10778 7828 10784 7840
rect 10836 7868 10842 7880
rect 11517 7871 11575 7877
rect 11517 7868 11529 7871
rect 10836 7840 11529 7868
rect 10836 7828 10842 7840
rect 11517 7837 11529 7840
rect 11563 7837 11575 7871
rect 12526 7868 12532 7880
rect 11517 7831 11575 7837
rect 11716 7840 12532 7868
rect 6914 7800 6920 7812
rect 6647 7772 6920 7800
rect 6914 7760 6920 7772
rect 6972 7760 6978 7812
rect 8294 7760 8300 7812
rect 8352 7800 8358 7812
rect 9401 7803 9459 7809
rect 9401 7800 9413 7803
rect 8352 7772 9413 7800
rect 8352 7760 8358 7772
rect 9401 7769 9413 7772
rect 9447 7800 9459 7803
rect 10870 7800 10876 7812
rect 9447 7772 10876 7800
rect 9447 7769 9459 7772
rect 9401 7763 9459 7769
rect 10870 7760 10876 7772
rect 10928 7760 10934 7812
rect 11057 7803 11115 7809
rect 11057 7769 11069 7803
rect 11103 7800 11115 7803
rect 11716 7800 11744 7840
rect 12526 7828 12532 7840
rect 12584 7828 12590 7880
rect 12986 7868 12992 7880
rect 12636 7840 12992 7868
rect 12636 7812 12664 7840
rect 12986 7828 12992 7840
rect 13044 7828 13050 7880
rect 13354 7868 13360 7880
rect 13315 7840 13360 7868
rect 13354 7828 13360 7840
rect 13412 7828 13418 7880
rect 14277 7871 14335 7877
rect 14277 7837 14289 7871
rect 14323 7868 14335 7871
rect 14458 7868 14464 7880
rect 14323 7840 14464 7868
rect 14323 7837 14335 7840
rect 14277 7831 14335 7837
rect 14458 7828 14464 7840
rect 14516 7828 14522 7880
rect 14642 7828 14648 7880
rect 14700 7868 14706 7880
rect 16945 7871 17003 7877
rect 14700 7840 16896 7868
rect 14700 7828 14706 7840
rect 11103 7772 11744 7800
rect 11784 7803 11842 7809
rect 11103 7769 11115 7772
rect 11057 7763 11115 7769
rect 11784 7769 11796 7803
rect 11830 7800 11842 7803
rect 12618 7800 12624 7812
rect 11830 7772 12624 7800
rect 11830 7769 11842 7772
rect 11784 7763 11842 7769
rect 12618 7760 12624 7772
rect 12676 7760 12682 7812
rect 12802 7760 12808 7812
rect 12860 7800 12866 7812
rect 14366 7800 14372 7812
rect 12860 7772 14372 7800
rect 12860 7760 12866 7772
rect 14366 7760 14372 7772
rect 14424 7760 14430 7812
rect 14737 7803 14795 7809
rect 14737 7769 14749 7803
rect 14783 7800 14795 7803
rect 16025 7803 16083 7809
rect 16025 7800 16037 7803
rect 14783 7772 16037 7800
rect 14783 7769 14795 7772
rect 14737 7763 14795 7769
rect 16025 7769 16037 7772
rect 16071 7769 16083 7803
rect 16025 7763 16083 7769
rect 16117 7803 16175 7809
rect 16117 7769 16129 7803
rect 16163 7800 16175 7803
rect 16206 7800 16212 7812
rect 16163 7772 16212 7800
rect 16163 7769 16175 7772
rect 16117 7763 16175 7769
rect 16206 7760 16212 7772
rect 16264 7760 16270 7812
rect 16868 7800 16896 7840
rect 16945 7837 16957 7871
rect 16991 7868 17003 7871
rect 17402 7868 17408 7880
rect 16991 7840 17408 7868
rect 16991 7837 17003 7840
rect 16945 7831 17003 7837
rect 17402 7828 17408 7840
rect 17460 7828 17466 7880
rect 17696 7868 17724 7899
rect 18598 7896 18604 7948
rect 18656 7936 18662 7948
rect 18877 7939 18935 7945
rect 18877 7936 18889 7939
rect 18656 7908 18889 7936
rect 18656 7896 18662 7908
rect 18877 7905 18889 7908
rect 18923 7905 18935 7939
rect 18877 7899 18935 7905
rect 19797 7939 19855 7945
rect 19797 7905 19809 7939
rect 19843 7936 19855 7939
rect 20622 7936 20628 7948
rect 19843 7908 20628 7936
rect 19843 7905 19855 7908
rect 19797 7899 19855 7905
rect 20622 7896 20628 7908
rect 20680 7896 20686 7948
rect 20717 7939 20775 7945
rect 20717 7905 20729 7939
rect 20763 7936 20775 7939
rect 20806 7936 20812 7948
rect 20763 7908 20812 7936
rect 20763 7905 20775 7908
rect 20717 7899 20775 7905
rect 20806 7896 20812 7908
rect 20864 7896 20870 7948
rect 21082 7936 21088 7948
rect 20916 7908 21088 7936
rect 18966 7868 18972 7880
rect 17696 7840 18972 7868
rect 18966 7828 18972 7840
rect 19024 7828 19030 7880
rect 19058 7828 19064 7880
rect 19116 7868 19122 7880
rect 19429 7871 19487 7877
rect 19429 7868 19441 7871
rect 19116 7840 19441 7868
rect 19116 7828 19122 7840
rect 19429 7837 19441 7840
rect 19475 7837 19487 7871
rect 19886 7868 19892 7880
rect 19847 7840 19892 7868
rect 19429 7831 19487 7837
rect 19886 7828 19892 7840
rect 19944 7828 19950 7880
rect 20916 7877 20944 7908
rect 21082 7896 21088 7908
rect 21140 7896 21146 7948
rect 19981 7871 20039 7877
rect 19981 7837 19993 7871
rect 20027 7868 20039 7871
rect 20901 7871 20959 7877
rect 20027 7840 20484 7868
rect 20027 7837 20039 7840
rect 19981 7831 20039 7837
rect 17773 7803 17831 7809
rect 17773 7800 17785 7803
rect 16868 7772 17785 7800
rect 17773 7769 17785 7772
rect 17819 7800 17831 7803
rect 18785 7803 18843 7809
rect 18785 7800 18797 7803
rect 17819 7772 18797 7800
rect 17819 7769 17831 7772
rect 17773 7763 17831 7769
rect 18785 7769 18797 7772
rect 18831 7800 18843 7803
rect 20456 7800 20484 7840
rect 20901 7837 20913 7871
rect 20947 7837 20959 7871
rect 20901 7831 20959 7837
rect 21361 7803 21419 7809
rect 21361 7800 21373 7803
rect 18831 7772 20024 7800
rect 20456 7772 21373 7800
rect 18831 7769 18843 7772
rect 18785 7763 18843 7769
rect 4706 7732 4712 7744
rect 4356 7704 4712 7732
rect 4157 7695 4215 7701
rect 4706 7692 4712 7704
rect 4764 7692 4770 7744
rect 4890 7732 4896 7744
rect 4851 7704 4896 7732
rect 4890 7692 4896 7704
rect 4948 7692 4954 7744
rect 5629 7735 5687 7741
rect 5629 7701 5641 7735
rect 5675 7732 5687 7735
rect 5810 7732 5816 7744
rect 5675 7704 5816 7732
rect 5675 7701 5687 7704
rect 5629 7695 5687 7701
rect 5810 7692 5816 7704
rect 5868 7692 5874 7744
rect 5902 7692 5908 7744
rect 5960 7732 5966 7744
rect 5997 7735 6055 7741
rect 5997 7732 6009 7735
rect 5960 7704 6009 7732
rect 5960 7692 5966 7704
rect 5997 7701 6009 7704
rect 6043 7701 6055 7735
rect 5997 7695 6055 7701
rect 6273 7735 6331 7741
rect 6273 7701 6285 7735
rect 6319 7732 6331 7735
rect 6638 7732 6644 7744
rect 6319 7704 6644 7732
rect 6319 7701 6331 7704
rect 6273 7695 6331 7701
rect 6638 7692 6644 7704
rect 6696 7692 6702 7744
rect 7742 7732 7748 7744
rect 7703 7704 7748 7732
rect 7742 7692 7748 7704
rect 7800 7692 7806 7744
rect 8110 7692 8116 7744
rect 8168 7732 8174 7744
rect 8570 7732 8576 7744
rect 8168 7704 8213 7732
rect 8531 7704 8576 7732
rect 8168 7692 8174 7704
rect 8570 7692 8576 7704
rect 8628 7692 8634 7744
rect 8662 7692 8668 7744
rect 8720 7732 8726 7744
rect 8941 7735 8999 7741
rect 8941 7732 8953 7735
rect 8720 7704 8953 7732
rect 8720 7692 8726 7704
rect 8941 7701 8953 7704
rect 8987 7701 8999 7735
rect 9766 7732 9772 7744
rect 9727 7704 9772 7732
rect 8941 7695 8999 7701
rect 9766 7692 9772 7704
rect 9824 7692 9830 7744
rect 10226 7692 10232 7744
rect 10284 7732 10290 7744
rect 10321 7735 10379 7741
rect 10321 7732 10333 7735
rect 10284 7704 10333 7732
rect 10284 7692 10290 7704
rect 10321 7701 10333 7704
rect 10367 7701 10379 7735
rect 10321 7695 10379 7701
rect 10965 7735 11023 7741
rect 10965 7701 10977 7735
rect 11011 7732 11023 7735
rect 11238 7732 11244 7744
rect 11011 7704 11244 7732
rect 11011 7701 11023 7704
rect 10965 7695 11023 7701
rect 11238 7692 11244 7704
rect 11296 7692 11302 7744
rect 11425 7735 11483 7741
rect 11425 7701 11437 7735
rect 11471 7732 11483 7735
rect 12250 7732 12256 7744
rect 11471 7704 12256 7732
rect 11471 7701 11483 7704
rect 11425 7695 11483 7701
rect 12250 7692 12256 7704
rect 12308 7692 12314 7744
rect 12986 7692 12992 7744
rect 13044 7732 13050 7744
rect 13449 7735 13507 7741
rect 13044 7704 13089 7732
rect 13044 7692 13050 7704
rect 13449 7701 13461 7735
rect 13495 7732 13507 7735
rect 13630 7732 13636 7744
rect 13495 7704 13636 7732
rect 13495 7701 13507 7704
rect 13449 7695 13507 7701
rect 13630 7692 13636 7704
rect 13688 7692 13694 7744
rect 14384 7732 14412 7760
rect 15105 7735 15163 7741
rect 15105 7732 15117 7735
rect 14384 7704 15117 7732
rect 15105 7701 15117 7704
rect 15151 7701 15163 7735
rect 15105 7695 15163 7701
rect 15197 7735 15255 7741
rect 15197 7701 15209 7735
rect 15243 7732 15255 7735
rect 15286 7732 15292 7744
rect 15243 7704 15292 7732
rect 15243 7701 15255 7704
rect 15197 7695 15255 7701
rect 15286 7692 15292 7704
rect 15344 7692 15350 7744
rect 15657 7735 15715 7741
rect 15657 7701 15669 7735
rect 15703 7732 15715 7735
rect 15930 7732 15936 7744
rect 15703 7704 15936 7732
rect 15703 7701 15715 7704
rect 15657 7695 15715 7701
rect 15930 7692 15936 7704
rect 15988 7692 15994 7744
rect 16224 7732 16252 7760
rect 17037 7735 17095 7741
rect 17037 7732 17049 7735
rect 16224 7704 17049 7732
rect 17037 7701 17049 7704
rect 17083 7701 17095 7735
rect 17037 7695 17095 7701
rect 17586 7692 17592 7744
rect 17644 7732 17650 7744
rect 17865 7735 17923 7741
rect 17865 7732 17877 7735
rect 17644 7704 17877 7732
rect 17644 7692 17650 7704
rect 17865 7701 17877 7704
rect 17911 7701 17923 7735
rect 17865 7695 17923 7701
rect 17954 7692 17960 7744
rect 18012 7732 18018 7744
rect 18693 7735 18751 7741
rect 18693 7732 18705 7735
rect 18012 7704 18705 7732
rect 18012 7692 18018 7704
rect 18693 7701 18705 7704
rect 18739 7732 18751 7735
rect 19334 7732 19340 7744
rect 18739 7704 19340 7732
rect 18739 7701 18751 7704
rect 18693 7695 18751 7701
rect 19334 7692 19340 7704
rect 19392 7692 19398 7744
rect 19996 7732 20024 7772
rect 21361 7769 21373 7772
rect 21407 7769 21419 7803
rect 21361 7763 21419 7769
rect 20714 7732 20720 7744
rect 19996 7704 20720 7732
rect 20714 7692 20720 7704
rect 20772 7692 20778 7744
rect 20809 7735 20867 7741
rect 20809 7701 20821 7735
rect 20855 7732 20867 7735
rect 21082 7732 21088 7744
rect 20855 7704 21088 7732
rect 20855 7701 20867 7704
rect 20809 7695 20867 7701
rect 21082 7692 21088 7704
rect 21140 7692 21146 7744
rect 1104 7642 22056 7664
rect 1104 7590 6148 7642
rect 6200 7590 6212 7642
rect 6264 7590 6276 7642
rect 6328 7590 6340 7642
rect 6392 7590 6404 7642
rect 6456 7590 11346 7642
rect 11398 7590 11410 7642
rect 11462 7590 11474 7642
rect 11526 7590 11538 7642
rect 11590 7590 11602 7642
rect 11654 7590 16544 7642
rect 16596 7590 16608 7642
rect 16660 7590 16672 7642
rect 16724 7590 16736 7642
rect 16788 7590 16800 7642
rect 16852 7590 21742 7642
rect 21794 7590 21806 7642
rect 21858 7590 21870 7642
rect 21922 7590 21934 7642
rect 21986 7590 21998 7642
rect 22050 7590 22056 7642
rect 1104 7568 22056 7590
rect 1578 7528 1584 7540
rect 1539 7500 1584 7528
rect 1578 7488 1584 7500
rect 1636 7488 1642 7540
rect 2406 7488 2412 7540
rect 2464 7528 2470 7540
rect 2590 7528 2596 7540
rect 2464 7500 2596 7528
rect 2464 7488 2470 7500
rect 2590 7488 2596 7500
rect 2648 7528 2654 7540
rect 4522 7528 4528 7540
rect 2648 7500 4528 7528
rect 2648 7488 2654 7500
rect 4522 7488 4528 7500
rect 4580 7488 4586 7540
rect 5166 7488 5172 7540
rect 5224 7528 5230 7540
rect 5994 7528 6000 7540
rect 5224 7500 6000 7528
rect 5224 7488 5230 7500
rect 5994 7488 6000 7500
rect 6052 7488 6058 7540
rect 6181 7531 6239 7537
rect 6181 7497 6193 7531
rect 6227 7528 6239 7531
rect 6822 7528 6828 7540
rect 6227 7500 6828 7528
rect 6227 7497 6239 7500
rect 6181 7491 6239 7497
rect 6822 7488 6828 7500
rect 6880 7488 6886 7540
rect 6914 7488 6920 7540
rect 6972 7488 6978 7540
rect 7561 7531 7619 7537
rect 7561 7497 7573 7531
rect 7607 7528 7619 7531
rect 8754 7528 8760 7540
rect 7607 7500 8760 7528
rect 7607 7497 7619 7500
rect 7561 7491 7619 7497
rect 8754 7488 8760 7500
rect 8812 7528 8818 7540
rect 10134 7528 10140 7540
rect 8812 7500 9076 7528
rect 10095 7500 10140 7528
rect 8812 7488 8818 7500
rect 2774 7420 2780 7472
rect 2832 7460 2838 7472
rect 2970 7463 3028 7469
rect 2970 7460 2982 7463
rect 2832 7432 2982 7460
rect 2832 7420 2838 7432
rect 2970 7429 2982 7432
rect 3016 7429 3028 7463
rect 4890 7460 4896 7472
rect 2970 7423 3028 7429
rect 3344 7432 4896 7460
rect 1394 7392 1400 7404
rect 1355 7364 1400 7392
rect 1394 7352 1400 7364
rect 1452 7352 1458 7404
rect 3344 7401 3372 7432
rect 4890 7420 4896 7432
rect 4948 7420 4954 7472
rect 5442 7420 5448 7472
rect 5500 7460 5506 7472
rect 6932 7460 6960 7488
rect 5500 7432 6960 7460
rect 5500 7420 5506 7432
rect 8386 7420 8392 7472
rect 8444 7460 8450 7472
rect 8444 7432 8984 7460
rect 8444 7420 8450 7432
rect 3237 7395 3295 7401
rect 3237 7361 3249 7395
rect 3283 7392 3295 7395
rect 3329 7395 3387 7401
rect 3329 7392 3341 7395
rect 3283 7364 3341 7392
rect 3283 7361 3295 7364
rect 3237 7355 3295 7361
rect 3329 7361 3341 7364
rect 3375 7361 3387 7395
rect 3329 7355 3387 7361
rect 3418 7352 3424 7404
rect 3476 7392 3482 7404
rect 3585 7395 3643 7401
rect 3585 7392 3597 7395
rect 3476 7364 3597 7392
rect 3476 7352 3482 7364
rect 3585 7361 3597 7364
rect 3631 7392 3643 7395
rect 4522 7392 4528 7404
rect 3631 7364 4528 7392
rect 3631 7361 3643 7364
rect 3585 7355 3643 7361
rect 4522 7352 4528 7364
rect 4580 7352 4586 7404
rect 4614 7352 4620 7404
rect 4672 7392 4678 7404
rect 5057 7395 5115 7401
rect 5057 7392 5069 7395
rect 4672 7364 5069 7392
rect 4672 7352 4678 7364
rect 5057 7361 5069 7364
rect 5103 7361 5115 7395
rect 5057 7355 5115 7361
rect 6733 7395 6791 7401
rect 6733 7361 6745 7395
rect 6779 7361 6791 7395
rect 6733 7355 6791 7361
rect 3436 7324 3464 7352
rect 4798 7324 4804 7336
rect 3353 7296 3464 7324
rect 4759 7296 4804 7324
rect 1857 7191 1915 7197
rect 1857 7157 1869 7191
rect 1903 7188 1915 7191
rect 3353 7188 3381 7296
rect 4798 7284 4804 7296
rect 4856 7284 4862 7336
rect 6457 7327 6515 7333
rect 6457 7293 6469 7327
rect 6503 7293 6515 7327
rect 6457 7287 6515 7293
rect 6641 7327 6699 7333
rect 6641 7293 6653 7327
rect 6687 7293 6699 7327
rect 6641 7287 6699 7293
rect 1903 7160 3381 7188
rect 1903 7157 1915 7160
rect 1857 7151 1915 7157
rect 4246 7148 4252 7200
rect 4304 7188 4310 7200
rect 4709 7191 4767 7197
rect 4709 7188 4721 7191
rect 4304 7160 4721 7188
rect 4304 7148 4310 7160
rect 4709 7157 4721 7160
rect 4755 7157 4767 7191
rect 4709 7151 4767 7157
rect 5166 7148 5172 7200
rect 5224 7188 5230 7200
rect 6472 7188 6500 7287
rect 6656 7200 6684 7287
rect 6748 7256 6776 7355
rect 6914 7352 6920 7404
rect 6972 7392 6978 7404
rect 7193 7395 7251 7401
rect 7193 7392 7205 7395
rect 6972 7364 7205 7392
rect 6972 7352 6978 7364
rect 7193 7361 7205 7364
rect 7239 7361 7251 7395
rect 7193 7355 7251 7361
rect 8294 7352 8300 7404
rect 8352 7392 8358 7404
rect 8674 7395 8732 7401
rect 8674 7392 8686 7395
rect 8352 7364 8686 7392
rect 8352 7352 8358 7364
rect 8674 7361 8686 7364
rect 8720 7392 8732 7395
rect 8846 7392 8852 7404
rect 8720 7364 8852 7392
rect 8720 7361 8732 7364
rect 8674 7355 8732 7361
rect 8846 7352 8852 7364
rect 8904 7352 8910 7404
rect 8956 7401 8984 7432
rect 9048 7401 9076 7500
rect 10134 7488 10140 7500
rect 10192 7488 10198 7540
rect 11238 7488 11244 7540
rect 11296 7528 11302 7540
rect 11793 7531 11851 7537
rect 11793 7528 11805 7531
rect 11296 7500 11805 7528
rect 11296 7488 11302 7500
rect 11793 7497 11805 7500
rect 11839 7497 11851 7531
rect 11793 7491 11851 7497
rect 12253 7531 12311 7537
rect 12253 7497 12265 7531
rect 12299 7528 12311 7531
rect 12986 7528 12992 7540
rect 12299 7500 12992 7528
rect 12299 7497 12311 7500
rect 12253 7491 12311 7497
rect 12986 7488 12992 7500
rect 13044 7488 13050 7540
rect 13630 7528 13636 7540
rect 13591 7500 13636 7528
rect 13630 7488 13636 7500
rect 13688 7488 13694 7540
rect 13725 7531 13783 7537
rect 13725 7497 13737 7531
rect 13771 7497 13783 7531
rect 13725 7491 13783 7497
rect 9674 7420 9680 7472
rect 9732 7460 9738 7472
rect 10045 7463 10103 7469
rect 10045 7460 10057 7463
rect 9732 7432 10057 7460
rect 9732 7420 9738 7432
rect 10045 7429 10057 7432
rect 10091 7460 10103 7463
rect 10318 7460 10324 7472
rect 10091 7432 10324 7460
rect 10091 7429 10103 7432
rect 10045 7423 10103 7429
rect 10318 7420 10324 7432
rect 10376 7420 10382 7472
rect 10870 7420 10876 7472
rect 10928 7460 10934 7472
rect 12161 7463 12219 7469
rect 10928 7432 11560 7460
rect 10928 7420 10934 7432
rect 8941 7395 8999 7401
rect 8941 7361 8953 7395
rect 8987 7361 8999 7395
rect 8941 7355 8999 7361
rect 9033 7395 9091 7401
rect 9033 7361 9045 7395
rect 9079 7392 9091 7395
rect 9490 7392 9496 7404
rect 9079 7364 9496 7392
rect 9079 7361 9091 7364
rect 9033 7355 9091 7361
rect 9490 7352 9496 7364
rect 9548 7352 9554 7404
rect 9858 7352 9864 7404
rect 9916 7392 9922 7404
rect 10962 7392 10968 7404
rect 9916 7364 10968 7392
rect 9916 7352 9922 7364
rect 10962 7352 10968 7364
rect 11020 7352 11026 7404
rect 11146 7392 11152 7404
rect 11107 7364 11152 7392
rect 11146 7352 11152 7364
rect 11204 7352 11210 7404
rect 11532 7401 11560 7432
rect 12161 7429 12173 7463
rect 12207 7460 12219 7463
rect 13740 7460 13768 7491
rect 14550 7488 14556 7540
rect 14608 7528 14614 7540
rect 14826 7528 14832 7540
rect 14608 7500 14832 7528
rect 14608 7488 14614 7500
rect 14826 7488 14832 7500
rect 14884 7488 14890 7540
rect 15010 7488 15016 7540
rect 15068 7528 15074 7540
rect 15286 7528 15292 7540
rect 15068 7500 15292 7528
rect 15068 7488 15074 7500
rect 15286 7488 15292 7500
rect 15344 7488 15350 7540
rect 15841 7531 15899 7537
rect 15841 7497 15853 7531
rect 15887 7528 15899 7531
rect 17129 7531 17187 7537
rect 17129 7528 17141 7531
rect 15887 7500 17141 7528
rect 15887 7497 15899 7500
rect 15841 7491 15899 7497
rect 17129 7497 17141 7500
rect 17175 7497 17187 7531
rect 17129 7491 17187 7497
rect 17865 7531 17923 7537
rect 17865 7497 17877 7531
rect 17911 7528 17923 7531
rect 18138 7528 18144 7540
rect 17911 7500 18144 7528
rect 17911 7497 17923 7500
rect 17865 7491 17923 7497
rect 18138 7488 18144 7500
rect 18196 7488 18202 7540
rect 18690 7528 18696 7540
rect 18340 7500 18696 7528
rect 12207 7432 13768 7460
rect 14016 7432 18276 7460
rect 12207 7429 12219 7432
rect 12161 7423 12219 7429
rect 11517 7395 11575 7401
rect 11517 7361 11529 7395
rect 11563 7361 11575 7395
rect 11974 7392 11980 7404
rect 11517 7355 11575 7361
rect 11624 7364 11980 7392
rect 7098 7284 7104 7336
rect 7156 7324 7162 7336
rect 7374 7324 7380 7336
rect 7156 7296 7380 7324
rect 7156 7284 7162 7296
rect 7374 7284 7380 7296
rect 7432 7284 7438 7336
rect 9306 7324 9312 7336
rect 9267 7296 9312 7324
rect 9306 7284 9312 7296
rect 9364 7284 9370 7336
rect 10597 7327 10655 7333
rect 10597 7324 10609 7327
rect 9508 7296 10609 7324
rect 6748 7228 8064 7256
rect 5224 7160 6500 7188
rect 5224 7148 5230 7160
rect 6638 7148 6644 7200
rect 6696 7148 6702 7200
rect 7098 7188 7104 7200
rect 7059 7160 7104 7188
rect 7098 7148 7104 7160
rect 7156 7148 7162 7200
rect 7377 7191 7435 7197
rect 7377 7157 7389 7191
rect 7423 7188 7435 7191
rect 7650 7188 7656 7200
rect 7423 7160 7656 7188
rect 7423 7157 7435 7160
rect 7377 7151 7435 7157
rect 7650 7148 7656 7160
rect 7708 7148 7714 7200
rect 8036 7188 8064 7228
rect 9214 7216 9220 7268
rect 9272 7256 9278 7268
rect 9508 7256 9536 7296
rect 10597 7293 10609 7296
rect 10643 7324 10655 7327
rect 11624 7324 11652 7364
rect 11974 7352 11980 7364
rect 12032 7352 12038 7404
rect 12066 7352 12072 7404
rect 12124 7392 12130 7404
rect 12250 7392 12256 7404
rect 12124 7364 12256 7392
rect 12124 7352 12130 7364
rect 12250 7352 12256 7364
rect 12308 7352 12314 7404
rect 12710 7392 12716 7404
rect 12671 7364 12716 7392
rect 12710 7352 12716 7364
rect 12768 7392 12774 7404
rect 13265 7395 13323 7401
rect 13265 7392 13277 7395
rect 12768 7364 13277 7392
rect 12768 7352 12774 7364
rect 13265 7361 13277 7364
rect 13311 7361 13323 7395
rect 13265 7355 13323 7361
rect 13538 7352 13544 7404
rect 13596 7392 13602 7404
rect 14016 7392 14044 7432
rect 13596 7364 14044 7392
rect 14093 7395 14151 7401
rect 13596 7352 13602 7364
rect 14093 7361 14105 7395
rect 14139 7392 14151 7395
rect 14550 7392 14556 7404
rect 14139 7364 14556 7392
rect 14139 7361 14151 7364
rect 14093 7355 14151 7361
rect 14550 7352 14556 7364
rect 14608 7352 14614 7404
rect 15013 7395 15071 7401
rect 15013 7361 15025 7395
rect 15059 7392 15071 7395
rect 15059 7364 15424 7392
rect 15059 7361 15071 7364
rect 15013 7355 15071 7361
rect 10643 7296 11652 7324
rect 10643 7293 10655 7296
rect 10597 7287 10655 7293
rect 11698 7284 11704 7336
rect 11756 7324 11762 7336
rect 12345 7327 12403 7333
rect 12345 7324 12357 7327
rect 11756 7296 12357 7324
rect 11756 7284 11762 7296
rect 12345 7293 12357 7296
rect 12391 7293 12403 7327
rect 12345 7287 12403 7293
rect 12618 7284 12624 7336
rect 12676 7324 12682 7336
rect 12989 7327 13047 7333
rect 12989 7324 13001 7327
rect 12676 7296 13001 7324
rect 12676 7284 12682 7296
rect 12989 7293 13001 7296
rect 13035 7293 13047 7327
rect 12989 7287 13047 7293
rect 13173 7327 13231 7333
rect 13173 7293 13185 7327
rect 13219 7293 13231 7327
rect 13173 7287 13231 7293
rect 9272 7228 9536 7256
rect 9272 7216 9278 7228
rect 9674 7216 9680 7268
rect 9732 7256 9738 7268
rect 10689 7259 10747 7265
rect 10689 7256 10701 7259
rect 9732 7228 10701 7256
rect 9732 7216 9738 7228
rect 10689 7225 10701 7228
rect 10735 7225 10747 7259
rect 10689 7219 10747 7225
rect 10870 7216 10876 7268
rect 10928 7256 10934 7268
rect 11238 7256 11244 7268
rect 10928 7228 11244 7256
rect 10928 7216 10934 7228
rect 11238 7216 11244 7228
rect 11296 7216 11302 7268
rect 11333 7259 11391 7265
rect 11333 7225 11345 7259
rect 11379 7256 11391 7259
rect 13188 7256 13216 7287
rect 13354 7284 13360 7336
rect 13412 7324 13418 7336
rect 14185 7327 14243 7333
rect 14185 7324 14197 7327
rect 13412 7296 14197 7324
rect 13412 7284 13418 7296
rect 14185 7293 14197 7296
rect 14231 7293 14243 7327
rect 14185 7287 14243 7293
rect 14277 7327 14335 7333
rect 14277 7293 14289 7327
rect 14323 7293 14335 7327
rect 14277 7287 14335 7293
rect 14829 7327 14887 7333
rect 14829 7293 14841 7327
rect 14875 7324 14887 7327
rect 14918 7324 14924 7336
rect 14875 7296 14924 7324
rect 14875 7293 14887 7296
rect 14829 7287 14887 7293
rect 13262 7256 13268 7268
rect 11379 7228 13032 7256
rect 13175 7228 13268 7256
rect 11379 7225 11391 7228
rect 11333 7219 11391 7225
rect 13004 7200 13032 7228
rect 13262 7216 13268 7228
rect 13320 7256 13326 7268
rect 13538 7256 13544 7268
rect 13320 7228 13544 7256
rect 13320 7216 13326 7228
rect 13538 7216 13544 7228
rect 13596 7216 13602 7268
rect 13722 7216 13728 7268
rect 13780 7256 13786 7268
rect 14292 7256 14320 7287
rect 14918 7284 14924 7296
rect 14976 7284 14982 7336
rect 15194 7324 15200 7336
rect 15155 7296 15200 7324
rect 15194 7284 15200 7296
rect 15252 7284 15258 7336
rect 15396 7333 15424 7364
rect 15470 7352 15476 7404
rect 15528 7392 15534 7404
rect 15528 7364 16068 7392
rect 15528 7352 15534 7364
rect 16040 7336 16068 7364
rect 16206 7352 16212 7404
rect 16264 7392 16270 7404
rect 16301 7395 16359 7401
rect 16301 7392 16313 7395
rect 16264 7364 16313 7392
rect 16264 7352 16270 7364
rect 16301 7361 16313 7364
rect 16347 7361 16359 7395
rect 16301 7355 16359 7361
rect 16390 7352 16396 7404
rect 16448 7392 16454 7404
rect 17037 7395 17095 7401
rect 17037 7392 17049 7395
rect 16448 7364 17049 7392
rect 16448 7352 16454 7364
rect 17037 7361 17049 7364
rect 17083 7361 17095 7395
rect 17037 7355 17095 7361
rect 15381 7327 15439 7333
rect 15381 7293 15393 7327
rect 15427 7324 15439 7327
rect 15838 7324 15844 7336
rect 15427 7296 15844 7324
rect 15427 7293 15439 7296
rect 15381 7287 15439 7293
rect 15838 7284 15844 7296
rect 15896 7284 15902 7336
rect 16022 7324 16028 7336
rect 15983 7296 16028 7324
rect 16022 7284 16028 7296
rect 16080 7284 16086 7336
rect 16482 7284 16488 7336
rect 16540 7324 16546 7336
rect 17221 7327 17279 7333
rect 17221 7324 17233 7327
rect 16540 7296 17233 7324
rect 16540 7284 16546 7296
rect 17221 7293 17233 7296
rect 17267 7293 17279 7327
rect 17221 7287 17279 7293
rect 17310 7284 17316 7336
rect 17368 7324 17374 7336
rect 17957 7327 18015 7333
rect 17957 7324 17969 7327
rect 17368 7296 17969 7324
rect 17368 7284 17374 7296
rect 17957 7293 17969 7296
rect 18003 7293 18015 7327
rect 18138 7324 18144 7336
rect 18099 7296 18144 7324
rect 17957 7287 18015 7293
rect 18138 7284 18144 7296
rect 18196 7284 18202 7336
rect 18248 7324 18276 7432
rect 18340 7401 18368 7500
rect 18690 7488 18696 7500
rect 18748 7488 18754 7540
rect 19705 7531 19763 7537
rect 19705 7497 19717 7531
rect 19751 7528 19763 7531
rect 19794 7528 19800 7540
rect 19751 7500 19800 7528
rect 19751 7497 19763 7500
rect 19705 7491 19763 7497
rect 19794 7488 19800 7500
rect 19852 7488 19858 7540
rect 19978 7488 19984 7540
rect 20036 7528 20042 7540
rect 20165 7531 20223 7537
rect 20165 7528 20177 7531
rect 20036 7500 20177 7528
rect 20036 7488 20042 7500
rect 20165 7497 20177 7500
rect 20211 7497 20223 7531
rect 21174 7528 21180 7540
rect 21135 7500 21180 7528
rect 20165 7491 20223 7497
rect 21174 7488 21180 7500
rect 21232 7488 21238 7540
rect 18598 7469 18604 7472
rect 18592 7460 18604 7469
rect 18559 7432 18604 7460
rect 18592 7423 18604 7432
rect 18598 7420 18604 7423
rect 18656 7420 18662 7472
rect 20254 7460 20260 7472
rect 19306 7432 20260 7460
rect 18325 7395 18383 7401
rect 18325 7361 18337 7395
rect 18371 7361 18383 7395
rect 19306 7392 19334 7432
rect 20254 7420 20260 7432
rect 20312 7420 20318 7472
rect 21450 7460 21456 7472
rect 21411 7432 21456 7460
rect 21450 7420 21456 7432
rect 21508 7420 21514 7472
rect 19978 7392 19984 7404
rect 18325 7355 18383 7361
rect 18441 7364 19334 7392
rect 19939 7364 19984 7392
rect 18441 7324 18469 7364
rect 19978 7352 19984 7364
rect 20036 7352 20042 7404
rect 20809 7395 20867 7401
rect 20809 7392 20821 7395
rect 20088 7364 20821 7392
rect 18248 7296 18469 7324
rect 19334 7284 19340 7336
rect 19392 7324 19398 7336
rect 20088 7324 20116 7364
rect 20809 7361 20821 7364
rect 20855 7392 20867 7395
rect 21082 7392 21088 7404
rect 20855 7364 21088 7392
rect 20855 7361 20867 7364
rect 20809 7355 20867 7361
rect 21082 7352 21088 7364
rect 21140 7352 21146 7404
rect 19392 7296 20116 7324
rect 20625 7327 20683 7333
rect 19392 7284 19398 7296
rect 20625 7293 20637 7327
rect 20671 7293 20683 7327
rect 20625 7287 20683 7293
rect 20717 7327 20775 7333
rect 20717 7293 20729 7327
rect 20763 7324 20775 7327
rect 20898 7324 20904 7336
rect 20763 7296 20904 7324
rect 20763 7293 20775 7296
rect 20717 7287 20775 7293
rect 13780 7228 14320 7256
rect 13780 7216 13786 7228
rect 15286 7216 15292 7268
rect 15344 7256 15350 7268
rect 16669 7259 16727 7265
rect 16669 7256 16681 7259
rect 15344 7228 16681 7256
rect 15344 7216 15350 7228
rect 16669 7225 16681 7228
rect 16715 7225 16727 7259
rect 17770 7256 17776 7268
rect 16669 7219 16727 7225
rect 17328 7228 17776 7256
rect 9858 7188 9864 7200
rect 8036 7160 9864 7188
rect 9858 7148 9864 7160
rect 9916 7148 9922 7200
rect 10413 7191 10471 7197
rect 10413 7157 10425 7191
rect 10459 7188 10471 7191
rect 10962 7188 10968 7200
rect 10459 7160 10968 7188
rect 10459 7157 10471 7160
rect 10413 7151 10471 7157
rect 10962 7148 10968 7160
rect 11020 7148 11026 7200
rect 11057 7191 11115 7197
rect 11057 7157 11069 7191
rect 11103 7188 11115 7191
rect 11606 7188 11612 7200
rect 11103 7160 11612 7188
rect 11103 7157 11115 7160
rect 11057 7151 11115 7157
rect 11606 7148 11612 7160
rect 11664 7148 11670 7200
rect 11701 7191 11759 7197
rect 11701 7157 11713 7191
rect 11747 7188 11759 7191
rect 12250 7188 12256 7200
rect 11747 7160 12256 7188
rect 11747 7157 11759 7160
rect 11701 7151 11759 7157
rect 12250 7148 12256 7160
rect 12308 7148 12314 7200
rect 12986 7148 12992 7200
rect 13044 7148 13050 7200
rect 14645 7191 14703 7197
rect 14645 7157 14657 7191
rect 14691 7188 14703 7191
rect 14826 7188 14832 7200
rect 14691 7160 14832 7188
rect 14691 7157 14703 7160
rect 14645 7151 14703 7157
rect 14826 7148 14832 7160
rect 14884 7188 14890 7200
rect 15378 7188 15384 7200
rect 14884 7160 15384 7188
rect 14884 7148 14890 7160
rect 15378 7148 15384 7160
rect 15436 7148 15442 7200
rect 16206 7188 16212 7200
rect 16167 7160 16212 7188
rect 16206 7148 16212 7160
rect 16264 7148 16270 7200
rect 16485 7191 16543 7197
rect 16485 7157 16497 7191
rect 16531 7188 16543 7191
rect 17328 7188 17356 7228
rect 17770 7216 17776 7228
rect 17828 7216 17834 7268
rect 20640 7256 20668 7287
rect 20898 7284 20904 7296
rect 20956 7324 20962 7336
rect 21174 7324 21180 7336
rect 20956 7296 21180 7324
rect 20956 7284 20962 7296
rect 21174 7284 21180 7296
rect 21232 7284 21238 7336
rect 20806 7256 20812 7268
rect 20640 7228 20812 7256
rect 20806 7216 20812 7228
rect 20864 7216 20870 7268
rect 17494 7188 17500 7200
rect 16531 7160 17356 7188
rect 17455 7160 17500 7188
rect 16531 7157 16543 7160
rect 16485 7151 16543 7157
rect 17494 7148 17500 7160
rect 17552 7148 17558 7200
rect 17678 7148 17684 7200
rect 17736 7188 17742 7200
rect 19797 7191 19855 7197
rect 19797 7188 19809 7191
rect 17736 7160 19809 7188
rect 17736 7148 17742 7160
rect 19797 7157 19809 7160
rect 19843 7157 19855 7191
rect 19797 7151 19855 7157
rect 20254 7148 20260 7200
rect 20312 7188 20318 7200
rect 21361 7191 21419 7197
rect 21361 7188 21373 7191
rect 20312 7160 21373 7188
rect 20312 7148 20318 7160
rect 21361 7157 21373 7160
rect 21407 7157 21419 7191
rect 21361 7151 21419 7157
rect 1104 7098 21896 7120
rect 1104 7046 3549 7098
rect 3601 7046 3613 7098
rect 3665 7046 3677 7098
rect 3729 7046 3741 7098
rect 3793 7046 3805 7098
rect 3857 7046 8747 7098
rect 8799 7046 8811 7098
rect 8863 7046 8875 7098
rect 8927 7046 8939 7098
rect 8991 7046 9003 7098
rect 9055 7046 13945 7098
rect 13997 7046 14009 7098
rect 14061 7046 14073 7098
rect 14125 7046 14137 7098
rect 14189 7046 14201 7098
rect 14253 7046 19143 7098
rect 19195 7046 19207 7098
rect 19259 7046 19271 7098
rect 19323 7046 19335 7098
rect 19387 7046 19399 7098
rect 19451 7046 21896 7098
rect 1104 7024 21896 7046
rect 3602 6984 3608 6996
rect 3563 6956 3608 6984
rect 3602 6944 3608 6956
rect 3660 6944 3666 6996
rect 3789 6987 3847 6993
rect 3789 6953 3801 6987
rect 3835 6984 3847 6987
rect 3970 6984 3976 6996
rect 3835 6956 3976 6984
rect 3835 6953 3847 6956
rect 3789 6947 3847 6953
rect 3970 6944 3976 6956
rect 4028 6944 4034 6996
rect 5074 6944 5080 6996
rect 5132 6984 5138 6996
rect 10226 6984 10232 6996
rect 5132 6956 10232 6984
rect 5132 6944 5138 6956
rect 10226 6944 10232 6956
rect 10284 6944 10290 6996
rect 10870 6944 10876 6996
rect 10928 6984 10934 6996
rect 12161 6987 12219 6993
rect 12161 6984 12173 6987
rect 10928 6956 12173 6984
rect 10928 6944 10934 6956
rect 12161 6953 12173 6956
rect 12207 6984 12219 6987
rect 12802 6984 12808 6996
rect 12207 6956 12808 6984
rect 12207 6953 12219 6956
rect 12161 6947 12219 6953
rect 12802 6944 12808 6956
rect 12860 6944 12866 6996
rect 13173 6987 13231 6993
rect 13173 6953 13185 6987
rect 13219 6984 13231 6987
rect 13354 6984 13360 6996
rect 13219 6956 13360 6984
rect 13219 6953 13231 6956
rect 13173 6947 13231 6953
rect 13354 6944 13360 6956
rect 13412 6944 13418 6996
rect 14458 6984 14464 6996
rect 13832 6956 14464 6984
rect 4522 6916 4528 6928
rect 4448 6888 4528 6916
rect 566 6808 572 6860
rect 624 6848 630 6860
rect 1486 6848 1492 6860
rect 624 6820 1492 6848
rect 624 6808 630 6820
rect 1486 6808 1492 6820
rect 1544 6808 1550 6860
rect 1949 6851 2007 6857
rect 1949 6817 1961 6851
rect 1995 6848 2007 6851
rect 2498 6848 2504 6860
rect 1995 6820 2504 6848
rect 1995 6817 2007 6820
rect 1949 6811 2007 6817
rect 2498 6808 2504 6820
rect 2556 6808 2562 6860
rect 2774 6808 2780 6860
rect 2832 6848 2838 6860
rect 2961 6851 3019 6857
rect 2961 6848 2973 6851
rect 2832 6820 2973 6848
rect 2832 6808 2838 6820
rect 2961 6817 2973 6820
rect 3007 6817 3019 6851
rect 2961 6811 3019 6817
rect 3602 6808 3608 6860
rect 3660 6848 3666 6860
rect 4448 6857 4476 6888
rect 4522 6876 4528 6888
rect 4580 6876 4586 6928
rect 4617 6919 4675 6925
rect 4617 6885 4629 6919
rect 4663 6885 4675 6919
rect 5902 6916 5908 6928
rect 4617 6879 4675 6885
rect 5552 6888 5908 6916
rect 4249 6851 4307 6857
rect 4249 6848 4261 6851
rect 3660 6820 4261 6848
rect 3660 6808 3666 6820
rect 4249 6817 4261 6820
rect 4295 6817 4307 6851
rect 4249 6811 4307 6817
rect 4433 6851 4491 6857
rect 4433 6817 4445 6851
rect 4479 6817 4491 6851
rect 4433 6811 4491 6817
rect 2130 6740 2136 6792
rect 2188 6780 2194 6792
rect 2225 6783 2283 6789
rect 2225 6780 2237 6783
rect 2188 6752 2237 6780
rect 2188 6740 2194 6752
rect 2225 6749 2237 6752
rect 2271 6780 2283 6783
rect 2866 6780 2872 6792
rect 2271 6752 2872 6780
rect 2271 6749 2283 6752
rect 2225 6743 2283 6749
rect 2866 6740 2872 6752
rect 2924 6740 2930 6792
rect 3142 6780 3148 6792
rect 3103 6752 3148 6780
rect 3142 6740 3148 6752
rect 3200 6740 3206 6792
rect 3234 6740 3240 6792
rect 3292 6780 3298 6792
rect 3418 6780 3424 6792
rect 3292 6752 3424 6780
rect 3292 6740 3298 6752
rect 3418 6740 3424 6752
rect 3476 6740 3482 6792
rect 14 6672 20 6724
rect 72 6712 78 6724
rect 934 6712 940 6724
rect 72 6684 940 6712
rect 72 6672 78 6684
rect 934 6672 940 6684
rect 992 6712 998 6724
rect 2409 6715 2467 6721
rect 2409 6712 2421 6715
rect 992 6684 2421 6712
rect 992 6672 998 6684
rect 2409 6681 2421 6684
rect 2455 6681 2467 6715
rect 2590 6712 2596 6724
rect 2551 6684 2596 6712
rect 2409 6675 2467 6681
rect 2590 6672 2596 6684
rect 2648 6672 2654 6724
rect 3878 6672 3884 6724
rect 3936 6712 3942 6724
rect 4062 6712 4068 6724
rect 3936 6684 4068 6712
rect 3936 6672 3942 6684
rect 4062 6672 4068 6684
rect 4120 6672 4126 6724
rect 4157 6715 4215 6721
rect 4157 6681 4169 6715
rect 4203 6712 4215 6715
rect 4632 6712 4660 6879
rect 5258 6848 5264 6860
rect 5219 6820 5264 6848
rect 5258 6808 5264 6820
rect 5316 6808 5322 6860
rect 5074 6740 5080 6792
rect 5132 6780 5138 6792
rect 5552 6780 5580 6888
rect 5902 6876 5908 6888
rect 5960 6876 5966 6928
rect 8294 6876 8300 6928
rect 8352 6916 8358 6928
rect 8757 6919 8815 6925
rect 8352 6888 8524 6916
rect 8352 6876 8358 6888
rect 5626 6808 5632 6860
rect 5684 6848 5690 6860
rect 5997 6851 6055 6857
rect 5997 6848 6009 6851
rect 5684 6820 6009 6848
rect 5684 6808 5690 6820
rect 5997 6817 6009 6820
rect 6043 6817 6055 6851
rect 7006 6848 7012 6860
rect 5997 6811 6055 6817
rect 6472 6820 7012 6848
rect 6472 6792 6500 6820
rect 7006 6808 7012 6820
rect 7064 6808 7070 6860
rect 8205 6851 8263 6857
rect 8205 6817 8217 6851
rect 8251 6848 8263 6851
rect 8386 6848 8392 6860
rect 8251 6820 8392 6848
rect 8251 6817 8263 6820
rect 8205 6811 8263 6817
rect 8386 6808 8392 6820
rect 8444 6808 8450 6860
rect 5905 6783 5963 6789
rect 5905 6780 5917 6783
rect 5132 6752 5917 6780
rect 5132 6740 5138 6752
rect 5905 6749 5917 6752
rect 5951 6749 5963 6783
rect 6454 6780 6460 6792
rect 6415 6752 6460 6780
rect 5905 6743 5963 6749
rect 6454 6740 6460 6752
rect 6512 6740 6518 6792
rect 6549 6783 6607 6789
rect 6549 6749 6561 6783
rect 6595 6749 6607 6783
rect 8496 6780 8524 6888
rect 8757 6885 8769 6919
rect 8803 6885 8815 6919
rect 10134 6916 10140 6928
rect 8757 6879 8815 6885
rect 9600 6888 10140 6916
rect 8772 6848 8800 6879
rect 8846 6848 8852 6860
rect 8772 6820 8852 6848
rect 8846 6808 8852 6820
rect 8904 6808 8910 6860
rect 9490 6848 9496 6860
rect 9451 6820 9496 6848
rect 9490 6808 9496 6820
rect 9548 6808 9554 6860
rect 6549 6743 6607 6749
rect 6840 6752 8524 6780
rect 6564 6712 6592 6743
rect 4203 6684 4660 6712
rect 4816 6684 6592 6712
rect 4203 6681 4215 6684
rect 4157 6675 4215 6681
rect 2130 6604 2136 6656
rect 2188 6644 2194 6656
rect 2685 6647 2743 6653
rect 2685 6644 2697 6647
rect 2188 6616 2697 6644
rect 2188 6604 2194 6616
rect 2685 6613 2697 6616
rect 2731 6644 2743 6647
rect 4816 6644 4844 6684
rect 4982 6644 4988 6656
rect 2731 6616 4844 6644
rect 4943 6616 4988 6644
rect 2731 6613 2743 6616
rect 2685 6607 2743 6613
rect 4982 6604 4988 6616
rect 5040 6604 5046 6656
rect 5074 6604 5080 6656
rect 5132 6644 5138 6656
rect 5132 6616 5177 6644
rect 5132 6604 5138 6616
rect 5258 6604 5264 6656
rect 5316 6644 5322 6656
rect 5445 6647 5503 6653
rect 5445 6644 5457 6647
rect 5316 6616 5457 6644
rect 5316 6604 5322 6616
rect 5445 6613 5457 6616
rect 5491 6613 5503 6647
rect 5810 6644 5816 6656
rect 5771 6616 5816 6644
rect 5445 6607 5503 6613
rect 5810 6604 5816 6616
rect 5868 6604 5874 6656
rect 6273 6647 6331 6653
rect 6273 6613 6285 6647
rect 6319 6644 6331 6647
rect 6546 6644 6552 6656
rect 6319 6616 6552 6644
rect 6319 6613 6331 6616
rect 6273 6607 6331 6613
rect 6546 6604 6552 6616
rect 6604 6604 6610 6656
rect 6638 6604 6644 6656
rect 6696 6644 6702 6656
rect 6840 6653 6868 6752
rect 8570 6740 8576 6792
rect 8628 6780 8634 6792
rect 9309 6783 9367 6789
rect 8628 6752 8721 6780
rect 8628 6740 8634 6752
rect 9309 6749 9321 6783
rect 9355 6780 9367 6783
rect 9600 6780 9628 6888
rect 10134 6876 10140 6888
rect 10192 6876 10198 6928
rect 11606 6876 11612 6928
rect 11664 6916 11670 6928
rect 11885 6919 11943 6925
rect 11664 6888 11836 6916
rect 11664 6876 11670 6888
rect 9355 6752 9628 6780
rect 9355 6749 9367 6752
rect 9309 6743 9367 6749
rect 10042 6740 10048 6792
rect 10100 6780 10106 6792
rect 10594 6780 10600 6792
rect 10100 6752 10600 6780
rect 10100 6740 10106 6752
rect 10594 6740 10600 6752
rect 10652 6780 10658 6792
rect 11241 6783 11299 6789
rect 11241 6780 11253 6783
rect 10652 6752 11253 6780
rect 10652 6740 10658 6752
rect 11241 6749 11253 6752
rect 11287 6749 11299 6783
rect 11241 6743 11299 6749
rect 11517 6783 11575 6789
rect 11517 6749 11529 6783
rect 11563 6780 11575 6783
rect 11563 6752 11597 6780
rect 11563 6749 11575 6752
rect 11517 6743 11575 6749
rect 7938 6715 7996 6721
rect 7938 6681 7950 6715
rect 7984 6681 7996 6715
rect 7938 6675 7996 6681
rect 6733 6647 6791 6653
rect 6733 6644 6745 6647
rect 6696 6616 6745 6644
rect 6696 6604 6702 6616
rect 6733 6613 6745 6616
rect 6779 6613 6791 6647
rect 6733 6607 6791 6613
rect 6825 6647 6883 6653
rect 6825 6613 6837 6647
rect 6871 6613 6883 6647
rect 6825 6607 6883 6613
rect 7282 6604 7288 6656
rect 7340 6644 7346 6656
rect 7558 6644 7564 6656
rect 7340 6616 7564 6644
rect 7340 6604 7346 6616
rect 7558 6604 7564 6616
rect 7616 6604 7622 6656
rect 7944 6644 7972 6675
rect 8110 6672 8116 6724
rect 8168 6712 8174 6724
rect 8297 6715 8355 6721
rect 8297 6712 8309 6715
rect 8168 6684 8309 6712
rect 8168 6672 8174 6684
rect 8297 6681 8309 6684
rect 8343 6681 8355 6715
rect 8297 6675 8355 6681
rect 8386 6672 8392 6724
rect 8444 6712 8450 6724
rect 8588 6712 8616 6740
rect 8444 6684 8616 6712
rect 8680 6684 9904 6712
rect 8444 6672 8450 6684
rect 8680 6644 8708 6684
rect 9876 6656 9904 6684
rect 10686 6672 10692 6724
rect 10744 6712 10750 6724
rect 10974 6715 11032 6721
rect 10974 6712 10986 6715
rect 10744 6684 10986 6712
rect 10744 6672 10750 6684
rect 10974 6681 10986 6684
rect 11020 6681 11032 6715
rect 11532 6712 11560 6743
rect 11808 6724 11836 6888
rect 11885 6885 11897 6919
rect 11931 6916 11943 6919
rect 11974 6916 11980 6928
rect 11931 6888 11980 6916
rect 11931 6885 11943 6888
rect 11885 6879 11943 6885
rect 11974 6876 11980 6888
rect 12032 6876 12038 6928
rect 13832 6916 13860 6956
rect 14458 6944 14464 6956
rect 14516 6944 14522 6996
rect 15102 6944 15108 6996
rect 15160 6984 15166 6996
rect 15160 6956 16712 6984
rect 15160 6944 15166 6956
rect 12452 6888 13860 6916
rect 11992 6848 12020 6876
rect 12158 6848 12164 6860
rect 11992 6820 12164 6848
rect 12158 6808 12164 6820
rect 12216 6808 12222 6860
rect 11609 6715 11667 6721
rect 11609 6712 11621 6715
rect 10974 6675 11032 6681
rect 11164 6684 11621 6712
rect 8938 6644 8944 6656
rect 7944 6616 8708 6644
rect 8899 6616 8944 6644
rect 8938 6604 8944 6616
rect 8996 6604 9002 6656
rect 9401 6647 9459 6653
rect 9401 6613 9413 6647
rect 9447 6644 9459 6647
rect 9582 6644 9588 6656
rect 9447 6616 9588 6644
rect 9447 6613 9459 6616
rect 9401 6607 9459 6613
rect 9582 6604 9588 6616
rect 9640 6604 9646 6656
rect 9858 6644 9864 6656
rect 9771 6616 9864 6644
rect 9858 6604 9864 6616
rect 9916 6604 9922 6656
rect 10410 6604 10416 6656
rect 10468 6644 10474 6656
rect 11164 6644 11192 6684
rect 11609 6681 11621 6684
rect 11655 6681 11667 6715
rect 11609 6675 11667 6681
rect 11790 6672 11796 6724
rect 11848 6672 11854 6724
rect 12069 6715 12127 6721
rect 12069 6681 12081 6715
rect 12115 6712 12127 6715
rect 12342 6712 12348 6724
rect 12115 6684 12348 6712
rect 12115 6681 12127 6684
rect 12069 6675 12127 6681
rect 12342 6672 12348 6684
rect 12400 6712 12406 6724
rect 12452 6712 12480 6888
rect 12618 6848 12624 6860
rect 12579 6820 12624 6848
rect 12618 6808 12624 6820
rect 12676 6808 12682 6860
rect 13078 6808 13084 6860
rect 13136 6848 13142 6860
rect 13633 6851 13691 6857
rect 13633 6848 13645 6851
rect 13136 6820 13645 6848
rect 13136 6808 13142 6820
rect 13633 6817 13645 6820
rect 13679 6817 13691 6851
rect 13633 6811 13691 6817
rect 15562 6808 15568 6860
rect 15620 6848 15626 6860
rect 16209 6851 16267 6857
rect 16209 6848 16221 6851
rect 15620 6820 16221 6848
rect 15620 6808 15626 6820
rect 16209 6817 16221 6820
rect 16255 6848 16267 6851
rect 16482 6848 16488 6860
rect 16255 6820 16488 6848
rect 16255 6817 16267 6820
rect 16209 6811 16267 6817
rect 16482 6808 16488 6820
rect 16540 6808 16546 6860
rect 12713 6783 12771 6789
rect 12713 6749 12725 6783
rect 12759 6780 12771 6783
rect 14090 6780 14096 6792
rect 12759 6752 13676 6780
rect 14051 6752 14096 6780
rect 12759 6749 12771 6752
rect 12713 6743 12771 6749
rect 13538 6712 13544 6724
rect 12400 6684 12480 6712
rect 13372 6684 13544 6712
rect 12400 6672 12406 6684
rect 13372 6656 13400 6684
rect 13538 6672 13544 6684
rect 13596 6672 13602 6724
rect 13648 6656 13676 6752
rect 14090 6740 14096 6752
rect 14148 6740 14154 6792
rect 15102 6740 15108 6792
rect 15160 6780 15166 6792
rect 16393 6783 16451 6789
rect 16393 6780 16405 6783
rect 15160 6752 16405 6780
rect 15160 6740 15166 6752
rect 16393 6749 16405 6752
rect 16439 6749 16451 6783
rect 16393 6743 16451 6749
rect 13814 6672 13820 6724
rect 13872 6712 13878 6724
rect 14338 6715 14396 6721
rect 14338 6712 14350 6715
rect 13872 6684 14350 6712
rect 13872 6672 13878 6684
rect 14338 6681 14350 6684
rect 14384 6712 14396 6715
rect 15194 6712 15200 6724
rect 14384 6684 15200 6712
rect 14384 6681 14396 6684
rect 14338 6675 14396 6681
rect 15194 6672 15200 6684
rect 15252 6672 15258 6724
rect 15930 6712 15936 6724
rect 15891 6684 15936 6712
rect 15930 6672 15936 6684
rect 15988 6672 15994 6724
rect 16684 6712 16712 6956
rect 18322 6944 18328 6996
rect 18380 6984 18386 6996
rect 19978 6984 19984 6996
rect 18380 6956 18920 6984
rect 19939 6956 19984 6984
rect 18380 6944 18386 6956
rect 17957 6851 18015 6857
rect 17957 6817 17969 6851
rect 18003 6848 18015 6851
rect 18322 6848 18328 6860
rect 18003 6820 18328 6848
rect 18003 6817 18015 6820
rect 17957 6811 18015 6817
rect 18322 6808 18328 6820
rect 18380 6808 18386 6860
rect 18417 6851 18475 6857
rect 18417 6817 18429 6851
rect 18463 6848 18475 6851
rect 18782 6848 18788 6860
rect 18463 6820 18788 6848
rect 18463 6817 18475 6820
rect 18417 6811 18475 6817
rect 18782 6808 18788 6820
rect 18840 6808 18846 6860
rect 18892 6848 18920 6956
rect 19978 6944 19984 6956
rect 20036 6944 20042 6996
rect 18966 6876 18972 6928
rect 19024 6916 19030 6928
rect 19024 6888 19932 6916
rect 19024 6876 19030 6888
rect 19150 6848 19156 6860
rect 18892 6820 19156 6848
rect 19150 6808 19156 6820
rect 19208 6808 19214 6860
rect 19429 6851 19487 6857
rect 19429 6817 19441 6851
rect 19475 6848 19487 6851
rect 19794 6848 19800 6860
rect 19475 6820 19800 6848
rect 19475 6817 19487 6820
rect 19429 6811 19487 6817
rect 19794 6808 19800 6820
rect 19852 6808 19858 6860
rect 19904 6848 19932 6888
rect 20898 6848 20904 6860
rect 19904 6820 20904 6848
rect 16942 6740 16948 6792
rect 17000 6780 17006 6792
rect 17690 6783 17748 6789
rect 17690 6780 17702 6783
rect 17000 6752 17702 6780
rect 17000 6740 17006 6752
rect 17690 6749 17702 6752
rect 17736 6749 17748 6783
rect 18233 6783 18291 6789
rect 18233 6780 18245 6783
rect 17690 6743 17748 6749
rect 17788 6752 18245 6780
rect 16684 6684 16988 6712
rect 11330 6644 11336 6656
rect 10468 6616 11192 6644
rect 11291 6616 11336 6644
rect 10468 6604 10474 6616
rect 11330 6604 11336 6616
rect 11388 6604 11394 6656
rect 12805 6647 12863 6653
rect 12805 6613 12817 6647
rect 12851 6644 12863 6647
rect 13078 6644 13084 6656
rect 12851 6616 13084 6644
rect 12851 6613 12863 6616
rect 12805 6607 12863 6613
rect 13078 6604 13084 6616
rect 13136 6604 13142 6656
rect 13354 6644 13360 6656
rect 13315 6616 13360 6644
rect 13354 6604 13360 6616
rect 13412 6604 13418 6656
rect 13449 6647 13507 6653
rect 13449 6613 13461 6647
rect 13495 6644 13507 6647
rect 13630 6644 13636 6656
rect 13495 6616 13636 6644
rect 13495 6613 13507 6616
rect 13449 6607 13507 6613
rect 13630 6604 13636 6616
rect 13688 6604 13694 6656
rect 13909 6647 13967 6653
rect 13909 6613 13921 6647
rect 13955 6644 13967 6647
rect 14182 6644 14188 6656
rect 13955 6616 14188 6644
rect 13955 6613 13967 6616
rect 13909 6607 13967 6613
rect 14182 6604 14188 6616
rect 14240 6604 14246 6656
rect 15470 6644 15476 6656
rect 15431 6616 15476 6644
rect 15470 6604 15476 6616
rect 15528 6604 15534 6656
rect 15562 6604 15568 6656
rect 15620 6644 15626 6656
rect 16022 6644 16028 6656
rect 15620 6616 15665 6644
rect 15983 6616 16028 6644
rect 15620 6604 15626 6616
rect 16022 6604 16028 6616
rect 16080 6604 16086 6656
rect 16577 6647 16635 6653
rect 16577 6613 16589 6647
rect 16623 6644 16635 6647
rect 16850 6644 16856 6656
rect 16623 6616 16856 6644
rect 16623 6613 16635 6616
rect 16577 6607 16635 6613
rect 16850 6604 16856 6616
rect 16908 6604 16914 6656
rect 16960 6644 16988 6684
rect 17788 6644 17816 6752
rect 18233 6749 18245 6752
rect 18279 6780 18291 6783
rect 18690 6780 18696 6792
rect 18279 6752 18696 6780
rect 18279 6749 18291 6752
rect 18233 6743 18291 6749
rect 18690 6740 18696 6752
rect 18748 6740 18754 6792
rect 20548 6789 20576 6820
rect 20898 6808 20904 6820
rect 20956 6808 20962 6860
rect 20349 6783 20407 6789
rect 20349 6780 20361 6783
rect 19306 6752 20361 6780
rect 18138 6672 18144 6724
rect 18196 6712 18202 6724
rect 19306 6712 19334 6752
rect 20349 6749 20361 6752
rect 20395 6749 20407 6783
rect 20349 6743 20407 6749
rect 20533 6783 20591 6789
rect 20533 6749 20545 6783
rect 20579 6749 20591 6783
rect 20533 6743 20591 6749
rect 20622 6740 20628 6792
rect 20680 6780 20686 6792
rect 20717 6783 20775 6789
rect 20717 6780 20729 6783
rect 20680 6752 20729 6780
rect 20680 6740 20686 6752
rect 20717 6749 20729 6752
rect 20763 6749 20775 6783
rect 20717 6743 20775 6749
rect 20993 6783 21051 6789
rect 20993 6749 21005 6783
rect 21039 6749 21051 6783
rect 20993 6743 21051 6749
rect 18196 6684 19334 6712
rect 19521 6715 19579 6721
rect 18196 6672 18202 6684
rect 19521 6681 19533 6715
rect 19567 6712 19579 6715
rect 19794 6712 19800 6724
rect 19567 6684 19800 6712
rect 19567 6681 19579 6684
rect 19521 6675 19579 6681
rect 19794 6672 19800 6684
rect 19852 6672 19858 6724
rect 20254 6672 20260 6724
rect 20312 6712 20318 6724
rect 21008 6712 21036 6743
rect 20312 6684 21036 6712
rect 20312 6672 20318 6684
rect 16960 6616 17816 6644
rect 17954 6604 17960 6656
rect 18012 6644 18018 6656
rect 18049 6647 18107 6653
rect 18049 6644 18061 6647
rect 18012 6616 18061 6644
rect 18012 6604 18018 6616
rect 18049 6613 18061 6616
rect 18095 6613 18107 6647
rect 18049 6607 18107 6613
rect 18322 6604 18328 6656
rect 18380 6644 18386 6656
rect 18601 6647 18659 6653
rect 18601 6644 18613 6647
rect 18380 6616 18613 6644
rect 18380 6604 18386 6616
rect 18601 6613 18613 6616
rect 18647 6613 18659 6647
rect 18601 6607 18659 6613
rect 18693 6647 18751 6653
rect 18693 6613 18705 6647
rect 18739 6644 18751 6647
rect 18966 6644 18972 6656
rect 18739 6616 18972 6644
rect 18739 6613 18751 6616
rect 18693 6607 18751 6613
rect 18966 6604 18972 6616
rect 19024 6604 19030 6656
rect 19061 6647 19119 6653
rect 19061 6613 19073 6647
rect 19107 6644 19119 6647
rect 19242 6644 19248 6656
rect 19107 6616 19248 6644
rect 19107 6613 19119 6616
rect 19061 6607 19119 6613
rect 19242 6604 19248 6616
rect 19300 6604 19306 6656
rect 19613 6647 19671 6653
rect 19613 6613 19625 6647
rect 19659 6644 19671 6647
rect 19702 6644 19708 6656
rect 19659 6616 19708 6644
rect 19659 6613 19671 6616
rect 19613 6607 19671 6613
rect 19702 6604 19708 6616
rect 19760 6604 19766 6656
rect 19886 6604 19892 6656
rect 19944 6644 19950 6656
rect 20073 6647 20131 6653
rect 20073 6644 20085 6647
rect 19944 6616 20085 6644
rect 19944 6604 19950 6616
rect 20073 6613 20085 6616
rect 20119 6613 20131 6647
rect 20073 6607 20131 6613
rect 1104 6554 22056 6576
rect 1104 6502 6148 6554
rect 6200 6502 6212 6554
rect 6264 6502 6276 6554
rect 6328 6502 6340 6554
rect 6392 6502 6404 6554
rect 6456 6502 11346 6554
rect 11398 6502 11410 6554
rect 11462 6502 11474 6554
rect 11526 6502 11538 6554
rect 11590 6502 11602 6554
rect 11654 6502 16544 6554
rect 16596 6502 16608 6554
rect 16660 6502 16672 6554
rect 16724 6502 16736 6554
rect 16788 6502 16800 6554
rect 16852 6502 21742 6554
rect 21794 6502 21806 6554
rect 21858 6502 21870 6554
rect 21922 6502 21934 6554
rect 21986 6502 21998 6554
rect 22050 6502 22056 6554
rect 1104 6480 22056 6502
rect 1857 6443 1915 6449
rect 1857 6409 1869 6443
rect 1903 6440 1915 6443
rect 1946 6440 1952 6452
rect 1903 6412 1952 6440
rect 1903 6409 1915 6412
rect 1857 6403 1915 6409
rect 1946 6400 1952 6412
rect 2004 6400 2010 6452
rect 2222 6440 2228 6452
rect 2183 6412 2228 6440
rect 2222 6400 2228 6412
rect 2280 6400 2286 6452
rect 2866 6400 2872 6452
rect 2924 6440 2930 6452
rect 4709 6443 4767 6449
rect 4709 6440 4721 6443
rect 2924 6412 4721 6440
rect 2924 6400 2930 6412
rect 4709 6409 4721 6412
rect 4755 6409 4767 6443
rect 4709 6403 4767 6409
rect 5813 6443 5871 6449
rect 5813 6409 5825 6443
rect 5859 6440 5871 6443
rect 6365 6443 6423 6449
rect 6365 6440 6377 6443
rect 5859 6412 6377 6440
rect 5859 6409 5871 6412
rect 5813 6403 5871 6409
rect 6365 6409 6377 6412
rect 6411 6409 6423 6443
rect 6365 6403 6423 6409
rect 6825 6443 6883 6449
rect 6825 6409 6837 6443
rect 6871 6440 6883 6443
rect 7282 6440 7288 6452
rect 6871 6412 7288 6440
rect 6871 6409 6883 6412
rect 6825 6403 6883 6409
rect 7282 6400 7288 6412
rect 7340 6400 7346 6452
rect 7561 6443 7619 6449
rect 7561 6409 7573 6443
rect 7607 6440 7619 6443
rect 8113 6443 8171 6449
rect 8113 6440 8125 6443
rect 7607 6412 8125 6440
rect 7607 6409 7619 6412
rect 7561 6403 7619 6409
rect 8113 6409 8125 6412
rect 8159 6409 8171 6443
rect 8113 6403 8171 6409
rect 8294 6400 8300 6452
rect 8352 6440 8358 6452
rect 8481 6443 8539 6449
rect 8481 6440 8493 6443
rect 8352 6412 8493 6440
rect 8352 6400 8358 6412
rect 8481 6409 8493 6412
rect 8527 6409 8539 6443
rect 8481 6403 8539 6409
rect 8573 6443 8631 6449
rect 8573 6409 8585 6443
rect 8619 6440 8631 6443
rect 8662 6440 8668 6452
rect 8619 6412 8668 6440
rect 8619 6409 8631 6412
rect 8573 6403 8631 6409
rect 8662 6400 8668 6412
rect 8720 6400 8726 6452
rect 8772 6412 10732 6440
rect 1486 6372 1492 6384
rect 1447 6344 1492 6372
rect 1486 6332 1492 6344
rect 1544 6332 1550 6384
rect 1673 6375 1731 6381
rect 1673 6341 1685 6375
rect 1719 6372 1731 6375
rect 1762 6372 1768 6384
rect 1719 6344 1768 6372
rect 1719 6341 1731 6344
rect 1673 6335 1731 6341
rect 1762 6332 1768 6344
rect 1820 6332 1826 6384
rect 3142 6372 3148 6384
rect 3103 6344 3148 6372
rect 3142 6332 3148 6344
rect 3200 6332 3206 6384
rect 3252 6344 4936 6372
rect 2774 6264 2780 6316
rect 2832 6304 2838 6316
rect 3252 6313 3280 6344
rect 4908 6316 4936 6344
rect 6546 6332 6552 6384
rect 6604 6372 6610 6384
rect 7653 6375 7711 6381
rect 6604 6344 7512 6372
rect 6604 6332 6610 6344
rect 3237 6307 3295 6313
rect 2832 6276 2877 6304
rect 2832 6264 2838 6276
rect 3237 6273 3249 6307
rect 3283 6273 3295 6307
rect 3493 6307 3551 6313
rect 3493 6304 3505 6307
rect 3237 6267 3295 6273
rect 3344 6276 3505 6304
rect 2317 6239 2375 6245
rect 2317 6205 2329 6239
rect 2363 6205 2375 6239
rect 2317 6199 2375 6205
rect 2501 6239 2559 6245
rect 2501 6205 2513 6239
rect 2547 6236 2559 6239
rect 2682 6236 2688 6248
rect 2547 6208 2688 6236
rect 2547 6205 2559 6208
rect 2501 6199 2559 6205
rect 2332 6100 2360 6199
rect 2682 6196 2688 6208
rect 2740 6196 2746 6248
rect 3344 6236 3372 6276
rect 3493 6273 3505 6276
rect 3539 6273 3551 6307
rect 3493 6267 3551 6273
rect 4246 6264 4252 6316
rect 4304 6304 4310 6316
rect 4522 6304 4528 6316
rect 4304 6276 4528 6304
rect 4304 6264 4310 6276
rect 4522 6264 4528 6276
rect 4580 6264 4586 6316
rect 4890 6304 4896 6316
rect 4851 6276 4896 6304
rect 4890 6264 4896 6276
rect 4948 6264 4954 6316
rect 4985 6307 5043 6313
rect 4985 6273 4997 6307
rect 5031 6304 5043 6307
rect 5350 6304 5356 6316
rect 5031 6276 5356 6304
rect 5031 6273 5043 6276
rect 4985 6267 5043 6273
rect 5350 6264 5356 6276
rect 5408 6264 5414 6316
rect 5721 6307 5779 6313
rect 5721 6273 5733 6307
rect 5767 6304 5779 6307
rect 6178 6304 6184 6316
rect 5767 6276 6184 6304
rect 5767 6273 5779 6276
rect 5721 6267 5779 6273
rect 6178 6264 6184 6276
rect 6236 6264 6242 6316
rect 6362 6264 6368 6316
rect 6420 6304 6426 6316
rect 6733 6307 6791 6313
rect 6733 6304 6745 6307
rect 6420 6276 6745 6304
rect 6420 6264 6426 6276
rect 6733 6273 6745 6276
rect 6779 6304 6791 6307
rect 7006 6304 7012 6316
rect 6779 6276 7012 6304
rect 6779 6273 6791 6276
rect 6733 6267 6791 6273
rect 7006 6264 7012 6276
rect 7064 6264 7070 6316
rect 3252 6208 3372 6236
rect 3252 6180 3280 6208
rect 4338 6196 4344 6248
rect 4396 6236 4402 6248
rect 4396 6208 5580 6236
rect 4396 6196 4402 6208
rect 2961 6171 3019 6177
rect 2961 6137 2973 6171
rect 3007 6168 3019 6171
rect 3142 6168 3148 6180
rect 3007 6140 3148 6168
rect 3007 6137 3019 6140
rect 2961 6131 3019 6137
rect 3142 6128 3148 6140
rect 3200 6128 3206 6180
rect 3234 6128 3240 6180
rect 3292 6128 3298 6180
rect 5074 6168 5080 6180
rect 4509 6140 5080 6168
rect 4509 6100 4537 6140
rect 5074 6128 5080 6140
rect 5132 6128 5138 6180
rect 5552 6168 5580 6208
rect 5626 6196 5632 6248
rect 5684 6236 5690 6248
rect 5905 6239 5963 6245
rect 5905 6236 5917 6239
rect 5684 6208 5917 6236
rect 5684 6196 5690 6208
rect 5905 6205 5917 6208
rect 5951 6205 5963 6239
rect 5905 6199 5963 6205
rect 6638 6196 6644 6248
rect 6696 6236 6702 6248
rect 6917 6239 6975 6245
rect 6917 6236 6929 6239
rect 6696 6208 6929 6236
rect 6696 6196 6702 6208
rect 6917 6205 6929 6208
rect 6963 6205 6975 6239
rect 7374 6236 7380 6248
rect 7335 6208 7380 6236
rect 6917 6199 6975 6205
rect 7374 6196 7380 6208
rect 7432 6196 7438 6248
rect 7484 6236 7512 6344
rect 7653 6341 7665 6375
rect 7699 6372 7711 6375
rect 8202 6372 8208 6384
rect 7699 6344 8208 6372
rect 7699 6341 7711 6344
rect 7653 6335 7711 6341
rect 8202 6332 8208 6344
rect 8260 6332 8266 6384
rect 8772 6304 8800 6412
rect 9582 6332 9588 6384
rect 9640 6372 9646 6384
rect 9640 6344 9996 6372
rect 9640 6332 9646 6344
rect 8404 6276 8800 6304
rect 8941 6307 8999 6313
rect 8404 6236 8432 6276
rect 8941 6273 8953 6307
rect 8987 6304 8999 6307
rect 9122 6304 9128 6316
rect 8987 6276 9128 6304
rect 8987 6273 8999 6276
rect 8941 6267 8999 6273
rect 9122 6264 9128 6276
rect 9180 6304 9186 6316
rect 9766 6304 9772 6316
rect 9180 6276 9772 6304
rect 9180 6264 9186 6276
rect 9766 6264 9772 6276
rect 9824 6264 9830 6316
rect 9968 6304 9996 6344
rect 10042 6332 10048 6384
rect 10100 6372 10106 6384
rect 10100 6344 10548 6372
rect 10100 6332 10106 6344
rect 10318 6304 10324 6316
rect 10376 6313 10382 6316
rect 9968 6276 10324 6304
rect 10318 6264 10324 6276
rect 10376 6267 10388 6313
rect 10376 6264 10382 6267
rect 7484 6208 8432 6236
rect 8757 6239 8815 6245
rect 8757 6205 8769 6239
rect 8803 6236 8815 6239
rect 9490 6236 9496 6248
rect 8803 6208 9496 6236
rect 8803 6205 8815 6208
rect 8757 6199 8815 6205
rect 9490 6196 9496 6208
rect 9548 6196 9554 6248
rect 10520 6236 10548 6344
rect 10594 6332 10600 6384
rect 10652 6332 10658 6384
rect 10704 6372 10732 6412
rect 11882 6400 11888 6452
rect 11940 6440 11946 6452
rect 12434 6440 12440 6452
rect 11940 6412 12440 6440
rect 11940 6400 11946 6412
rect 12434 6400 12440 6412
rect 12492 6400 12498 6452
rect 13357 6443 13415 6449
rect 13357 6409 13369 6443
rect 13403 6440 13415 6443
rect 16022 6440 16028 6452
rect 13403 6412 16028 6440
rect 13403 6409 13415 6412
rect 13357 6403 13415 6409
rect 16022 6400 16028 6412
rect 16080 6400 16086 6452
rect 16574 6440 16580 6452
rect 16132 6412 16580 6440
rect 12989 6375 13047 6381
rect 12989 6372 13001 6375
rect 10704 6344 13001 6372
rect 12989 6341 13001 6344
rect 13035 6341 13047 6375
rect 12989 6335 13047 6341
rect 13814 6332 13820 6384
rect 13872 6332 13878 6384
rect 16132 6372 16160 6412
rect 16574 6400 16580 6412
rect 16632 6440 16638 6452
rect 16669 6443 16727 6449
rect 16669 6440 16681 6443
rect 16632 6412 16681 6440
rect 16632 6400 16638 6412
rect 16669 6409 16681 6412
rect 16715 6409 16727 6443
rect 16669 6403 16727 6409
rect 17034 6400 17040 6452
rect 17092 6440 17098 6452
rect 17092 6412 18552 6440
rect 17092 6400 17098 6412
rect 14476 6344 16160 6372
rect 10612 6304 10640 6332
rect 10689 6307 10747 6313
rect 10689 6304 10701 6307
rect 10612 6276 10701 6304
rect 10689 6273 10701 6276
rect 10735 6273 10747 6307
rect 10689 6267 10747 6273
rect 11333 6307 11391 6313
rect 11333 6273 11345 6307
rect 11379 6304 11391 6307
rect 11885 6307 11943 6313
rect 11885 6304 11897 6307
rect 11379 6276 11897 6304
rect 11379 6273 11391 6276
rect 11333 6267 11391 6273
rect 11885 6273 11897 6276
rect 11931 6273 11943 6307
rect 13832 6304 13860 6332
rect 13998 6304 14004 6316
rect 11885 6267 11943 6273
rect 12728 6276 13860 6304
rect 13959 6276 14004 6304
rect 10597 6239 10655 6245
rect 10597 6236 10609 6239
rect 10520 6208 10609 6236
rect 10597 6205 10609 6208
rect 10643 6205 10655 6239
rect 10597 6199 10655 6205
rect 11057 6239 11115 6245
rect 11057 6205 11069 6239
rect 11103 6236 11115 6239
rect 11974 6236 11980 6248
rect 11103 6208 11980 6236
rect 11103 6205 11115 6208
rect 11057 6199 11115 6205
rect 11974 6196 11980 6208
rect 12032 6196 12038 6248
rect 12728 6245 12756 6276
rect 13998 6264 14004 6276
rect 14056 6264 14062 6316
rect 14090 6264 14096 6316
rect 14148 6304 14154 6316
rect 14476 6313 14504 6344
rect 14461 6307 14519 6313
rect 14461 6304 14473 6307
rect 14148 6276 14473 6304
rect 14148 6264 14154 6276
rect 14461 6273 14473 6276
rect 14507 6273 14519 6307
rect 14461 6267 14519 6273
rect 14728 6307 14786 6313
rect 14728 6273 14740 6307
rect 14774 6304 14786 6307
rect 15470 6304 15476 6316
rect 14774 6276 15476 6304
rect 14774 6273 14786 6276
rect 14728 6267 14786 6273
rect 15470 6264 15476 6276
rect 15528 6264 15534 6316
rect 15838 6264 15844 6316
rect 15896 6304 15902 6316
rect 16022 6304 16028 6316
rect 15896 6276 16028 6304
rect 15896 6264 15902 6276
rect 16022 6264 16028 6276
rect 16080 6264 16086 6316
rect 16132 6313 16160 6344
rect 16298 6332 16304 6384
rect 16356 6372 16362 6384
rect 16758 6372 16764 6384
rect 16356 6344 16764 6372
rect 16356 6332 16362 6344
rect 16758 6332 16764 6344
rect 16816 6332 16822 6384
rect 18414 6372 18420 6384
rect 16868 6344 18420 6372
rect 16868 6313 16896 6344
rect 16117 6307 16175 6313
rect 16117 6273 16129 6307
rect 16163 6273 16175 6307
rect 16117 6267 16175 6273
rect 16485 6307 16543 6313
rect 16485 6273 16497 6307
rect 16531 6273 16543 6307
rect 16485 6267 16543 6273
rect 16853 6307 16911 6313
rect 16853 6273 16865 6307
rect 16899 6273 16911 6307
rect 17034 6304 17040 6316
rect 16995 6276 17040 6304
rect 16853 6267 16911 6273
rect 12069 6239 12127 6245
rect 12069 6205 12081 6239
rect 12115 6205 12127 6239
rect 12069 6199 12127 6205
rect 12713 6239 12771 6245
rect 12713 6205 12725 6239
rect 12759 6205 12771 6239
rect 12894 6236 12900 6248
rect 12855 6208 12900 6236
rect 12713 6199 12771 6205
rect 5718 6168 5724 6180
rect 5552 6140 5724 6168
rect 5718 6128 5724 6140
rect 5776 6128 5782 6180
rect 7834 6168 7840 6180
rect 5828 6140 7840 6168
rect 2332 6072 4537 6100
rect 4614 6060 4620 6112
rect 4672 6100 4678 6112
rect 4672 6072 4717 6100
rect 4672 6060 4678 6072
rect 4890 6060 4896 6112
rect 4948 6100 4954 6112
rect 5169 6103 5227 6109
rect 5169 6100 5181 6103
rect 4948 6072 5181 6100
rect 4948 6060 4954 6072
rect 5169 6069 5181 6072
rect 5215 6069 5227 6103
rect 5350 6100 5356 6112
rect 5311 6072 5356 6100
rect 5169 6063 5227 6069
rect 5350 6060 5356 6072
rect 5408 6060 5414 6112
rect 5442 6060 5448 6112
rect 5500 6100 5506 6112
rect 5828 6100 5856 6140
rect 7834 6128 7840 6140
rect 7892 6128 7898 6180
rect 8202 6128 8208 6180
rect 8260 6168 8266 6180
rect 8938 6168 8944 6180
rect 8260 6140 8944 6168
rect 8260 6128 8266 6140
rect 8938 6128 8944 6140
rect 8996 6128 9002 6180
rect 9125 6171 9183 6177
rect 9125 6137 9137 6171
rect 9171 6168 9183 6171
rect 9398 6168 9404 6180
rect 9171 6140 9404 6168
rect 9171 6137 9183 6140
rect 9125 6131 9183 6137
rect 9398 6128 9404 6140
rect 9456 6128 9462 6180
rect 10778 6128 10784 6180
rect 10836 6168 10842 6180
rect 11517 6171 11575 6177
rect 11517 6168 11529 6171
rect 10836 6140 11529 6168
rect 10836 6128 10842 6140
rect 11517 6137 11529 6140
rect 11563 6137 11575 6171
rect 11517 6131 11575 6137
rect 11606 6128 11612 6180
rect 11664 6168 11670 6180
rect 12084 6168 12112 6199
rect 12894 6196 12900 6208
rect 12952 6196 12958 6248
rect 13725 6239 13783 6245
rect 13725 6205 13737 6239
rect 13771 6205 13783 6239
rect 13725 6199 13783 6205
rect 11664 6140 12112 6168
rect 13740 6168 13768 6199
rect 13814 6196 13820 6248
rect 13872 6236 13878 6248
rect 13909 6239 13967 6245
rect 13909 6236 13921 6239
rect 13872 6208 13921 6236
rect 13872 6196 13878 6208
rect 13909 6205 13921 6208
rect 13955 6205 13967 6239
rect 13909 6199 13967 6205
rect 15746 6196 15752 6248
rect 15804 6236 15810 6248
rect 16500 6236 16528 6267
rect 17034 6264 17040 6276
rect 17092 6264 17098 6316
rect 17328 6313 17356 6344
rect 18414 6332 18420 6344
rect 18472 6332 18478 6384
rect 18524 6372 18552 6412
rect 18598 6400 18604 6452
rect 18656 6440 18662 6452
rect 18693 6443 18751 6449
rect 18693 6440 18705 6443
rect 18656 6412 18705 6440
rect 18656 6400 18662 6412
rect 18693 6409 18705 6412
rect 18739 6409 18751 6443
rect 19242 6440 19248 6452
rect 19203 6412 19248 6440
rect 18693 6403 18751 6409
rect 19242 6400 19248 6412
rect 19300 6400 19306 6452
rect 19702 6440 19708 6452
rect 19663 6412 19708 6440
rect 19702 6400 19708 6412
rect 19760 6400 19766 6452
rect 19794 6400 19800 6452
rect 19852 6440 19858 6452
rect 19852 6412 19897 6440
rect 19852 6400 19858 6412
rect 20714 6400 20720 6452
rect 20772 6440 20778 6452
rect 20993 6443 21051 6449
rect 20993 6440 21005 6443
rect 20772 6412 21005 6440
rect 20772 6400 20778 6412
rect 20993 6409 21005 6412
rect 21039 6409 21051 6443
rect 21358 6440 21364 6452
rect 21319 6412 21364 6440
rect 20993 6403 21051 6409
rect 21358 6400 21364 6412
rect 21416 6400 21422 6452
rect 21450 6400 21456 6452
rect 21508 6440 21514 6452
rect 21726 6440 21732 6452
rect 21508 6412 21732 6440
rect 21508 6400 21514 6412
rect 21726 6400 21732 6412
rect 21784 6400 21790 6452
rect 18524 6344 21588 6372
rect 17586 6313 17592 6316
rect 17313 6307 17371 6313
rect 17313 6273 17325 6307
rect 17359 6273 17371 6307
rect 17580 6304 17592 6313
rect 17499 6276 17592 6304
rect 17313 6267 17371 6273
rect 17580 6267 17592 6276
rect 17644 6304 17650 6316
rect 18782 6304 18788 6316
rect 17644 6276 18788 6304
rect 17586 6264 17592 6267
rect 17644 6264 17650 6276
rect 18782 6264 18788 6276
rect 18840 6264 18846 6316
rect 19337 6307 19395 6313
rect 19337 6273 19349 6307
rect 19383 6304 19395 6307
rect 19518 6304 19524 6316
rect 19383 6276 19524 6304
rect 19383 6273 19395 6276
rect 19337 6267 19395 6273
rect 19518 6264 19524 6276
rect 19576 6264 19582 6316
rect 20162 6304 20168 6316
rect 20123 6276 20168 6304
rect 20162 6264 20168 6276
rect 20220 6264 20226 6316
rect 20714 6264 20720 6316
rect 20772 6304 20778 6316
rect 20901 6307 20959 6313
rect 20901 6304 20913 6307
rect 20772 6276 20913 6304
rect 20772 6264 20778 6276
rect 20901 6273 20913 6276
rect 20947 6273 20959 6307
rect 20901 6267 20959 6273
rect 15804 6208 16436 6236
rect 16500 6208 17356 6236
rect 15804 6196 15810 6208
rect 14458 6168 14464 6180
rect 13740 6140 14464 6168
rect 11664 6128 11670 6140
rect 14458 6128 14464 6140
rect 14516 6128 14522 6180
rect 15841 6171 15899 6177
rect 15841 6137 15853 6171
rect 15887 6168 15899 6171
rect 16206 6168 16212 6180
rect 15887 6140 16212 6168
rect 15887 6137 15899 6140
rect 15841 6131 15899 6137
rect 16206 6128 16212 6140
rect 16264 6128 16270 6180
rect 16408 6168 16436 6208
rect 17034 6168 17040 6180
rect 16408 6140 17040 6168
rect 17034 6128 17040 6140
rect 17092 6128 17098 6180
rect 17126 6128 17132 6180
rect 17184 6168 17190 6180
rect 17221 6171 17279 6177
rect 17221 6168 17233 6171
rect 17184 6140 17233 6168
rect 17184 6128 17190 6140
rect 17221 6137 17233 6140
rect 17267 6137 17279 6171
rect 17221 6131 17279 6137
rect 5500 6072 5856 6100
rect 5500 6060 5506 6072
rect 5902 6060 5908 6112
rect 5960 6100 5966 6112
rect 6270 6100 6276 6112
rect 5960 6072 6276 6100
rect 5960 6060 5966 6072
rect 6270 6060 6276 6072
rect 6328 6060 6334 6112
rect 8021 6103 8079 6109
rect 8021 6069 8033 6103
rect 8067 6100 8079 6103
rect 8294 6100 8300 6112
rect 8067 6072 8300 6100
rect 8067 6069 8079 6072
rect 8021 6063 8079 6069
rect 8294 6060 8300 6072
rect 8352 6060 8358 6112
rect 9217 6103 9275 6109
rect 9217 6069 9229 6103
rect 9263 6100 9275 6103
rect 9674 6100 9680 6112
rect 9263 6072 9680 6100
rect 9263 6069 9275 6072
rect 9217 6063 9275 6069
rect 9674 6060 9680 6072
rect 9732 6100 9738 6112
rect 10686 6100 10692 6112
rect 9732 6072 10692 6100
rect 9732 6060 9738 6072
rect 10686 6060 10692 6072
rect 10744 6060 10750 6112
rect 10870 6100 10876 6112
rect 10831 6072 10876 6100
rect 10870 6060 10876 6072
rect 10928 6060 10934 6112
rect 11238 6060 11244 6112
rect 11296 6100 11302 6112
rect 12437 6103 12495 6109
rect 12437 6100 12449 6103
rect 11296 6072 12449 6100
rect 11296 6060 11302 6072
rect 12437 6069 12449 6072
rect 12483 6100 12495 6103
rect 12986 6100 12992 6112
rect 12483 6072 12992 6100
rect 12483 6069 12495 6072
rect 12437 6063 12495 6069
rect 12986 6060 12992 6072
rect 13044 6060 13050 6112
rect 13538 6100 13544 6112
rect 13499 6072 13544 6100
rect 13538 6060 13544 6072
rect 13596 6100 13602 6112
rect 13998 6100 14004 6112
rect 13596 6072 14004 6100
rect 13596 6060 13602 6072
rect 13998 6060 14004 6072
rect 14056 6060 14062 6112
rect 14366 6100 14372 6112
rect 14327 6072 14372 6100
rect 14366 6060 14372 6072
rect 14424 6060 14430 6112
rect 14826 6060 14832 6112
rect 14884 6100 14890 6112
rect 15933 6103 15991 6109
rect 15933 6100 15945 6103
rect 14884 6072 15945 6100
rect 14884 6060 14890 6072
rect 15933 6069 15945 6072
rect 15979 6069 15991 6103
rect 15933 6063 15991 6069
rect 16114 6060 16120 6112
rect 16172 6100 16178 6112
rect 16301 6103 16359 6109
rect 16301 6100 16313 6103
rect 16172 6072 16313 6100
rect 16172 6060 16178 6072
rect 16301 6069 16313 6072
rect 16347 6069 16359 6103
rect 17328 6100 17356 6208
rect 18598 6196 18604 6248
rect 18656 6236 18662 6248
rect 19061 6239 19119 6245
rect 19061 6236 19073 6239
rect 18656 6208 19073 6236
rect 18656 6196 18662 6208
rect 19061 6205 19073 6208
rect 19107 6236 19119 6239
rect 20254 6236 20260 6248
rect 19107 6208 19334 6236
rect 20215 6208 20260 6236
rect 19107 6205 19119 6208
rect 19061 6199 19119 6205
rect 19306 6168 19334 6208
rect 20254 6196 20260 6208
rect 20312 6196 20318 6248
rect 20349 6239 20407 6245
rect 20349 6205 20361 6239
rect 20395 6205 20407 6239
rect 20806 6236 20812 6248
rect 20767 6208 20812 6236
rect 20349 6199 20407 6205
rect 20364 6168 20392 6199
rect 20806 6196 20812 6208
rect 20864 6196 20870 6248
rect 19306 6140 20392 6168
rect 21560 6112 21588 6344
rect 18877 6103 18935 6109
rect 18877 6100 18889 6103
rect 17328 6072 18889 6100
rect 16301 6063 16359 6069
rect 18877 6069 18889 6072
rect 18923 6100 18935 6103
rect 18966 6100 18972 6112
rect 18923 6072 18972 6100
rect 18923 6069 18935 6072
rect 18877 6063 18935 6069
rect 18966 6060 18972 6072
rect 19024 6060 19030 6112
rect 21542 6100 21548 6112
rect 21503 6072 21548 6100
rect 21542 6060 21548 6072
rect 21600 6060 21606 6112
rect 1104 6010 21896 6032
rect 1104 5958 3549 6010
rect 3601 5958 3613 6010
rect 3665 5958 3677 6010
rect 3729 5958 3741 6010
rect 3793 5958 3805 6010
rect 3857 5958 8747 6010
rect 8799 5958 8811 6010
rect 8863 5958 8875 6010
rect 8927 5958 8939 6010
rect 8991 5958 9003 6010
rect 9055 5958 13945 6010
rect 13997 5958 14009 6010
rect 14061 5958 14073 6010
rect 14125 5958 14137 6010
rect 14189 5958 14201 6010
rect 14253 5958 19143 6010
rect 19195 5958 19207 6010
rect 19259 5958 19271 6010
rect 19323 5958 19335 6010
rect 19387 5958 19399 6010
rect 19451 5958 21896 6010
rect 1104 5936 21896 5958
rect 3605 5899 3663 5905
rect 3605 5865 3617 5899
rect 3651 5896 3663 5899
rect 3878 5896 3884 5908
rect 3651 5868 3884 5896
rect 3651 5865 3663 5868
rect 3605 5859 3663 5865
rect 3878 5856 3884 5868
rect 3936 5856 3942 5908
rect 4982 5896 4988 5908
rect 4172 5868 4988 5896
rect 2777 5763 2835 5769
rect 2777 5729 2789 5763
rect 2823 5760 2835 5763
rect 2866 5760 2872 5772
rect 2823 5732 2872 5760
rect 2823 5729 2835 5732
rect 2777 5723 2835 5729
rect 2866 5720 2872 5732
rect 2924 5720 2930 5772
rect 3053 5763 3111 5769
rect 3053 5729 3065 5763
rect 3099 5760 3111 5763
rect 3878 5760 3884 5772
rect 3099 5732 3884 5760
rect 3099 5729 3111 5732
rect 3053 5723 3111 5729
rect 3878 5720 3884 5732
rect 3936 5720 3942 5772
rect 3973 5695 4031 5701
rect 2608 5664 3924 5692
rect 2608 5636 2636 5664
rect 2590 5633 2596 5636
rect 2532 5627 2596 5633
rect 2532 5593 2544 5627
rect 2578 5593 2596 5627
rect 2532 5587 2596 5593
rect 2590 5584 2596 5587
rect 2648 5584 2654 5636
rect 2682 5584 2688 5636
rect 2740 5624 2746 5636
rect 3237 5627 3295 5633
rect 3237 5624 3249 5627
rect 2740 5596 3249 5624
rect 2740 5584 2746 5596
rect 3237 5593 3249 5596
rect 3283 5593 3295 5627
rect 3237 5587 3295 5593
rect 1397 5559 1455 5565
rect 1397 5525 1409 5559
rect 1443 5556 1455 5559
rect 2130 5556 2136 5568
rect 1443 5528 2136 5556
rect 1443 5525 1455 5528
rect 1397 5519 1455 5525
rect 2130 5516 2136 5528
rect 2188 5516 2194 5568
rect 3142 5556 3148 5568
rect 3103 5528 3148 5556
rect 3142 5516 3148 5528
rect 3200 5516 3206 5568
rect 3896 5556 3924 5664
rect 3973 5661 3985 5695
rect 4019 5692 4031 5695
rect 4172 5692 4200 5868
rect 4982 5856 4988 5868
rect 5040 5856 5046 5908
rect 5902 5896 5908 5908
rect 5863 5868 5908 5896
rect 5902 5856 5908 5868
rect 5960 5856 5966 5908
rect 6178 5896 6184 5908
rect 6139 5868 6184 5896
rect 6178 5856 6184 5868
rect 6236 5856 6242 5908
rect 6546 5856 6552 5908
rect 6604 5896 6610 5908
rect 10594 5896 10600 5908
rect 6604 5868 10600 5896
rect 6604 5856 6610 5868
rect 10594 5856 10600 5868
rect 10652 5856 10658 5908
rect 10870 5856 10876 5908
rect 10928 5896 10934 5908
rect 13909 5899 13967 5905
rect 10928 5868 11652 5896
rect 10928 5856 10934 5868
rect 4246 5788 4252 5840
rect 4304 5788 4310 5840
rect 6089 5831 6147 5837
rect 6089 5797 6101 5831
rect 6135 5828 6147 5831
rect 6270 5828 6276 5840
rect 6135 5800 6276 5828
rect 6135 5797 6147 5800
rect 6089 5791 6147 5797
rect 6270 5788 6276 5800
rect 6328 5788 6334 5840
rect 6362 5788 6368 5840
rect 6420 5828 6426 5840
rect 7282 5828 7288 5840
rect 6420 5800 7288 5828
rect 6420 5788 6426 5800
rect 7282 5788 7288 5800
rect 7340 5788 7346 5840
rect 7926 5788 7932 5840
rect 7984 5828 7990 5840
rect 8110 5828 8116 5840
rect 7984 5800 8116 5828
rect 7984 5788 7990 5800
rect 8110 5788 8116 5800
rect 8168 5788 8174 5840
rect 9582 5828 9588 5840
rect 8772 5800 9588 5828
rect 4264 5701 4292 5788
rect 8772 5772 8800 5800
rect 9582 5788 9588 5800
rect 9640 5788 9646 5840
rect 10962 5788 10968 5840
rect 11020 5828 11026 5840
rect 11333 5831 11391 5837
rect 11333 5828 11345 5831
rect 11020 5800 11345 5828
rect 11020 5788 11026 5800
rect 11333 5797 11345 5800
rect 11379 5797 11391 5831
rect 11624 5828 11652 5868
rect 13909 5865 13921 5899
rect 13955 5896 13967 5899
rect 14642 5896 14648 5908
rect 13955 5868 14648 5896
rect 13955 5865 13967 5868
rect 13909 5859 13967 5865
rect 14642 5856 14648 5868
rect 14700 5856 14706 5908
rect 15105 5899 15163 5905
rect 15105 5865 15117 5899
rect 15151 5896 15163 5899
rect 18322 5896 18328 5908
rect 15151 5868 18328 5896
rect 15151 5865 15163 5868
rect 15105 5859 15163 5865
rect 18322 5856 18328 5868
rect 18380 5856 18386 5908
rect 18414 5856 18420 5908
rect 18472 5896 18478 5908
rect 19518 5896 19524 5908
rect 18472 5868 18736 5896
rect 19479 5868 19524 5896
rect 18472 5856 18478 5868
rect 15470 5828 15476 5840
rect 11624 5800 15476 5828
rect 11333 5791 11391 5797
rect 15470 5788 15476 5800
rect 15528 5788 15534 5840
rect 16945 5831 17003 5837
rect 16945 5797 16957 5831
rect 16991 5797 17003 5831
rect 17310 5828 17316 5840
rect 17223 5800 17316 5828
rect 16945 5791 17003 5797
rect 6638 5720 6644 5772
rect 6696 5760 6702 5772
rect 6733 5763 6791 5769
rect 6733 5760 6745 5763
rect 6696 5732 6745 5760
rect 6696 5720 6702 5732
rect 6733 5729 6745 5732
rect 6779 5729 6791 5763
rect 7374 5760 7380 5772
rect 7335 5732 7380 5760
rect 6733 5723 6791 5729
rect 7374 5720 7380 5732
rect 7432 5720 7438 5772
rect 8205 5763 8263 5769
rect 8205 5729 8217 5763
rect 8251 5760 8263 5763
rect 8754 5760 8760 5772
rect 8251 5732 8760 5760
rect 8251 5729 8263 5732
rect 8205 5723 8263 5729
rect 8754 5720 8760 5732
rect 8812 5720 8818 5772
rect 9125 5763 9183 5769
rect 9125 5729 9137 5763
rect 9171 5760 9183 5763
rect 9674 5760 9680 5772
rect 9171 5732 9680 5760
rect 9171 5729 9183 5732
rect 9125 5723 9183 5729
rect 9674 5720 9680 5732
rect 9732 5720 9738 5772
rect 9858 5760 9864 5772
rect 9819 5732 9864 5760
rect 9858 5720 9864 5732
rect 9916 5720 9922 5772
rect 10781 5763 10839 5769
rect 10781 5729 10793 5763
rect 10827 5760 10839 5763
rect 10870 5760 10876 5772
rect 10827 5732 10876 5760
rect 10827 5729 10839 5732
rect 10781 5723 10839 5729
rect 10870 5720 10876 5732
rect 10928 5760 10934 5772
rect 11517 5763 11575 5769
rect 11517 5760 11529 5763
rect 10928 5732 11529 5760
rect 10928 5720 10934 5732
rect 11517 5729 11529 5732
rect 11563 5729 11575 5763
rect 13170 5760 13176 5772
rect 11517 5723 11575 5729
rect 11808 5732 12480 5760
rect 13131 5732 13176 5760
rect 4019 5664 4200 5692
rect 4249 5695 4307 5701
rect 4019 5661 4031 5664
rect 3973 5655 4031 5661
rect 4249 5661 4261 5695
rect 4295 5661 4307 5695
rect 5718 5692 5724 5704
rect 5631 5664 5724 5692
rect 4249 5655 4307 5661
rect 5718 5652 5724 5664
rect 5776 5692 5782 5704
rect 7466 5692 7472 5704
rect 5776 5664 7472 5692
rect 5776 5652 5782 5664
rect 7466 5652 7472 5664
rect 7524 5652 7530 5704
rect 7561 5695 7619 5701
rect 7561 5661 7573 5695
rect 7607 5692 7619 5695
rect 7742 5692 7748 5704
rect 7607 5664 7748 5692
rect 7607 5661 7619 5664
rect 7561 5655 7619 5661
rect 7742 5652 7748 5664
rect 7800 5652 7806 5704
rect 9217 5695 9275 5701
rect 9217 5661 9229 5695
rect 9263 5692 9275 5695
rect 10594 5692 10600 5704
rect 9263 5664 10600 5692
rect 9263 5661 9275 5664
rect 9217 5655 9275 5661
rect 10594 5652 10600 5664
rect 10652 5652 10658 5704
rect 11532 5692 11560 5723
rect 11532 5688 11744 5692
rect 11808 5688 11836 5732
rect 12158 5692 12164 5704
rect 11532 5664 11836 5688
rect 11716 5660 11836 5664
rect 11900 5664 12164 5692
rect 4154 5624 4160 5636
rect 4115 5596 4160 5624
rect 4154 5584 4160 5596
rect 4212 5584 4218 5636
rect 4516 5627 4574 5633
rect 4516 5593 4528 5627
rect 4562 5593 4574 5627
rect 4982 5624 4988 5636
rect 4516 5587 4574 5593
rect 4724 5596 4988 5624
rect 4246 5556 4252 5568
rect 3896 5528 4252 5556
rect 4246 5516 4252 5528
rect 4304 5516 4310 5568
rect 4531 5556 4559 5587
rect 4724 5556 4752 5596
rect 4982 5584 4988 5596
rect 5040 5584 5046 5636
rect 6822 5624 6828 5636
rect 6735 5596 6828 5624
rect 5626 5556 5632 5568
rect 4531 5528 4752 5556
rect 5587 5528 5632 5556
rect 5626 5516 5632 5528
rect 5684 5516 5690 5568
rect 5718 5516 5724 5568
rect 5776 5556 5782 5568
rect 6362 5556 6368 5568
rect 5776 5528 6368 5556
rect 5776 5516 5782 5528
rect 6362 5516 6368 5528
rect 6420 5516 6426 5568
rect 6454 5516 6460 5568
rect 6512 5556 6518 5568
rect 6549 5559 6607 5565
rect 6549 5556 6561 5559
rect 6512 5528 6561 5556
rect 6512 5516 6518 5528
rect 6549 5525 6561 5528
rect 6595 5525 6607 5559
rect 6549 5519 6607 5525
rect 6641 5559 6699 5565
rect 6641 5525 6653 5559
rect 6687 5556 6699 5559
rect 6748 5556 6776 5596
rect 6822 5584 6828 5596
rect 6880 5624 6886 5636
rect 8202 5624 8208 5636
rect 6880 5596 8208 5624
rect 6880 5584 6886 5596
rect 8202 5584 8208 5596
rect 8260 5584 8266 5636
rect 8297 5627 8355 5633
rect 8297 5593 8309 5627
rect 8343 5624 8355 5627
rect 8662 5624 8668 5636
rect 8343 5596 8668 5624
rect 8343 5593 8355 5596
rect 8297 5587 8355 5593
rect 8662 5584 8668 5596
rect 8720 5584 8726 5636
rect 9309 5627 9367 5633
rect 9309 5624 9321 5627
rect 8772 5596 9321 5624
rect 6687 5528 6776 5556
rect 6687 5525 6699 5528
rect 6641 5519 6699 5525
rect 6914 5516 6920 5568
rect 6972 5556 6978 5568
rect 7009 5559 7067 5565
rect 7009 5556 7021 5559
rect 6972 5528 7021 5556
rect 6972 5516 6978 5528
rect 7009 5525 7021 5528
rect 7055 5525 7067 5559
rect 7466 5556 7472 5568
rect 7427 5528 7472 5556
rect 7009 5519 7067 5525
rect 7466 5516 7472 5528
rect 7524 5516 7530 5568
rect 7926 5556 7932 5568
rect 7887 5528 7932 5556
rect 7926 5516 7932 5528
rect 7984 5516 7990 5568
rect 8389 5559 8447 5565
rect 8389 5525 8401 5559
rect 8435 5556 8447 5559
rect 8570 5556 8576 5568
rect 8435 5528 8576 5556
rect 8435 5525 8447 5528
rect 8389 5519 8447 5525
rect 8570 5516 8576 5528
rect 8628 5516 8634 5568
rect 8772 5565 8800 5596
rect 9309 5593 9321 5596
rect 9355 5593 9367 5627
rect 9309 5587 9367 5593
rect 9398 5584 9404 5636
rect 9456 5624 9462 5636
rect 9858 5624 9864 5636
rect 9456 5596 9864 5624
rect 9456 5584 9462 5596
rect 9858 5584 9864 5596
rect 9916 5584 9922 5636
rect 10965 5627 11023 5633
rect 10965 5593 10977 5627
rect 11011 5624 11023 5627
rect 11330 5624 11336 5636
rect 11011 5596 11336 5624
rect 11011 5593 11023 5596
rect 10965 5587 11023 5593
rect 11330 5584 11336 5596
rect 11388 5584 11394 5636
rect 8757 5559 8815 5565
rect 8757 5525 8769 5559
rect 8803 5525 8815 5559
rect 8757 5519 8815 5525
rect 9677 5559 9735 5565
rect 9677 5525 9689 5559
rect 9723 5556 9735 5559
rect 10045 5559 10103 5565
rect 10045 5556 10057 5559
rect 9723 5528 10057 5556
rect 9723 5525 9735 5528
rect 9677 5519 9735 5525
rect 10045 5525 10057 5528
rect 10091 5525 10103 5559
rect 10045 5519 10103 5525
rect 10134 5516 10140 5568
rect 10192 5556 10198 5568
rect 10502 5556 10508 5568
rect 10192 5528 10237 5556
rect 10463 5528 10508 5556
rect 10192 5516 10198 5528
rect 10502 5516 10508 5528
rect 10560 5516 10566 5568
rect 10873 5559 10931 5565
rect 10873 5525 10885 5559
rect 10919 5556 10931 5559
rect 11238 5556 11244 5568
rect 10919 5528 11244 5556
rect 10919 5525 10931 5528
rect 10873 5519 10931 5525
rect 11238 5516 11244 5528
rect 11296 5516 11302 5568
rect 11606 5516 11612 5568
rect 11664 5556 11670 5568
rect 11701 5559 11759 5565
rect 11701 5556 11713 5559
rect 11664 5528 11713 5556
rect 11664 5516 11670 5528
rect 11701 5525 11713 5528
rect 11747 5525 11759 5559
rect 11701 5519 11759 5525
rect 11793 5559 11851 5565
rect 11793 5525 11805 5559
rect 11839 5556 11851 5559
rect 11900 5556 11928 5664
rect 12158 5652 12164 5664
rect 12216 5652 12222 5704
rect 12452 5701 12480 5732
rect 13170 5720 13176 5732
rect 13228 5720 13234 5772
rect 13357 5763 13415 5769
rect 13357 5729 13369 5763
rect 13403 5760 13415 5763
rect 13630 5760 13636 5772
rect 13403 5732 13636 5760
rect 13403 5729 13415 5732
rect 13357 5723 13415 5729
rect 13630 5720 13636 5732
rect 13688 5720 13694 5772
rect 14274 5760 14280 5772
rect 13740 5732 14280 5760
rect 12437 5695 12495 5701
rect 12437 5661 12449 5695
rect 12483 5661 12495 5695
rect 13078 5692 13084 5704
rect 13039 5664 13084 5692
rect 12437 5655 12495 5661
rect 13078 5652 13084 5664
rect 13136 5652 13142 5704
rect 13740 5701 13768 5732
rect 14274 5720 14280 5732
rect 14332 5720 14338 5772
rect 14458 5760 14464 5772
rect 14419 5732 14464 5760
rect 14458 5720 14464 5732
rect 14516 5760 14522 5772
rect 16574 5760 16580 5772
rect 14516 5732 15608 5760
rect 16535 5732 16580 5760
rect 14516 5720 14522 5732
rect 13725 5695 13783 5701
rect 13725 5661 13737 5695
rect 13771 5661 13783 5695
rect 13725 5655 13783 5661
rect 14093 5695 14151 5701
rect 14093 5661 14105 5695
rect 14139 5692 14151 5695
rect 14918 5692 14924 5704
rect 14139 5664 14924 5692
rect 14139 5661 14151 5664
rect 14093 5655 14151 5661
rect 14918 5652 14924 5664
rect 14976 5652 14982 5704
rect 15378 5692 15384 5704
rect 15120 5664 15384 5692
rect 11974 5584 11980 5636
rect 12032 5624 12038 5636
rect 12253 5627 12311 5633
rect 12253 5624 12265 5627
rect 12032 5596 12265 5624
rect 12032 5584 12038 5596
rect 12253 5593 12265 5596
rect 12299 5593 12311 5627
rect 12253 5587 12311 5593
rect 13906 5584 13912 5636
rect 13964 5624 13970 5636
rect 14645 5627 14703 5633
rect 14645 5624 14657 5627
rect 13964 5596 14657 5624
rect 13964 5584 13970 5596
rect 14645 5593 14657 5596
rect 14691 5593 14703 5627
rect 14645 5587 14703 5593
rect 12158 5556 12164 5568
rect 11839 5528 11928 5556
rect 12119 5528 12164 5556
rect 11839 5525 11851 5528
rect 11793 5519 11851 5525
rect 12158 5516 12164 5528
rect 12216 5516 12222 5568
rect 12710 5556 12716 5568
rect 12671 5528 12716 5556
rect 12710 5516 12716 5528
rect 12768 5516 12774 5568
rect 13538 5556 13544 5568
rect 13499 5528 13544 5556
rect 13538 5516 13544 5528
rect 13596 5556 13602 5568
rect 13814 5556 13820 5568
rect 13596 5528 13820 5556
rect 13596 5516 13602 5528
rect 13814 5516 13820 5528
rect 13872 5516 13878 5568
rect 14182 5516 14188 5568
rect 14240 5556 14246 5568
rect 14277 5559 14335 5565
rect 14277 5556 14289 5559
rect 14240 5528 14289 5556
rect 14240 5516 14246 5528
rect 14277 5525 14289 5528
rect 14323 5525 14335 5559
rect 14277 5519 14335 5525
rect 14458 5516 14464 5568
rect 14516 5556 14522 5568
rect 14737 5559 14795 5565
rect 14737 5556 14749 5559
rect 14516 5528 14749 5556
rect 14516 5516 14522 5528
rect 14737 5525 14749 5528
rect 14783 5556 14795 5559
rect 15120 5556 15148 5664
rect 15378 5652 15384 5664
rect 15436 5652 15442 5704
rect 15580 5692 15608 5732
rect 16574 5720 16580 5732
rect 16632 5720 16638 5772
rect 16960 5760 16988 5791
rect 17310 5788 17316 5800
rect 17368 5828 17374 5840
rect 17586 5828 17592 5840
rect 17368 5800 17592 5828
rect 17368 5788 17374 5800
rect 17586 5788 17592 5800
rect 17644 5788 17650 5840
rect 18708 5769 18736 5868
rect 19518 5856 19524 5868
rect 19576 5856 19582 5908
rect 20162 5856 20168 5908
rect 20220 5896 20226 5908
rect 20349 5899 20407 5905
rect 20349 5896 20361 5899
rect 20220 5868 20361 5896
rect 20220 5856 20226 5868
rect 20349 5865 20361 5868
rect 20395 5865 20407 5899
rect 20349 5859 20407 5865
rect 20990 5856 20996 5908
rect 21048 5896 21054 5908
rect 21361 5899 21419 5905
rect 21361 5896 21373 5899
rect 21048 5868 21373 5896
rect 21048 5856 21054 5868
rect 21361 5865 21373 5868
rect 21407 5865 21419 5899
rect 21361 5859 21419 5865
rect 19429 5831 19487 5837
rect 19429 5797 19441 5831
rect 19475 5828 19487 5831
rect 21266 5828 21272 5840
rect 19475 5800 21272 5828
rect 19475 5797 19487 5800
rect 19429 5791 19487 5797
rect 21266 5788 21272 5800
rect 21324 5788 21330 5840
rect 18693 5763 18751 5769
rect 16960 5732 17724 5760
rect 16758 5692 16764 5704
rect 15580 5664 16620 5692
rect 16719 5664 16764 5692
rect 16298 5584 16304 5636
rect 16356 5633 16362 5636
rect 16356 5624 16368 5633
rect 16592 5624 16620 5664
rect 16758 5652 16764 5664
rect 16816 5652 16822 5704
rect 17034 5692 17040 5704
rect 16995 5664 17040 5692
rect 17034 5652 17040 5664
rect 17092 5652 17098 5704
rect 17696 5692 17724 5732
rect 18693 5729 18705 5763
rect 18739 5729 18751 5763
rect 18693 5723 18751 5729
rect 18782 5720 18788 5772
rect 18840 5760 18846 5772
rect 20165 5763 20223 5769
rect 20165 5760 20177 5763
rect 18840 5732 20177 5760
rect 18840 5720 18846 5732
rect 20165 5729 20177 5732
rect 20211 5729 20223 5763
rect 20165 5723 20223 5729
rect 17862 5692 17868 5704
rect 17696 5664 17868 5692
rect 17862 5652 17868 5664
rect 17920 5652 17926 5704
rect 18874 5652 18880 5704
rect 18932 5692 18938 5704
rect 18969 5695 19027 5701
rect 18969 5692 18981 5695
rect 18932 5664 18981 5692
rect 18932 5652 18938 5664
rect 18969 5661 18981 5664
rect 19015 5661 19027 5695
rect 18969 5655 19027 5661
rect 19058 5652 19064 5704
rect 19116 5692 19122 5704
rect 19245 5695 19303 5701
rect 19245 5692 19257 5695
rect 19116 5664 19257 5692
rect 19116 5652 19122 5664
rect 19245 5661 19257 5664
rect 19291 5661 19303 5695
rect 19886 5692 19892 5704
rect 19847 5664 19892 5692
rect 19245 5655 19303 5661
rect 19886 5652 19892 5664
rect 19944 5652 19950 5704
rect 20180 5692 20208 5723
rect 20438 5720 20444 5772
rect 20496 5760 20502 5772
rect 20809 5763 20867 5769
rect 20809 5760 20821 5763
rect 20496 5732 20821 5760
rect 20496 5720 20502 5732
rect 20809 5729 20821 5732
rect 20855 5729 20867 5763
rect 20809 5723 20867 5729
rect 20901 5763 20959 5769
rect 20901 5729 20913 5763
rect 20947 5729 20959 5763
rect 20901 5723 20959 5729
rect 20916 5692 20944 5723
rect 20180 5664 20944 5692
rect 21266 5652 21272 5704
rect 21324 5692 21330 5704
rect 22554 5692 22560 5704
rect 21324 5664 22560 5692
rect 21324 5652 21330 5664
rect 22554 5652 22560 5664
rect 22612 5652 22618 5704
rect 18138 5624 18144 5636
rect 16356 5596 16401 5624
rect 16592 5596 18144 5624
rect 16356 5587 16368 5596
rect 16356 5584 16362 5587
rect 18138 5584 18144 5596
rect 18196 5624 18202 5636
rect 18426 5627 18484 5633
rect 18426 5624 18438 5627
rect 18196 5596 18438 5624
rect 18196 5584 18202 5596
rect 18426 5593 18438 5596
rect 18472 5593 18484 5627
rect 18782 5624 18788 5636
rect 18743 5596 18788 5624
rect 18426 5587 18484 5593
rect 18782 5584 18788 5596
rect 18840 5584 18846 5636
rect 19702 5584 19708 5636
rect 19760 5624 19766 5636
rect 19981 5627 20039 5633
rect 19981 5624 19993 5627
rect 19760 5596 19993 5624
rect 19760 5584 19766 5596
rect 19981 5593 19993 5596
rect 20027 5593 20039 5627
rect 19981 5587 20039 5593
rect 21453 5627 21511 5633
rect 21453 5593 21465 5627
rect 21499 5624 21511 5627
rect 21726 5624 21732 5636
rect 21499 5596 21732 5624
rect 21499 5593 21511 5596
rect 21453 5587 21511 5593
rect 21726 5584 21732 5596
rect 21784 5584 21790 5636
rect 14783 5528 15148 5556
rect 15197 5559 15255 5565
rect 14783 5525 14795 5528
rect 14737 5519 14795 5525
rect 15197 5525 15209 5559
rect 15243 5556 15255 5559
rect 15378 5556 15384 5568
rect 15243 5528 15384 5556
rect 15243 5525 15255 5528
rect 15197 5519 15255 5525
rect 15378 5516 15384 5528
rect 15436 5516 15442 5568
rect 16758 5516 16764 5568
rect 16816 5556 16822 5568
rect 17126 5556 17132 5568
rect 16816 5528 17132 5556
rect 16816 5516 16822 5528
rect 17126 5516 17132 5528
rect 17184 5516 17190 5568
rect 17221 5559 17279 5565
rect 17221 5525 17233 5559
rect 17267 5556 17279 5559
rect 17862 5556 17868 5568
rect 17267 5528 17868 5556
rect 17267 5525 17279 5528
rect 17221 5519 17279 5525
rect 17862 5516 17868 5528
rect 17920 5516 17926 5568
rect 20714 5556 20720 5568
rect 20675 5528 20720 5556
rect 20714 5516 20720 5528
rect 20772 5516 20778 5568
rect 382 5448 388 5500
rect 440 5488 446 5500
rect 934 5488 940 5500
rect 440 5460 940 5488
rect 440 5448 446 5460
rect 934 5448 940 5460
rect 992 5448 998 5500
rect 1104 5466 22056 5488
rect 1104 5414 6148 5466
rect 6200 5414 6212 5466
rect 6264 5414 6276 5466
rect 6328 5414 6340 5466
rect 6392 5414 6404 5466
rect 6456 5414 11346 5466
rect 11398 5414 11410 5466
rect 11462 5414 11474 5466
rect 11526 5414 11538 5466
rect 11590 5414 11602 5466
rect 11654 5414 16544 5466
rect 16596 5414 16608 5466
rect 16660 5414 16672 5466
rect 16724 5414 16736 5466
rect 16788 5414 16800 5466
rect 16852 5414 21742 5466
rect 21794 5414 21806 5466
rect 21858 5414 21870 5466
rect 21922 5414 21934 5466
rect 21986 5414 21998 5466
rect 22050 5414 22056 5466
rect 1104 5392 22056 5414
rect 3326 5352 3332 5364
rect 3287 5324 3332 5352
rect 3326 5312 3332 5324
rect 3384 5312 3390 5364
rect 4062 5352 4068 5364
rect 4023 5324 4068 5352
rect 4062 5312 4068 5324
rect 4120 5312 4126 5364
rect 4157 5355 4215 5361
rect 4157 5321 4169 5355
rect 4203 5352 4215 5355
rect 4430 5352 4436 5364
rect 4203 5324 4436 5352
rect 4203 5321 4215 5324
rect 4157 5315 4215 5321
rect 4430 5312 4436 5324
rect 4488 5352 4494 5364
rect 4488 5324 5672 5352
rect 4488 5312 4494 5324
rect 198 5244 204 5296
rect 256 5284 262 5296
rect 1026 5284 1032 5296
rect 256 5256 1032 5284
rect 256 5244 262 5256
rect 1026 5244 1032 5256
rect 1084 5284 1090 5296
rect 2409 5287 2467 5293
rect 2409 5284 2421 5287
rect 1084 5256 2421 5284
rect 1084 5244 1090 5256
rect 2409 5253 2421 5256
rect 2455 5253 2467 5287
rect 2409 5247 2467 5253
rect 3237 5287 3295 5293
rect 3237 5253 3249 5287
rect 3283 5284 3295 5287
rect 3510 5284 3516 5296
rect 3283 5256 3516 5284
rect 3283 5253 3295 5256
rect 3237 5247 3295 5253
rect 3510 5244 3516 5256
rect 3568 5244 3574 5296
rect 5534 5284 5540 5296
rect 4356 5256 5540 5284
rect 1949 5219 2007 5225
rect 1949 5185 1961 5219
rect 1995 5216 2007 5219
rect 2038 5216 2044 5228
rect 1995 5188 2044 5216
rect 1995 5185 2007 5188
rect 1949 5179 2007 5185
rect 2038 5176 2044 5188
rect 2096 5176 2102 5228
rect 2777 5219 2835 5225
rect 2777 5185 2789 5219
rect 2823 5216 2835 5219
rect 3326 5216 3332 5228
rect 2823 5188 3332 5216
rect 2823 5185 2835 5188
rect 2777 5179 2835 5185
rect 3326 5176 3332 5188
rect 3384 5176 3390 5228
rect 3878 5176 3884 5228
rect 3936 5216 3942 5228
rect 4154 5216 4160 5228
rect 3936 5188 4160 5216
rect 3936 5176 3942 5188
rect 4154 5176 4160 5188
rect 4212 5176 4218 5228
rect 1762 5108 1768 5160
rect 1820 5148 1826 5160
rect 2225 5151 2283 5157
rect 2225 5148 2237 5151
rect 1820 5120 2237 5148
rect 1820 5108 1826 5120
rect 2225 5117 2237 5120
rect 2271 5148 2283 5151
rect 3050 5148 3056 5160
rect 2271 5120 3056 5148
rect 2271 5117 2283 5120
rect 2225 5111 2283 5117
rect 3050 5108 3056 5120
rect 3108 5108 3114 5160
rect 4356 5157 4384 5256
rect 5534 5244 5540 5256
rect 5592 5244 5598 5296
rect 4525 5219 4583 5225
rect 4525 5185 4537 5219
rect 4571 5216 4583 5219
rect 4982 5216 4988 5228
rect 4571 5188 4988 5216
rect 4571 5185 4583 5188
rect 4525 5179 4583 5185
rect 3513 5151 3571 5157
rect 3513 5117 3525 5151
rect 3559 5117 3571 5151
rect 3513 5111 3571 5117
rect 4341 5151 4399 5157
rect 4341 5117 4353 5151
rect 4387 5117 4399 5151
rect 4341 5111 4399 5117
rect 3528 5080 3556 5111
rect 4154 5080 4160 5092
rect 3528 5052 4160 5080
rect 4154 5040 4160 5052
rect 4212 5080 4218 5092
rect 4540 5080 4568 5179
rect 4982 5176 4988 5188
rect 5040 5176 5046 5228
rect 4801 5151 4859 5157
rect 4801 5117 4813 5151
rect 4847 5117 4859 5151
rect 5644 5148 5672 5324
rect 5718 5312 5724 5364
rect 5776 5352 5782 5364
rect 5813 5355 5871 5361
rect 5813 5352 5825 5355
rect 5776 5324 5825 5352
rect 5776 5312 5782 5324
rect 5813 5321 5825 5324
rect 5859 5321 5871 5355
rect 5813 5315 5871 5321
rect 5902 5312 5908 5364
rect 5960 5352 5966 5364
rect 6825 5355 6883 5361
rect 6825 5352 6837 5355
rect 5960 5324 6837 5352
rect 5960 5312 5966 5324
rect 6825 5321 6837 5324
rect 6871 5321 6883 5355
rect 6825 5315 6883 5321
rect 7466 5312 7472 5364
rect 7524 5352 7530 5364
rect 7837 5355 7895 5361
rect 7837 5352 7849 5355
rect 7524 5324 7849 5352
rect 7524 5312 7530 5324
rect 7837 5321 7849 5324
rect 7883 5321 7895 5355
rect 7837 5315 7895 5321
rect 8018 5312 8024 5364
rect 8076 5352 8082 5364
rect 8297 5355 8355 5361
rect 8297 5352 8309 5355
rect 8076 5324 8309 5352
rect 8076 5312 8082 5324
rect 8297 5321 8309 5324
rect 8343 5321 8355 5355
rect 8297 5315 8355 5321
rect 8665 5355 8723 5361
rect 8665 5321 8677 5355
rect 8711 5352 8723 5355
rect 8754 5352 8760 5364
rect 8711 5324 8760 5352
rect 8711 5321 8723 5324
rect 8665 5315 8723 5321
rect 8754 5312 8760 5324
rect 8812 5312 8818 5364
rect 10134 5312 10140 5364
rect 10192 5352 10198 5364
rect 10413 5355 10471 5361
rect 10413 5352 10425 5355
rect 10192 5324 10425 5352
rect 10192 5312 10198 5324
rect 10413 5321 10425 5324
rect 10459 5321 10471 5355
rect 10778 5352 10784 5364
rect 10739 5324 10784 5352
rect 10413 5315 10471 5321
rect 10778 5312 10784 5324
rect 10836 5312 10842 5364
rect 10873 5355 10931 5361
rect 10873 5321 10885 5355
rect 10919 5352 10931 5355
rect 11517 5355 11575 5361
rect 11517 5352 11529 5355
rect 10919 5324 11529 5352
rect 10919 5321 10931 5324
rect 10873 5315 10931 5321
rect 11517 5321 11529 5324
rect 11563 5321 11575 5355
rect 11517 5315 11575 5321
rect 11606 5312 11612 5364
rect 11664 5352 11670 5364
rect 11882 5352 11888 5364
rect 11664 5324 11888 5352
rect 11664 5312 11670 5324
rect 11882 5312 11888 5324
rect 11940 5312 11946 5364
rect 11977 5355 12035 5361
rect 11977 5321 11989 5355
rect 12023 5352 12035 5355
rect 12158 5352 12164 5364
rect 12023 5324 12164 5352
rect 12023 5321 12035 5324
rect 11977 5315 12035 5321
rect 12158 5312 12164 5324
rect 12216 5312 12222 5364
rect 12250 5312 12256 5364
rect 12308 5352 12314 5364
rect 12618 5352 12624 5364
rect 12308 5324 12624 5352
rect 12308 5312 12314 5324
rect 12618 5312 12624 5324
rect 12676 5312 12682 5364
rect 14366 5312 14372 5364
rect 14424 5352 14430 5364
rect 17037 5355 17095 5361
rect 17037 5352 17049 5355
rect 14424 5324 17049 5352
rect 14424 5312 14430 5324
rect 17037 5321 17049 5324
rect 17083 5321 17095 5355
rect 17037 5315 17095 5321
rect 17129 5355 17187 5361
rect 17129 5321 17141 5355
rect 17175 5352 17187 5355
rect 17494 5352 17500 5364
rect 17175 5324 17500 5352
rect 17175 5321 17187 5324
rect 17129 5315 17187 5321
rect 17494 5312 17500 5324
rect 17552 5312 17558 5364
rect 17773 5355 17831 5361
rect 17773 5321 17785 5355
rect 17819 5352 17831 5355
rect 19426 5352 19432 5364
rect 17819 5324 19432 5352
rect 17819 5321 17831 5324
rect 17773 5315 17831 5321
rect 19426 5312 19432 5324
rect 19484 5312 19490 5364
rect 19521 5355 19579 5361
rect 19521 5321 19533 5355
rect 19567 5352 19579 5355
rect 19567 5324 19901 5352
rect 19567 5321 19579 5324
rect 19521 5315 19579 5321
rect 19628 5296 19656 5324
rect 7282 5284 7288 5296
rect 5920 5256 7288 5284
rect 5920 5225 5948 5256
rect 7282 5244 7288 5256
rect 7340 5244 7346 5296
rect 7484 5256 8524 5284
rect 5905 5219 5963 5225
rect 5905 5185 5917 5219
rect 5951 5185 5963 5219
rect 6270 5216 6276 5228
rect 5905 5179 5963 5185
rect 6012 5188 6276 5216
rect 6012 5148 6040 5188
rect 6270 5176 6276 5188
rect 6328 5176 6334 5228
rect 6733 5219 6791 5225
rect 6733 5185 6745 5219
rect 6779 5216 6791 5219
rect 7006 5216 7012 5228
rect 6779 5188 7012 5216
rect 6779 5185 6791 5188
rect 6733 5179 6791 5185
rect 7006 5176 7012 5188
rect 7064 5176 7070 5228
rect 7484 5225 7512 5256
rect 7469 5219 7527 5225
rect 7469 5185 7481 5219
rect 7515 5216 7527 5219
rect 7745 5219 7803 5225
rect 7515 5188 7696 5216
rect 7515 5185 7527 5188
rect 7469 5179 7527 5185
rect 5644 5120 6040 5148
rect 6089 5151 6147 5157
rect 4801 5111 4859 5117
rect 6089 5117 6101 5151
rect 6135 5148 6147 5151
rect 6638 5148 6644 5160
rect 6135 5120 6644 5148
rect 6135 5117 6147 5120
rect 6089 5111 6147 5117
rect 4212 5052 4568 5080
rect 4816 5080 4844 5111
rect 6104 5080 6132 5111
rect 6638 5108 6644 5120
rect 6696 5148 6702 5160
rect 6917 5151 6975 5157
rect 6917 5148 6929 5151
rect 6696 5120 6929 5148
rect 6696 5108 6702 5120
rect 6917 5117 6929 5120
rect 6963 5117 6975 5151
rect 6917 5111 6975 5117
rect 4816 5052 6132 5080
rect 4212 5040 4218 5052
rect 7006 5040 7012 5092
rect 7064 5080 7070 5092
rect 7668 5080 7696 5188
rect 7745 5185 7757 5219
rect 7791 5216 7803 5219
rect 8018 5216 8024 5228
rect 7791 5188 8024 5216
rect 7791 5185 7803 5188
rect 7745 5179 7803 5185
rect 8018 5176 8024 5188
rect 8076 5176 8082 5228
rect 8205 5219 8263 5225
rect 8205 5185 8217 5219
rect 8251 5185 8263 5219
rect 8205 5179 8263 5185
rect 8496 5216 8524 5256
rect 9674 5244 9680 5296
rect 9732 5284 9738 5296
rect 9800 5287 9858 5293
rect 9800 5284 9812 5287
rect 9732 5256 9812 5284
rect 9732 5244 9738 5256
rect 9800 5253 9812 5256
rect 9846 5284 9858 5287
rect 9846 5256 12020 5284
rect 9846 5253 9858 5256
rect 9800 5247 9858 5253
rect 11992 5228 12020 5256
rect 13722 5244 13728 5296
rect 13780 5284 13786 5296
rect 14676 5287 14734 5293
rect 14676 5284 14688 5287
rect 13780 5256 14688 5284
rect 13780 5244 13786 5256
rect 14676 5253 14688 5256
rect 14722 5284 14734 5287
rect 16117 5287 16175 5293
rect 16117 5284 16129 5287
rect 14722 5256 16129 5284
rect 14722 5253 14734 5256
rect 14676 5247 14734 5253
rect 16117 5253 16129 5256
rect 16163 5253 16175 5287
rect 16117 5247 16175 5253
rect 16301 5287 16359 5293
rect 16301 5253 16313 5287
rect 16347 5284 16359 5287
rect 16942 5284 16948 5296
rect 16347 5256 16948 5284
rect 16347 5253 16359 5256
rect 16301 5247 16359 5253
rect 16942 5244 16948 5256
rect 17000 5244 17006 5296
rect 17218 5244 17224 5296
rect 17276 5284 17282 5296
rect 17276 5256 17908 5284
rect 17276 5244 17282 5256
rect 9306 5216 9312 5228
rect 8496 5188 9312 5216
rect 7834 5108 7840 5160
rect 7892 5148 7898 5160
rect 8220 5148 8248 5179
rect 8496 5157 8524 5188
rect 9306 5176 9312 5188
rect 9364 5176 9370 5228
rect 10042 5216 10048 5228
rect 10003 5188 10048 5216
rect 10042 5176 10048 5188
rect 10100 5176 10106 5228
rect 10137 5219 10195 5225
rect 10137 5185 10149 5219
rect 10183 5216 10195 5219
rect 10502 5216 10508 5228
rect 10183 5188 10508 5216
rect 10183 5185 10195 5188
rect 10137 5179 10195 5185
rect 10502 5176 10508 5188
rect 10560 5176 10566 5228
rect 11333 5219 11391 5225
rect 11333 5185 11345 5219
rect 11379 5216 11391 5219
rect 11606 5216 11612 5228
rect 11379 5188 11612 5216
rect 11379 5185 11391 5188
rect 11333 5179 11391 5185
rect 11606 5176 11612 5188
rect 11664 5176 11670 5228
rect 11882 5216 11888 5228
rect 11843 5188 11888 5216
rect 11882 5176 11888 5188
rect 11940 5176 11946 5228
rect 11974 5176 11980 5228
rect 12032 5176 12038 5228
rect 12250 5176 12256 5228
rect 12308 5216 12314 5228
rect 12345 5219 12403 5225
rect 12345 5216 12357 5219
rect 12308 5188 12357 5216
rect 12308 5176 12314 5188
rect 12345 5185 12357 5188
rect 12391 5185 12403 5219
rect 12345 5179 12403 5185
rect 12710 5176 12716 5228
rect 12768 5216 12774 5228
rect 12897 5219 12955 5225
rect 12897 5216 12909 5219
rect 12768 5188 12909 5216
rect 12768 5176 12774 5188
rect 12897 5185 12909 5188
rect 12943 5185 12955 5219
rect 12897 5179 12955 5185
rect 12989 5219 13047 5225
rect 12989 5185 13001 5219
rect 13035 5216 13047 5219
rect 13078 5216 13084 5228
rect 13035 5188 13084 5216
rect 13035 5185 13047 5188
rect 12989 5179 13047 5185
rect 13078 5176 13084 5188
rect 13136 5176 13142 5228
rect 14826 5176 14832 5228
rect 14884 5216 14890 5228
rect 14921 5219 14979 5225
rect 14921 5216 14933 5219
rect 14884 5188 14933 5216
rect 14884 5176 14890 5188
rect 14921 5185 14933 5188
rect 14967 5185 14979 5219
rect 14921 5179 14979 5185
rect 15013 5219 15071 5225
rect 15013 5185 15025 5219
rect 15059 5216 15071 5219
rect 15102 5216 15108 5228
rect 15059 5188 15108 5216
rect 15059 5185 15071 5188
rect 15013 5179 15071 5185
rect 15102 5176 15108 5188
rect 15160 5176 15166 5228
rect 15654 5216 15660 5228
rect 15615 5188 15660 5216
rect 15654 5176 15660 5188
rect 15712 5176 15718 5228
rect 17586 5216 17592 5228
rect 17547 5188 17592 5216
rect 17586 5176 17592 5188
rect 17644 5176 17650 5228
rect 17880 5225 17908 5256
rect 18064 5256 19334 5284
rect 17865 5219 17923 5225
rect 17865 5185 17877 5219
rect 17911 5185 17923 5219
rect 17865 5179 17923 5185
rect 7892 5120 8248 5148
rect 8481 5151 8539 5157
rect 7892 5108 7898 5120
rect 8481 5117 8493 5151
rect 8527 5117 8539 5151
rect 8481 5111 8539 5117
rect 10686 5108 10692 5160
rect 10744 5148 10750 5160
rect 10965 5151 11023 5157
rect 10965 5148 10977 5151
rect 10744 5120 10977 5148
rect 10744 5108 10750 5120
rect 10965 5117 10977 5120
rect 11011 5117 11023 5151
rect 10965 5111 11023 5117
rect 11146 5108 11152 5160
rect 11204 5148 11210 5160
rect 12069 5151 12127 5157
rect 12069 5148 12081 5151
rect 11204 5120 12081 5148
rect 11204 5108 11210 5120
rect 12069 5117 12081 5120
rect 12115 5117 12127 5151
rect 12069 5111 12127 5117
rect 12805 5151 12863 5157
rect 12805 5117 12817 5151
rect 12851 5148 12863 5151
rect 12851 5120 13584 5148
rect 12851 5117 12863 5120
rect 12805 5111 12863 5117
rect 7742 5080 7748 5092
rect 7064 5052 7604 5080
rect 7668 5052 7748 5080
rect 7064 5040 7070 5052
rect 2498 5012 2504 5024
rect 2459 4984 2504 5012
rect 2498 4972 2504 4984
rect 2556 4972 2562 5024
rect 2866 4972 2872 5024
rect 2924 5012 2930 5024
rect 2924 4984 2969 5012
rect 2924 4972 2930 4984
rect 3326 4972 3332 5024
rect 3384 5012 3390 5024
rect 3697 5015 3755 5021
rect 3697 5012 3709 5015
rect 3384 4984 3709 5012
rect 3384 4972 3390 4984
rect 3697 4981 3709 4984
rect 3743 4981 3755 5015
rect 3697 4975 3755 4981
rect 4246 4972 4252 5024
rect 4304 5012 4310 5024
rect 4430 5012 4436 5024
rect 4304 4984 4436 5012
rect 4304 4972 4310 4984
rect 4430 4972 4436 4984
rect 4488 4972 4494 5024
rect 5445 5015 5503 5021
rect 5445 4981 5457 5015
rect 5491 5012 5503 5015
rect 5718 5012 5724 5024
rect 5491 4984 5724 5012
rect 5491 4981 5503 4984
rect 5445 4975 5503 4981
rect 5718 4972 5724 4984
rect 5776 4972 5782 5024
rect 6362 5012 6368 5024
rect 6323 4984 6368 5012
rect 6362 4972 6368 4984
rect 6420 4972 6426 5024
rect 7282 5012 7288 5024
rect 7243 4984 7288 5012
rect 7282 4972 7288 4984
rect 7340 4972 7346 5024
rect 7576 5021 7604 5052
rect 7742 5040 7748 5052
rect 7800 5040 7806 5092
rect 13556 5024 13584 5120
rect 15194 5108 15200 5160
rect 15252 5148 15258 5160
rect 15381 5151 15439 5157
rect 15381 5148 15393 5151
rect 15252 5120 15393 5148
rect 15252 5108 15258 5120
rect 15381 5117 15393 5120
rect 15427 5117 15439 5151
rect 15381 5111 15439 5117
rect 15565 5151 15623 5157
rect 15565 5117 15577 5151
rect 15611 5148 15623 5151
rect 16482 5148 16488 5160
rect 15611 5120 16488 5148
rect 15611 5117 15623 5120
rect 15565 5111 15623 5117
rect 16482 5108 16488 5120
rect 16540 5108 16546 5160
rect 16945 5151 17003 5157
rect 16945 5117 16957 5151
rect 16991 5148 17003 5151
rect 17310 5148 17316 5160
rect 16991 5120 17316 5148
rect 16991 5117 17003 5120
rect 16945 5111 17003 5117
rect 17310 5108 17316 5120
rect 17368 5108 17374 5160
rect 18064 5148 18092 5256
rect 18141 5219 18199 5225
rect 18141 5185 18153 5219
rect 18187 5216 18199 5219
rect 18230 5216 18236 5228
rect 18187 5188 18236 5216
rect 18187 5185 18199 5188
rect 18141 5179 18199 5185
rect 18230 5176 18236 5188
rect 18288 5176 18294 5228
rect 18414 5225 18420 5228
rect 18408 5179 18420 5225
rect 18472 5216 18478 5228
rect 19306 5216 19334 5256
rect 19610 5244 19616 5296
rect 19668 5244 19674 5296
rect 19873 5293 19901 5324
rect 20898 5312 20904 5364
rect 20956 5352 20962 5364
rect 20993 5355 21051 5361
rect 20993 5352 21005 5355
rect 20956 5324 21005 5352
rect 20956 5312 20962 5324
rect 20993 5321 21005 5324
rect 21039 5321 21051 5355
rect 21358 5352 21364 5364
rect 21319 5324 21364 5352
rect 20993 5315 21051 5321
rect 21358 5312 21364 5324
rect 21416 5312 21422 5364
rect 21726 5312 21732 5364
rect 21784 5352 21790 5364
rect 22462 5352 22468 5364
rect 21784 5324 22468 5352
rect 21784 5312 21790 5324
rect 22462 5312 22468 5324
rect 22520 5312 22526 5364
rect 19858 5287 19916 5293
rect 19858 5253 19870 5287
rect 19904 5253 19916 5287
rect 21450 5284 21456 5296
rect 21411 5256 21456 5284
rect 19858 5247 19916 5253
rect 21450 5244 21456 5256
rect 21508 5244 21514 5296
rect 20254 5216 20260 5228
rect 18472 5188 18508 5216
rect 19306 5188 20260 5216
rect 18414 5176 18420 5179
rect 18472 5176 18478 5188
rect 20254 5176 20260 5188
rect 20312 5176 20318 5228
rect 21177 5219 21235 5225
rect 21177 5185 21189 5219
rect 21223 5216 21235 5219
rect 21358 5216 21364 5228
rect 21223 5188 21364 5216
rect 21223 5185 21235 5188
rect 21177 5179 21235 5185
rect 21358 5176 21364 5188
rect 21416 5216 21422 5228
rect 22738 5216 22744 5228
rect 21416 5188 22744 5216
rect 21416 5176 21422 5188
rect 22738 5176 22744 5188
rect 22796 5176 22802 5228
rect 17512 5120 18092 5148
rect 19613 5151 19671 5157
rect 16025 5083 16083 5089
rect 16025 5049 16037 5083
rect 16071 5080 16083 5083
rect 16390 5080 16396 5092
rect 16071 5052 16396 5080
rect 16071 5049 16083 5052
rect 16025 5043 16083 5049
rect 16390 5040 16396 5052
rect 16448 5040 16454 5092
rect 17512 5089 17540 5120
rect 19613 5117 19625 5151
rect 19659 5117 19671 5151
rect 19613 5111 19671 5117
rect 17497 5083 17555 5089
rect 17497 5049 17509 5083
rect 17543 5049 17555 5083
rect 17497 5043 17555 5049
rect 7561 5015 7619 5021
rect 7561 4981 7573 5015
rect 7607 4981 7619 5015
rect 7561 4975 7619 4981
rect 8938 4972 8944 5024
rect 8996 5012 9002 5024
rect 10134 5012 10140 5024
rect 8996 4984 10140 5012
rect 8996 4972 9002 4984
rect 10134 4972 10140 4984
rect 10192 4972 10198 5024
rect 10318 5012 10324 5024
rect 10279 4984 10324 5012
rect 10318 4972 10324 4984
rect 10376 4972 10382 5024
rect 11882 4972 11888 5024
rect 11940 5012 11946 5024
rect 12342 5012 12348 5024
rect 11940 4984 12348 5012
rect 11940 4972 11946 4984
rect 12342 4972 12348 4984
rect 12400 4972 12406 5024
rect 12529 5015 12587 5021
rect 12529 4981 12541 5015
rect 12575 5012 12587 5015
rect 13262 5012 13268 5024
rect 12575 4984 13268 5012
rect 12575 4981 12587 4984
rect 12529 4975 12587 4981
rect 13262 4972 13268 4984
rect 13320 4972 13326 5024
rect 13357 5015 13415 5021
rect 13357 4981 13369 5015
rect 13403 5012 13415 5015
rect 13446 5012 13452 5024
rect 13403 4984 13452 5012
rect 13403 4981 13415 4984
rect 13357 4975 13415 4981
rect 13446 4972 13452 4984
rect 13504 4972 13510 5024
rect 13538 4972 13544 5024
rect 13596 5012 13602 5024
rect 15194 5012 15200 5024
rect 13596 4984 13641 5012
rect 15155 4984 15200 5012
rect 13596 4972 13602 4984
rect 15194 4972 15200 4984
rect 15252 4972 15258 5024
rect 18049 5015 18107 5021
rect 18049 4981 18061 5015
rect 18095 5012 18107 5015
rect 18506 5012 18512 5024
rect 18095 4984 18512 5012
rect 18095 4981 18107 4984
rect 18049 4975 18107 4981
rect 18506 4972 18512 4984
rect 18564 4972 18570 5024
rect 18874 4972 18880 5024
rect 18932 5012 18938 5024
rect 19628 5012 19656 5111
rect 20806 5108 20812 5160
rect 20864 5148 20870 5160
rect 21450 5148 21456 5160
rect 20864 5120 21456 5148
rect 20864 5108 20870 5120
rect 21450 5108 21456 5120
rect 21508 5108 21514 5160
rect 18932 4984 19656 5012
rect 18932 4972 18938 4984
rect 1104 4922 21896 4944
rect 1104 4870 3549 4922
rect 3601 4870 3613 4922
rect 3665 4870 3677 4922
rect 3729 4870 3741 4922
rect 3793 4870 3805 4922
rect 3857 4870 8747 4922
rect 8799 4870 8811 4922
rect 8863 4870 8875 4922
rect 8927 4870 8939 4922
rect 8991 4870 9003 4922
rect 9055 4870 13945 4922
rect 13997 4870 14009 4922
rect 14061 4870 14073 4922
rect 14125 4870 14137 4922
rect 14189 4870 14201 4922
rect 14253 4870 19143 4922
rect 19195 4870 19207 4922
rect 19259 4870 19271 4922
rect 19323 4870 19335 4922
rect 19387 4870 19399 4922
rect 19451 4870 21896 4922
rect 1104 4848 21896 4870
rect 2130 4768 2136 4820
rect 2188 4808 2194 4820
rect 2188 4780 3096 4808
rect 2188 4768 2194 4780
rect 2866 4740 2872 4752
rect 2516 4712 2872 4740
rect 1946 4672 1952 4684
rect 1907 4644 1952 4672
rect 1946 4632 1952 4644
rect 2004 4632 2010 4684
rect 2516 4681 2544 4712
rect 2866 4700 2872 4712
rect 2924 4700 2930 4752
rect 3068 4740 3096 4780
rect 3142 4768 3148 4820
rect 3200 4808 3206 4820
rect 4157 4811 4215 4817
rect 4157 4808 4169 4811
rect 3200 4780 4169 4808
rect 3200 4768 3206 4780
rect 4157 4777 4169 4780
rect 4203 4777 4215 4811
rect 4157 4771 4215 4777
rect 5626 4768 5632 4820
rect 5684 4808 5690 4820
rect 5810 4808 5816 4820
rect 5684 4780 5816 4808
rect 5684 4768 5690 4780
rect 5810 4768 5816 4780
rect 5868 4768 5874 4820
rect 6270 4808 6276 4820
rect 6231 4780 6276 4808
rect 6270 4768 6276 4780
rect 6328 4768 6334 4820
rect 7469 4811 7527 4817
rect 7469 4777 7481 4811
rect 7515 4808 7527 4811
rect 7558 4808 7564 4820
rect 7515 4780 7564 4808
rect 7515 4777 7527 4780
rect 7469 4771 7527 4777
rect 7558 4768 7564 4780
rect 7616 4768 7622 4820
rect 8662 4768 8668 4820
rect 8720 4808 8726 4820
rect 8941 4811 8999 4817
rect 8941 4808 8953 4811
rect 8720 4780 8953 4808
rect 8720 4768 8726 4780
rect 8941 4777 8953 4780
rect 8987 4777 8999 4811
rect 8941 4771 8999 4777
rect 9030 4768 9036 4820
rect 9088 4808 9094 4820
rect 9769 4811 9827 4817
rect 9088 4780 9674 4808
rect 9088 4768 9094 4780
rect 3234 4740 3240 4752
rect 3068 4712 3240 4740
rect 3234 4700 3240 4712
rect 3292 4740 3298 4752
rect 3292 4712 4752 4740
rect 3292 4700 3298 4712
rect 2501 4675 2559 4681
rect 2501 4641 2513 4675
rect 2547 4641 2559 4675
rect 2501 4635 2559 4641
rect 2590 4632 2596 4684
rect 2648 4672 2654 4684
rect 3326 4672 3332 4684
rect 2648 4644 2693 4672
rect 3287 4644 3332 4672
rect 2648 4632 2654 4644
rect 3326 4632 3332 4644
rect 3384 4632 3390 4684
rect 3513 4675 3571 4681
rect 3513 4641 3525 4675
rect 3559 4672 3571 4675
rect 4062 4672 4068 4684
rect 3559 4644 4068 4672
rect 3559 4641 3571 4644
rect 3513 4635 3571 4641
rect 4062 4632 4068 4644
rect 4120 4632 4126 4684
rect 4724 4681 4752 4712
rect 4798 4700 4804 4752
rect 4856 4740 4862 4752
rect 5350 4740 5356 4752
rect 4856 4712 5356 4740
rect 4856 4700 4862 4712
rect 5350 4700 5356 4712
rect 5408 4700 5414 4752
rect 5552 4712 8432 4740
rect 4709 4675 4767 4681
rect 4709 4641 4721 4675
rect 4755 4641 4767 4675
rect 5552 4672 5580 4712
rect 5718 4672 5724 4684
rect 4709 4635 4767 4641
rect 4908 4644 5580 4672
rect 5679 4644 5724 4672
rect 934 4564 940 4616
rect 992 4604 998 4616
rect 1489 4607 1547 4613
rect 1489 4604 1501 4607
rect 992 4576 1501 4604
rect 992 4564 998 4576
rect 1489 4573 1501 4576
rect 1535 4573 1547 4607
rect 2406 4604 2412 4616
rect 2367 4576 2412 4604
rect 1489 4567 1547 4573
rect 2406 4564 2412 4576
rect 2464 4564 2470 4616
rect 3973 4607 4031 4613
rect 3973 4573 3985 4607
rect 4019 4604 4031 4607
rect 4908 4604 4936 4644
rect 5718 4632 5724 4644
rect 5776 4632 5782 4684
rect 5810 4632 5816 4684
rect 5868 4672 5874 4684
rect 6457 4675 6515 4681
rect 5868 4644 5913 4672
rect 5868 4632 5874 4644
rect 6457 4641 6469 4675
rect 6503 4672 6515 4675
rect 6822 4672 6828 4684
rect 6503 4644 6828 4672
rect 6503 4641 6515 4644
rect 6457 4635 6515 4641
rect 6822 4632 6828 4644
rect 6880 4672 6886 4684
rect 7466 4672 7472 4684
rect 6880 4644 7472 4672
rect 6880 4632 6886 4644
rect 7466 4632 7472 4644
rect 7524 4632 7530 4684
rect 7745 4675 7803 4681
rect 7745 4641 7757 4675
rect 7791 4672 7803 4675
rect 8202 4672 8208 4684
rect 7791 4644 8208 4672
rect 7791 4641 7803 4644
rect 7745 4635 7803 4641
rect 8202 4632 8208 4644
rect 8260 4632 8266 4684
rect 8404 4672 8432 4712
rect 8478 4700 8484 4752
rect 8536 4740 8542 4752
rect 8757 4743 8815 4749
rect 8757 4740 8769 4743
rect 8536 4712 8769 4740
rect 8536 4700 8542 4712
rect 8757 4709 8769 4712
rect 8803 4709 8815 4743
rect 9646 4740 9674 4780
rect 9769 4777 9781 4811
rect 9815 4808 9827 4811
rect 9950 4808 9956 4820
rect 9815 4780 9956 4808
rect 9815 4777 9827 4780
rect 9769 4771 9827 4777
rect 9950 4768 9956 4780
rect 10008 4768 10014 4820
rect 10594 4808 10600 4820
rect 10555 4780 10600 4808
rect 10594 4768 10600 4780
rect 10652 4768 10658 4820
rect 10778 4768 10784 4820
rect 10836 4808 10842 4820
rect 12434 4808 12440 4820
rect 10836 4780 12440 4808
rect 10836 4768 10842 4780
rect 12434 4768 12440 4780
rect 12492 4768 12498 4820
rect 12986 4768 12992 4820
rect 13044 4808 13050 4820
rect 17678 4808 17684 4820
rect 13044 4780 13676 4808
rect 13044 4768 13050 4780
rect 9646 4712 11560 4740
rect 8757 4703 8815 4709
rect 9585 4675 9643 4681
rect 8404 4644 9536 4672
rect 4019 4576 4936 4604
rect 4985 4607 5043 4613
rect 4019 4573 4031 4576
rect 3973 4567 4031 4573
rect 4985 4573 4997 4607
rect 5031 4604 5043 4607
rect 5074 4604 5080 4616
rect 5031 4576 5080 4604
rect 5031 4573 5043 4576
rect 4985 4567 5043 4573
rect 5074 4564 5080 4576
rect 5132 4564 5138 4616
rect 5629 4607 5687 4613
rect 5629 4573 5641 4607
rect 5675 4604 5687 4607
rect 6362 4604 6368 4616
rect 5675 4576 6368 4604
rect 5675 4573 5687 4576
rect 5629 4567 5687 4573
rect 6362 4564 6368 4576
rect 6420 4564 6426 4616
rect 6638 4564 6644 4616
rect 6696 4604 6702 4616
rect 6733 4607 6791 4613
rect 6733 4604 6745 4607
rect 6696 4576 6745 4604
rect 6696 4564 6702 4576
rect 6733 4573 6745 4576
rect 6779 4573 6791 4607
rect 8573 4607 8631 4613
rect 6733 4567 6791 4573
rect 7024 4600 8524 4604
rect 8573 4600 8585 4607
rect 7024 4576 8585 4600
rect 1673 4539 1731 4545
rect 1673 4505 1685 4539
rect 1719 4536 1731 4539
rect 1762 4536 1768 4548
rect 1719 4508 1768 4536
rect 1719 4505 1731 4508
rect 1673 4499 1731 4505
rect 1762 4496 1768 4508
rect 1820 4496 1826 4548
rect 2222 4496 2228 4548
rect 2280 4536 2286 4548
rect 2590 4536 2596 4548
rect 2280 4508 2596 4536
rect 2280 4496 2286 4508
rect 2590 4496 2596 4508
rect 2648 4496 2654 4548
rect 3237 4539 3295 4545
rect 3237 4505 3249 4539
rect 3283 4536 3295 4539
rect 4430 4536 4436 4548
rect 3283 4508 4436 4536
rect 3283 4505 3295 4508
rect 3237 4499 3295 4505
rect 4430 4496 4436 4508
rect 4488 4496 4494 4548
rect 4525 4539 4583 4545
rect 4525 4505 4537 4539
rect 4571 4536 4583 4539
rect 4571 4508 5304 4536
rect 4571 4505 4583 4508
rect 4525 4499 4583 4505
rect 1026 4428 1032 4480
rect 1084 4468 1090 4480
rect 1394 4468 1400 4480
rect 1084 4440 1400 4468
rect 1084 4428 1090 4440
rect 1394 4428 1400 4440
rect 1452 4428 1458 4480
rect 2038 4428 2044 4480
rect 2096 4468 2102 4480
rect 2096 4440 2141 4468
rect 2096 4428 2102 4440
rect 2406 4428 2412 4480
rect 2464 4468 2470 4480
rect 2869 4471 2927 4477
rect 2869 4468 2881 4471
rect 2464 4440 2881 4468
rect 2464 4428 2470 4440
rect 2869 4437 2881 4440
rect 2915 4437 2927 4471
rect 2869 4431 2927 4437
rect 4617 4471 4675 4477
rect 4617 4437 4629 4471
rect 4663 4468 4675 4471
rect 4798 4468 4804 4480
rect 4663 4440 4804 4468
rect 4663 4437 4675 4440
rect 4617 4431 4675 4437
rect 4798 4428 4804 4440
rect 4856 4428 4862 4480
rect 5074 4428 5080 4480
rect 5132 4468 5138 4480
rect 5276 4477 5304 4508
rect 5902 4496 5908 4548
rect 5960 4536 5966 4548
rect 6178 4536 6184 4548
rect 5960 4508 6184 4536
rect 5960 4496 5966 4508
rect 6178 4496 6184 4508
rect 6236 4496 6242 4548
rect 5169 4471 5227 4477
rect 5169 4468 5181 4471
rect 5132 4440 5181 4468
rect 5132 4428 5138 4440
rect 5169 4437 5181 4440
rect 5215 4437 5227 4471
rect 5169 4431 5227 4437
rect 5261 4471 5319 4477
rect 5261 4437 5273 4471
rect 5307 4437 5319 4471
rect 5261 4431 5319 4437
rect 5626 4428 5632 4480
rect 5684 4468 5690 4480
rect 7024 4468 7052 4576
rect 8496 4573 8585 4576
rect 8619 4600 8631 4607
rect 8662 4600 8668 4616
rect 8619 4573 8668 4600
rect 8496 4572 8668 4573
rect 8573 4567 8631 4572
rect 8662 4564 8668 4572
rect 8720 4564 8726 4616
rect 9508 4604 9536 4644
rect 9585 4641 9597 4675
rect 9631 4672 9643 4675
rect 9674 4672 9680 4684
rect 9631 4644 9680 4672
rect 9631 4641 9643 4644
rect 9585 4635 9643 4641
rect 9674 4632 9680 4644
rect 9732 4632 9738 4684
rect 9766 4632 9772 4684
rect 9824 4672 9830 4684
rect 10321 4675 10379 4681
rect 10321 4672 10333 4675
rect 9824 4644 10333 4672
rect 9824 4632 9830 4644
rect 10321 4641 10333 4644
rect 10367 4641 10379 4675
rect 11146 4672 11152 4684
rect 11107 4644 11152 4672
rect 10321 4635 10379 4641
rect 11146 4632 11152 4644
rect 11204 4632 11210 4684
rect 10137 4607 10195 4613
rect 10137 4604 10149 4607
rect 9508 4576 10149 4604
rect 10137 4573 10149 4576
rect 10183 4573 10195 4607
rect 10137 4567 10195 4573
rect 10226 4564 10232 4616
rect 10284 4604 10290 4616
rect 10962 4604 10968 4616
rect 10284 4576 10329 4604
rect 10923 4576 10968 4604
rect 10284 4564 10290 4576
rect 10962 4564 10968 4576
rect 11020 4564 11026 4616
rect 7650 4496 7656 4548
rect 7708 4536 7714 4548
rect 9309 4539 9367 4545
rect 9309 4536 9321 4539
rect 7708 4508 9321 4536
rect 7708 4496 7714 4508
rect 9309 4505 9321 4508
rect 9355 4505 9367 4539
rect 9309 4499 9367 4505
rect 7834 4468 7840 4480
rect 5684 4440 7052 4468
rect 7795 4440 7840 4468
rect 5684 4428 5690 4440
rect 7834 4428 7840 4440
rect 7892 4428 7898 4480
rect 7926 4428 7932 4480
rect 7984 4468 7990 4480
rect 8297 4471 8355 4477
rect 7984 4440 8029 4468
rect 7984 4428 7990 4440
rect 8297 4437 8309 4471
rect 8343 4468 8355 4471
rect 8938 4468 8944 4480
rect 8343 4440 8944 4468
rect 8343 4437 8355 4440
rect 8297 4431 8355 4437
rect 8938 4428 8944 4440
rect 8996 4428 9002 4480
rect 9214 4428 9220 4480
rect 9272 4468 9278 4480
rect 9401 4471 9459 4477
rect 9401 4468 9413 4471
rect 9272 4440 9413 4468
rect 9272 4428 9278 4440
rect 9401 4437 9413 4440
rect 9447 4437 9459 4471
rect 9401 4431 9459 4437
rect 11057 4471 11115 4477
rect 11057 4437 11069 4471
rect 11103 4468 11115 4471
rect 11425 4471 11483 4477
rect 11425 4468 11437 4471
rect 11103 4440 11437 4468
rect 11103 4437 11115 4440
rect 11057 4431 11115 4437
rect 11425 4437 11437 4440
rect 11471 4437 11483 4471
rect 11532 4468 11560 4712
rect 13078 4700 13084 4752
rect 13136 4740 13142 4752
rect 13136 4712 13181 4740
rect 13136 4700 13142 4712
rect 11974 4672 11980 4684
rect 11935 4644 11980 4672
rect 11974 4632 11980 4644
rect 12032 4632 12038 4684
rect 12529 4675 12587 4681
rect 12529 4641 12541 4675
rect 12575 4672 12587 4675
rect 12710 4672 12716 4684
rect 12575 4644 12716 4672
rect 12575 4641 12587 4644
rect 12529 4635 12587 4641
rect 12710 4632 12716 4644
rect 12768 4632 12774 4684
rect 12986 4632 12992 4684
rect 13044 4672 13050 4684
rect 13354 4672 13360 4684
rect 13044 4644 13360 4672
rect 13044 4632 13050 4644
rect 13354 4632 13360 4644
rect 13412 4632 13418 4684
rect 13648 4681 13676 4780
rect 14292 4780 17684 4808
rect 13633 4675 13691 4681
rect 13633 4641 13645 4675
rect 13679 4641 13691 4675
rect 13633 4635 13691 4641
rect 13722 4632 13728 4684
rect 13780 4672 13786 4684
rect 14292 4681 14320 4780
rect 17678 4768 17684 4780
rect 17736 4768 17742 4820
rect 18230 4768 18236 4820
rect 18288 4808 18294 4820
rect 18874 4808 18880 4820
rect 18288 4780 18880 4808
rect 18288 4768 18294 4780
rect 18874 4768 18880 4780
rect 18932 4768 18938 4820
rect 14921 4743 14979 4749
rect 14921 4709 14933 4743
rect 14967 4740 14979 4743
rect 14967 4712 18828 4740
rect 14967 4709 14979 4712
rect 14921 4703 14979 4709
rect 14277 4675 14335 4681
rect 13780 4644 13825 4672
rect 13780 4632 13786 4644
rect 14277 4641 14289 4675
rect 14323 4641 14335 4675
rect 14458 4672 14464 4684
rect 14419 4644 14464 4672
rect 14277 4635 14335 4641
rect 14458 4632 14464 4644
rect 14516 4632 14522 4684
rect 15197 4675 15255 4681
rect 15197 4641 15209 4675
rect 15243 4672 15255 4675
rect 16298 4672 16304 4684
rect 15243 4644 16304 4672
rect 15243 4641 15255 4644
rect 15197 4635 15255 4641
rect 16298 4632 16304 4644
rect 16356 4632 16362 4684
rect 16485 4675 16543 4681
rect 16485 4641 16497 4675
rect 16531 4672 16543 4675
rect 16942 4672 16948 4684
rect 16531 4644 16948 4672
rect 16531 4641 16543 4644
rect 16485 4635 16543 4641
rect 16942 4632 16948 4644
rect 17000 4672 17006 4684
rect 17221 4675 17279 4681
rect 17221 4672 17233 4675
rect 17000 4644 17233 4672
rect 17000 4632 17006 4644
rect 17221 4641 17233 4644
rect 17267 4641 17279 4675
rect 17678 4672 17684 4684
rect 17639 4644 17684 4672
rect 17221 4635 17279 4641
rect 17678 4632 17684 4644
rect 17736 4632 17742 4684
rect 17773 4675 17831 4681
rect 17773 4641 17785 4675
rect 17819 4672 17831 4675
rect 18046 4672 18052 4684
rect 17819 4644 18052 4672
rect 17819 4641 17831 4644
rect 17773 4635 17831 4641
rect 18046 4632 18052 4644
rect 18104 4632 18110 4684
rect 18800 4681 18828 4712
rect 22002 4700 22008 4752
rect 22060 4740 22066 4752
rect 22646 4740 22652 4752
rect 22060 4712 22652 4740
rect 22060 4700 22066 4712
rect 22646 4700 22652 4712
rect 22704 4700 22710 4752
rect 18785 4675 18843 4681
rect 18785 4641 18797 4675
rect 18831 4641 18843 4675
rect 18785 4635 18843 4641
rect 18874 4632 18880 4684
rect 18932 4672 18938 4684
rect 19429 4675 19487 4681
rect 18932 4644 18977 4672
rect 18932 4632 18938 4644
rect 19429 4641 19441 4675
rect 19475 4672 19487 4675
rect 19610 4672 19616 4684
rect 19475 4644 19616 4672
rect 19475 4641 19487 4644
rect 19429 4635 19487 4641
rect 19610 4632 19616 4644
rect 19668 4632 19674 4684
rect 20717 4675 20775 4681
rect 20717 4641 20729 4675
rect 20763 4672 20775 4675
rect 21910 4672 21916 4684
rect 20763 4644 21916 4672
rect 20763 4641 20775 4644
rect 20717 4635 20775 4641
rect 21910 4632 21916 4644
rect 21968 4632 21974 4684
rect 11793 4607 11851 4613
rect 11793 4573 11805 4607
rect 11839 4604 11851 4607
rect 12894 4604 12900 4616
rect 11839 4576 12900 4604
rect 11839 4573 11851 4576
rect 11793 4567 11851 4573
rect 12894 4564 12900 4576
rect 12952 4564 12958 4616
rect 13078 4564 13084 4616
rect 13136 4604 13142 4616
rect 13541 4607 13599 4613
rect 13541 4604 13553 4607
rect 13136 4576 13553 4604
rect 13136 4564 13142 4576
rect 13541 4573 13553 4576
rect 13587 4573 13599 4607
rect 13541 4567 13599 4573
rect 14550 4564 14556 4616
rect 14608 4564 14614 4616
rect 15286 4604 15292 4616
rect 15247 4576 15292 4604
rect 15286 4564 15292 4576
rect 15344 4564 15350 4616
rect 15381 4607 15439 4613
rect 15381 4573 15393 4607
rect 15427 4604 15439 4607
rect 15562 4604 15568 4616
rect 15427 4576 15568 4604
rect 15427 4573 15439 4576
rect 15381 4567 15439 4573
rect 15562 4564 15568 4576
rect 15620 4564 15626 4616
rect 16209 4607 16267 4613
rect 16209 4573 16221 4607
rect 16255 4604 16267 4607
rect 16390 4604 16396 4616
rect 16255 4576 16396 4604
rect 16255 4573 16267 4576
rect 16209 4567 16267 4573
rect 16390 4564 16396 4576
rect 16448 4564 16454 4616
rect 16574 4564 16580 4616
rect 16632 4604 16638 4616
rect 20349 4607 20407 4613
rect 20349 4604 20361 4607
rect 16632 4576 20361 4604
rect 16632 4564 16638 4576
rect 20349 4573 20361 4576
rect 20395 4573 20407 4607
rect 20990 4604 20996 4616
rect 20951 4576 20996 4604
rect 20349 4567 20407 4573
rect 20990 4564 20996 4576
rect 21048 4564 21054 4616
rect 12526 4496 12532 4548
rect 12584 4536 12590 4548
rect 12621 4539 12679 4545
rect 12621 4536 12633 4539
rect 12584 4508 12633 4536
rect 12584 4496 12590 4508
rect 12621 4505 12633 4508
rect 12667 4505 12679 4539
rect 12621 4499 12679 4505
rect 12710 4496 12716 4548
rect 12768 4536 12774 4548
rect 14568 4536 14596 4564
rect 12768 4508 14596 4536
rect 12768 4496 12774 4508
rect 15102 4496 15108 4548
rect 15160 4536 15166 4548
rect 15160 4508 15884 4536
rect 15160 4496 15166 4508
rect 11885 4471 11943 4477
rect 11885 4468 11897 4471
rect 11532 4440 11897 4468
rect 11425 4431 11483 4437
rect 11885 4437 11897 4440
rect 11931 4468 11943 4471
rect 11974 4468 11980 4480
rect 11931 4440 11980 4468
rect 11931 4437 11943 4440
rect 11885 4431 11943 4437
rect 11974 4428 11980 4440
rect 12032 4428 12038 4480
rect 13170 4468 13176 4480
rect 13131 4440 13176 4468
rect 13170 4428 13176 4440
rect 13228 4428 13234 4480
rect 14550 4468 14556 4480
rect 14511 4440 14556 4468
rect 14550 4428 14556 4440
rect 14608 4428 14614 4480
rect 15746 4468 15752 4480
rect 15707 4440 15752 4468
rect 15746 4428 15752 4440
rect 15804 4428 15810 4480
rect 15856 4477 15884 4508
rect 16114 4496 16120 4548
rect 16172 4536 16178 4548
rect 16301 4539 16359 4545
rect 16301 4536 16313 4539
rect 16172 4508 16313 4536
rect 16172 4496 16178 4508
rect 16301 4505 16313 4508
rect 16347 4505 16359 4539
rect 16301 4499 16359 4505
rect 16942 4496 16948 4548
rect 17000 4536 17006 4548
rect 17037 4539 17095 4545
rect 17037 4536 17049 4539
rect 17000 4508 17049 4536
rect 17000 4496 17006 4508
rect 17037 4505 17049 4508
rect 17083 4536 17095 4539
rect 17218 4536 17224 4548
rect 17083 4508 17224 4536
rect 17083 4505 17095 4508
rect 17037 4499 17095 4505
rect 17218 4496 17224 4508
rect 17276 4496 17282 4548
rect 17770 4496 17776 4548
rect 17828 4536 17834 4548
rect 17865 4539 17923 4545
rect 17865 4536 17877 4539
rect 17828 4508 17877 4536
rect 17828 4496 17834 4508
rect 17865 4505 17877 4508
rect 17911 4505 17923 4539
rect 18693 4539 18751 4545
rect 18693 4536 18705 4539
rect 17865 4499 17923 4505
rect 18248 4508 18705 4536
rect 15841 4471 15899 4477
rect 15841 4437 15853 4471
rect 15887 4437 15899 4471
rect 15841 4431 15899 4437
rect 16390 4428 16396 4480
rect 16448 4468 16454 4480
rect 16669 4471 16727 4477
rect 16669 4468 16681 4471
rect 16448 4440 16681 4468
rect 16448 4428 16454 4440
rect 16669 4437 16681 4440
rect 16715 4437 16727 4471
rect 16669 4431 16727 4437
rect 16758 4428 16764 4480
rect 16816 4468 16822 4480
rect 17129 4471 17187 4477
rect 17129 4468 17141 4471
rect 16816 4440 17141 4468
rect 16816 4428 16822 4440
rect 17129 4437 17141 4440
rect 17175 4468 17187 4471
rect 17954 4468 17960 4480
rect 17175 4440 17960 4468
rect 17175 4437 17187 4440
rect 17129 4431 17187 4437
rect 17954 4428 17960 4440
rect 18012 4428 18018 4480
rect 18248 4477 18276 4508
rect 18693 4505 18705 4508
rect 18739 4505 18751 4539
rect 20533 4539 20591 4545
rect 20533 4536 20545 4539
rect 18693 4499 18751 4505
rect 19306 4508 20545 4536
rect 18233 4471 18291 4477
rect 18233 4437 18245 4471
rect 18279 4437 18291 4471
rect 18233 4431 18291 4437
rect 18322 4428 18328 4480
rect 18380 4468 18386 4480
rect 18380 4440 18425 4468
rect 18380 4428 18386 4440
rect 18598 4428 18604 4480
rect 18656 4468 18662 4480
rect 19306 4468 19334 4508
rect 20533 4505 20545 4508
rect 20579 4505 20591 4539
rect 20533 4499 20591 4505
rect 19518 4468 19524 4480
rect 18656 4440 19334 4468
rect 19479 4440 19524 4468
rect 18656 4428 18662 4440
rect 19518 4428 19524 4440
rect 19576 4428 19582 4480
rect 19610 4428 19616 4480
rect 19668 4468 19674 4480
rect 19978 4468 19984 4480
rect 19668 4440 19713 4468
rect 19939 4440 19984 4468
rect 19668 4428 19674 4440
rect 19978 4428 19984 4440
rect 20036 4428 20042 4480
rect 20070 4428 20076 4480
rect 20128 4468 20134 4480
rect 20128 4440 20173 4468
rect 20128 4428 20134 4440
rect 1104 4378 22056 4400
rect 1104 4326 6148 4378
rect 6200 4326 6212 4378
rect 6264 4326 6276 4378
rect 6328 4326 6340 4378
rect 6392 4326 6404 4378
rect 6456 4326 11346 4378
rect 11398 4326 11410 4378
rect 11462 4326 11474 4378
rect 11526 4326 11538 4378
rect 11590 4326 11602 4378
rect 11654 4326 16544 4378
rect 16596 4326 16608 4378
rect 16660 4326 16672 4378
rect 16724 4326 16736 4378
rect 16788 4326 16800 4378
rect 16852 4326 21742 4378
rect 21794 4326 21806 4378
rect 21858 4326 21870 4378
rect 21922 4326 21934 4378
rect 21986 4326 21998 4378
rect 22050 4326 22056 4378
rect 1104 4304 22056 4326
rect 2038 4224 2044 4276
rect 2096 4264 2102 4276
rect 2225 4267 2283 4273
rect 2225 4264 2237 4267
rect 2096 4236 2237 4264
rect 2096 4224 2102 4236
rect 2225 4233 2237 4236
rect 2271 4233 2283 4267
rect 4154 4264 4160 4276
rect 4115 4236 4160 4264
rect 2225 4227 2283 4233
rect 4154 4224 4160 4236
rect 4212 4224 4218 4276
rect 4430 4224 4436 4276
rect 4488 4264 4494 4276
rect 5445 4267 5503 4273
rect 5445 4264 5457 4267
rect 4488 4236 5457 4264
rect 4488 4224 4494 4236
rect 5445 4233 5457 4236
rect 5491 4233 5503 4267
rect 5810 4264 5816 4276
rect 5771 4236 5816 4264
rect 5445 4227 5503 4233
rect 5810 4224 5816 4236
rect 5868 4224 5874 4276
rect 5905 4267 5963 4273
rect 5905 4233 5917 4267
rect 5951 4264 5963 4267
rect 6086 4264 6092 4276
rect 5951 4236 6092 4264
rect 5951 4233 5963 4236
rect 5905 4227 5963 4233
rect 6086 4224 6092 4236
rect 6144 4224 6150 4276
rect 6914 4264 6920 4276
rect 6748 4236 6920 4264
rect 2317 4199 2375 4205
rect 2317 4165 2329 4199
rect 2363 4196 2375 4199
rect 5258 4196 5264 4208
rect 2363 4168 5264 4196
rect 2363 4165 2375 4168
rect 2317 4159 2375 4165
rect 5258 4156 5264 4168
rect 5316 4156 5322 4208
rect 5350 4156 5356 4208
rect 5408 4196 5414 4208
rect 6748 4196 6776 4236
rect 6914 4224 6920 4236
rect 6972 4224 6978 4276
rect 7098 4224 7104 4276
rect 7156 4264 7162 4276
rect 10965 4267 11023 4273
rect 10965 4264 10977 4267
rect 7156 4236 10977 4264
rect 7156 4224 7162 4236
rect 10965 4233 10977 4236
rect 11011 4233 11023 4267
rect 10965 4227 11023 4233
rect 11793 4267 11851 4273
rect 11793 4233 11805 4267
rect 11839 4264 11851 4267
rect 11974 4264 11980 4276
rect 11839 4236 11980 4264
rect 11839 4233 11851 4236
rect 11793 4227 11851 4233
rect 11974 4224 11980 4236
rect 12032 4224 12038 4276
rect 12526 4264 12532 4276
rect 12084 4236 12532 4264
rect 7190 4196 7196 4208
rect 5408 4168 6776 4196
rect 6840 4168 7196 4196
rect 5408 4156 5414 4168
rect 1397 4131 1455 4137
rect 1397 4097 1409 4131
rect 1443 4128 1455 4131
rect 1486 4128 1492 4140
rect 1443 4100 1492 4128
rect 1443 4097 1455 4100
rect 1397 4091 1455 4097
rect 1486 4088 1492 4100
rect 1544 4088 1550 4140
rect 1857 4131 1915 4137
rect 1857 4097 1869 4131
rect 1903 4097 1915 4131
rect 1857 4091 1915 4097
rect 1670 3992 1676 4004
rect 1631 3964 1676 3992
rect 1670 3952 1676 3964
rect 1728 3952 1734 4004
rect 1581 3927 1639 3933
rect 1581 3893 1593 3927
rect 1627 3924 1639 3927
rect 1872 3924 1900 4091
rect 2774 4088 2780 4140
rect 2832 4128 2838 4140
rect 3044 4131 3102 4137
rect 2832 4100 2877 4128
rect 2832 4088 2838 4100
rect 3044 4097 3056 4131
rect 3090 4128 3102 4131
rect 3326 4128 3332 4140
rect 3090 4100 3332 4128
rect 3090 4097 3102 4100
rect 3044 4091 3102 4097
rect 3326 4088 3332 4100
rect 3384 4088 3390 4140
rect 4246 4128 4252 4140
rect 4207 4100 4252 4128
rect 4246 4088 4252 4100
rect 4304 4088 4310 4140
rect 4982 4128 4988 4140
rect 4943 4100 4988 4128
rect 4982 4088 4988 4100
rect 5040 4088 5046 4140
rect 6362 4128 6368 4140
rect 5184 4100 6132 4128
rect 6323 4100 6368 4128
rect 2130 4060 2136 4072
rect 2091 4032 2136 4060
rect 2130 4020 2136 4032
rect 2188 4020 2194 4072
rect 5074 4060 5080 4072
rect 5035 4032 5080 4060
rect 5074 4020 5080 4032
rect 5132 4020 5138 4072
rect 2682 3992 2688 4004
rect 2643 3964 2688 3992
rect 2682 3952 2688 3964
rect 2740 3952 2746 4004
rect 4246 3952 4252 4004
rect 4304 3992 4310 4004
rect 4433 3995 4491 4001
rect 4433 3992 4445 3995
rect 4304 3964 4445 3992
rect 4304 3952 4310 3964
rect 4433 3961 4445 3964
rect 4479 3961 4491 3995
rect 4433 3955 4491 3961
rect 4890 3952 4896 4004
rect 4948 3992 4954 4004
rect 5184 3992 5212 4100
rect 5261 4063 5319 4069
rect 5261 4029 5273 4063
rect 5307 4029 5319 4063
rect 5994 4060 6000 4072
rect 5955 4032 6000 4060
rect 5261 4023 5319 4029
rect 4948 3964 5212 3992
rect 5276 3992 5304 4023
rect 5994 4020 6000 4032
rect 6052 4020 6058 4072
rect 6104 4060 6132 4100
rect 6362 4088 6368 4100
rect 6420 4088 6426 4140
rect 6641 4131 6699 4137
rect 6641 4097 6653 4131
rect 6687 4128 6699 4131
rect 6730 4128 6736 4140
rect 6687 4100 6736 4128
rect 6687 4097 6699 4100
rect 6641 4091 6699 4097
rect 6730 4088 6736 4100
rect 6788 4088 6794 4140
rect 6840 4137 6868 4168
rect 7190 4156 7196 4168
rect 7248 4156 7254 4208
rect 7374 4156 7380 4208
rect 7432 4156 7438 4208
rect 7466 4156 7472 4208
rect 7524 4196 7530 4208
rect 7926 4196 7932 4208
rect 7524 4168 7932 4196
rect 7524 4156 7530 4168
rect 7926 4156 7932 4168
rect 7984 4156 7990 4208
rect 8110 4156 8116 4208
rect 8168 4196 8174 4208
rect 8941 4199 8999 4205
rect 8941 4196 8953 4199
rect 8168 4168 8953 4196
rect 8168 4156 8174 4168
rect 8941 4165 8953 4168
rect 8987 4165 8999 4199
rect 8941 4159 8999 4165
rect 9030 4156 9036 4208
rect 9088 4196 9094 4208
rect 9088 4168 9133 4196
rect 9088 4156 9094 4168
rect 11238 4156 11244 4208
rect 11296 4196 11302 4208
rect 12084 4196 12112 4236
rect 12526 4224 12532 4236
rect 12584 4224 12590 4276
rect 13170 4224 13176 4276
rect 13228 4264 13234 4276
rect 13357 4267 13415 4273
rect 13357 4264 13369 4267
rect 13228 4236 13369 4264
rect 13228 4224 13234 4236
rect 13357 4233 13369 4236
rect 13403 4233 13415 4267
rect 13357 4227 13415 4233
rect 13446 4224 13452 4276
rect 13504 4264 13510 4276
rect 14277 4267 14335 4273
rect 14277 4264 14289 4267
rect 13504 4236 14289 4264
rect 13504 4224 13510 4236
rect 14277 4233 14289 4236
rect 14323 4233 14335 4267
rect 14277 4227 14335 4233
rect 14737 4267 14795 4273
rect 14737 4233 14749 4267
rect 14783 4233 14795 4267
rect 14737 4227 14795 4233
rect 11296 4168 12112 4196
rect 11296 4156 11302 4168
rect 12434 4156 12440 4208
rect 12492 4196 12498 4208
rect 12492 4168 13492 4196
rect 12492 4156 12498 4168
rect 6825 4131 6883 4137
rect 6825 4097 6837 4131
rect 6871 4097 6883 4131
rect 6825 4091 6883 4097
rect 7276 4131 7334 4137
rect 7276 4097 7288 4131
rect 7322 4128 7334 4131
rect 7392 4128 7420 4156
rect 7322 4100 7420 4128
rect 7322 4097 7334 4100
rect 7276 4091 7334 4097
rect 7558 4088 7564 4140
rect 7616 4128 7622 4140
rect 8386 4128 8392 4140
rect 7616 4100 8392 4128
rect 7616 4088 7622 4100
rect 8386 4088 8392 4100
rect 8444 4088 8450 4140
rect 9582 4128 9588 4140
rect 9543 4100 9588 4128
rect 9582 4088 9588 4100
rect 9640 4088 9646 4140
rect 9861 4131 9919 4137
rect 9861 4097 9873 4131
rect 9907 4128 9919 4131
rect 9907 4100 10272 4128
rect 9907 4097 9919 4100
rect 9861 4091 9919 4097
rect 10244 4072 10272 4100
rect 10318 4088 10324 4140
rect 10376 4128 10382 4140
rect 11606 4128 11612 4140
rect 10376 4100 11468 4128
rect 11567 4100 11612 4128
rect 10376 4088 10382 4100
rect 7006 4060 7012 4072
rect 6104 4032 7012 4060
rect 7006 4020 7012 4032
rect 7064 4020 7070 4072
rect 9217 4063 9275 4069
rect 9217 4029 9229 4063
rect 9263 4060 9275 4063
rect 9674 4060 9680 4072
rect 9263 4032 9680 4060
rect 9263 4029 9275 4032
rect 9217 4023 9275 4029
rect 9674 4020 9680 4032
rect 9732 4020 9738 4072
rect 10226 4060 10232 4072
rect 10187 4032 10232 4060
rect 10226 4020 10232 4032
rect 10284 4020 10290 4072
rect 11057 4063 11115 4069
rect 11057 4060 11069 4063
rect 10336 4032 11069 4060
rect 5534 3992 5540 4004
rect 5276 3964 5540 3992
rect 4948 3952 4954 3964
rect 5534 3952 5540 3964
rect 5592 3992 5598 4004
rect 6638 3992 6644 4004
rect 5592 3964 6644 3992
rect 5592 3952 5598 3964
rect 6638 3952 6644 3964
rect 6696 3952 6702 4004
rect 8202 3952 8208 4004
rect 8260 3992 8266 4004
rect 8389 3995 8447 4001
rect 8389 3992 8401 3995
rect 8260 3964 8401 3992
rect 8260 3952 8266 3964
rect 8389 3961 8401 3964
rect 8435 3961 8447 3995
rect 8570 3992 8576 4004
rect 8531 3964 8576 3992
rect 8389 3955 8447 3961
rect 8570 3952 8576 3964
rect 8628 3952 8634 4004
rect 10336 3992 10364 4032
rect 11057 4029 11069 4032
rect 11103 4029 11115 4063
rect 11057 4023 11115 4029
rect 11149 4063 11207 4069
rect 11149 4029 11161 4063
rect 11195 4029 11207 4063
rect 11440 4060 11468 4100
rect 11606 4088 11612 4100
rect 11664 4088 11670 4140
rect 11885 4131 11943 4137
rect 11885 4128 11897 4131
rect 11716 4100 11897 4128
rect 11716 4060 11744 4100
rect 11885 4097 11897 4100
rect 11931 4097 11943 4131
rect 11885 4091 11943 4097
rect 12066 4088 12072 4140
rect 12124 4128 12130 4140
rect 12161 4131 12219 4137
rect 12161 4128 12173 4131
rect 12124 4100 12173 4128
rect 12124 4088 12130 4100
rect 12161 4097 12173 4100
rect 12207 4097 12219 4131
rect 12161 4091 12219 4097
rect 12621 4131 12679 4137
rect 12621 4097 12633 4131
rect 12667 4128 12679 4131
rect 13262 4128 13268 4140
rect 12667 4100 13268 4128
rect 12667 4097 12679 4100
rect 12621 4091 12679 4097
rect 13262 4088 13268 4100
rect 13320 4088 13326 4140
rect 13464 4137 13492 4168
rect 13449 4131 13507 4137
rect 13449 4097 13461 4131
rect 13495 4128 13507 4131
rect 14185 4131 14243 4137
rect 14743 4132 14771 4227
rect 15102 4224 15108 4276
rect 15160 4264 15166 4276
rect 15197 4267 15255 4273
rect 15197 4264 15209 4267
rect 15160 4236 15209 4264
rect 15160 4224 15166 4236
rect 15197 4233 15209 4236
rect 15243 4233 15255 4267
rect 15930 4264 15936 4276
rect 15891 4236 15936 4264
rect 15197 4227 15255 4233
rect 15930 4224 15936 4236
rect 15988 4224 15994 4276
rect 17678 4264 17684 4276
rect 16684 4236 17684 4264
rect 16390 4196 16396 4208
rect 15120 4168 16396 4196
rect 15120 4137 15148 4168
rect 16390 4156 16396 4168
rect 16448 4156 16454 4208
rect 16684 4137 16712 4236
rect 17678 4224 17684 4236
rect 17736 4224 17742 4276
rect 18325 4267 18383 4273
rect 18325 4233 18337 4267
rect 18371 4264 18383 4267
rect 18414 4264 18420 4276
rect 18371 4236 18420 4264
rect 18371 4233 18383 4236
rect 18325 4227 18383 4233
rect 18414 4224 18420 4236
rect 18472 4224 18478 4276
rect 18785 4267 18843 4273
rect 18785 4233 18797 4267
rect 18831 4264 18843 4267
rect 19245 4267 19303 4273
rect 19245 4264 19257 4267
rect 18831 4236 19257 4264
rect 18831 4233 18843 4236
rect 18785 4227 18843 4233
rect 19245 4233 19257 4236
rect 19291 4233 19303 4267
rect 19245 4227 19303 4233
rect 19613 4267 19671 4273
rect 19613 4233 19625 4267
rect 19659 4264 19671 4267
rect 20070 4264 20076 4276
rect 19659 4236 20076 4264
rect 19659 4233 19671 4236
rect 19613 4227 19671 4233
rect 20070 4224 20076 4236
rect 20128 4224 20134 4276
rect 17034 4196 17040 4208
rect 16947 4168 17040 4196
rect 16960 4137 16988 4168
rect 17034 4156 17040 4168
rect 17092 4196 17098 4208
rect 18230 4196 18236 4208
rect 17092 4168 18236 4196
rect 17092 4156 17098 4168
rect 18230 4156 18236 4168
rect 18288 4156 18294 4208
rect 19794 4156 19800 4208
rect 19852 4196 19858 4208
rect 19852 4168 19932 4196
rect 19852 4156 19858 4168
rect 17218 4137 17224 4140
rect 13495 4100 14044 4128
rect 13495 4097 13507 4100
rect 13449 4091 13507 4097
rect 12986 4060 12992 4072
rect 11440 4032 11744 4060
rect 11799 4032 12992 4060
rect 11149 4023 11207 4029
rect 8671 3964 10364 3992
rect 1627 3896 1900 3924
rect 1627 3893 1639 3896
rect 1581 3887 1639 3893
rect 4614 3884 4620 3936
rect 4672 3924 4678 3936
rect 6546 3924 6552 3936
rect 4672 3896 4717 3924
rect 6507 3896 6552 3924
rect 4672 3884 4678 3896
rect 6546 3884 6552 3896
rect 6604 3884 6610 3936
rect 6730 3884 6736 3936
rect 6788 3924 6794 3936
rect 8671 3924 8699 3964
rect 10502 3952 10508 4004
rect 10560 3992 10566 4004
rect 11164 3992 11192 4023
rect 11799 3992 11827 4032
rect 12986 4020 12992 4032
rect 13044 4020 13050 4072
rect 13170 4060 13176 4072
rect 13131 4032 13176 4060
rect 13170 4020 13176 4032
rect 13228 4060 13234 4072
rect 13538 4060 13544 4072
rect 13228 4032 13544 4060
rect 13228 4020 13234 4032
rect 13538 4020 13544 4032
rect 13596 4020 13602 4072
rect 10560 3964 11192 3992
rect 11716 3964 11827 3992
rect 12805 3995 12863 4001
rect 10560 3952 10566 3964
rect 6788 3896 8699 3924
rect 6788 3884 6794 3896
rect 8938 3884 8944 3936
rect 8996 3924 9002 3936
rect 9214 3924 9220 3936
rect 8996 3896 9220 3924
rect 8996 3884 9002 3896
rect 9214 3884 9220 3896
rect 9272 3884 9278 3936
rect 9490 3924 9496 3936
rect 9451 3896 9496 3924
rect 9490 3884 9496 3896
rect 9548 3884 9554 3936
rect 9674 3884 9680 3936
rect 9732 3924 9738 3936
rect 10597 3927 10655 3933
rect 10597 3924 10609 3927
rect 9732 3896 10609 3924
rect 9732 3884 9738 3896
rect 10597 3893 10609 3896
rect 10643 3893 10655 3927
rect 10597 3887 10655 3893
rect 10686 3884 10692 3936
rect 10744 3924 10750 3936
rect 11716 3924 11744 3964
rect 12805 3961 12817 3995
rect 12851 3992 12863 3995
rect 13722 3992 13728 4004
rect 12851 3964 13728 3992
rect 12851 3961 12863 3964
rect 12805 3955 12863 3961
rect 13722 3952 13728 3964
rect 13780 3952 13786 4004
rect 14016 3992 14044 4100
rect 14185 4097 14197 4131
rect 14231 4128 14243 4131
rect 14691 4128 14771 4132
rect 14231 4104 14771 4128
rect 15105 4131 15163 4137
rect 14231 4100 14719 4104
rect 14231 4097 14243 4100
rect 14185 4091 14243 4097
rect 15105 4097 15117 4131
rect 15151 4097 15163 4131
rect 16669 4131 16727 4137
rect 16669 4128 16681 4131
rect 15105 4091 15163 4097
rect 15764 4100 16681 4128
rect 14093 4063 14151 4069
rect 14093 4029 14105 4063
rect 14139 4060 14151 4063
rect 14274 4060 14280 4072
rect 14139 4032 14280 4060
rect 14139 4029 14151 4032
rect 14093 4023 14151 4029
rect 14274 4020 14280 4032
rect 14332 4020 14338 4072
rect 15286 4060 15292 4072
rect 15247 4032 15292 4060
rect 15286 4020 15292 4032
rect 15344 4020 15350 4072
rect 15764 4069 15792 4100
rect 16669 4097 16681 4100
rect 16715 4097 16727 4131
rect 16669 4091 16727 4097
rect 16945 4131 17003 4137
rect 16945 4097 16957 4131
rect 16991 4097 17003 4131
rect 17212 4128 17224 4137
rect 17179 4100 17224 4128
rect 16945 4091 17003 4097
rect 17212 4091 17224 4100
rect 17218 4088 17224 4091
rect 17276 4088 17282 4140
rect 18874 4088 18880 4140
rect 18932 4128 18938 4140
rect 18932 4100 19840 4128
rect 18932 4088 18938 4100
rect 15749 4063 15807 4069
rect 15749 4029 15761 4063
rect 15795 4029 15807 4063
rect 15749 4023 15807 4029
rect 15838 4020 15844 4072
rect 15896 4060 15902 4072
rect 16390 4060 16396 4072
rect 15896 4032 15941 4060
rect 16351 4032 16396 4060
rect 15896 4020 15902 4032
rect 16390 4020 16396 4032
rect 16448 4020 16454 4072
rect 18414 4020 18420 4072
rect 18472 4060 18478 4072
rect 18509 4063 18567 4069
rect 18509 4060 18521 4063
rect 18472 4032 18521 4060
rect 18472 4020 18478 4032
rect 18509 4029 18521 4032
rect 18555 4029 18567 4063
rect 18690 4060 18696 4072
rect 18651 4032 18696 4060
rect 18509 4023 18567 4029
rect 18690 4020 18696 4032
rect 18748 4020 18754 4072
rect 19058 4020 19064 4072
rect 19116 4020 19122 4072
rect 19812 4069 19840 4100
rect 19705 4063 19763 4069
rect 19705 4029 19717 4063
rect 19751 4029 19763 4063
rect 19705 4023 19763 4029
rect 19797 4063 19855 4069
rect 19797 4029 19809 4063
rect 19843 4029 19855 4063
rect 19904 4060 19932 4168
rect 19978 4088 19984 4140
rect 20036 4128 20042 4140
rect 20257 4131 20315 4137
rect 20257 4128 20269 4131
rect 20036 4100 20269 4128
rect 20036 4088 20042 4100
rect 20257 4097 20269 4100
rect 20303 4097 20315 4131
rect 20257 4091 20315 4097
rect 20346 4088 20352 4140
rect 20404 4128 20410 4140
rect 20533 4131 20591 4137
rect 20533 4128 20545 4131
rect 20404 4100 20545 4128
rect 20404 4088 20410 4100
rect 20533 4097 20545 4100
rect 20579 4097 20591 4131
rect 20993 4131 21051 4137
rect 20993 4128 21005 4131
rect 20533 4091 20591 4097
rect 20640 4100 21005 4128
rect 20640 4060 20668 4100
rect 20993 4097 21005 4100
rect 21039 4097 21051 4131
rect 20993 4091 21051 4097
rect 19904 4032 20668 4060
rect 20717 4063 20775 4069
rect 19797 4023 19855 4029
rect 20717 4029 20729 4063
rect 20763 4060 20775 4063
rect 20806 4060 20812 4072
rect 20763 4032 20812 4060
rect 20763 4029 20775 4032
rect 20717 4023 20775 4029
rect 15010 3992 15016 4004
rect 14016 3964 15016 3992
rect 15010 3952 15016 3964
rect 15068 3952 15074 4004
rect 12066 3924 12072 3936
rect 10744 3896 11744 3924
rect 12027 3896 12072 3924
rect 10744 3884 10750 3896
rect 12066 3884 12072 3896
rect 12124 3884 12130 3936
rect 12342 3924 12348 3936
rect 12303 3896 12348 3924
rect 12342 3884 12348 3896
rect 12400 3884 12406 3936
rect 12986 3924 12992 3936
rect 12947 3896 12992 3924
rect 12986 3884 12992 3896
rect 13044 3884 13050 3936
rect 13817 3927 13875 3933
rect 13817 3893 13829 3927
rect 13863 3924 13875 3927
rect 14458 3924 14464 3936
rect 13863 3896 14464 3924
rect 13863 3893 13875 3896
rect 13817 3887 13875 3893
rect 14458 3884 14464 3896
rect 14516 3884 14522 3936
rect 14550 3884 14556 3936
rect 14608 3924 14614 3936
rect 14645 3927 14703 3933
rect 14645 3924 14657 3927
rect 14608 3896 14657 3924
rect 14608 3884 14614 3896
rect 14645 3893 14657 3896
rect 14691 3893 14703 3927
rect 16298 3924 16304 3936
rect 16259 3896 16304 3924
rect 14645 3887 14703 3893
rect 16298 3884 16304 3896
rect 16356 3884 16362 3936
rect 16850 3924 16856 3936
rect 16811 3896 16856 3924
rect 16850 3884 16856 3896
rect 16908 3884 16914 3936
rect 19076 3924 19104 4020
rect 19153 3995 19211 4001
rect 19153 3961 19165 3995
rect 19199 3992 19211 3995
rect 19610 3992 19616 4004
rect 19199 3964 19616 3992
rect 19199 3961 19211 3964
rect 19153 3955 19211 3961
rect 19610 3952 19616 3964
rect 19668 3952 19674 4004
rect 19720 3992 19748 4023
rect 20806 4020 20812 4032
rect 20864 4020 20870 4072
rect 19978 3992 19984 4004
rect 19720 3964 19984 3992
rect 19978 3952 19984 3964
rect 20036 3952 20042 4004
rect 20073 3927 20131 3933
rect 20073 3924 20085 3927
rect 19076 3896 20085 3924
rect 20073 3893 20085 3896
rect 20119 3893 20131 3927
rect 20073 3887 20131 3893
rect 20349 3927 20407 3933
rect 20349 3893 20361 3927
rect 20395 3924 20407 3927
rect 20438 3924 20444 3936
rect 20395 3896 20444 3924
rect 20395 3893 20407 3896
rect 20349 3887 20407 3893
rect 20438 3884 20444 3896
rect 20496 3884 20502 3936
rect 1104 3834 21896 3856
rect 1104 3782 3549 3834
rect 3601 3782 3613 3834
rect 3665 3782 3677 3834
rect 3729 3782 3741 3834
rect 3793 3782 3805 3834
rect 3857 3782 8747 3834
rect 8799 3782 8811 3834
rect 8863 3782 8875 3834
rect 8927 3782 8939 3834
rect 8991 3782 9003 3834
rect 9055 3782 13945 3834
rect 13997 3782 14009 3834
rect 14061 3782 14073 3834
rect 14125 3782 14137 3834
rect 14189 3782 14201 3834
rect 14253 3782 19143 3834
rect 19195 3782 19207 3834
rect 19259 3782 19271 3834
rect 19323 3782 19335 3834
rect 19387 3782 19399 3834
rect 19451 3782 21896 3834
rect 1104 3760 21896 3782
rect 1857 3723 1915 3729
rect 1857 3689 1869 3723
rect 1903 3720 1915 3723
rect 1903 3692 3464 3720
rect 1903 3689 1915 3692
rect 1857 3683 1915 3689
rect 750 3612 756 3664
rect 808 3652 814 3664
rect 1946 3652 1952 3664
rect 808 3624 1952 3652
rect 808 3612 814 3624
rect 1946 3612 1952 3624
rect 2004 3612 2010 3664
rect 3326 3652 3332 3664
rect 3239 3624 3332 3652
rect 3326 3612 3332 3624
rect 3384 3612 3390 3664
rect 3436 3652 3464 3692
rect 3510 3680 3516 3732
rect 3568 3720 3574 3732
rect 5166 3720 5172 3732
rect 3568 3692 5172 3720
rect 3568 3680 3574 3692
rect 5166 3680 5172 3692
rect 5224 3680 5230 3732
rect 5902 3680 5908 3732
rect 5960 3720 5966 3732
rect 6365 3723 6423 3729
rect 5960 3692 6224 3720
rect 5960 3680 5966 3692
rect 3786 3652 3792 3664
rect 3436 3624 3792 3652
rect 3786 3612 3792 3624
rect 3844 3612 3850 3664
rect 5537 3655 5595 3661
rect 5537 3621 5549 3655
rect 5583 3652 5595 3655
rect 5994 3652 6000 3664
rect 5583 3624 6000 3652
rect 5583 3621 5595 3624
rect 5537 3615 5595 3621
rect 5994 3612 6000 3624
rect 6052 3612 6058 3664
rect 6196 3652 6224 3692
rect 6365 3689 6377 3723
rect 6411 3720 6423 3723
rect 7834 3720 7840 3732
rect 6411 3692 7840 3720
rect 6411 3689 6423 3692
rect 6365 3683 6423 3689
rect 7834 3680 7840 3692
rect 7892 3680 7898 3732
rect 7926 3680 7932 3732
rect 7984 3720 7990 3732
rect 10318 3720 10324 3732
rect 7984 3692 10324 3720
rect 7984 3680 7990 3692
rect 10318 3680 10324 3692
rect 10376 3680 10382 3732
rect 10505 3723 10563 3729
rect 10505 3689 10517 3723
rect 10551 3720 10563 3723
rect 11606 3720 11612 3732
rect 10551 3692 11612 3720
rect 10551 3689 10563 3692
rect 10505 3683 10563 3689
rect 11606 3680 11612 3692
rect 11664 3720 11670 3732
rect 12158 3720 12164 3732
rect 11664 3692 12164 3720
rect 11664 3680 11670 3692
rect 12158 3680 12164 3692
rect 12216 3680 12222 3732
rect 13262 3680 13268 3732
rect 13320 3720 13326 3732
rect 14093 3723 14151 3729
rect 14093 3720 14105 3723
rect 13320 3692 14105 3720
rect 13320 3680 13326 3692
rect 14093 3689 14105 3692
rect 14139 3689 14151 3723
rect 14093 3683 14151 3689
rect 15565 3723 15623 3729
rect 15565 3689 15577 3723
rect 15611 3720 15623 3723
rect 16114 3720 16120 3732
rect 15611 3692 16120 3720
rect 15611 3689 15623 3692
rect 15565 3683 15623 3689
rect 16114 3680 16120 3692
rect 16172 3680 16178 3732
rect 16298 3680 16304 3732
rect 16356 3720 16362 3732
rect 17957 3723 18015 3729
rect 16356 3692 17448 3720
rect 16356 3680 16362 3692
rect 6822 3652 6828 3664
rect 6196 3624 6828 3652
rect 6822 3612 6828 3624
rect 6880 3612 6886 3664
rect 8202 3652 8208 3664
rect 8128 3624 8208 3652
rect 3344 3584 3372 3612
rect 5813 3587 5871 3593
rect 3344 3556 3924 3584
rect 1394 3516 1400 3528
rect 1355 3488 1400 3516
rect 1394 3476 1400 3488
rect 1452 3476 1458 3528
rect 1673 3519 1731 3525
rect 1673 3485 1685 3519
rect 1719 3485 1731 3519
rect 1673 3479 1731 3485
rect 1949 3519 2007 3525
rect 1949 3485 1961 3519
rect 1995 3516 2007 3519
rect 2774 3516 2780 3528
rect 1995 3488 2780 3516
rect 1995 3485 2007 3488
rect 1949 3479 2007 3485
rect 1210 3408 1216 3460
rect 1268 3448 1274 3460
rect 1688 3448 1716 3479
rect 2774 3476 2780 3488
rect 2832 3476 2838 3528
rect 3418 3516 3424 3528
rect 3379 3488 3424 3516
rect 3418 3476 3424 3488
rect 3476 3476 3482 3528
rect 3789 3519 3847 3525
rect 3789 3485 3801 3519
rect 3835 3485 3847 3519
rect 3896 3516 3924 3556
rect 5813 3553 5825 3587
rect 5859 3584 5871 3587
rect 6270 3584 6276 3596
rect 5859 3556 6276 3584
rect 5859 3553 5871 3556
rect 5813 3547 5871 3553
rect 6270 3544 6276 3556
rect 6328 3544 6334 3596
rect 8128 3593 8156 3624
rect 8202 3612 8208 3624
rect 8260 3652 8266 3664
rect 10597 3655 10655 3661
rect 8260 3624 8984 3652
rect 8260 3612 8266 3624
rect 8113 3587 8171 3593
rect 8113 3553 8125 3587
rect 8159 3553 8171 3587
rect 8294 3584 8300 3596
rect 8255 3556 8300 3584
rect 8113 3547 8171 3553
rect 8294 3544 8300 3556
rect 8352 3544 8358 3596
rect 8956 3584 8984 3624
rect 10597 3621 10609 3655
rect 10643 3652 10655 3655
rect 10870 3652 10876 3664
rect 10643 3624 10876 3652
rect 10643 3621 10655 3624
rect 10597 3615 10655 3621
rect 10870 3612 10876 3624
rect 10928 3612 10934 3664
rect 12253 3655 12311 3661
rect 12253 3652 12265 3655
rect 11992 3624 12265 3652
rect 11992 3593 12020 3624
rect 12253 3621 12265 3624
rect 12299 3621 12311 3655
rect 12253 3615 12311 3621
rect 12434 3612 12440 3664
rect 12492 3612 12498 3664
rect 13538 3612 13544 3664
rect 13596 3652 13602 3664
rect 15105 3655 15163 3661
rect 13596 3624 14688 3652
rect 13596 3612 13602 3624
rect 11977 3587 12035 3593
rect 8956 3556 9076 3584
rect 7834 3516 7840 3528
rect 3896 3488 7696 3516
rect 7795 3488 7840 3516
rect 3789 3479 3847 3485
rect 1268 3420 1716 3448
rect 1268 3408 1274 3420
rect 1578 3380 1584 3392
rect 1539 3352 1584 3380
rect 1578 3340 1584 3352
rect 1636 3340 1642 3392
rect 1688 3380 1716 3420
rect 2216 3451 2274 3457
rect 2216 3417 2228 3451
rect 2262 3448 2274 3451
rect 2498 3448 2504 3460
rect 2262 3420 2504 3448
rect 2262 3417 2274 3420
rect 2216 3411 2274 3417
rect 2498 3408 2504 3420
rect 2556 3408 2562 3460
rect 2792 3448 2820 3476
rect 3804 3448 3832 3479
rect 2792 3420 3832 3448
rect 4056 3451 4114 3457
rect 4056 3417 4068 3451
rect 4102 3448 4114 3451
rect 4154 3448 4160 3460
rect 4102 3420 4160 3448
rect 4102 3417 4114 3420
rect 4056 3411 4114 3417
rect 4154 3408 4160 3420
rect 4212 3448 4218 3460
rect 4706 3448 4712 3460
rect 4212 3420 4712 3448
rect 4212 3408 4218 3420
rect 4706 3408 4712 3420
rect 4764 3408 4770 3460
rect 5350 3448 5356 3460
rect 5311 3420 5356 3448
rect 5350 3408 5356 3420
rect 5408 3408 5414 3460
rect 5442 3408 5448 3460
rect 5500 3448 5506 3460
rect 6638 3448 6644 3460
rect 5500 3420 6644 3448
rect 5500 3408 5506 3420
rect 6638 3408 6644 3420
rect 6696 3408 6702 3460
rect 7570 3451 7628 3457
rect 7570 3417 7582 3451
rect 7616 3417 7628 3451
rect 7668 3448 7696 3488
rect 7834 3476 7840 3488
rect 7892 3476 7898 3528
rect 8018 3476 8024 3528
rect 8076 3516 8082 3528
rect 8938 3516 8944 3528
rect 8076 3488 8944 3516
rect 8076 3476 8082 3488
rect 8938 3476 8944 3488
rect 8996 3476 9002 3528
rect 9048 3516 9076 3556
rect 11977 3553 11989 3587
rect 12023 3553 12035 3587
rect 11977 3547 12035 3553
rect 12161 3587 12219 3593
rect 12161 3553 12173 3587
rect 12207 3584 12219 3587
rect 12452 3584 12480 3612
rect 14550 3584 14556 3596
rect 12207 3556 12480 3584
rect 14511 3556 14556 3584
rect 12207 3553 12219 3556
rect 12161 3547 12219 3553
rect 9197 3519 9255 3525
rect 9197 3516 9209 3519
rect 9048 3488 9209 3516
rect 9197 3485 9209 3488
rect 9243 3485 9255 3519
rect 10502 3516 10508 3528
rect 9197 3479 9255 3485
rect 9646 3488 10508 3516
rect 9646 3448 9674 3488
rect 10502 3476 10508 3488
rect 10560 3476 10566 3528
rect 10870 3476 10876 3528
rect 10928 3516 10934 3528
rect 11992 3516 12020 3547
rect 14550 3544 14556 3556
rect 14608 3544 14614 3596
rect 14660 3593 14688 3624
rect 15105 3621 15117 3655
rect 15151 3652 15163 3655
rect 15286 3652 15292 3664
rect 15151 3624 15292 3652
rect 15151 3621 15163 3624
rect 15105 3615 15163 3621
rect 15286 3612 15292 3624
rect 15344 3612 15350 3664
rect 14645 3587 14703 3593
rect 14645 3553 14657 3587
rect 14691 3553 14703 3587
rect 17218 3584 17224 3596
rect 14645 3547 14703 3553
rect 16960 3556 17224 3584
rect 10928 3488 12020 3516
rect 12437 3519 12495 3525
rect 10928 3476 10934 3488
rect 12437 3485 12449 3519
rect 12483 3516 12495 3519
rect 12529 3519 12587 3525
rect 12529 3516 12541 3519
rect 12483 3488 12541 3516
rect 12483 3485 12495 3488
rect 12437 3479 12495 3485
rect 12529 3485 12541 3488
rect 12575 3516 12587 3519
rect 13262 3516 13268 3528
rect 12575 3488 13268 3516
rect 12575 3485 12587 3488
rect 12529 3479 12587 3485
rect 13262 3476 13268 3488
rect 13320 3476 13326 3528
rect 13630 3476 13636 3528
rect 13688 3516 13694 3528
rect 13688 3488 14320 3516
rect 13688 3476 13694 3488
rect 7668 3420 9674 3448
rect 7570 3411 7628 3417
rect 3050 3380 3056 3392
rect 1688 3352 3056 3380
rect 3050 3340 3056 3352
rect 3108 3340 3114 3392
rect 3605 3383 3663 3389
rect 3605 3349 3617 3383
rect 3651 3380 3663 3383
rect 3878 3380 3884 3392
rect 3651 3352 3884 3380
rect 3651 3349 3663 3352
rect 3605 3343 3663 3349
rect 3878 3340 3884 3352
rect 3936 3340 3942 3392
rect 4246 3340 4252 3392
rect 4304 3380 4310 3392
rect 5258 3380 5264 3392
rect 4304 3352 5264 3380
rect 4304 3340 4310 3352
rect 5258 3340 5264 3352
rect 5316 3340 5322 3392
rect 5902 3380 5908 3392
rect 5863 3352 5908 3380
rect 5902 3340 5908 3352
rect 5960 3340 5966 3392
rect 5994 3340 6000 3392
rect 6052 3380 6058 3392
rect 6052 3352 6097 3380
rect 6052 3340 6058 3352
rect 6270 3340 6276 3392
rect 6328 3380 6334 3392
rect 6457 3383 6515 3389
rect 6457 3380 6469 3383
rect 6328 3352 6469 3380
rect 6328 3340 6334 3352
rect 6457 3349 6469 3352
rect 6503 3380 6515 3383
rect 7374 3380 7380 3392
rect 6503 3352 7380 3380
rect 6503 3349 6515 3352
rect 6457 3343 6515 3349
rect 7374 3340 7380 3352
rect 7432 3340 7438 3392
rect 7585 3380 7613 3411
rect 10134 3408 10140 3460
rect 10192 3448 10198 3460
rect 10686 3448 10692 3460
rect 10192 3420 10692 3448
rect 10192 3408 10198 3420
rect 10686 3408 10692 3420
rect 10744 3408 10750 3460
rect 11732 3451 11790 3457
rect 11732 3417 11744 3451
rect 11778 3448 11790 3451
rect 12796 3451 12854 3457
rect 11778 3420 12434 3448
rect 11778 3417 11790 3420
rect 11732 3411 11790 3417
rect 7742 3380 7748 3392
rect 7585 3352 7748 3380
rect 7742 3340 7748 3352
rect 7800 3380 7806 3392
rect 8018 3380 8024 3392
rect 7800 3352 8024 3380
rect 7800 3340 7806 3352
rect 8018 3340 8024 3352
rect 8076 3340 8082 3392
rect 8386 3380 8392 3392
rect 8347 3352 8392 3380
rect 8386 3340 8392 3352
rect 8444 3340 8450 3392
rect 8757 3383 8815 3389
rect 8757 3349 8769 3383
rect 8803 3380 8815 3383
rect 9398 3380 9404 3392
rect 8803 3352 9404 3380
rect 8803 3349 8815 3352
rect 8757 3343 8815 3349
rect 9398 3340 9404 3352
rect 9456 3340 9462 3392
rect 10226 3340 10232 3392
rect 10284 3380 10290 3392
rect 10321 3383 10379 3389
rect 10321 3380 10333 3383
rect 10284 3352 10333 3380
rect 10284 3340 10290 3352
rect 10321 3349 10333 3352
rect 10367 3349 10379 3383
rect 12406 3380 12434 3420
rect 12796 3417 12808 3451
rect 12842 3448 12854 3451
rect 13170 3448 13176 3460
rect 12842 3420 13176 3448
rect 12842 3417 12854 3420
rect 12796 3411 12854 3417
rect 13170 3408 13176 3420
rect 13228 3408 13234 3460
rect 14292 3448 14320 3488
rect 14734 3476 14740 3528
rect 14792 3516 14798 3528
rect 14921 3519 14979 3525
rect 14921 3516 14933 3519
rect 14792 3488 14933 3516
rect 14792 3476 14798 3488
rect 14921 3485 14933 3488
rect 14967 3485 14979 3519
rect 16960 3516 16988 3556
rect 17218 3544 17224 3556
rect 17276 3584 17282 3596
rect 17313 3587 17371 3593
rect 17313 3584 17325 3587
rect 17276 3556 17325 3584
rect 17276 3544 17282 3556
rect 17313 3553 17325 3556
rect 17359 3553 17371 3587
rect 17420 3584 17448 3692
rect 17957 3689 17969 3723
rect 18003 3720 18015 3723
rect 18690 3720 18696 3732
rect 18003 3692 18696 3720
rect 18003 3689 18015 3692
rect 17957 3683 18015 3689
rect 18690 3680 18696 3692
rect 18748 3680 18754 3732
rect 20441 3723 20499 3729
rect 20441 3689 20453 3723
rect 20487 3720 20499 3723
rect 20714 3720 20720 3732
rect 20487 3692 20720 3720
rect 20487 3689 20499 3692
rect 20441 3683 20499 3689
rect 20714 3680 20720 3692
rect 20772 3680 20778 3732
rect 18414 3652 18420 3664
rect 18156 3624 18420 3652
rect 18156 3593 18184 3624
rect 18414 3612 18420 3624
rect 18472 3612 18478 3664
rect 18782 3612 18788 3664
rect 18840 3652 18846 3664
rect 19337 3655 19395 3661
rect 19337 3652 19349 3655
rect 18840 3624 19349 3652
rect 18840 3612 18846 3624
rect 19337 3621 19349 3624
rect 19383 3621 19395 3655
rect 19337 3615 19395 3621
rect 19613 3655 19671 3661
rect 19613 3621 19625 3655
rect 19659 3621 19671 3655
rect 20254 3652 20260 3664
rect 19613 3615 19671 3621
rect 20088 3624 20260 3652
rect 17497 3587 17555 3593
rect 17497 3584 17509 3587
rect 17420 3556 17509 3584
rect 17313 3547 17371 3553
rect 17497 3553 17509 3556
rect 17543 3553 17555 3587
rect 17497 3547 17555 3553
rect 18141 3587 18199 3593
rect 18141 3553 18153 3587
rect 18187 3553 18199 3587
rect 18322 3584 18328 3596
rect 18283 3556 18328 3584
rect 18141 3547 18199 3553
rect 14921 3479 14979 3485
rect 15672 3488 16988 3516
rect 15010 3448 15016 3460
rect 14292 3420 15016 3448
rect 15010 3408 15016 3420
rect 15068 3408 15074 3460
rect 13538 3380 13544 3392
rect 12406 3352 13544 3380
rect 10321 3343 10379 3349
rect 13538 3340 13544 3352
rect 13596 3340 13602 3392
rect 13906 3380 13912 3392
rect 13819 3352 13912 3380
rect 13906 3340 13912 3352
rect 13964 3380 13970 3392
rect 14182 3380 14188 3392
rect 13964 3352 14188 3380
rect 13964 3340 13970 3352
rect 14182 3340 14188 3352
rect 14240 3340 14246 3392
rect 14274 3340 14280 3392
rect 14332 3380 14338 3392
rect 14461 3383 14519 3389
rect 14461 3380 14473 3383
rect 14332 3352 14473 3380
rect 14332 3340 14338 3352
rect 14461 3349 14473 3352
rect 14507 3349 14519 3383
rect 14461 3343 14519 3349
rect 15194 3340 15200 3392
rect 15252 3380 15258 3392
rect 15672 3389 15700 3488
rect 17034 3476 17040 3528
rect 17092 3516 17098 3528
rect 17328 3516 17356 3547
rect 18322 3544 18328 3556
rect 18380 3544 18386 3596
rect 19628 3584 19656 3615
rect 18432 3556 19656 3584
rect 17092 3488 17137 3516
rect 17328 3488 18184 3516
rect 17092 3476 17098 3488
rect 16022 3408 16028 3460
rect 16080 3448 16086 3460
rect 16390 3448 16396 3460
rect 16080 3420 16396 3448
rect 16080 3408 16086 3420
rect 16390 3408 16396 3420
rect 16448 3408 16454 3460
rect 16850 3457 16856 3460
rect 16792 3451 16856 3457
rect 16792 3448 16804 3451
rect 16763 3420 16804 3448
rect 16792 3417 16804 3420
rect 16838 3417 16856 3451
rect 16792 3411 16856 3417
rect 16850 3408 16856 3411
rect 16908 3448 16914 3460
rect 17862 3448 17868 3460
rect 16908 3420 17868 3448
rect 16908 3408 16914 3420
rect 17862 3408 17868 3420
rect 17920 3408 17926 3460
rect 18156 3448 18184 3488
rect 18230 3476 18236 3528
rect 18288 3516 18294 3528
rect 18432 3516 18460 3556
rect 18874 3516 18880 3528
rect 18288 3488 18460 3516
rect 18708 3488 18880 3516
rect 18288 3476 18294 3488
rect 18708 3460 18736 3488
rect 18874 3476 18880 3488
rect 18932 3476 18938 3528
rect 19058 3516 19064 3528
rect 19019 3488 19064 3516
rect 19058 3476 19064 3488
rect 19116 3476 19122 3528
rect 19521 3519 19579 3525
rect 19521 3485 19533 3519
rect 19567 3485 19579 3519
rect 19521 3479 19579 3485
rect 19797 3519 19855 3525
rect 19797 3485 19809 3519
rect 19843 3516 19855 3519
rect 19886 3516 19892 3528
rect 19843 3488 19892 3516
rect 19843 3485 19855 3488
rect 19797 3479 19855 3485
rect 18690 3448 18696 3460
rect 18156 3420 18696 3448
rect 18690 3408 18696 3420
rect 18748 3408 18754 3460
rect 19426 3448 19432 3460
rect 18800 3420 19432 3448
rect 15657 3383 15715 3389
rect 15252 3352 15297 3380
rect 15252 3340 15258 3352
rect 15657 3349 15669 3383
rect 15703 3349 15715 3383
rect 15657 3343 15715 3349
rect 15746 3340 15752 3392
rect 15804 3380 15810 3392
rect 16298 3380 16304 3392
rect 15804 3352 16304 3380
rect 15804 3340 15810 3352
rect 16298 3340 16304 3352
rect 16356 3340 16362 3392
rect 17126 3340 17132 3392
rect 17184 3380 17190 3392
rect 17494 3380 17500 3392
rect 17184 3352 17500 3380
rect 17184 3340 17190 3352
rect 17494 3340 17500 3352
rect 17552 3340 17558 3392
rect 17589 3383 17647 3389
rect 17589 3349 17601 3383
rect 17635 3380 17647 3383
rect 17678 3380 17684 3392
rect 17635 3352 17684 3380
rect 17635 3349 17647 3352
rect 17589 3343 17647 3349
rect 17678 3340 17684 3352
rect 17736 3340 17742 3392
rect 18138 3340 18144 3392
rect 18196 3380 18202 3392
rect 18800 3389 18828 3420
rect 19426 3408 19432 3420
rect 19484 3408 19490 3460
rect 19536 3448 19564 3479
rect 19886 3476 19892 3488
rect 19944 3476 19950 3528
rect 20088 3525 20116 3624
rect 20254 3612 20260 3624
rect 20312 3652 20318 3664
rect 21358 3652 21364 3664
rect 20312 3624 21364 3652
rect 20312 3612 20318 3624
rect 21358 3612 21364 3624
rect 21416 3612 21422 3664
rect 20898 3544 20904 3596
rect 20956 3584 20962 3596
rect 20993 3587 21051 3593
rect 20993 3584 21005 3587
rect 20956 3556 21005 3584
rect 20956 3544 20962 3556
rect 20993 3553 21005 3556
rect 21039 3553 21051 3587
rect 20993 3547 21051 3553
rect 20073 3519 20131 3525
rect 20073 3485 20085 3519
rect 20119 3485 20131 3519
rect 20346 3516 20352 3528
rect 20307 3488 20352 3516
rect 20073 3479 20131 3485
rect 20346 3476 20352 3488
rect 20404 3476 20410 3528
rect 21453 3519 21511 3525
rect 21453 3485 21465 3519
rect 21499 3516 21511 3519
rect 22094 3516 22100 3528
rect 21499 3488 22100 3516
rect 21499 3485 21511 3488
rect 21453 3479 21511 3485
rect 22094 3476 22100 3488
rect 22152 3476 22158 3528
rect 20806 3448 20812 3460
rect 19536 3420 20208 3448
rect 20767 3420 20812 3448
rect 18417 3383 18475 3389
rect 18417 3380 18429 3383
rect 18196 3352 18429 3380
rect 18196 3340 18202 3352
rect 18417 3349 18429 3352
rect 18463 3349 18475 3383
rect 18417 3343 18475 3349
rect 18785 3383 18843 3389
rect 18785 3349 18797 3383
rect 18831 3349 18843 3383
rect 18785 3343 18843 3349
rect 18874 3340 18880 3392
rect 18932 3380 18938 3392
rect 19886 3380 19892 3392
rect 18932 3352 18977 3380
rect 19847 3352 19892 3380
rect 18932 3340 18938 3352
rect 19886 3340 19892 3352
rect 19944 3340 19950 3392
rect 20180 3389 20208 3420
rect 20806 3408 20812 3420
rect 20864 3408 20870 3460
rect 20901 3451 20959 3457
rect 20901 3417 20913 3451
rect 20947 3448 20959 3451
rect 21082 3448 21088 3460
rect 20947 3420 21088 3448
rect 20947 3417 20959 3420
rect 20901 3411 20959 3417
rect 21082 3408 21088 3420
rect 21140 3408 21146 3460
rect 20165 3383 20223 3389
rect 20165 3349 20177 3383
rect 20211 3349 20223 3383
rect 20165 3343 20223 3349
rect 20714 3340 20720 3392
rect 20772 3380 20778 3392
rect 21361 3383 21419 3389
rect 21361 3380 21373 3383
rect 20772 3352 21373 3380
rect 20772 3340 20778 3352
rect 21361 3349 21373 3352
rect 21407 3349 21419 3383
rect 21361 3343 21419 3349
rect 1104 3290 22056 3312
rect 1104 3238 6148 3290
rect 6200 3238 6212 3290
rect 6264 3238 6276 3290
rect 6328 3238 6340 3290
rect 6392 3238 6404 3290
rect 6456 3238 11346 3290
rect 11398 3238 11410 3290
rect 11462 3238 11474 3290
rect 11526 3238 11538 3290
rect 11590 3238 11602 3290
rect 11654 3238 16544 3290
rect 16596 3238 16608 3290
rect 16660 3238 16672 3290
rect 16724 3238 16736 3290
rect 16788 3238 16800 3290
rect 16852 3238 21742 3290
rect 21794 3238 21806 3290
rect 21858 3238 21870 3290
rect 21922 3238 21934 3290
rect 21986 3238 21998 3290
rect 22050 3238 22056 3290
rect 1104 3216 22056 3238
rect 2406 3176 2412 3188
rect 2367 3148 2412 3176
rect 2406 3136 2412 3148
rect 2464 3136 2470 3188
rect 2501 3179 2559 3185
rect 2501 3145 2513 3179
rect 2547 3176 2559 3179
rect 2961 3179 3019 3185
rect 2961 3176 2973 3179
rect 2547 3148 2973 3176
rect 2547 3145 2559 3148
rect 2501 3139 2559 3145
rect 2961 3145 2973 3148
rect 3007 3145 3019 3179
rect 2961 3139 3019 3145
rect 3421 3179 3479 3185
rect 3421 3145 3433 3179
rect 3467 3176 3479 3179
rect 4614 3176 4620 3188
rect 3467 3148 4620 3176
rect 3467 3145 3479 3148
rect 3421 3139 3479 3145
rect 4614 3136 4620 3148
rect 4672 3136 4678 3188
rect 4706 3136 4712 3188
rect 4764 3176 4770 3188
rect 5810 3176 5816 3188
rect 4764 3148 5816 3176
rect 4764 3136 4770 3148
rect 5810 3136 5816 3148
rect 5868 3136 5874 3188
rect 5902 3136 5908 3188
rect 5960 3176 5966 3188
rect 6457 3179 6515 3185
rect 6457 3176 6469 3179
rect 5960 3148 6469 3176
rect 5960 3136 5966 3148
rect 6457 3145 6469 3148
rect 6503 3145 6515 3179
rect 6457 3139 6515 3145
rect 6546 3136 6552 3188
rect 6604 3176 6610 3188
rect 6822 3176 6828 3188
rect 6604 3148 6828 3176
rect 6604 3136 6610 3148
rect 6822 3136 6828 3148
rect 6880 3176 6886 3188
rect 6917 3179 6975 3185
rect 6917 3176 6929 3179
rect 6880 3148 6929 3176
rect 6880 3136 6886 3148
rect 6917 3145 6929 3148
rect 6963 3145 6975 3179
rect 6917 3139 6975 3145
rect 7006 3136 7012 3188
rect 7064 3176 7070 3188
rect 7834 3176 7840 3188
rect 7064 3148 7840 3176
rect 7064 3136 7070 3148
rect 7834 3136 7840 3148
rect 7892 3136 7898 3188
rect 7926 3136 7932 3188
rect 7984 3176 7990 3188
rect 9398 3176 9404 3188
rect 7984 3148 8892 3176
rect 9359 3148 9404 3176
rect 7984 3136 7990 3148
rect 1118 3068 1124 3120
rect 1176 3108 1182 3120
rect 4062 3108 4068 3120
rect 1176 3080 4068 3108
rect 1176 3068 1182 3080
rect 1596 3049 1624 3080
rect 4062 3068 4068 3080
rect 4120 3068 4126 3120
rect 5068 3111 5126 3117
rect 4540 3080 5028 3108
rect 1581 3043 1639 3049
rect 1581 3009 1593 3043
rect 1627 3009 1639 3043
rect 1581 3003 1639 3009
rect 1857 3043 1915 3049
rect 1857 3009 1869 3043
rect 1903 3040 1915 3043
rect 2682 3040 2688 3052
rect 1903 3012 2688 3040
rect 1903 3009 1915 3012
rect 1857 3003 1915 3009
rect 2682 3000 2688 3012
rect 2740 3000 2746 3052
rect 3326 3040 3332 3052
rect 3287 3012 3332 3040
rect 3326 3000 3332 3012
rect 3384 3000 3390 3052
rect 4540 3040 4568 3080
rect 4264 3012 4568 3040
rect 4617 3043 4675 3049
rect 2317 2975 2375 2981
rect 2317 2941 2329 2975
rect 2363 2972 2375 2975
rect 2498 2972 2504 2984
rect 2363 2944 2504 2972
rect 2363 2941 2375 2944
rect 2317 2935 2375 2941
rect 2498 2932 2504 2944
rect 2556 2972 2562 2984
rect 3510 2972 3516 2984
rect 2556 2944 3516 2972
rect 2556 2932 2562 2944
rect 3510 2932 3516 2944
rect 3568 2932 3574 2984
rect 3605 2975 3663 2981
rect 3605 2941 3617 2975
rect 3651 2972 3663 2975
rect 4154 2972 4160 2984
rect 3651 2944 4160 2972
rect 3651 2941 3663 2944
rect 3605 2935 3663 2941
rect 4154 2932 4160 2944
rect 4212 2932 4218 2984
rect 1489 2907 1547 2913
rect 1489 2873 1501 2907
rect 1535 2904 1547 2907
rect 1854 2904 1860 2916
rect 1535 2876 1860 2904
rect 1535 2873 1547 2876
rect 1489 2867 1547 2873
rect 1854 2864 1860 2876
rect 1912 2864 1918 2916
rect 2869 2907 2927 2913
rect 2148 2876 2774 2904
rect 2148 2848 2176 2876
rect 1762 2836 1768 2848
rect 1723 2808 1768 2836
rect 1762 2796 1768 2808
rect 1820 2796 1826 2848
rect 2038 2836 2044 2848
rect 1999 2808 2044 2836
rect 2038 2796 2044 2808
rect 2096 2796 2102 2848
rect 2130 2796 2136 2848
rect 2188 2796 2194 2848
rect 2746 2836 2774 2876
rect 2869 2873 2881 2907
rect 2915 2904 2927 2907
rect 4264 2904 4292 3012
rect 4617 3009 4629 3043
rect 4663 3009 4675 3043
rect 4617 3003 4675 3009
rect 4801 3043 4859 3049
rect 4801 3009 4813 3043
rect 4847 3040 4859 3043
rect 4890 3040 4896 3052
rect 4847 3012 4896 3040
rect 4847 3009 4859 3012
rect 4801 3003 4859 3009
rect 4341 2975 4399 2981
rect 4341 2941 4353 2975
rect 4387 2941 4399 2975
rect 4341 2935 4399 2941
rect 2915 2876 4292 2904
rect 2915 2873 2927 2876
rect 2869 2867 2927 2873
rect 4246 2836 4252 2848
rect 2746 2808 4252 2836
rect 4246 2796 4252 2808
rect 4304 2796 4310 2848
rect 4356 2836 4384 2935
rect 4632 2916 4660 3003
rect 4890 3000 4896 3012
rect 4948 3000 4954 3052
rect 5000 3040 5028 3080
rect 5068 3077 5080 3111
rect 5114 3108 5126 3111
rect 5442 3108 5448 3120
rect 5114 3080 5448 3108
rect 5114 3077 5126 3080
rect 5068 3071 5126 3077
rect 5442 3068 5448 3080
rect 5500 3068 5506 3120
rect 7392 3080 8800 3108
rect 6730 3040 6736 3052
rect 5000 3012 6736 3040
rect 6730 3000 6736 3012
rect 6788 3000 6794 3052
rect 6825 3043 6883 3049
rect 6825 3009 6837 3043
rect 6871 3040 6883 3043
rect 6914 3040 6920 3052
rect 6871 3012 6920 3040
rect 6871 3009 6883 3012
rect 6825 3003 6883 3009
rect 6914 3000 6920 3012
rect 6972 3000 6978 3052
rect 7101 2975 7159 2981
rect 7101 2941 7113 2975
rect 7147 2972 7159 2975
rect 7282 2972 7288 2984
rect 7147 2944 7288 2972
rect 7147 2941 7159 2944
rect 7101 2935 7159 2941
rect 7282 2932 7288 2944
rect 7340 2972 7346 2984
rect 7392 2981 7420 3080
rect 7650 3040 7656 3052
rect 7611 3012 7656 3040
rect 7650 3000 7656 3012
rect 7708 3000 7714 3052
rect 8481 3043 8539 3049
rect 8481 3009 8493 3043
rect 8527 3009 8539 3043
rect 8481 3003 8539 3009
rect 7377 2975 7435 2981
rect 7377 2972 7389 2975
rect 7340 2944 7389 2972
rect 7340 2932 7346 2944
rect 7377 2941 7389 2944
rect 7423 2941 7435 2975
rect 7377 2935 7435 2941
rect 7466 2932 7472 2984
rect 7524 2972 7530 2984
rect 7561 2975 7619 2981
rect 7561 2972 7573 2975
rect 7524 2944 7573 2972
rect 7524 2932 7530 2944
rect 7561 2941 7573 2944
rect 7607 2941 7619 2975
rect 7561 2935 7619 2941
rect 8294 2932 8300 2984
rect 8352 2972 8358 2984
rect 8496 2972 8524 3003
rect 8352 2944 8524 2972
rect 8352 2932 8358 2944
rect 8570 2932 8576 2984
rect 8628 2972 8634 2984
rect 8772 2981 8800 3080
rect 8864 3040 8892 3148
rect 9398 3136 9404 3148
rect 9456 3136 9462 3188
rect 9861 3179 9919 3185
rect 9861 3145 9873 3179
rect 9907 3176 9919 3179
rect 10318 3176 10324 3188
rect 9907 3148 10324 3176
rect 9907 3145 9919 3148
rect 9861 3139 9919 3145
rect 10318 3136 10324 3148
rect 10376 3136 10382 3188
rect 12342 3176 12348 3188
rect 12084 3148 12348 3176
rect 9214 3068 9220 3120
rect 9272 3108 9278 3120
rect 9309 3111 9367 3117
rect 9309 3108 9321 3111
rect 9272 3080 9321 3108
rect 9272 3068 9278 3080
rect 9309 3077 9321 3080
rect 9355 3077 9367 3111
rect 9766 3108 9772 3120
rect 9309 3071 9367 3077
rect 9416 3080 9772 3108
rect 9416 3040 9444 3080
rect 9766 3068 9772 3080
rect 9824 3068 9830 3120
rect 11977 3111 12035 3117
rect 11977 3077 11989 3111
rect 12023 3108 12035 3111
rect 12084 3108 12112 3148
rect 12342 3136 12348 3148
rect 12400 3136 12406 3188
rect 12805 3179 12863 3185
rect 12805 3145 12817 3179
rect 12851 3176 12863 3179
rect 13538 3176 13544 3188
rect 12851 3148 13544 3176
rect 12851 3145 12863 3148
rect 12805 3139 12863 3145
rect 13538 3136 13544 3148
rect 13596 3136 13602 3188
rect 14274 3176 14280 3188
rect 14235 3148 14280 3176
rect 14274 3136 14280 3148
rect 14332 3136 14338 3188
rect 14458 3136 14464 3188
rect 14516 3176 14522 3188
rect 14737 3179 14795 3185
rect 14737 3176 14749 3179
rect 14516 3148 14749 3176
rect 14516 3136 14522 3148
rect 14737 3145 14749 3148
rect 14783 3145 14795 3179
rect 14737 3139 14795 3145
rect 16390 3136 16396 3188
rect 16448 3176 16454 3188
rect 16448 3148 17540 3176
rect 16448 3136 16454 3148
rect 12526 3108 12532 3120
rect 12023 3080 12112 3108
rect 12023 3077 12035 3080
rect 11977 3071 12035 3077
rect 10226 3049 10232 3052
rect 9876 3040 9996 3044
rect 10209 3043 10232 3049
rect 10209 3040 10221 3043
rect 8864 3012 9444 3040
rect 9600 3016 10221 3040
rect 9600 3012 9904 3016
rect 9968 3012 10221 3016
rect 8757 2975 8815 2981
rect 8628 2944 8673 2972
rect 8628 2932 8634 2944
rect 8757 2941 8769 2975
rect 8803 2941 8815 2975
rect 8757 2935 8815 2941
rect 8938 2932 8944 2984
rect 8996 2972 9002 2984
rect 9600 2981 9628 3012
rect 10209 3009 10221 3012
rect 10284 3040 10290 3052
rect 11885 3043 11943 3049
rect 10284 3012 10357 3040
rect 11885 3036 11897 3043
rect 11931 3036 11943 3043
rect 10209 3003 10232 3009
rect 10226 3000 10232 3003
rect 10284 3000 10290 3012
rect 11882 2984 11888 3036
rect 11940 2984 11946 3036
rect 9585 2975 9643 2981
rect 8996 2944 9536 2972
rect 8996 2932 9002 2944
rect 4614 2864 4620 2916
rect 4672 2864 4678 2916
rect 5810 2864 5816 2916
rect 5868 2904 5874 2916
rect 6181 2907 6239 2913
rect 6181 2904 6193 2907
rect 5868 2876 6193 2904
rect 5868 2864 5874 2876
rect 6181 2873 6193 2876
rect 6227 2904 6239 2907
rect 7926 2904 7932 2916
rect 6227 2876 7932 2904
rect 6227 2873 6239 2876
rect 6181 2867 6239 2873
rect 7926 2864 7932 2876
rect 7984 2864 7990 2916
rect 8021 2907 8079 2913
rect 8021 2873 8033 2907
rect 8067 2904 8079 2907
rect 8202 2904 8208 2916
rect 8067 2876 8208 2904
rect 8067 2873 8079 2876
rect 8021 2867 8079 2873
rect 8202 2864 8208 2876
rect 8260 2864 8266 2916
rect 8588 2904 8616 2932
rect 9508 2904 9536 2944
rect 9585 2941 9597 2975
rect 9631 2941 9643 2975
rect 9585 2935 9643 2941
rect 9858 2932 9864 2984
rect 9916 2972 9922 2984
rect 9953 2975 10011 2981
rect 9953 2972 9965 2975
rect 9916 2944 9965 2972
rect 9916 2932 9922 2944
rect 9953 2941 9965 2944
rect 9999 2941 10011 2975
rect 9953 2935 10011 2941
rect 11054 2932 11060 2984
rect 11112 2972 11118 2984
rect 11112 2944 11836 2972
rect 11112 2932 11118 2944
rect 9876 2904 9904 2932
rect 8588 2876 9076 2904
rect 9508 2876 9904 2904
rect 5534 2836 5540 2848
rect 4356 2808 5540 2836
rect 5534 2796 5540 2808
rect 5592 2796 5598 2848
rect 7190 2796 7196 2848
rect 7248 2836 7254 2848
rect 7834 2836 7840 2848
rect 7248 2808 7840 2836
rect 7248 2796 7254 2808
rect 7834 2796 7840 2808
rect 7892 2796 7898 2848
rect 8110 2796 8116 2848
rect 8168 2836 8174 2848
rect 8168 2808 8213 2836
rect 8168 2796 8174 2808
rect 8294 2796 8300 2848
rect 8352 2836 8358 2848
rect 8941 2839 8999 2845
rect 8941 2836 8953 2839
rect 8352 2808 8953 2836
rect 8352 2796 8358 2808
rect 8941 2805 8953 2808
rect 8987 2805 8999 2839
rect 9048 2836 9076 2876
rect 10962 2864 10968 2916
rect 11020 2904 11026 2916
rect 11517 2907 11575 2913
rect 11517 2904 11529 2907
rect 11020 2876 11529 2904
rect 11020 2864 11026 2876
rect 11517 2873 11529 2876
rect 11563 2873 11575 2907
rect 11808 2904 11836 2944
rect 12084 2904 12112 3080
rect 12185 3080 12532 3108
rect 12185 2981 12213 3080
rect 12526 3068 12532 3080
rect 12584 3108 12590 3120
rect 14826 3108 14832 3120
rect 12584 3080 12940 3108
rect 12584 3068 12590 3080
rect 12342 3040 12348 3052
rect 12303 3012 12348 3040
rect 12342 3000 12348 3012
rect 12400 3000 12406 3052
rect 12161 2975 12219 2981
rect 12161 2941 12173 2975
rect 12207 2941 12219 2975
rect 12802 2972 12808 2984
rect 12161 2935 12219 2941
rect 12406 2944 12808 2972
rect 11808 2876 12112 2904
rect 11517 2867 11575 2873
rect 11238 2836 11244 2848
rect 9048 2808 11244 2836
rect 8941 2799 8999 2805
rect 11238 2796 11244 2808
rect 11296 2796 11302 2848
rect 11333 2839 11391 2845
rect 11333 2805 11345 2839
rect 11379 2836 11391 2839
rect 12406 2836 12434 2944
rect 12802 2932 12808 2944
rect 12860 2932 12866 2984
rect 12526 2836 12532 2848
rect 11379 2808 12434 2836
rect 12487 2808 12532 2836
rect 11379 2805 11391 2808
rect 11333 2799 11391 2805
rect 12526 2796 12532 2808
rect 12584 2796 12590 2848
rect 12912 2836 12940 3080
rect 14108 3080 14832 3108
rect 13906 3000 13912 3052
rect 13964 3049 13970 3052
rect 13964 3043 13987 3049
rect 13975 3009 13987 3043
rect 13964 3003 13987 3009
rect 13964 3000 13970 3003
rect 14108 2972 14136 3080
rect 14826 3068 14832 3080
rect 14884 3068 14890 3120
rect 15654 3108 15660 3120
rect 15396 3080 15660 3108
rect 14642 3040 14648 3052
rect 14603 3012 14648 3040
rect 14642 3000 14648 3012
rect 14700 3000 14706 3052
rect 15396 3049 15424 3080
rect 15654 3068 15660 3080
rect 15712 3068 15718 3120
rect 15381 3043 15439 3049
rect 15381 3009 15393 3043
rect 15427 3009 15439 3043
rect 15381 3003 15439 3009
rect 15470 3000 15476 3052
rect 15528 3040 15534 3052
rect 15565 3043 15623 3049
rect 15565 3040 15577 3043
rect 15528 3012 15577 3040
rect 15528 3000 15534 3012
rect 15565 3009 15577 3012
rect 15611 3009 15623 3043
rect 16114 3040 16120 3052
rect 16075 3012 16120 3040
rect 15565 3003 15623 3009
rect 16114 3000 16120 3012
rect 16172 3000 16178 3052
rect 16393 3043 16451 3049
rect 16393 3009 16405 3043
rect 16439 3009 16451 3043
rect 16393 3003 16451 3009
rect 14185 2975 14243 2981
rect 14185 2972 14197 2975
rect 14108 2944 14197 2972
rect 14185 2941 14197 2944
rect 14231 2941 14243 2975
rect 14185 2935 14243 2941
rect 14274 2932 14280 2984
rect 14332 2972 14338 2984
rect 14829 2975 14887 2981
rect 14829 2972 14841 2975
rect 14332 2944 14841 2972
rect 14332 2932 14338 2944
rect 14829 2941 14841 2944
rect 14875 2941 14887 2975
rect 14829 2935 14887 2941
rect 15010 2932 15016 2984
rect 15068 2972 15074 2984
rect 16408 2972 16436 3003
rect 16482 3000 16488 3052
rect 16540 3040 16546 3052
rect 16853 3043 16911 3049
rect 16853 3040 16865 3043
rect 16540 3012 16865 3040
rect 16540 3000 16546 3012
rect 16853 3009 16865 3012
rect 16899 3009 16911 3043
rect 16853 3003 16911 3009
rect 16942 3000 16948 3052
rect 17000 3040 17006 3052
rect 17000 3012 17045 3040
rect 17000 3000 17006 3012
rect 17310 3000 17316 3052
rect 17368 3040 17374 3052
rect 17512 3049 17540 3148
rect 17586 3136 17592 3188
rect 17644 3176 17650 3188
rect 17681 3179 17739 3185
rect 17681 3176 17693 3179
rect 17644 3148 17693 3176
rect 17644 3136 17650 3148
rect 17681 3145 17693 3148
rect 17727 3145 17739 3179
rect 18138 3176 18144 3188
rect 18099 3148 18144 3176
rect 17681 3139 17739 3145
rect 18138 3136 18144 3148
rect 18196 3136 18202 3188
rect 18509 3179 18567 3185
rect 18509 3145 18521 3179
rect 18555 3176 18567 3179
rect 18969 3179 19027 3185
rect 18969 3176 18981 3179
rect 18555 3148 18981 3176
rect 18555 3145 18567 3148
rect 18509 3139 18567 3145
rect 18969 3145 18981 3148
rect 19015 3145 19027 3179
rect 18969 3139 19027 3145
rect 19429 3179 19487 3185
rect 19429 3145 19441 3179
rect 19475 3176 19487 3179
rect 22186 3176 22192 3188
rect 19475 3148 19932 3176
rect 19475 3145 19487 3148
rect 19429 3139 19487 3145
rect 17954 3068 17960 3120
rect 18012 3108 18018 3120
rect 18874 3108 18880 3120
rect 18012 3080 18880 3108
rect 18012 3068 18018 3080
rect 18874 3068 18880 3080
rect 18932 3068 18938 3120
rect 19337 3111 19395 3117
rect 19337 3077 19349 3111
rect 19383 3108 19395 3111
rect 19518 3108 19524 3120
rect 19383 3080 19524 3108
rect 19383 3077 19395 3080
rect 19337 3071 19395 3077
rect 19518 3068 19524 3080
rect 19576 3068 19582 3120
rect 17405 3043 17463 3049
rect 17405 3040 17417 3043
rect 17368 3012 17417 3040
rect 17368 3000 17374 3012
rect 17405 3009 17417 3012
rect 17451 3009 17463 3043
rect 17405 3003 17463 3009
rect 17497 3043 17555 3049
rect 17497 3009 17509 3043
rect 17543 3009 17555 3043
rect 17497 3003 17555 3009
rect 17773 3043 17831 3049
rect 17773 3009 17785 3043
rect 17819 3009 17831 3043
rect 17773 3003 17831 3009
rect 15068 2944 16436 2972
rect 15068 2932 15074 2944
rect 16758 2932 16764 2984
rect 16816 2972 16822 2984
rect 17788 2972 17816 3003
rect 17862 3000 17868 3052
rect 17920 3040 17926 3052
rect 17920 3012 19564 3040
rect 17920 3000 17926 3012
rect 18598 2972 18604 2984
rect 16816 2944 17816 2972
rect 18559 2944 18604 2972
rect 16816 2932 16822 2944
rect 18598 2932 18604 2944
rect 18656 2932 18662 2984
rect 18690 2932 18696 2984
rect 18748 2972 18754 2984
rect 19536 2981 19564 3012
rect 19521 2975 19579 2981
rect 18748 2944 18793 2972
rect 18748 2932 18754 2944
rect 19521 2941 19533 2975
rect 19567 2972 19579 2975
rect 19794 2972 19800 2984
rect 19567 2944 19800 2972
rect 19567 2941 19579 2944
rect 19521 2935 19579 2941
rect 19794 2932 19800 2944
rect 19852 2932 19858 2984
rect 19904 2972 19932 3148
rect 20548 3148 22192 3176
rect 20070 3040 20076 3052
rect 20031 3012 20076 3040
rect 20070 3000 20076 3012
rect 20128 3000 20134 3052
rect 20438 3040 20444 3052
rect 20399 3012 20444 3040
rect 20438 3000 20444 3012
rect 20496 3000 20502 3052
rect 20548 3049 20576 3148
rect 22186 3136 22192 3148
rect 22244 3136 22250 3188
rect 22278 3108 22284 3120
rect 20916 3080 22284 3108
rect 20916 3049 20944 3080
rect 22278 3068 22284 3080
rect 22336 3068 22342 3120
rect 20533 3043 20591 3049
rect 20533 3009 20545 3043
rect 20579 3009 20591 3043
rect 20533 3003 20591 3009
rect 20901 3043 20959 3049
rect 20901 3009 20913 3043
rect 20947 3009 20959 3043
rect 20901 3003 20959 3009
rect 21269 3043 21327 3049
rect 21269 3009 21281 3043
rect 21315 3040 21327 3043
rect 22370 3040 22376 3052
rect 21315 3012 22376 3040
rect 21315 3009 21327 3012
rect 21269 3003 21327 3009
rect 22370 3000 22376 3012
rect 22428 3000 22434 3052
rect 21174 2972 21180 2984
rect 19904 2944 21180 2972
rect 21174 2932 21180 2944
rect 21232 2932 21238 2984
rect 15378 2904 15384 2916
rect 14200 2876 15384 2904
rect 14200 2836 14228 2876
rect 15378 2864 15384 2876
rect 15436 2864 15442 2916
rect 15654 2864 15660 2916
rect 15712 2904 15718 2916
rect 17129 2907 17187 2913
rect 15712 2876 16252 2904
rect 15712 2864 15718 2876
rect 12912 2808 14228 2836
rect 14366 2796 14372 2848
rect 14424 2836 14430 2848
rect 15197 2839 15255 2845
rect 15197 2836 15209 2839
rect 14424 2808 15209 2836
rect 14424 2796 14430 2808
rect 15197 2805 15209 2808
rect 15243 2805 15255 2839
rect 15197 2799 15255 2805
rect 15470 2796 15476 2848
rect 15528 2836 15534 2848
rect 15749 2839 15807 2845
rect 15749 2836 15761 2839
rect 15528 2808 15761 2836
rect 15528 2796 15534 2808
rect 15749 2805 15761 2808
rect 15795 2805 15807 2839
rect 15930 2836 15936 2848
rect 15891 2808 15936 2836
rect 15749 2799 15807 2805
rect 15930 2796 15936 2808
rect 15988 2796 15994 2848
rect 16224 2845 16252 2876
rect 17129 2873 17141 2907
rect 17175 2904 17187 2907
rect 17175 2876 19012 2904
rect 17175 2873 17187 2876
rect 17129 2867 17187 2873
rect 18984 2848 19012 2876
rect 19610 2864 19616 2916
rect 19668 2904 19674 2916
rect 20257 2907 20315 2913
rect 20257 2904 20269 2907
rect 19668 2876 20269 2904
rect 19668 2864 19674 2876
rect 20257 2873 20269 2876
rect 20303 2873 20315 2907
rect 20257 2867 20315 2873
rect 20622 2864 20628 2916
rect 20680 2904 20686 2916
rect 21085 2907 21143 2913
rect 21085 2904 21097 2907
rect 20680 2876 21097 2904
rect 20680 2864 20686 2876
rect 21085 2873 21097 2876
rect 21131 2873 21143 2907
rect 21085 2867 21143 2873
rect 16209 2839 16267 2845
rect 16209 2805 16221 2839
rect 16255 2805 16267 2839
rect 16666 2836 16672 2848
rect 16627 2808 16672 2836
rect 16209 2799 16267 2805
rect 16666 2796 16672 2808
rect 16724 2796 16730 2848
rect 17218 2796 17224 2848
rect 17276 2836 17282 2848
rect 17957 2839 18015 2845
rect 17276 2808 17321 2836
rect 17276 2796 17282 2808
rect 17957 2805 17969 2839
rect 18003 2836 18015 2839
rect 18046 2836 18052 2848
rect 18003 2808 18052 2836
rect 18003 2805 18015 2808
rect 17957 2799 18015 2805
rect 18046 2796 18052 2808
rect 18104 2796 18110 2848
rect 18690 2796 18696 2848
rect 18748 2836 18754 2848
rect 18874 2836 18880 2848
rect 18748 2808 18880 2836
rect 18748 2796 18754 2808
rect 18874 2796 18880 2808
rect 18932 2796 18938 2848
rect 18966 2796 18972 2848
rect 19024 2796 19030 2848
rect 19058 2796 19064 2848
rect 19116 2836 19122 2848
rect 19889 2839 19947 2845
rect 19889 2836 19901 2839
rect 19116 2808 19901 2836
rect 19116 2796 19122 2808
rect 19889 2805 19901 2808
rect 19935 2805 19947 2839
rect 19889 2799 19947 2805
rect 20346 2796 20352 2848
rect 20404 2836 20410 2848
rect 20717 2839 20775 2845
rect 20717 2836 20729 2839
rect 20404 2808 20729 2836
rect 20404 2796 20410 2808
rect 20717 2805 20729 2808
rect 20763 2805 20775 2839
rect 20717 2799 20775 2805
rect 21358 2796 21364 2848
rect 21416 2836 21422 2848
rect 21453 2839 21511 2845
rect 21453 2836 21465 2839
rect 21416 2808 21465 2836
rect 21416 2796 21422 2808
rect 21453 2805 21465 2808
rect 21499 2805 21511 2839
rect 21453 2799 21511 2805
rect 1104 2746 21896 2768
rect 1104 2694 3549 2746
rect 3601 2694 3613 2746
rect 3665 2694 3677 2746
rect 3729 2694 3741 2746
rect 3793 2694 3805 2746
rect 3857 2694 8747 2746
rect 8799 2694 8811 2746
rect 8863 2694 8875 2746
rect 8927 2694 8939 2746
rect 8991 2694 9003 2746
rect 9055 2694 13945 2746
rect 13997 2694 14009 2746
rect 14061 2694 14073 2746
rect 14125 2694 14137 2746
rect 14189 2694 14201 2746
rect 14253 2694 19143 2746
rect 19195 2694 19207 2746
rect 19259 2694 19271 2746
rect 19323 2694 19335 2746
rect 19387 2694 19399 2746
rect 19451 2694 21896 2746
rect 1104 2672 21896 2694
rect 2774 2592 2780 2644
rect 2832 2632 2838 2644
rect 4246 2632 4252 2644
rect 2832 2604 4252 2632
rect 2832 2592 2838 2604
rect 4246 2592 4252 2604
rect 4304 2592 4310 2644
rect 5626 2632 5632 2644
rect 5587 2604 5632 2632
rect 5626 2592 5632 2604
rect 5684 2592 5690 2644
rect 5813 2635 5871 2641
rect 5813 2601 5825 2635
rect 5859 2632 5871 2635
rect 6822 2632 6828 2644
rect 5859 2604 6828 2632
rect 5859 2601 5871 2604
rect 5813 2595 5871 2601
rect 6822 2592 6828 2604
rect 6880 2592 6886 2644
rect 7466 2632 7472 2644
rect 7427 2604 7472 2632
rect 7466 2592 7472 2604
rect 7524 2592 7530 2644
rect 7650 2632 7656 2644
rect 7611 2604 7656 2632
rect 7650 2592 7656 2604
rect 7708 2592 7714 2644
rect 8018 2592 8024 2644
rect 8076 2632 8082 2644
rect 8076 2604 8432 2632
rect 8076 2592 8082 2604
rect 3234 2564 3240 2576
rect 1964 2536 3240 2564
rect 1964 2505 1992 2536
rect 3234 2524 3240 2536
rect 3292 2524 3298 2576
rect 3602 2564 3608 2576
rect 3563 2536 3608 2564
rect 3602 2524 3608 2536
rect 3660 2524 3666 2576
rect 3694 2524 3700 2576
rect 3752 2564 3758 2576
rect 3970 2564 3976 2576
rect 3752 2536 3976 2564
rect 3752 2524 3758 2536
rect 3970 2524 3976 2536
rect 4028 2524 4034 2576
rect 4154 2564 4160 2576
rect 4115 2536 4160 2564
rect 4154 2524 4160 2536
rect 4212 2524 4218 2576
rect 5534 2524 5540 2576
rect 5592 2564 5598 2576
rect 5902 2564 5908 2576
rect 5592 2536 5908 2564
rect 5592 2524 5598 2536
rect 5902 2524 5908 2536
rect 5960 2524 5966 2576
rect 8294 2564 8300 2576
rect 7300 2536 8300 2564
rect 1949 2499 2007 2505
rect 1949 2465 1961 2499
rect 1995 2465 2007 2499
rect 1949 2459 2007 2465
rect 2038 2456 2044 2508
rect 2096 2496 2102 2508
rect 2096 2468 4108 2496
rect 2096 2456 2102 2468
rect 2225 2431 2283 2437
rect 2225 2397 2237 2431
rect 2271 2428 2283 2431
rect 2774 2428 2780 2440
rect 2271 2400 2780 2428
rect 2271 2397 2283 2400
rect 2225 2391 2283 2397
rect 2774 2388 2780 2400
rect 2832 2388 2838 2440
rect 3145 2431 3203 2437
rect 3145 2397 3157 2431
rect 3191 2397 3203 2431
rect 3145 2391 3203 2397
rect 2682 2320 2688 2372
rect 2740 2360 2746 2372
rect 3160 2360 3188 2391
rect 2740 2332 3188 2360
rect 3421 2363 3479 2369
rect 2740 2320 2746 2332
rect 3421 2329 3433 2363
rect 3467 2360 3479 2363
rect 3602 2360 3608 2372
rect 3467 2332 3608 2360
rect 3467 2329 3479 2332
rect 3421 2323 3479 2329
rect 3602 2320 3608 2332
rect 3660 2320 3666 2372
rect 3970 2360 3976 2372
rect 3931 2332 3976 2360
rect 3970 2320 3976 2332
rect 4028 2320 4034 2372
rect 4080 2360 4108 2468
rect 5258 2456 5264 2508
rect 5316 2496 5322 2508
rect 6917 2499 6975 2505
rect 5316 2468 6132 2496
rect 5316 2456 5322 2468
rect 4249 2431 4307 2437
rect 4249 2397 4261 2431
rect 4295 2428 4307 2431
rect 4890 2428 4896 2440
rect 4295 2400 4896 2428
rect 4295 2397 4307 2400
rect 4249 2391 4307 2397
rect 4890 2388 4896 2400
rect 4948 2388 4954 2440
rect 5994 2388 6000 2440
rect 6052 2388 6058 2440
rect 6104 2428 6132 2468
rect 6917 2465 6929 2499
rect 6963 2496 6975 2499
rect 7098 2496 7104 2508
rect 6963 2468 7104 2496
rect 6963 2465 6975 2468
rect 6917 2459 6975 2465
rect 7098 2456 7104 2468
rect 7156 2456 7162 2508
rect 7300 2437 7328 2536
rect 8294 2524 8300 2536
rect 8352 2524 8358 2576
rect 7374 2456 7380 2508
rect 7432 2496 7438 2508
rect 8021 2499 8079 2505
rect 8021 2496 8033 2499
rect 7432 2468 8033 2496
rect 7432 2456 7438 2468
rect 8021 2465 8033 2468
rect 8067 2465 8079 2499
rect 8202 2496 8208 2508
rect 8163 2468 8208 2496
rect 8021 2459 8079 2465
rect 8202 2456 8208 2468
rect 8260 2456 8266 2508
rect 8404 2496 8432 2604
rect 9858 2592 9864 2644
rect 9916 2632 9922 2644
rect 10870 2632 10876 2644
rect 9916 2604 10876 2632
rect 9916 2592 9922 2604
rect 10870 2592 10876 2604
rect 10928 2592 10934 2644
rect 11146 2592 11152 2644
rect 11204 2632 11210 2644
rect 11701 2635 11759 2641
rect 11701 2632 11713 2635
rect 11204 2604 11713 2632
rect 11204 2592 11210 2604
rect 11701 2601 11713 2604
rect 11747 2601 11759 2635
rect 11701 2595 11759 2601
rect 14642 2592 14648 2644
rect 14700 2632 14706 2644
rect 14829 2635 14887 2641
rect 14829 2632 14841 2635
rect 14700 2604 14841 2632
rect 14700 2592 14706 2604
rect 14829 2601 14841 2604
rect 14875 2601 14887 2635
rect 14829 2595 14887 2601
rect 15838 2592 15844 2644
rect 15896 2632 15902 2644
rect 16761 2635 16819 2641
rect 16761 2632 16773 2635
rect 15896 2604 16773 2632
rect 15896 2592 15902 2604
rect 16761 2601 16773 2604
rect 16807 2601 16819 2635
rect 16761 2595 16819 2601
rect 17678 2592 17684 2644
rect 17736 2632 17742 2644
rect 18693 2635 18751 2641
rect 18693 2632 18705 2635
rect 17736 2604 18705 2632
rect 17736 2592 17742 2604
rect 18693 2601 18705 2604
rect 18739 2601 18751 2635
rect 18693 2595 18751 2601
rect 20070 2592 20076 2644
rect 20128 2632 20134 2644
rect 20441 2635 20499 2641
rect 20441 2632 20453 2635
rect 20128 2604 20453 2632
rect 20128 2592 20134 2604
rect 20441 2601 20453 2604
rect 20487 2601 20499 2635
rect 20441 2595 20499 2601
rect 8662 2564 8668 2576
rect 8623 2536 8668 2564
rect 8662 2524 8668 2536
rect 8720 2524 8726 2576
rect 9766 2524 9772 2576
rect 9824 2564 9830 2576
rect 12342 2564 12348 2576
rect 9824 2536 9996 2564
rect 12303 2536 12348 2564
rect 9824 2524 9830 2536
rect 9493 2499 9551 2505
rect 9493 2496 9505 2499
rect 8404 2468 9505 2496
rect 9493 2465 9505 2468
rect 9539 2465 9551 2499
rect 9493 2459 9551 2465
rect 9861 2499 9919 2505
rect 9861 2465 9873 2499
rect 9907 2465 9919 2499
rect 9968 2496 9996 2536
rect 12342 2524 12348 2536
rect 12400 2524 12406 2576
rect 13630 2524 13636 2576
rect 13688 2564 13694 2576
rect 15013 2567 15071 2573
rect 15013 2564 15025 2567
rect 13688 2536 15025 2564
rect 13688 2524 13694 2536
rect 15013 2533 15025 2536
rect 15059 2533 15071 2567
rect 15013 2527 15071 2533
rect 15102 2524 15108 2576
rect 15160 2564 15166 2576
rect 16117 2567 16175 2573
rect 16117 2564 16129 2567
rect 15160 2536 16129 2564
rect 15160 2524 15166 2536
rect 16117 2533 16129 2536
rect 16163 2533 16175 2567
rect 16117 2527 16175 2533
rect 16206 2524 16212 2576
rect 16264 2564 16270 2576
rect 17129 2567 17187 2573
rect 17129 2564 17141 2567
rect 16264 2536 17141 2564
rect 16264 2524 16270 2536
rect 17129 2533 17141 2536
rect 17175 2533 17187 2567
rect 17129 2527 17187 2533
rect 17310 2524 17316 2576
rect 17368 2564 17374 2576
rect 18233 2567 18291 2573
rect 18233 2564 18245 2567
rect 17368 2536 18245 2564
rect 17368 2524 17374 2536
rect 18233 2533 18245 2536
rect 18279 2533 18291 2567
rect 18233 2527 18291 2533
rect 18414 2524 18420 2576
rect 18472 2524 18478 2576
rect 18598 2524 18604 2576
rect 18656 2564 18662 2576
rect 19245 2567 19303 2573
rect 19245 2564 19257 2567
rect 18656 2536 19257 2564
rect 18656 2524 18662 2536
rect 19245 2533 19257 2536
rect 19291 2533 19303 2567
rect 20257 2567 20315 2573
rect 20257 2564 20269 2567
rect 19245 2527 19303 2533
rect 19352 2536 20269 2564
rect 11149 2499 11207 2505
rect 11149 2496 11161 2499
rect 9968 2468 11161 2496
rect 9861 2459 9919 2465
rect 11149 2465 11161 2468
rect 11195 2465 11207 2499
rect 11149 2459 11207 2465
rect 7193 2431 7251 2437
rect 7193 2428 7205 2431
rect 6104 2400 7205 2428
rect 7193 2397 7205 2400
rect 7239 2397 7251 2431
rect 7193 2391 7251 2397
rect 7285 2431 7343 2437
rect 7285 2397 7297 2431
rect 7331 2397 7343 2431
rect 7285 2391 7343 2397
rect 7392 2400 7880 2428
rect 4494 2363 4552 2369
rect 4494 2360 4506 2363
rect 4080 2332 4506 2360
rect 4494 2329 4506 2332
rect 4540 2329 4552 2363
rect 4494 2323 4552 2329
rect 4614 2320 4620 2372
rect 4672 2360 4678 2372
rect 5905 2363 5963 2369
rect 5905 2360 5917 2363
rect 4672 2332 5917 2360
rect 4672 2320 4678 2332
rect 5905 2329 5917 2332
rect 5951 2329 5963 2363
rect 5905 2323 5963 2329
rect 2915 2295 2973 2301
rect 2915 2261 2927 2295
rect 2961 2292 2973 2295
rect 5810 2292 5816 2304
rect 2961 2264 5816 2292
rect 2961 2261 2973 2264
rect 2915 2255 2973 2261
rect 5810 2252 5816 2264
rect 5868 2252 5874 2304
rect 6012 2292 6040 2388
rect 6089 2363 6147 2369
rect 6089 2329 6101 2363
rect 6135 2360 6147 2363
rect 6638 2360 6644 2372
rect 6135 2332 6644 2360
rect 6135 2329 6147 2332
rect 6089 2323 6147 2329
rect 6638 2320 6644 2332
rect 6696 2320 6702 2372
rect 6730 2320 6736 2372
rect 6788 2360 6794 2372
rect 7392 2360 7420 2400
rect 6788 2332 7420 2360
rect 6788 2320 6794 2332
rect 7650 2320 7656 2372
rect 7708 2360 7714 2372
rect 7745 2363 7803 2369
rect 7745 2360 7757 2363
rect 7708 2332 7757 2360
rect 7708 2320 7714 2332
rect 7745 2329 7757 2332
rect 7791 2329 7803 2363
rect 7852 2360 7880 2400
rect 8110 2388 8116 2440
rect 8168 2428 8174 2440
rect 8297 2431 8355 2437
rect 8297 2428 8309 2431
rect 8168 2400 8309 2428
rect 8168 2388 8174 2400
rect 8297 2397 8309 2400
rect 8343 2397 8355 2431
rect 8297 2391 8355 2397
rect 8386 2388 8392 2440
rect 8444 2428 8450 2440
rect 8662 2428 8668 2440
rect 8444 2400 8668 2428
rect 8444 2388 8450 2400
rect 8662 2388 8668 2400
rect 8720 2388 8726 2440
rect 9398 2428 9404 2440
rect 9359 2400 9404 2428
rect 9398 2388 9404 2400
rect 9456 2388 9462 2440
rect 9876 2360 9904 2459
rect 12066 2456 12072 2508
rect 12124 2496 12130 2508
rect 12124 2468 13032 2496
rect 12124 2456 12130 2468
rect 9950 2388 9956 2440
rect 10008 2428 10014 2440
rect 10965 2431 11023 2437
rect 10965 2428 10977 2431
rect 10008 2400 10977 2428
rect 10008 2388 10014 2400
rect 10965 2397 10977 2400
rect 11011 2397 11023 2431
rect 10965 2391 11023 2397
rect 11609 2431 11667 2437
rect 11609 2397 11621 2431
rect 11655 2428 11667 2431
rect 11698 2428 11704 2440
rect 11655 2400 11704 2428
rect 11655 2397 11667 2400
rect 11609 2391 11667 2397
rect 11698 2388 11704 2400
rect 11756 2388 11762 2440
rect 11882 2428 11888 2440
rect 11843 2400 11888 2428
rect 11882 2388 11888 2400
rect 11940 2388 11946 2440
rect 12342 2388 12348 2440
rect 12400 2428 12406 2440
rect 13004 2437 13032 2468
rect 13170 2456 13176 2508
rect 13228 2496 13234 2508
rect 14185 2499 14243 2505
rect 14185 2496 14197 2499
rect 13228 2468 14197 2496
rect 13228 2456 13234 2468
rect 14185 2465 14197 2468
rect 14231 2465 14243 2499
rect 15930 2496 15936 2508
rect 14185 2459 14243 2465
rect 15212 2468 15936 2496
rect 12529 2431 12587 2437
rect 12529 2428 12541 2431
rect 12400 2400 12541 2428
rect 12400 2388 12406 2400
rect 12529 2397 12541 2400
rect 12575 2397 12587 2431
rect 12529 2391 12587 2397
rect 12897 2431 12955 2437
rect 12897 2397 12909 2431
rect 12943 2397 12955 2431
rect 12897 2391 12955 2397
rect 12989 2431 13047 2437
rect 12989 2397 13001 2431
rect 13035 2397 13047 2431
rect 13354 2428 13360 2440
rect 13315 2400 13360 2428
rect 12989 2391 13047 2397
rect 10137 2363 10195 2369
rect 10137 2360 10149 2363
rect 7852 2332 9904 2360
rect 9968 2332 10149 2360
rect 7745 2323 7803 2329
rect 8941 2295 8999 2301
rect 8941 2292 8953 2295
rect 6012 2264 8953 2292
rect 8941 2261 8953 2264
rect 8987 2261 8999 2295
rect 9306 2292 9312 2304
rect 9267 2264 9312 2292
rect 8941 2255 8999 2261
rect 9306 2252 9312 2264
rect 9364 2252 9370 2304
rect 9490 2252 9496 2304
rect 9548 2292 9554 2304
rect 9968 2292 9996 2332
rect 10137 2329 10149 2332
rect 10183 2329 10195 2363
rect 11057 2363 11115 2369
rect 11057 2360 11069 2363
rect 10137 2323 10195 2329
rect 10520 2332 11069 2360
rect 9548 2264 9996 2292
rect 10045 2295 10103 2301
rect 9548 2252 9554 2264
rect 10045 2261 10057 2295
rect 10091 2292 10103 2295
rect 10226 2292 10232 2304
rect 10091 2264 10232 2292
rect 10091 2261 10103 2264
rect 10045 2255 10103 2261
rect 10226 2252 10232 2264
rect 10284 2252 10290 2304
rect 10520 2301 10548 2332
rect 11057 2329 11069 2332
rect 11103 2329 11115 2363
rect 12912 2360 12940 2391
rect 13354 2388 13360 2400
rect 13412 2388 13418 2440
rect 13722 2388 13728 2440
rect 13780 2428 13786 2440
rect 13909 2431 13967 2437
rect 13909 2428 13921 2431
rect 13780 2400 13921 2428
rect 13780 2388 13786 2400
rect 13909 2397 13921 2400
rect 13955 2397 13967 2431
rect 13909 2391 13967 2397
rect 14461 2431 14519 2437
rect 14461 2397 14473 2431
rect 14507 2428 14519 2431
rect 15010 2428 15016 2440
rect 14507 2400 15016 2428
rect 14507 2397 14519 2400
rect 14461 2391 14519 2397
rect 15010 2388 15016 2400
rect 15068 2388 15074 2440
rect 15212 2437 15240 2468
rect 15930 2456 15936 2468
rect 15988 2456 15994 2508
rect 18138 2496 18144 2508
rect 17328 2468 18144 2496
rect 15197 2431 15255 2437
rect 15197 2397 15209 2431
rect 15243 2397 15255 2431
rect 15197 2391 15255 2397
rect 15286 2388 15292 2440
rect 15344 2428 15350 2440
rect 15654 2428 15660 2440
rect 15344 2400 15389 2428
rect 15615 2400 15660 2428
rect 15344 2388 15350 2400
rect 15654 2388 15660 2400
rect 15712 2388 15718 2440
rect 16301 2431 16359 2437
rect 16301 2397 16313 2431
rect 16347 2428 16359 2431
rect 16666 2428 16672 2440
rect 16347 2400 16672 2428
rect 16347 2397 16359 2400
rect 16301 2391 16359 2397
rect 16666 2388 16672 2400
rect 16724 2388 16730 2440
rect 16945 2431 17003 2437
rect 16945 2397 16957 2431
rect 16991 2428 17003 2431
rect 17218 2428 17224 2440
rect 16991 2400 17224 2428
rect 16991 2397 17003 2400
rect 16945 2391 17003 2397
rect 17218 2388 17224 2400
rect 17276 2388 17282 2440
rect 17328 2437 17356 2468
rect 18138 2456 18144 2468
rect 18196 2456 18202 2508
rect 18432 2496 18460 2524
rect 19352 2496 19380 2536
rect 20257 2533 20269 2536
rect 20303 2533 20315 2567
rect 20257 2527 20315 2533
rect 19794 2496 19800 2508
rect 18432 2468 19380 2496
rect 19755 2468 19800 2496
rect 19794 2456 19800 2468
rect 19852 2456 19858 2508
rect 20993 2499 21051 2505
rect 20993 2465 21005 2499
rect 21039 2496 21051 2499
rect 22922 2496 22928 2508
rect 21039 2468 22928 2496
rect 21039 2465 21051 2468
rect 20993 2459 21051 2465
rect 22922 2456 22928 2468
rect 22980 2456 22986 2508
rect 17313 2431 17371 2437
rect 17313 2397 17325 2431
rect 17359 2397 17371 2431
rect 17313 2391 17371 2397
rect 17681 2431 17739 2437
rect 17681 2397 17693 2431
rect 17727 2428 17739 2431
rect 17954 2428 17960 2440
rect 17727 2400 17960 2428
rect 17727 2397 17739 2400
rect 17681 2391 17739 2397
rect 17954 2388 17960 2400
rect 18012 2388 18018 2440
rect 18049 2431 18107 2437
rect 18049 2397 18061 2431
rect 18095 2397 18107 2431
rect 18049 2391 18107 2397
rect 12912 2332 13768 2360
rect 11057 2323 11115 2329
rect 10505 2295 10563 2301
rect 10505 2261 10517 2295
rect 10551 2261 10563 2295
rect 10505 2255 10563 2261
rect 10594 2252 10600 2304
rect 10652 2292 10658 2304
rect 12066 2292 12072 2304
rect 10652 2264 10697 2292
rect 12027 2264 12072 2292
rect 10652 2252 10658 2264
rect 12066 2252 12072 2264
rect 12124 2252 12130 2304
rect 12526 2252 12532 2304
rect 12584 2292 12590 2304
rect 12713 2295 12771 2301
rect 12713 2292 12725 2295
rect 12584 2264 12725 2292
rect 12584 2252 12590 2264
rect 12713 2261 12725 2264
rect 12759 2261 12771 2295
rect 12713 2255 12771 2261
rect 12894 2252 12900 2304
rect 12952 2292 12958 2304
rect 13173 2295 13231 2301
rect 13173 2292 13185 2295
rect 12952 2264 13185 2292
rect 12952 2252 12958 2264
rect 13173 2261 13185 2264
rect 13219 2261 13231 2295
rect 13173 2255 13231 2261
rect 13262 2252 13268 2304
rect 13320 2292 13326 2304
rect 13740 2301 13768 2332
rect 13998 2320 14004 2372
rect 14056 2360 14062 2372
rect 14056 2332 14688 2360
rect 14056 2320 14062 2332
rect 13541 2295 13599 2301
rect 13541 2292 13553 2295
rect 13320 2264 13553 2292
rect 13320 2252 13326 2264
rect 13541 2261 13553 2264
rect 13587 2261 13599 2295
rect 13541 2255 13599 2261
rect 13725 2295 13783 2301
rect 13725 2261 13737 2295
rect 13771 2261 13783 2295
rect 13725 2255 13783 2261
rect 13814 2252 13820 2304
rect 13872 2292 13878 2304
rect 14369 2295 14427 2301
rect 14369 2292 14381 2295
rect 13872 2264 14381 2292
rect 13872 2252 13878 2264
rect 14369 2261 14381 2264
rect 14415 2292 14427 2295
rect 14458 2292 14464 2304
rect 14415 2264 14464 2292
rect 14415 2261 14427 2264
rect 14369 2255 14427 2261
rect 14458 2252 14464 2264
rect 14516 2252 14522 2304
rect 14660 2292 14688 2332
rect 14734 2320 14740 2372
rect 14792 2360 14798 2372
rect 14792 2332 15884 2360
rect 14792 2320 14798 2332
rect 15856 2301 15884 2332
rect 17034 2320 17040 2372
rect 17092 2360 17098 2372
rect 18064 2360 18092 2391
rect 18322 2388 18328 2440
rect 18380 2428 18386 2440
rect 18417 2431 18475 2437
rect 18417 2428 18429 2431
rect 18380 2400 18429 2428
rect 18380 2388 18386 2400
rect 18417 2397 18429 2400
rect 18463 2397 18475 2431
rect 18417 2391 18475 2397
rect 18506 2388 18512 2440
rect 18564 2428 18570 2440
rect 18564 2400 18609 2428
rect 18564 2388 18570 2400
rect 18966 2388 18972 2440
rect 19024 2428 19030 2440
rect 19061 2431 19119 2437
rect 19061 2428 19073 2431
rect 19024 2400 19073 2428
rect 19024 2388 19030 2400
rect 19061 2397 19073 2400
rect 19107 2397 19119 2431
rect 19061 2391 19119 2397
rect 19702 2388 19708 2440
rect 19760 2428 19766 2440
rect 20073 2431 20131 2437
rect 20073 2428 20085 2431
rect 19760 2400 20085 2428
rect 19760 2388 19766 2400
rect 20073 2397 20085 2400
rect 20119 2397 20131 2431
rect 20073 2391 20131 2397
rect 20530 2388 20536 2440
rect 20588 2428 20594 2440
rect 20625 2431 20683 2437
rect 20625 2428 20637 2431
rect 20588 2400 20637 2428
rect 20588 2388 20594 2400
rect 20625 2397 20637 2400
rect 20671 2397 20683 2431
rect 20625 2391 20683 2397
rect 20714 2388 20720 2440
rect 20772 2428 20778 2440
rect 21542 2428 21548 2440
rect 20772 2400 21548 2428
rect 20772 2388 20778 2400
rect 21542 2388 21548 2400
rect 21600 2388 21606 2440
rect 19613 2363 19671 2369
rect 17092 2332 17908 2360
rect 18064 2332 18920 2360
rect 17092 2320 17098 2332
rect 15473 2295 15531 2301
rect 15473 2292 15485 2295
rect 14660 2264 15485 2292
rect 15473 2261 15485 2264
rect 15519 2261 15531 2295
rect 15473 2255 15531 2261
rect 15841 2295 15899 2301
rect 15841 2261 15853 2295
rect 15887 2261 15899 2295
rect 16390 2292 16396 2304
rect 16351 2264 16396 2292
rect 15841 2255 15899 2261
rect 16390 2252 16396 2264
rect 16448 2252 16454 2304
rect 16942 2252 16948 2304
rect 17000 2292 17006 2304
rect 17880 2301 17908 2332
rect 18892 2301 18920 2332
rect 19613 2329 19625 2363
rect 19659 2360 19671 2363
rect 20162 2360 20168 2372
rect 19659 2332 20168 2360
rect 19659 2329 19671 2332
rect 19613 2323 19671 2329
rect 20162 2320 20168 2332
rect 20220 2320 20226 2372
rect 17497 2295 17555 2301
rect 17497 2292 17509 2295
rect 17000 2264 17509 2292
rect 17000 2252 17006 2264
rect 17497 2261 17509 2264
rect 17543 2261 17555 2295
rect 17497 2255 17555 2261
rect 17865 2295 17923 2301
rect 17865 2261 17877 2295
rect 17911 2261 17923 2295
rect 17865 2255 17923 2261
rect 18877 2295 18935 2301
rect 18877 2261 18889 2295
rect 18923 2261 18935 2295
rect 18877 2255 18935 2261
rect 19705 2295 19763 2301
rect 19705 2261 19717 2295
rect 19751 2292 19763 2295
rect 21266 2292 21272 2304
rect 19751 2264 21272 2292
rect 19751 2261 19763 2264
rect 19705 2255 19763 2261
rect 21266 2252 21272 2264
rect 21324 2252 21330 2304
rect 1104 2202 22056 2224
rect 1104 2150 6148 2202
rect 6200 2150 6212 2202
rect 6264 2150 6276 2202
rect 6328 2150 6340 2202
rect 6392 2150 6404 2202
rect 6456 2150 11346 2202
rect 11398 2150 11410 2202
rect 11462 2150 11474 2202
rect 11526 2150 11538 2202
rect 11590 2150 11602 2202
rect 11654 2150 16544 2202
rect 16596 2150 16608 2202
rect 16660 2150 16672 2202
rect 16724 2150 16736 2202
rect 16788 2150 16800 2202
rect 16852 2150 21742 2202
rect 21794 2150 21806 2202
rect 21858 2150 21870 2202
rect 21922 2150 21934 2202
rect 21986 2150 21998 2202
rect 22050 2150 22056 2202
rect 1104 2128 22056 2150
rect 3970 2048 3976 2100
rect 4028 2088 4034 2100
rect 4028 2060 5488 2088
rect 4028 2048 4034 2060
rect 1302 1980 1308 2032
rect 1360 2020 1366 2032
rect 5258 2020 5264 2032
rect 1360 1992 5264 2020
rect 1360 1980 1366 1992
rect 5258 1980 5264 1992
rect 5316 1980 5322 2032
rect 5460 2020 5488 2060
rect 5534 2048 5540 2100
rect 5592 2088 5598 2100
rect 10226 2088 10232 2100
rect 5592 2060 10232 2088
rect 5592 2048 5598 2060
rect 10226 2048 10232 2060
rect 10284 2048 10290 2100
rect 11054 2048 11060 2100
rect 11112 2088 11118 2100
rect 12342 2088 12348 2100
rect 11112 2060 12348 2088
rect 11112 2048 11118 2060
rect 12342 2048 12348 2060
rect 12400 2088 12406 2100
rect 16390 2088 16396 2100
rect 12400 2060 16396 2088
rect 12400 2048 12406 2060
rect 16390 2048 16396 2060
rect 16448 2048 16454 2100
rect 18322 2048 18328 2100
rect 18380 2088 18386 2100
rect 19886 2088 19892 2100
rect 18380 2060 19892 2088
rect 18380 2048 18386 2060
rect 19886 2048 19892 2060
rect 19944 2048 19950 2100
rect 7374 2020 7380 2032
rect 5460 1992 7380 2020
rect 7374 1980 7380 1992
rect 7432 1980 7438 2032
rect 7466 1980 7472 2032
rect 7524 2020 7530 2032
rect 12250 2020 12256 2032
rect 7524 1992 12256 2020
rect 7524 1980 7530 1992
rect 12250 1980 12256 1992
rect 12308 1980 12314 2032
rect 12618 1980 12624 2032
rect 12676 2020 12682 2032
rect 15654 2020 15660 2032
rect 12676 1992 15660 2020
rect 12676 1980 12682 1992
rect 15654 1980 15660 1992
rect 15712 1980 15718 2032
rect 17494 1980 17500 2032
rect 17552 2020 17558 2032
rect 19794 2020 19800 2032
rect 17552 1992 19800 2020
rect 17552 1980 17558 1992
rect 19794 1980 19800 1992
rect 19852 1980 19858 2032
rect 1854 1912 1860 1964
rect 1912 1952 1918 1964
rect 5442 1952 5448 1964
rect 1912 1924 5448 1952
rect 1912 1912 1918 1924
rect 5442 1912 5448 1924
rect 5500 1912 5506 1964
rect 5810 1912 5816 1964
rect 5868 1952 5874 1964
rect 8570 1952 8576 1964
rect 5868 1924 8576 1952
rect 5868 1912 5874 1924
rect 8570 1912 8576 1924
rect 8628 1912 8634 1964
rect 14550 1912 14556 1964
rect 14608 1952 14614 1964
rect 19242 1952 19248 1964
rect 14608 1924 19248 1952
rect 14608 1912 14614 1924
rect 19242 1912 19248 1924
rect 19300 1912 19306 1964
rect 6638 1844 6644 1896
rect 6696 1884 6702 1896
rect 8846 1884 8852 1896
rect 6696 1856 8852 1884
rect 6696 1844 6702 1856
rect 8846 1844 8852 1856
rect 8904 1884 8910 1896
rect 10778 1884 10784 1896
rect 8904 1856 10784 1884
rect 8904 1844 8910 1856
rect 10778 1844 10784 1856
rect 10836 1844 10842 1896
rect 14918 1844 14924 1896
rect 14976 1884 14982 1896
rect 19150 1884 19156 1896
rect 14976 1856 19156 1884
rect 14976 1844 14982 1856
rect 19150 1844 19156 1856
rect 19208 1844 19214 1896
rect 3786 1776 3792 1828
rect 3844 1816 3850 1828
rect 7558 1816 7564 1828
rect 3844 1788 7564 1816
rect 3844 1776 3850 1788
rect 7558 1776 7564 1788
rect 7616 1776 7622 1828
rect 14458 1776 14464 1828
rect 14516 1816 14522 1828
rect 19978 1816 19984 1828
rect 14516 1788 19984 1816
rect 14516 1776 14522 1788
rect 19978 1776 19984 1788
rect 20036 1776 20042 1828
rect 3602 1708 3608 1760
rect 3660 1748 3666 1760
rect 6730 1748 6736 1760
rect 3660 1720 6736 1748
rect 3660 1708 3666 1720
rect 6730 1708 6736 1720
rect 6788 1708 6794 1760
rect 1486 1640 1492 1692
rect 1544 1680 1550 1692
rect 9674 1680 9680 1692
rect 1544 1652 9680 1680
rect 1544 1640 1550 1652
rect 9674 1640 9680 1652
rect 9732 1640 9738 1692
rect 8110 1300 8116 1352
rect 8168 1340 8174 1352
rect 10594 1340 10600 1352
rect 8168 1312 10600 1340
rect 8168 1300 8174 1312
rect 10594 1300 10600 1312
rect 10652 1300 10658 1352
rect 17126 1340 17132 1352
rect 10796 1312 17132 1340
rect 5074 1164 5080 1216
rect 5132 1204 5138 1216
rect 10796 1204 10824 1312
rect 17126 1300 17132 1312
rect 17184 1300 17190 1352
rect 16114 1272 16120 1284
rect 5132 1176 10824 1204
rect 12406 1244 16120 1272
rect 5132 1164 5138 1176
rect 5718 1096 5724 1148
rect 5776 1136 5782 1148
rect 12406 1136 12434 1244
rect 16114 1232 16120 1244
rect 16172 1232 16178 1284
rect 5776 1108 12434 1136
rect 5776 1096 5782 1108
rect 7466 76 7472 128
rect 7524 116 7530 128
rect 22830 116 22836 128
rect 7524 88 22836 116
rect 7524 76 7530 88
rect 22830 76 22836 88
rect 22888 76 22894 128
rect 3970 8 3976 60
rect 4028 48 4034 60
rect 20438 48 20444 60
rect 4028 20 20444 48
rect 4028 8 4034 20
rect 20438 8 20444 20
rect 20496 8 20502 60
<< via1 >>
rect 1032 21224 1084 21276
rect 14648 21224 14700 21276
rect 1216 21156 1268 21208
rect 14280 21156 14332 21208
rect 1584 21088 1636 21140
rect 2044 21088 2096 21140
rect 2412 21088 2464 21140
rect 15936 21088 15988 21140
rect 2044 20952 2096 21004
rect 16120 20952 16172 21004
rect 3884 20884 3936 20936
rect 9128 20884 9180 20936
rect 1952 20748 2004 20800
rect 4068 20748 4120 20800
rect 7380 20748 7432 20800
rect 17684 20748 17736 20800
rect 18052 20748 18104 20800
rect 19708 20748 19760 20800
rect 6148 20646 6200 20698
rect 6212 20646 6264 20698
rect 6276 20646 6328 20698
rect 6340 20646 6392 20698
rect 6404 20646 6456 20698
rect 11346 20646 11398 20698
rect 11410 20646 11462 20698
rect 11474 20646 11526 20698
rect 11538 20646 11590 20698
rect 11602 20646 11654 20698
rect 16544 20646 16596 20698
rect 16608 20646 16660 20698
rect 16672 20646 16724 20698
rect 16736 20646 16788 20698
rect 16800 20646 16852 20698
rect 21742 20646 21794 20698
rect 21806 20646 21858 20698
rect 21870 20646 21922 20698
rect 21934 20646 21986 20698
rect 21998 20646 22050 20698
rect 1860 20587 1912 20596
rect 1860 20553 1869 20587
rect 1869 20553 1903 20587
rect 1903 20553 1912 20587
rect 1860 20544 1912 20553
rect 3884 20587 3936 20596
rect 3884 20553 3893 20587
rect 3893 20553 3927 20587
rect 3927 20553 3936 20587
rect 3884 20544 3936 20553
rect 2872 20519 2924 20528
rect 2872 20485 2881 20519
rect 2881 20485 2915 20519
rect 2915 20485 2924 20519
rect 2872 20476 2924 20485
rect 4160 20476 4212 20528
rect 9772 20544 9824 20596
rect 10876 20544 10928 20596
rect 11704 20544 11756 20596
rect 11980 20544 12032 20596
rect 12440 20544 12492 20596
rect 12716 20544 12768 20596
rect 13084 20544 13136 20596
rect 13452 20544 13504 20596
rect 13820 20544 13872 20596
rect 14556 20544 14608 20596
rect 15200 20544 15252 20596
rect 15384 20544 15436 20596
rect 15752 20544 15804 20596
rect 16580 20544 16632 20596
rect 17500 20544 17552 20596
rect 19524 20587 19576 20596
rect 1952 20408 2004 20460
rect 2044 20451 2096 20460
rect 2044 20417 2053 20451
rect 2053 20417 2087 20451
rect 2087 20417 2096 20451
rect 2044 20408 2096 20417
rect 2596 20408 2648 20460
rect 2688 20451 2740 20460
rect 2688 20417 2697 20451
rect 2697 20417 2731 20451
rect 2731 20417 2740 20451
rect 2688 20408 2740 20417
rect 2964 20408 3016 20460
rect 3332 20408 3384 20460
rect 4712 20408 4764 20460
rect 7104 20408 7156 20460
rect 7288 20408 7340 20460
rect 3976 20383 4028 20392
rect 3976 20349 3985 20383
rect 3985 20349 4019 20383
rect 4019 20349 4028 20383
rect 3976 20340 4028 20349
rect 5908 20383 5960 20392
rect 5908 20349 5917 20383
rect 5917 20349 5951 20383
rect 5951 20349 5960 20383
rect 5908 20340 5960 20349
rect 10600 20476 10652 20528
rect 3424 20272 3476 20324
rect 1492 20247 1544 20256
rect 1492 20213 1501 20247
rect 1501 20213 1535 20247
rect 1535 20213 1544 20247
rect 1492 20204 1544 20213
rect 2136 20204 2188 20256
rect 3884 20204 3936 20256
rect 8392 20340 8444 20392
rect 8668 20408 8720 20460
rect 9128 20451 9180 20460
rect 9128 20417 9137 20451
rect 9137 20417 9171 20451
rect 9171 20417 9180 20451
rect 9128 20408 9180 20417
rect 10140 20451 10192 20460
rect 9496 20340 9548 20392
rect 10140 20417 10149 20451
rect 10149 20417 10183 20451
rect 10183 20417 10192 20451
rect 10140 20408 10192 20417
rect 10508 20451 10560 20460
rect 10508 20417 10517 20451
rect 10517 20417 10551 20451
rect 10551 20417 10560 20451
rect 10508 20408 10560 20417
rect 10692 20408 10744 20460
rect 11796 20408 11848 20460
rect 13084 20451 13136 20460
rect 13084 20417 13093 20451
rect 13093 20417 13127 20451
rect 13127 20417 13136 20451
rect 13084 20408 13136 20417
rect 14372 20451 14424 20460
rect 10416 20340 10468 20392
rect 10784 20383 10836 20392
rect 10784 20349 10793 20383
rect 10793 20349 10827 20383
rect 10827 20349 10836 20383
rect 10784 20340 10836 20349
rect 11888 20340 11940 20392
rect 14372 20417 14381 20451
rect 14381 20417 14415 20451
rect 14415 20417 14424 20451
rect 14372 20408 14424 20417
rect 14740 20451 14792 20460
rect 14740 20417 14749 20451
rect 14749 20417 14783 20451
rect 14783 20417 14792 20451
rect 14740 20408 14792 20417
rect 16304 20476 16356 20528
rect 19524 20553 19533 20587
rect 19533 20553 19567 20587
rect 19567 20553 19576 20587
rect 19524 20544 19576 20553
rect 19984 20587 20036 20596
rect 19984 20553 19993 20587
rect 19993 20553 20027 20587
rect 20027 20553 20036 20587
rect 19984 20544 20036 20553
rect 21180 20544 21232 20596
rect 15476 20451 15528 20460
rect 15476 20417 15485 20451
rect 15485 20417 15519 20451
rect 15519 20417 15528 20451
rect 15476 20408 15528 20417
rect 15844 20451 15896 20460
rect 15844 20417 15853 20451
rect 15853 20417 15887 20451
rect 15887 20417 15896 20451
rect 15844 20408 15896 20417
rect 16212 20451 16264 20460
rect 16212 20417 16221 20451
rect 16221 20417 16255 20451
rect 16255 20417 16264 20451
rect 16212 20408 16264 20417
rect 15568 20340 15620 20392
rect 17040 20408 17092 20460
rect 17132 20408 17184 20460
rect 17408 20451 17460 20460
rect 17408 20417 17417 20451
rect 17417 20417 17451 20451
rect 17451 20417 17460 20451
rect 17408 20408 17460 20417
rect 17592 20408 17644 20460
rect 18144 20451 18196 20460
rect 18144 20417 18153 20451
rect 18153 20417 18187 20451
rect 18187 20417 18196 20451
rect 18144 20408 18196 20417
rect 18328 20408 18380 20460
rect 5356 20247 5408 20256
rect 5356 20213 5365 20247
rect 5365 20213 5399 20247
rect 5399 20213 5408 20247
rect 5356 20204 5408 20213
rect 5540 20204 5592 20256
rect 6828 20204 6880 20256
rect 7748 20247 7800 20256
rect 7748 20213 7757 20247
rect 7757 20213 7791 20247
rect 7791 20213 7800 20247
rect 7748 20204 7800 20213
rect 8300 20204 8352 20256
rect 9312 20204 9364 20256
rect 10232 20272 10284 20324
rect 10968 20272 11020 20324
rect 14188 20272 14240 20324
rect 16028 20272 16080 20324
rect 16948 20272 17000 20324
rect 17960 20340 18012 20392
rect 18972 20408 19024 20460
rect 19708 20451 19760 20460
rect 19708 20417 19717 20451
rect 19717 20417 19751 20451
rect 19751 20417 19760 20451
rect 19708 20408 19760 20417
rect 19800 20451 19852 20460
rect 19800 20417 19809 20451
rect 19809 20417 19843 20451
rect 19843 20417 19852 20451
rect 19800 20408 19852 20417
rect 19064 20340 19116 20392
rect 11152 20204 11204 20256
rect 13820 20204 13872 20256
rect 15660 20204 15712 20256
rect 16120 20204 16172 20256
rect 17224 20204 17276 20256
rect 18880 20272 18932 20324
rect 20720 20408 20772 20460
rect 21364 20408 21416 20460
rect 21548 20272 21600 20324
rect 20168 20204 20220 20256
rect 20352 20247 20404 20256
rect 20352 20213 20361 20247
rect 20361 20213 20395 20247
rect 20395 20213 20404 20247
rect 20352 20204 20404 20213
rect 21088 20247 21140 20256
rect 21088 20213 21097 20247
rect 21097 20213 21131 20247
rect 21131 20213 21140 20247
rect 21088 20204 21140 20213
rect 3549 20102 3601 20154
rect 3613 20102 3665 20154
rect 3677 20102 3729 20154
rect 3741 20102 3793 20154
rect 3805 20102 3857 20154
rect 8747 20102 8799 20154
rect 8811 20102 8863 20154
rect 8875 20102 8927 20154
rect 8939 20102 8991 20154
rect 9003 20102 9055 20154
rect 13945 20102 13997 20154
rect 14009 20102 14061 20154
rect 14073 20102 14125 20154
rect 14137 20102 14189 20154
rect 14201 20102 14253 20154
rect 19143 20102 19195 20154
rect 19207 20102 19259 20154
rect 19271 20102 19323 20154
rect 19335 20102 19387 20154
rect 19399 20102 19451 20154
rect 2228 20043 2280 20052
rect 2228 20009 2237 20043
rect 2237 20009 2271 20043
rect 2271 20009 2280 20043
rect 2228 20000 2280 20009
rect 2320 20000 2372 20052
rect 4252 19864 4304 19916
rect 4896 19864 4948 19916
rect 6736 20000 6788 20052
rect 7932 20000 7984 20052
rect 11244 20000 11296 20052
rect 12440 19932 12492 19984
rect 14372 19932 14424 19984
rect 1952 19796 2004 19848
rect 2320 19796 2372 19848
rect 2412 19839 2464 19848
rect 2412 19805 2421 19839
rect 2421 19805 2455 19839
rect 2455 19805 2464 19839
rect 2412 19796 2464 19805
rect 3148 19796 3200 19848
rect 3884 19796 3936 19848
rect 4620 19839 4672 19848
rect 3056 19728 3108 19780
rect 4252 19728 4304 19780
rect 1492 19703 1544 19712
rect 1492 19669 1501 19703
rect 1501 19669 1535 19703
rect 1535 19669 1544 19703
rect 1492 19660 1544 19669
rect 1860 19703 1912 19712
rect 1860 19669 1869 19703
rect 1869 19669 1903 19703
rect 1903 19669 1912 19703
rect 1860 19660 1912 19669
rect 3148 19703 3200 19712
rect 3148 19669 3157 19703
rect 3157 19669 3191 19703
rect 3191 19669 3200 19703
rect 3148 19660 3200 19669
rect 4068 19660 4120 19712
rect 4620 19805 4629 19839
rect 4629 19805 4663 19839
rect 4663 19805 4672 19839
rect 4620 19796 4672 19805
rect 4436 19728 4488 19780
rect 4804 19796 4856 19848
rect 6828 19839 6880 19848
rect 6828 19805 6837 19839
rect 6837 19805 6871 19839
rect 6871 19805 6880 19839
rect 6828 19796 6880 19805
rect 7472 19796 7524 19848
rect 5448 19728 5500 19780
rect 5724 19728 5776 19780
rect 8300 19864 8352 19916
rect 8392 19864 8444 19916
rect 11060 19864 11112 19916
rect 4528 19660 4580 19712
rect 5080 19660 5132 19712
rect 7748 19660 7800 19712
rect 8392 19728 8444 19780
rect 8300 19703 8352 19712
rect 8300 19669 8309 19703
rect 8309 19669 8343 19703
rect 8343 19669 8352 19703
rect 8576 19703 8628 19712
rect 8300 19660 8352 19669
rect 8576 19669 8585 19703
rect 8585 19669 8619 19703
rect 8619 19669 8628 19703
rect 8576 19660 8628 19669
rect 8760 19660 8812 19712
rect 10876 19839 10928 19848
rect 10876 19805 10885 19839
rect 10885 19805 10919 19839
rect 10919 19805 10928 19839
rect 10876 19796 10928 19805
rect 11244 19796 11296 19848
rect 12992 19796 13044 19848
rect 14188 19839 14240 19848
rect 10968 19728 11020 19780
rect 13176 19728 13228 19780
rect 14188 19805 14197 19839
rect 14197 19805 14231 19839
rect 14231 19805 14240 19839
rect 14188 19796 14240 19805
rect 15568 20000 15620 20052
rect 16212 20000 16264 20052
rect 17132 20043 17184 20052
rect 17132 20009 17141 20043
rect 17141 20009 17175 20043
rect 17175 20009 17184 20043
rect 17132 20000 17184 20009
rect 17592 20043 17644 20052
rect 17592 20009 17601 20043
rect 17601 20009 17635 20043
rect 17635 20009 17644 20043
rect 17592 20000 17644 20009
rect 17684 20043 17736 20052
rect 17684 20009 17693 20043
rect 17693 20009 17727 20043
rect 17727 20009 17736 20043
rect 17684 20000 17736 20009
rect 18236 20000 18288 20052
rect 18696 20000 18748 20052
rect 19340 20000 19392 20052
rect 20076 20000 20128 20052
rect 15844 19932 15896 19984
rect 17960 19975 18012 19984
rect 17960 19941 17969 19975
rect 17969 19941 18003 19975
rect 18003 19941 18012 19975
rect 17960 19932 18012 19941
rect 18788 19932 18840 19984
rect 19064 19932 19116 19984
rect 15752 19864 15804 19916
rect 15660 19839 15712 19848
rect 15660 19805 15669 19839
rect 15669 19805 15703 19839
rect 15703 19805 15712 19839
rect 15660 19796 15712 19805
rect 16396 19864 16448 19916
rect 11704 19660 11756 19712
rect 13544 19660 13596 19712
rect 13820 19703 13872 19712
rect 13820 19669 13829 19703
rect 13829 19669 13863 19703
rect 13863 19669 13872 19703
rect 13820 19660 13872 19669
rect 13912 19660 13964 19712
rect 15200 19660 15252 19712
rect 16396 19728 16448 19780
rect 16948 19796 17000 19848
rect 17224 19796 17276 19848
rect 17684 19864 17736 19916
rect 19616 19907 19668 19916
rect 19616 19873 19625 19907
rect 19625 19873 19659 19907
rect 19659 19873 19668 19907
rect 20260 19907 20312 19916
rect 19616 19864 19668 19873
rect 17132 19728 17184 19780
rect 18420 19796 18472 19848
rect 18788 19796 18840 19848
rect 19524 19796 19576 19848
rect 19616 19728 19668 19780
rect 20260 19873 20269 19907
rect 20269 19873 20303 19907
rect 20303 19873 20312 19907
rect 20260 19864 20312 19873
rect 20444 19796 20496 19848
rect 21180 19796 21232 19848
rect 20260 19728 20312 19780
rect 20812 19728 20864 19780
rect 16304 19703 16356 19712
rect 16304 19669 16313 19703
rect 16313 19669 16347 19703
rect 16347 19669 16356 19703
rect 16304 19660 16356 19669
rect 21548 19660 21600 19712
rect 6148 19558 6200 19610
rect 6212 19558 6264 19610
rect 6276 19558 6328 19610
rect 6340 19558 6392 19610
rect 6404 19558 6456 19610
rect 11346 19558 11398 19610
rect 11410 19558 11462 19610
rect 11474 19558 11526 19610
rect 11538 19558 11590 19610
rect 11602 19558 11654 19610
rect 16544 19558 16596 19610
rect 16608 19558 16660 19610
rect 16672 19558 16724 19610
rect 16736 19558 16788 19610
rect 16800 19558 16852 19610
rect 21742 19558 21794 19610
rect 21806 19558 21858 19610
rect 21870 19558 21922 19610
rect 21934 19558 21986 19610
rect 21998 19558 22050 19610
rect 1768 19456 1820 19508
rect 20 19388 72 19440
rect 940 19388 992 19440
rect 1400 19320 1452 19372
rect 2044 19363 2096 19372
rect 2044 19329 2053 19363
rect 2053 19329 2087 19363
rect 2087 19329 2096 19363
rect 2044 19320 2096 19329
rect 2136 19320 2188 19372
rect 3056 19388 3108 19440
rect 5356 19388 5408 19440
rect 5540 19456 5592 19508
rect 8208 19456 8260 19508
rect 6736 19431 6788 19440
rect 6736 19397 6745 19431
rect 6745 19397 6779 19431
rect 6779 19397 6788 19431
rect 6736 19388 6788 19397
rect 7932 19388 7984 19440
rect 8668 19388 8720 19440
rect 10232 19456 10284 19508
rect 11888 19456 11940 19508
rect 12992 19499 13044 19508
rect 12992 19465 13001 19499
rect 13001 19465 13035 19499
rect 13035 19465 13044 19499
rect 12992 19456 13044 19465
rect 13084 19456 13136 19508
rect 14188 19456 14240 19508
rect 10416 19388 10468 19440
rect 10876 19388 10928 19440
rect 3424 19184 3476 19236
rect 3608 19320 3660 19372
rect 4804 19363 4856 19372
rect 4528 19252 4580 19304
rect 4804 19329 4813 19363
rect 4813 19329 4847 19363
rect 4847 19329 4856 19363
rect 4804 19320 4856 19329
rect 7104 19320 7156 19372
rect 7288 19363 7340 19372
rect 7288 19329 7297 19363
rect 7297 19329 7331 19363
rect 7331 19329 7340 19363
rect 7288 19320 7340 19329
rect 8484 19320 8536 19372
rect 6276 19252 6328 19304
rect 7012 19252 7064 19304
rect 7564 19295 7616 19304
rect 7564 19261 7573 19295
rect 7573 19261 7607 19295
rect 7607 19261 7616 19295
rect 7564 19252 7616 19261
rect 7748 19252 7800 19304
rect 7932 19252 7984 19304
rect 9128 19320 9180 19372
rect 11060 19363 11112 19372
rect 11060 19329 11069 19363
rect 11069 19329 11103 19363
rect 11103 19329 11112 19363
rect 11060 19320 11112 19329
rect 12164 19388 12216 19440
rect 13912 19388 13964 19440
rect 14740 19456 14792 19508
rect 15844 19456 15896 19508
rect 13360 19363 13412 19372
rect 8760 19295 8812 19304
rect 8760 19261 8769 19295
rect 8769 19261 8803 19295
rect 8803 19261 8812 19295
rect 8760 19252 8812 19261
rect 13360 19329 13369 19363
rect 13369 19329 13403 19363
rect 13403 19329 13412 19363
rect 13360 19320 13412 19329
rect 14096 19320 14148 19372
rect 12900 19252 12952 19304
rect 13544 19295 13596 19304
rect 13544 19261 13553 19295
rect 13553 19261 13587 19295
rect 13587 19261 13596 19295
rect 13544 19252 13596 19261
rect 15752 19320 15804 19372
rect 17408 19456 17460 19508
rect 18328 19456 18380 19508
rect 18788 19499 18840 19508
rect 18788 19465 18797 19499
rect 18797 19465 18831 19499
rect 18831 19465 18840 19499
rect 18788 19456 18840 19465
rect 18972 19456 19024 19508
rect 19064 19499 19116 19508
rect 19064 19465 19073 19499
rect 19073 19465 19107 19499
rect 19107 19465 19116 19499
rect 19064 19456 19116 19465
rect 16856 19363 16908 19372
rect 16856 19329 16865 19363
rect 16865 19329 16899 19363
rect 16899 19329 16908 19363
rect 16856 19320 16908 19329
rect 16120 19252 16172 19304
rect 1492 19159 1544 19168
rect 1492 19125 1501 19159
rect 1501 19125 1535 19159
rect 1535 19125 1544 19159
rect 1492 19116 1544 19125
rect 2228 19159 2280 19168
rect 2228 19125 2237 19159
rect 2237 19125 2271 19159
rect 2271 19125 2280 19159
rect 2228 19116 2280 19125
rect 3056 19159 3108 19168
rect 3056 19125 3065 19159
rect 3065 19125 3099 19159
rect 3099 19125 3108 19159
rect 3056 19116 3108 19125
rect 3332 19116 3384 19168
rect 3608 19116 3660 19168
rect 3884 19159 3936 19168
rect 3884 19125 3893 19159
rect 3893 19125 3927 19159
rect 3927 19125 3936 19159
rect 3884 19116 3936 19125
rect 4988 19116 5040 19168
rect 5080 19116 5132 19168
rect 8392 19184 8444 19236
rect 8852 19184 8904 19236
rect 6552 19116 6604 19168
rect 6736 19116 6788 19168
rect 6920 19159 6972 19168
rect 6920 19125 6929 19159
rect 6929 19125 6963 19159
rect 6963 19125 6972 19159
rect 6920 19116 6972 19125
rect 7012 19116 7064 19168
rect 7656 19116 7708 19168
rect 9588 19116 9640 19168
rect 9680 19159 9732 19168
rect 9680 19125 9689 19159
rect 9689 19125 9723 19159
rect 9723 19125 9732 19159
rect 11060 19184 11112 19236
rect 15936 19184 15988 19236
rect 9680 19116 9732 19125
rect 12808 19116 12860 19168
rect 13176 19116 13228 19168
rect 15660 19116 15712 19168
rect 18144 19388 18196 19440
rect 20076 19456 20128 19508
rect 20536 19499 20588 19508
rect 20536 19465 20545 19499
rect 20545 19465 20579 19499
rect 20579 19465 20588 19499
rect 20536 19456 20588 19465
rect 21456 19499 21508 19508
rect 21456 19465 21465 19499
rect 21465 19465 21499 19499
rect 21499 19465 21508 19499
rect 21456 19456 21508 19465
rect 17776 19363 17828 19372
rect 17776 19329 17785 19363
rect 17785 19329 17819 19363
rect 17819 19329 17828 19363
rect 17776 19320 17828 19329
rect 18236 19320 18288 19372
rect 18696 19363 18748 19372
rect 17316 19227 17368 19236
rect 17316 19193 17325 19227
rect 17325 19193 17359 19227
rect 17359 19193 17368 19227
rect 17316 19184 17368 19193
rect 17408 19159 17460 19168
rect 17408 19125 17417 19159
rect 17417 19125 17451 19159
rect 17451 19125 17460 19159
rect 17408 19116 17460 19125
rect 17684 19159 17736 19168
rect 17684 19125 17693 19159
rect 17693 19125 17727 19159
rect 17727 19125 17736 19159
rect 17684 19116 17736 19125
rect 18696 19329 18705 19363
rect 18705 19329 18739 19363
rect 18739 19329 18748 19363
rect 18696 19320 18748 19329
rect 19156 19320 19208 19372
rect 20168 19388 20220 19440
rect 20260 19388 20312 19440
rect 18604 19252 18656 19304
rect 19432 19320 19484 19372
rect 19892 19320 19944 19372
rect 20444 19320 20496 19372
rect 20996 19363 21048 19372
rect 20996 19329 21005 19363
rect 21005 19329 21039 19363
rect 21039 19329 21048 19363
rect 20996 19320 21048 19329
rect 21272 19363 21324 19372
rect 21272 19329 21281 19363
rect 21281 19329 21315 19363
rect 21315 19329 21324 19363
rect 21272 19320 21324 19329
rect 20628 19252 20680 19304
rect 20260 19184 20312 19236
rect 18972 19116 19024 19168
rect 3549 19014 3601 19066
rect 3613 19014 3665 19066
rect 3677 19014 3729 19066
rect 3741 19014 3793 19066
rect 3805 19014 3857 19066
rect 8747 19014 8799 19066
rect 8811 19014 8863 19066
rect 8875 19014 8927 19066
rect 8939 19014 8991 19066
rect 9003 19014 9055 19066
rect 13945 19014 13997 19066
rect 14009 19014 14061 19066
rect 14073 19014 14125 19066
rect 14137 19014 14189 19066
rect 14201 19014 14253 19066
rect 19143 19014 19195 19066
rect 19207 19014 19259 19066
rect 19271 19014 19323 19066
rect 19335 19014 19387 19066
rect 19399 19014 19451 19066
rect 3148 18912 3200 18964
rect 2228 18844 2280 18896
rect 6276 18912 6328 18964
rect 6736 18912 6788 18964
rect 7932 18912 7984 18964
rect 8484 18955 8536 18964
rect 8484 18921 8493 18955
rect 8493 18921 8527 18955
rect 8527 18921 8536 18955
rect 8484 18912 8536 18921
rect 8668 18912 8720 18964
rect 10600 18912 10652 18964
rect 11796 18912 11848 18964
rect 12900 18912 12952 18964
rect 13360 18912 13412 18964
rect 15476 18955 15528 18964
rect 15476 18921 15485 18955
rect 15485 18921 15519 18955
rect 15519 18921 15528 18955
rect 15476 18912 15528 18921
rect 17040 18912 17092 18964
rect 18052 18912 18104 18964
rect 18512 18955 18564 18964
rect 18512 18921 18521 18955
rect 18521 18921 18555 18955
rect 18555 18921 18564 18955
rect 18512 18912 18564 18921
rect 5356 18887 5408 18896
rect 5356 18853 5365 18887
rect 5365 18853 5399 18887
rect 5399 18853 5408 18887
rect 5356 18844 5408 18853
rect 3332 18819 3384 18828
rect 3332 18785 3341 18819
rect 3341 18785 3375 18819
rect 3375 18785 3384 18819
rect 3332 18776 3384 18785
rect 3424 18819 3476 18828
rect 3424 18785 3433 18819
rect 3433 18785 3467 18819
rect 3467 18785 3476 18819
rect 3424 18776 3476 18785
rect 3884 18776 3936 18828
rect 4436 18819 4488 18828
rect 4436 18785 4445 18819
rect 4445 18785 4479 18819
rect 4479 18785 4488 18819
rect 4436 18776 4488 18785
rect 4712 18819 4764 18828
rect 4712 18785 4721 18819
rect 4721 18785 4755 18819
rect 4755 18785 4764 18819
rect 4712 18776 4764 18785
rect 2228 18708 2280 18760
rect 2596 18708 2648 18760
rect 3976 18708 4028 18760
rect 4068 18708 4120 18760
rect 5632 18776 5684 18828
rect 8116 18844 8168 18896
rect 6276 18751 6328 18760
rect 6276 18717 6285 18751
rect 6285 18717 6319 18751
rect 6319 18717 6328 18751
rect 6276 18708 6328 18717
rect 7564 18776 7616 18828
rect 9588 18776 9640 18828
rect 16948 18844 17000 18896
rect 7748 18708 7800 18760
rect 6644 18683 6696 18692
rect 6644 18649 6653 18683
rect 6653 18649 6687 18683
rect 6687 18649 6696 18683
rect 6644 18640 6696 18649
rect 6920 18640 6972 18692
rect 1492 18615 1544 18624
rect 1492 18581 1501 18615
rect 1501 18581 1535 18615
rect 1535 18581 1544 18615
rect 1492 18572 1544 18581
rect 2044 18572 2096 18624
rect 2504 18572 2556 18624
rect 2688 18572 2740 18624
rect 3148 18572 3200 18624
rect 3332 18572 3384 18624
rect 4252 18572 4304 18624
rect 4896 18615 4948 18624
rect 4896 18581 4905 18615
rect 4905 18581 4939 18615
rect 4939 18581 4948 18615
rect 4896 18572 4948 18581
rect 4988 18615 5040 18624
rect 4988 18581 4997 18615
rect 4997 18581 5031 18615
rect 5031 18581 5040 18615
rect 4988 18572 5040 18581
rect 5356 18572 5408 18624
rect 5816 18615 5868 18624
rect 5816 18581 5825 18615
rect 5825 18581 5859 18615
rect 5859 18581 5868 18615
rect 5816 18572 5868 18581
rect 5908 18615 5960 18624
rect 5908 18581 5917 18615
rect 5917 18581 5951 18615
rect 5951 18581 5960 18615
rect 5908 18572 5960 18581
rect 7656 18572 7708 18624
rect 7748 18572 7800 18624
rect 9772 18708 9824 18760
rect 10232 18751 10284 18760
rect 8208 18640 8260 18692
rect 9864 18640 9916 18692
rect 10232 18717 10241 18751
rect 10241 18717 10275 18751
rect 10275 18717 10284 18751
rect 10232 18708 10284 18717
rect 10600 18751 10652 18760
rect 10600 18717 10609 18751
rect 10609 18717 10643 18751
rect 10643 18717 10652 18751
rect 10600 18708 10652 18717
rect 10784 18751 10836 18760
rect 10784 18717 10793 18751
rect 10793 18717 10827 18751
rect 10827 18717 10836 18751
rect 10784 18708 10836 18717
rect 11888 18776 11940 18828
rect 12164 18776 12216 18828
rect 12348 18776 12400 18828
rect 12900 18776 12952 18828
rect 13176 18819 13228 18828
rect 13176 18785 13185 18819
rect 13185 18785 13219 18819
rect 13219 18785 13228 18819
rect 13176 18776 13228 18785
rect 11980 18708 12032 18760
rect 8024 18615 8076 18624
rect 8024 18581 8033 18615
rect 8033 18581 8067 18615
rect 8067 18581 8076 18615
rect 8024 18572 8076 18581
rect 8116 18615 8168 18624
rect 8116 18581 8125 18615
rect 8125 18581 8159 18615
rect 8159 18581 8168 18615
rect 8116 18572 8168 18581
rect 8300 18572 8352 18624
rect 8484 18572 8536 18624
rect 8760 18615 8812 18624
rect 8760 18581 8769 18615
rect 8769 18581 8803 18615
rect 8803 18581 8812 18615
rect 8760 18572 8812 18581
rect 9312 18615 9364 18624
rect 9312 18581 9321 18615
rect 9321 18581 9355 18615
rect 9355 18581 9364 18615
rect 9312 18572 9364 18581
rect 9404 18615 9456 18624
rect 9404 18581 9413 18615
rect 9413 18581 9447 18615
rect 9447 18581 9456 18615
rect 9404 18572 9456 18581
rect 9772 18572 9824 18624
rect 12072 18572 12124 18624
rect 12532 18615 12584 18624
rect 12532 18581 12541 18615
rect 12541 18581 12575 18615
rect 12575 18581 12584 18615
rect 13452 18640 13504 18692
rect 16028 18776 16080 18828
rect 17408 18776 17460 18828
rect 15016 18751 15068 18760
rect 15016 18717 15025 18751
rect 15025 18717 15059 18751
rect 15059 18717 15068 18751
rect 15016 18708 15068 18717
rect 15108 18708 15160 18760
rect 15568 18751 15620 18760
rect 15568 18717 15577 18751
rect 15577 18717 15611 18751
rect 15611 18717 15620 18751
rect 15568 18708 15620 18717
rect 18052 18751 18104 18760
rect 18052 18717 18061 18751
rect 18061 18717 18095 18751
rect 18095 18717 18104 18751
rect 18052 18708 18104 18717
rect 19294 18776 19346 18828
rect 19432 18776 19484 18828
rect 18420 18708 18472 18760
rect 18788 18708 18840 18760
rect 18972 18708 19024 18760
rect 19984 18751 20036 18760
rect 19984 18717 19993 18751
rect 19993 18717 20027 18751
rect 20027 18717 20036 18751
rect 19984 18708 20036 18717
rect 22284 18912 22336 18964
rect 20720 18844 20772 18896
rect 20536 18776 20588 18828
rect 12532 18572 12584 18581
rect 13268 18615 13320 18624
rect 13268 18581 13277 18615
rect 13277 18581 13311 18615
rect 13311 18581 13320 18615
rect 13268 18572 13320 18581
rect 13728 18572 13780 18624
rect 14280 18572 14332 18624
rect 14648 18572 14700 18624
rect 19616 18640 19668 18692
rect 20536 18640 20588 18692
rect 20904 18683 20956 18692
rect 20904 18649 20913 18683
rect 20913 18649 20947 18683
rect 20947 18649 20956 18683
rect 20904 18640 20956 18649
rect 15660 18572 15712 18624
rect 16120 18572 16172 18624
rect 16396 18615 16448 18624
rect 16396 18581 16405 18615
rect 16405 18581 16439 18615
rect 16439 18581 16448 18615
rect 16396 18572 16448 18581
rect 17224 18615 17276 18624
rect 17224 18581 17233 18615
rect 17233 18581 17267 18615
rect 17267 18581 17276 18615
rect 17224 18572 17276 18581
rect 18880 18572 18932 18624
rect 19156 18572 19208 18624
rect 19340 18572 19392 18624
rect 19524 18572 19576 18624
rect 20628 18572 20680 18624
rect 21456 18615 21508 18624
rect 21456 18581 21465 18615
rect 21465 18581 21499 18615
rect 21499 18581 21508 18615
rect 21456 18572 21508 18581
rect 6148 18470 6200 18522
rect 6212 18470 6264 18522
rect 6276 18470 6328 18522
rect 6340 18470 6392 18522
rect 6404 18470 6456 18522
rect 11346 18470 11398 18522
rect 11410 18470 11462 18522
rect 11474 18470 11526 18522
rect 11538 18470 11590 18522
rect 11602 18470 11654 18522
rect 16544 18470 16596 18522
rect 16608 18470 16660 18522
rect 16672 18470 16724 18522
rect 16736 18470 16788 18522
rect 16800 18470 16852 18522
rect 21742 18470 21794 18522
rect 21806 18470 21858 18522
rect 21870 18470 21922 18522
rect 21934 18470 21986 18522
rect 21998 18470 22050 18522
rect 3056 18411 3108 18420
rect 3056 18377 3065 18411
rect 3065 18377 3099 18411
rect 3099 18377 3108 18411
rect 3056 18368 3108 18377
rect 3148 18411 3200 18420
rect 3148 18377 3157 18411
rect 3157 18377 3191 18411
rect 3191 18377 3200 18411
rect 3148 18368 3200 18377
rect 4068 18368 4120 18420
rect 5080 18368 5132 18420
rect 3332 18300 3384 18352
rect 2044 18275 2096 18284
rect 2044 18241 2053 18275
rect 2053 18241 2087 18275
rect 2087 18241 2096 18275
rect 2044 18232 2096 18241
rect 2412 18232 2464 18284
rect 2504 18232 2556 18284
rect 3056 18232 3108 18284
rect 4712 18275 4764 18284
rect 4712 18241 4730 18275
rect 4730 18241 4764 18275
rect 4712 18232 4764 18241
rect 2964 18207 3016 18216
rect 2964 18173 2973 18207
rect 2973 18173 3007 18207
rect 3007 18173 3016 18207
rect 2964 18164 3016 18173
rect 1860 18139 1912 18148
rect 1860 18105 1869 18139
rect 1869 18105 1903 18139
rect 1903 18105 1912 18139
rect 1860 18096 1912 18105
rect 3976 18096 4028 18148
rect 1492 18071 1544 18080
rect 1492 18037 1501 18071
rect 1501 18037 1535 18071
rect 1535 18037 1544 18071
rect 1492 18028 1544 18037
rect 2412 18071 2464 18080
rect 2412 18037 2421 18071
rect 2421 18037 2455 18071
rect 2455 18037 2464 18071
rect 2412 18028 2464 18037
rect 4068 18028 4120 18080
rect 5264 18275 5316 18284
rect 5264 18241 5273 18275
rect 5273 18241 5307 18275
rect 5307 18241 5316 18275
rect 5264 18232 5316 18241
rect 5448 18232 5500 18284
rect 5540 18207 5592 18216
rect 5540 18173 5549 18207
rect 5549 18173 5583 18207
rect 5583 18173 5592 18207
rect 5540 18164 5592 18173
rect 5816 18368 5868 18420
rect 5908 18368 5960 18420
rect 7288 18368 7340 18420
rect 7840 18368 7892 18420
rect 8300 18368 8352 18420
rect 9312 18411 9364 18420
rect 9312 18377 9321 18411
rect 9321 18377 9355 18411
rect 9355 18377 9364 18411
rect 9312 18368 9364 18377
rect 10140 18411 10192 18420
rect 10140 18377 10149 18411
rect 10149 18377 10183 18411
rect 10183 18377 10192 18411
rect 10140 18368 10192 18377
rect 6920 18300 6972 18352
rect 7196 18300 7248 18352
rect 7472 18343 7524 18352
rect 7472 18309 7481 18343
rect 7481 18309 7515 18343
rect 7515 18309 7524 18343
rect 7472 18300 7524 18309
rect 7656 18300 7708 18352
rect 5816 18275 5868 18284
rect 5816 18241 5825 18275
rect 5825 18241 5859 18275
rect 5859 18241 5868 18275
rect 5816 18232 5868 18241
rect 6552 18232 6604 18284
rect 8760 18300 8812 18352
rect 6184 18164 6236 18216
rect 6368 18164 6420 18216
rect 6828 18096 6880 18148
rect 7104 18096 7156 18148
rect 5264 18028 5316 18080
rect 6000 18028 6052 18080
rect 6276 18028 6328 18080
rect 7748 18028 7800 18080
rect 8300 18207 8352 18216
rect 8300 18173 8309 18207
rect 8309 18173 8343 18207
rect 8343 18173 8352 18207
rect 8300 18164 8352 18173
rect 8576 18164 8628 18216
rect 8760 18164 8812 18216
rect 9496 18232 9548 18284
rect 9864 18275 9916 18284
rect 9864 18241 9873 18275
rect 9873 18241 9907 18275
rect 9907 18241 9916 18275
rect 9864 18232 9916 18241
rect 10416 18275 10468 18284
rect 10416 18241 10425 18275
rect 10425 18241 10459 18275
rect 10459 18241 10468 18275
rect 10692 18368 10744 18420
rect 11244 18411 11296 18420
rect 11244 18377 11253 18411
rect 11253 18377 11287 18411
rect 11287 18377 11296 18411
rect 11244 18368 11296 18377
rect 11888 18411 11940 18420
rect 11888 18377 11897 18411
rect 11897 18377 11931 18411
rect 11931 18377 11940 18411
rect 11888 18368 11940 18377
rect 11980 18368 12032 18420
rect 12348 18300 12400 18352
rect 12532 18368 12584 18420
rect 13636 18368 13688 18420
rect 14648 18411 14700 18420
rect 14648 18377 14657 18411
rect 14657 18377 14691 18411
rect 14691 18377 14700 18411
rect 14648 18368 14700 18377
rect 15384 18411 15436 18420
rect 15384 18377 15393 18411
rect 15393 18377 15427 18411
rect 15427 18377 15436 18411
rect 15384 18368 15436 18377
rect 18604 18368 18656 18420
rect 19616 18368 19668 18420
rect 19800 18411 19852 18420
rect 19800 18377 19809 18411
rect 19809 18377 19843 18411
rect 19843 18377 19852 18411
rect 19800 18368 19852 18377
rect 19892 18368 19944 18420
rect 14280 18300 14332 18352
rect 18512 18300 18564 18352
rect 10416 18232 10468 18241
rect 9956 18164 10008 18216
rect 11704 18232 11756 18284
rect 12164 18232 12216 18284
rect 13084 18275 13136 18284
rect 8392 18096 8444 18148
rect 11244 18164 11296 18216
rect 13084 18241 13093 18275
rect 13093 18241 13127 18275
rect 13127 18241 13136 18275
rect 13084 18232 13136 18241
rect 15476 18232 15528 18284
rect 13176 18207 13228 18216
rect 9312 18028 9364 18080
rect 9680 18071 9732 18080
rect 9680 18037 9689 18071
rect 9689 18037 9723 18071
rect 9723 18037 9732 18071
rect 10784 18096 10836 18148
rect 9680 18028 9732 18037
rect 11244 18028 11296 18080
rect 11888 18028 11940 18080
rect 12072 18096 12124 18148
rect 13176 18173 13185 18207
rect 13185 18173 13219 18207
rect 13219 18173 13228 18207
rect 13176 18164 13228 18173
rect 14924 18164 14976 18216
rect 13636 18096 13688 18148
rect 16120 18164 16172 18216
rect 19340 18232 19392 18284
rect 20168 18232 20220 18284
rect 20628 18368 20680 18420
rect 21272 18368 21324 18420
rect 20812 18232 20864 18284
rect 20996 18232 21048 18284
rect 21088 18232 21140 18284
rect 21272 18275 21324 18284
rect 21272 18241 21281 18275
rect 21281 18241 21315 18275
rect 21315 18241 21324 18275
rect 21272 18232 21324 18241
rect 16212 18096 16264 18148
rect 18420 18096 18472 18148
rect 19248 18096 19300 18148
rect 20168 18096 20220 18148
rect 20628 18096 20680 18148
rect 21088 18139 21140 18148
rect 21088 18105 21097 18139
rect 21097 18105 21131 18139
rect 21131 18105 21140 18139
rect 21088 18096 21140 18105
rect 12256 18028 12308 18080
rect 12440 18028 12492 18080
rect 15292 18071 15344 18080
rect 15292 18037 15301 18071
rect 15301 18037 15335 18071
rect 15335 18037 15344 18071
rect 15292 18028 15344 18037
rect 15568 18071 15620 18080
rect 15568 18037 15577 18071
rect 15577 18037 15611 18071
rect 15611 18037 15620 18071
rect 15568 18028 15620 18037
rect 22192 18096 22244 18148
rect 21456 18071 21508 18080
rect 21456 18037 21465 18071
rect 21465 18037 21499 18071
rect 21499 18037 21508 18071
rect 21456 18028 21508 18037
rect 3549 17926 3601 17978
rect 3613 17926 3665 17978
rect 3677 17926 3729 17978
rect 3741 17926 3793 17978
rect 3805 17926 3857 17978
rect 8747 17926 8799 17978
rect 8811 17926 8863 17978
rect 8875 17926 8927 17978
rect 8939 17926 8991 17978
rect 9003 17926 9055 17978
rect 13945 17926 13997 17978
rect 14009 17926 14061 17978
rect 14073 17926 14125 17978
rect 14137 17926 14189 17978
rect 14201 17926 14253 17978
rect 19143 17926 19195 17978
rect 19207 17926 19259 17978
rect 19271 17926 19323 17978
rect 19335 17926 19387 17978
rect 19399 17926 19451 17978
rect 1584 17824 1636 17876
rect 2228 17824 2280 17876
rect 5264 17824 5316 17876
rect 5540 17824 5592 17876
rect 7288 17824 7340 17876
rect 8116 17824 8168 17876
rect 9404 17824 9456 17876
rect 9772 17824 9824 17876
rect 10232 17824 10284 17876
rect 10692 17824 10744 17876
rect 1584 17688 1636 17740
rect 1676 17663 1728 17672
rect 1676 17629 1685 17663
rect 1685 17629 1719 17663
rect 1719 17629 1728 17663
rect 1676 17620 1728 17629
rect 1492 17527 1544 17536
rect 1492 17493 1501 17527
rect 1501 17493 1535 17527
rect 1535 17493 1544 17527
rect 1492 17484 1544 17493
rect 1860 17527 1912 17536
rect 1860 17493 1869 17527
rect 1869 17493 1903 17527
rect 1903 17493 1912 17527
rect 1860 17484 1912 17493
rect 2228 17620 2280 17672
rect 3332 17756 3384 17808
rect 3240 17688 3292 17740
rect 3700 17688 3752 17740
rect 3884 17620 3936 17672
rect 4344 17620 4396 17672
rect 4804 17620 4856 17672
rect 6000 17756 6052 17808
rect 5908 17731 5960 17740
rect 5908 17697 5917 17731
rect 5917 17697 5951 17731
rect 5951 17697 5960 17731
rect 5908 17688 5960 17697
rect 8392 17756 8444 17808
rect 3332 17552 3384 17604
rect 3608 17552 3660 17604
rect 3700 17552 3752 17604
rect 5264 17552 5316 17604
rect 5632 17595 5684 17604
rect 5632 17561 5650 17595
rect 5650 17561 5684 17595
rect 6092 17620 6144 17672
rect 6368 17663 6420 17672
rect 6368 17629 6377 17663
rect 6377 17629 6411 17663
rect 6411 17629 6420 17663
rect 6368 17620 6420 17629
rect 8116 17688 8168 17740
rect 8576 17731 8628 17740
rect 8576 17697 8585 17731
rect 8585 17697 8619 17731
rect 8619 17697 8628 17731
rect 8576 17688 8628 17697
rect 8944 17688 8996 17740
rect 5632 17552 5684 17561
rect 6276 17552 6328 17604
rect 6920 17552 6972 17604
rect 9772 17552 9824 17604
rect 3148 17527 3200 17536
rect 3148 17493 3157 17527
rect 3157 17493 3191 17527
rect 3191 17493 3200 17527
rect 3148 17484 3200 17493
rect 3240 17527 3292 17536
rect 3240 17493 3249 17527
rect 3249 17493 3283 17527
rect 3283 17493 3292 17527
rect 3792 17527 3844 17536
rect 3240 17484 3292 17493
rect 3792 17493 3801 17527
rect 3801 17493 3835 17527
rect 3835 17493 3844 17527
rect 3792 17484 3844 17493
rect 4068 17484 4120 17536
rect 4436 17484 4488 17536
rect 4712 17484 4764 17536
rect 5448 17484 5500 17536
rect 6184 17484 6236 17536
rect 7196 17484 7248 17536
rect 7564 17527 7616 17536
rect 7564 17493 7573 17527
rect 7573 17493 7607 17527
rect 7607 17493 7616 17527
rect 7564 17484 7616 17493
rect 8208 17484 8260 17536
rect 8484 17527 8536 17536
rect 8484 17493 8493 17527
rect 8493 17493 8527 17527
rect 8527 17493 8536 17527
rect 8484 17484 8536 17493
rect 8852 17484 8904 17536
rect 13176 17824 13228 17876
rect 15016 17824 15068 17876
rect 15752 17824 15804 17876
rect 13452 17756 13504 17808
rect 10324 17595 10376 17604
rect 10324 17561 10358 17595
rect 10358 17561 10376 17595
rect 10324 17552 10376 17561
rect 10416 17552 10468 17604
rect 11980 17688 12032 17740
rect 12808 17688 12860 17740
rect 14280 17731 14332 17740
rect 14280 17697 14289 17731
rect 14289 17697 14323 17731
rect 14323 17697 14332 17731
rect 14280 17688 14332 17697
rect 17040 17824 17092 17876
rect 17776 17824 17828 17876
rect 18788 17824 18840 17876
rect 19616 17824 19668 17876
rect 20444 17824 20496 17876
rect 20996 17867 21048 17876
rect 20996 17833 21005 17867
rect 21005 17833 21039 17867
rect 21039 17833 21048 17867
rect 20996 17824 21048 17833
rect 19708 17756 19760 17808
rect 19984 17688 20036 17740
rect 21364 17756 21416 17808
rect 21548 17756 21600 17808
rect 22284 17688 22336 17740
rect 11888 17620 11940 17672
rect 11520 17552 11572 17604
rect 12624 17620 12676 17672
rect 13452 17620 13504 17672
rect 15200 17620 15252 17672
rect 15660 17620 15712 17672
rect 20076 17663 20128 17672
rect 20076 17629 20085 17663
rect 20085 17629 20119 17663
rect 20119 17629 20128 17663
rect 20076 17620 20128 17629
rect 20260 17620 20312 17672
rect 20720 17663 20772 17672
rect 20720 17629 20729 17663
rect 20729 17629 20763 17663
rect 20763 17629 20772 17663
rect 20720 17620 20772 17629
rect 21180 17663 21232 17672
rect 21180 17629 21189 17663
rect 21189 17629 21223 17663
rect 21223 17629 21232 17663
rect 21180 17620 21232 17629
rect 13820 17595 13872 17604
rect 13820 17561 13829 17595
rect 13829 17561 13863 17595
rect 13863 17561 13872 17595
rect 13820 17552 13872 17561
rect 15752 17552 15804 17604
rect 16948 17552 17000 17604
rect 19708 17595 19760 17604
rect 19708 17561 19717 17595
rect 19717 17561 19751 17595
rect 19751 17561 19760 17595
rect 19708 17552 19760 17561
rect 20536 17552 20588 17604
rect 12440 17484 12492 17536
rect 13360 17484 13412 17536
rect 14924 17484 14976 17536
rect 15108 17527 15160 17536
rect 15108 17493 15117 17527
rect 15117 17493 15151 17527
rect 15151 17493 15160 17527
rect 15108 17484 15160 17493
rect 20168 17484 20220 17536
rect 20720 17484 20772 17536
rect 22376 17552 22428 17604
rect 6148 17382 6200 17434
rect 6212 17382 6264 17434
rect 6276 17382 6328 17434
rect 6340 17382 6392 17434
rect 6404 17382 6456 17434
rect 11346 17382 11398 17434
rect 11410 17382 11462 17434
rect 11474 17382 11526 17434
rect 11538 17382 11590 17434
rect 11602 17382 11654 17434
rect 16544 17382 16596 17434
rect 16608 17382 16660 17434
rect 16672 17382 16724 17434
rect 16736 17382 16788 17434
rect 16800 17382 16852 17434
rect 21742 17382 21794 17434
rect 21806 17382 21858 17434
rect 21870 17382 21922 17434
rect 21934 17382 21986 17434
rect 21998 17382 22050 17434
rect 1400 17280 1452 17332
rect 3424 17255 3476 17264
rect 2964 17144 3016 17196
rect 3424 17221 3436 17255
rect 3436 17221 3476 17255
rect 3424 17212 3476 17221
rect 3608 17212 3660 17264
rect 4068 17212 4120 17264
rect 4988 17280 5040 17332
rect 5540 17280 5592 17332
rect 6276 17280 6328 17332
rect 8024 17323 8076 17332
rect 1400 16983 1452 16992
rect 1400 16949 1409 16983
rect 1409 16949 1443 16983
rect 1443 16949 1452 16983
rect 1400 16940 1452 16949
rect 2136 16940 2188 16992
rect 2688 16940 2740 16992
rect 4804 17144 4856 17196
rect 4988 17187 5040 17196
rect 4988 17153 4997 17187
rect 4997 17153 5031 17187
rect 5031 17153 5040 17187
rect 4988 17144 5040 17153
rect 4252 17076 4304 17128
rect 5448 17076 5500 17128
rect 5172 17008 5224 17060
rect 5908 17144 5960 17196
rect 6644 17212 6696 17264
rect 6920 17212 6972 17264
rect 8024 17289 8033 17323
rect 8033 17289 8067 17323
rect 8067 17289 8076 17323
rect 8024 17280 8076 17289
rect 8208 17280 8260 17332
rect 8852 17323 8904 17332
rect 6828 17144 6880 17196
rect 6184 17076 6236 17128
rect 6644 17076 6696 17128
rect 7472 17144 7524 17196
rect 8484 17212 8536 17264
rect 7932 17144 7984 17196
rect 8852 17289 8861 17323
rect 8861 17289 8895 17323
rect 8895 17289 8904 17323
rect 8852 17280 8904 17289
rect 8668 17212 8720 17264
rect 11060 17280 11112 17332
rect 11244 17280 11296 17332
rect 9036 17212 9088 17264
rect 9956 17212 10008 17264
rect 9864 17144 9916 17196
rect 10140 17187 10192 17196
rect 10140 17153 10158 17187
rect 10158 17153 10192 17187
rect 10140 17144 10192 17153
rect 10600 17187 10652 17196
rect 10600 17153 10609 17187
rect 10609 17153 10643 17187
rect 10643 17153 10652 17187
rect 11888 17280 11940 17332
rect 12440 17280 12492 17332
rect 13636 17280 13688 17332
rect 14924 17323 14976 17332
rect 14924 17289 14933 17323
rect 14933 17289 14967 17323
rect 14967 17289 14976 17323
rect 14924 17280 14976 17289
rect 15016 17280 15068 17332
rect 11980 17212 12032 17264
rect 12900 17212 12952 17264
rect 17040 17323 17092 17332
rect 17040 17289 17049 17323
rect 17049 17289 17083 17323
rect 17083 17289 17092 17323
rect 17040 17280 17092 17289
rect 19616 17280 19668 17332
rect 21272 17280 21324 17332
rect 10600 17144 10652 17153
rect 13452 17187 13504 17196
rect 13452 17153 13461 17187
rect 13461 17153 13495 17187
rect 13495 17153 13504 17187
rect 13452 17144 13504 17153
rect 15108 17144 15160 17196
rect 15292 17187 15344 17196
rect 15292 17153 15301 17187
rect 15301 17153 15335 17187
rect 15335 17153 15344 17187
rect 15292 17144 15344 17153
rect 7288 17119 7340 17128
rect 7288 17085 7297 17119
rect 7297 17085 7331 17119
rect 7331 17085 7340 17119
rect 7288 17076 7340 17085
rect 8300 17076 8352 17128
rect 8944 17076 8996 17128
rect 10416 17119 10468 17128
rect 10416 17085 10425 17119
rect 10425 17085 10459 17119
rect 10459 17085 10468 17119
rect 10416 17076 10468 17085
rect 4620 16940 4672 16992
rect 6000 16940 6052 16992
rect 6644 16983 6696 16992
rect 6644 16949 6653 16983
rect 6653 16949 6687 16983
rect 6687 16949 6696 16983
rect 6644 16940 6696 16949
rect 7012 17008 7064 17060
rect 8392 17008 8444 17060
rect 9036 17051 9088 17060
rect 9036 17017 9045 17051
rect 9045 17017 9079 17051
rect 9079 17017 9088 17051
rect 9036 17008 9088 17017
rect 12532 17008 12584 17060
rect 10692 16940 10744 16992
rect 11704 16940 11756 16992
rect 13176 16983 13228 16992
rect 13176 16949 13185 16983
rect 13185 16949 13219 16983
rect 13219 16949 13228 16983
rect 13176 16940 13228 16949
rect 13728 16940 13780 16992
rect 15016 17076 15068 17128
rect 15384 17119 15436 17128
rect 15384 17085 15393 17119
rect 15393 17085 15427 17119
rect 15427 17085 15436 17119
rect 15384 17076 15436 17085
rect 16212 17119 16264 17128
rect 15200 17008 15252 17060
rect 16212 17085 16221 17119
rect 16221 17085 16255 17119
rect 16255 17085 16264 17119
rect 16212 17076 16264 17085
rect 18972 17144 19024 17196
rect 21272 17187 21324 17196
rect 21272 17153 21281 17187
rect 21281 17153 21315 17187
rect 21315 17153 21324 17187
rect 21272 17144 21324 17153
rect 17132 17119 17184 17128
rect 17132 17085 17141 17119
rect 17141 17085 17175 17119
rect 17175 17085 17184 17119
rect 17132 17076 17184 17085
rect 17224 17119 17276 17128
rect 17224 17085 17233 17119
rect 17233 17085 17267 17119
rect 17267 17085 17276 17119
rect 17224 17076 17276 17085
rect 15752 17051 15804 17060
rect 15752 17017 15761 17051
rect 15761 17017 15795 17051
rect 15795 17017 15804 17051
rect 15752 17008 15804 17017
rect 16396 17008 16448 17060
rect 20628 17076 20680 17128
rect 21180 17051 21232 17060
rect 21180 17017 21189 17051
rect 21189 17017 21223 17051
rect 21223 17017 21232 17051
rect 21180 17008 21232 17017
rect 22928 17008 22980 17060
rect 15108 16940 15160 16992
rect 17224 16940 17276 16992
rect 17500 16983 17552 16992
rect 17500 16949 17509 16983
rect 17509 16949 17543 16983
rect 17543 16949 17552 16983
rect 17500 16940 17552 16949
rect 19616 16940 19668 16992
rect 20812 16940 20864 16992
rect 21456 16983 21508 16992
rect 21456 16949 21465 16983
rect 21465 16949 21499 16983
rect 21499 16949 21508 16983
rect 21456 16940 21508 16949
rect 3549 16838 3601 16890
rect 3613 16838 3665 16890
rect 3677 16838 3729 16890
rect 3741 16838 3793 16890
rect 3805 16838 3857 16890
rect 8747 16838 8799 16890
rect 8811 16838 8863 16890
rect 8875 16838 8927 16890
rect 8939 16838 8991 16890
rect 9003 16838 9055 16890
rect 13945 16838 13997 16890
rect 14009 16838 14061 16890
rect 14073 16838 14125 16890
rect 14137 16838 14189 16890
rect 14201 16838 14253 16890
rect 19143 16838 19195 16890
rect 19207 16838 19259 16890
rect 19271 16838 19323 16890
rect 19335 16838 19387 16890
rect 19399 16838 19451 16890
rect 1124 16668 1176 16720
rect 1308 16600 1360 16652
rect 2596 16736 2648 16788
rect 3148 16736 3200 16788
rect 5816 16736 5868 16788
rect 6276 16736 6328 16788
rect 7748 16779 7800 16788
rect 3424 16668 3476 16720
rect 3884 16668 3936 16720
rect 6000 16668 6052 16720
rect 6920 16668 6972 16720
rect 1400 16575 1452 16584
rect 1400 16541 1409 16575
rect 1409 16541 1443 16575
rect 1443 16541 1452 16575
rect 1400 16532 1452 16541
rect 2044 16575 2096 16584
rect 2044 16541 2053 16575
rect 2053 16541 2087 16575
rect 2087 16541 2096 16575
rect 2044 16532 2096 16541
rect 5356 16643 5408 16652
rect 5356 16609 5365 16643
rect 5365 16609 5399 16643
rect 5399 16609 5408 16643
rect 5356 16600 5408 16609
rect 5448 16643 5500 16652
rect 5448 16609 5457 16643
rect 5457 16609 5491 16643
rect 5491 16609 5500 16643
rect 5448 16600 5500 16609
rect 5632 16600 5684 16652
rect 6184 16600 6236 16652
rect 7748 16745 7757 16779
rect 7757 16745 7791 16779
rect 7791 16745 7800 16779
rect 7748 16736 7800 16745
rect 9496 16736 9548 16788
rect 9864 16736 9916 16788
rect 10600 16736 10652 16788
rect 11152 16736 11204 16788
rect 11796 16736 11848 16788
rect 12348 16779 12400 16788
rect 12348 16745 12357 16779
rect 12357 16745 12391 16779
rect 12391 16745 12400 16779
rect 12348 16736 12400 16745
rect 12992 16736 13044 16788
rect 14280 16736 14332 16788
rect 15292 16736 15344 16788
rect 17132 16736 17184 16788
rect 7288 16600 7340 16652
rect 7932 16643 7984 16652
rect 7932 16609 7941 16643
rect 7941 16609 7975 16643
rect 7975 16609 7984 16643
rect 7932 16600 7984 16609
rect 8392 16668 8444 16720
rect 8668 16668 8720 16720
rect 11060 16668 11112 16720
rect 9772 16600 9824 16652
rect 9956 16643 10008 16652
rect 9956 16609 9965 16643
rect 9965 16609 9999 16643
rect 9999 16609 10008 16643
rect 9956 16600 10008 16609
rect 10140 16643 10192 16652
rect 10140 16609 10149 16643
rect 10149 16609 10183 16643
rect 10183 16609 10192 16643
rect 10140 16600 10192 16609
rect 3976 16532 4028 16584
rect 4712 16532 4764 16584
rect 6644 16532 6696 16584
rect 7748 16532 7800 16584
rect 8116 16532 8168 16584
rect 10416 16532 10468 16584
rect 10600 16532 10652 16584
rect 11152 16600 11204 16652
rect 11704 16643 11756 16652
rect 11704 16609 11713 16643
rect 11713 16609 11747 16643
rect 11747 16609 11756 16643
rect 11704 16600 11756 16609
rect 12440 16668 12492 16720
rect 12716 16668 12768 16720
rect 15660 16668 15712 16720
rect 12900 16643 12952 16652
rect 12900 16609 12909 16643
rect 12909 16609 12943 16643
rect 12943 16609 12952 16643
rect 12900 16600 12952 16609
rect 12716 16532 12768 16584
rect 12808 16575 12860 16584
rect 12808 16541 12817 16575
rect 12817 16541 12851 16575
rect 12851 16541 12860 16575
rect 13360 16575 13412 16584
rect 12808 16532 12860 16541
rect 13360 16541 13369 16575
rect 13369 16541 13403 16575
rect 13403 16541 13412 16575
rect 13360 16532 13412 16541
rect 15200 16575 15252 16584
rect 15200 16541 15218 16575
rect 15218 16541 15252 16575
rect 15200 16532 15252 16541
rect 2228 16464 2280 16516
rect 4344 16464 4396 16516
rect 1584 16439 1636 16448
rect 1584 16405 1593 16439
rect 1593 16405 1627 16439
rect 1627 16405 1636 16439
rect 1584 16396 1636 16405
rect 1860 16439 1912 16448
rect 1860 16405 1869 16439
rect 1869 16405 1903 16439
rect 1903 16405 1912 16439
rect 1860 16396 1912 16405
rect 4160 16439 4212 16448
rect 4160 16405 4169 16439
rect 4169 16405 4203 16439
rect 4203 16405 4212 16439
rect 4160 16396 4212 16405
rect 4896 16439 4948 16448
rect 4896 16405 4905 16439
rect 4905 16405 4939 16439
rect 4939 16405 4948 16439
rect 5908 16464 5960 16516
rect 7196 16464 7248 16516
rect 4896 16396 4948 16405
rect 6828 16396 6880 16448
rect 6920 16439 6972 16448
rect 6920 16405 6929 16439
rect 6929 16405 6963 16439
rect 6963 16405 6972 16439
rect 7380 16439 7432 16448
rect 6920 16396 6972 16405
rect 7380 16405 7389 16439
rect 7389 16405 7423 16439
rect 7423 16405 7432 16439
rect 7380 16396 7432 16405
rect 8852 16396 8904 16448
rect 8944 16439 8996 16448
rect 8944 16405 8953 16439
rect 8953 16405 8987 16439
rect 8987 16405 8996 16439
rect 9588 16464 9640 16516
rect 11060 16464 11112 16516
rect 8944 16396 8996 16405
rect 9864 16439 9916 16448
rect 9864 16405 9873 16439
rect 9873 16405 9907 16439
rect 9907 16405 9916 16439
rect 9864 16396 9916 16405
rect 11244 16439 11296 16448
rect 11244 16405 11253 16439
rect 11253 16405 11287 16439
rect 11287 16405 11296 16439
rect 11244 16396 11296 16405
rect 11980 16396 12032 16448
rect 13268 16464 13320 16516
rect 16212 16643 16264 16652
rect 16212 16609 16221 16643
rect 16221 16609 16255 16643
rect 16255 16609 16264 16643
rect 16212 16600 16264 16609
rect 17224 16600 17276 16652
rect 16396 16532 16448 16584
rect 19524 16736 19576 16788
rect 19984 16736 20036 16788
rect 20536 16779 20588 16788
rect 20536 16745 20545 16779
rect 20545 16745 20579 16779
rect 20579 16745 20588 16779
rect 20536 16736 20588 16745
rect 21272 16736 21324 16788
rect 17776 16643 17828 16652
rect 17776 16609 17785 16643
rect 17785 16609 17819 16643
rect 17819 16609 17828 16643
rect 17776 16600 17828 16609
rect 16948 16464 17000 16516
rect 19800 16600 19852 16652
rect 20260 16600 20312 16652
rect 20812 16600 20864 16652
rect 18052 16532 18104 16584
rect 20628 16575 20680 16584
rect 20628 16541 20637 16575
rect 20637 16541 20671 16575
rect 20671 16541 20680 16575
rect 20628 16532 20680 16541
rect 12532 16396 12584 16448
rect 12992 16396 13044 16448
rect 13176 16439 13228 16448
rect 13176 16405 13185 16439
rect 13185 16405 13219 16439
rect 13219 16405 13228 16439
rect 13176 16396 13228 16405
rect 15476 16396 15528 16448
rect 15936 16439 15988 16448
rect 15936 16405 15945 16439
rect 15945 16405 15979 16439
rect 15979 16405 15988 16439
rect 15936 16396 15988 16405
rect 16120 16396 16172 16448
rect 20444 16464 20496 16516
rect 21088 16532 21140 16584
rect 17500 16396 17552 16448
rect 20076 16439 20128 16448
rect 20076 16405 20085 16439
rect 20085 16405 20119 16439
rect 20119 16405 20128 16439
rect 20076 16396 20128 16405
rect 20168 16396 20220 16448
rect 21456 16439 21508 16448
rect 21456 16405 21465 16439
rect 21465 16405 21499 16439
rect 21499 16405 21508 16439
rect 21456 16396 21508 16405
rect 20 16260 72 16312
rect 940 16260 992 16312
rect 6148 16294 6200 16346
rect 6212 16294 6264 16346
rect 6276 16294 6328 16346
rect 6340 16294 6392 16346
rect 6404 16294 6456 16346
rect 11346 16294 11398 16346
rect 11410 16294 11462 16346
rect 11474 16294 11526 16346
rect 11538 16294 11590 16346
rect 11602 16294 11654 16346
rect 16544 16294 16596 16346
rect 16608 16294 16660 16346
rect 16672 16294 16724 16346
rect 16736 16294 16788 16346
rect 16800 16294 16852 16346
rect 21742 16294 21794 16346
rect 21806 16294 21858 16346
rect 21870 16294 21922 16346
rect 21934 16294 21986 16346
rect 21998 16294 22050 16346
rect 2044 16192 2096 16244
rect 5632 16192 5684 16244
rect 4620 16167 4672 16176
rect 2136 16056 2188 16108
rect 2228 16031 2280 16040
rect 2228 15997 2237 16031
rect 2237 15997 2271 16031
rect 2271 15997 2280 16031
rect 2228 15988 2280 15997
rect 2412 16031 2464 16040
rect 2412 15997 2421 16031
rect 2421 15997 2455 16031
rect 2455 15997 2464 16031
rect 2412 15988 2464 15997
rect 3240 15988 3292 16040
rect 3884 15988 3936 16040
rect 112 15920 164 15972
rect 1492 15895 1544 15904
rect 1492 15861 1501 15895
rect 1501 15861 1535 15895
rect 1535 15861 1544 15895
rect 1492 15852 1544 15861
rect 3148 15920 3200 15972
rect 4620 16133 4654 16167
rect 4654 16133 4672 16167
rect 4620 16124 4672 16133
rect 5264 16124 5316 16176
rect 6000 16192 6052 16244
rect 6184 16124 6236 16176
rect 7012 16124 7064 16176
rect 10140 16192 10192 16244
rect 11336 16192 11388 16244
rect 12164 16235 12216 16244
rect 12164 16201 12173 16235
rect 12173 16201 12207 16235
rect 12207 16201 12216 16235
rect 12164 16192 12216 16201
rect 12716 16192 12768 16244
rect 15384 16192 15436 16244
rect 15752 16192 15804 16244
rect 4436 16056 4488 16108
rect 6000 16056 6052 16108
rect 7196 16056 7248 16108
rect 7840 16056 7892 16108
rect 8116 16099 8168 16108
rect 8116 16065 8125 16099
rect 8125 16065 8159 16099
rect 8159 16065 8168 16099
rect 8116 16056 8168 16065
rect 8760 16056 8812 16108
rect 9404 16056 9456 16108
rect 6368 16031 6420 16040
rect 4252 15852 4304 15904
rect 6368 15997 6377 16031
rect 6377 15997 6411 16031
rect 6411 15997 6420 16031
rect 6368 15988 6420 15997
rect 5448 15852 5500 15904
rect 6552 15852 6604 15904
rect 9680 15988 9732 16040
rect 9588 15920 9640 15972
rect 10140 16056 10192 16108
rect 10784 15988 10836 16040
rect 10968 16031 11020 16040
rect 10968 15997 10977 16031
rect 10977 15997 11011 16031
rect 11011 15997 11020 16031
rect 10968 15988 11020 15997
rect 12072 16124 12124 16176
rect 13360 16124 13412 16176
rect 14280 16124 14332 16176
rect 11612 16056 11664 16108
rect 11796 16056 11848 16108
rect 13176 16056 13228 16108
rect 15936 16124 15988 16176
rect 17868 16124 17920 16176
rect 17960 16124 18012 16176
rect 19708 16124 19760 16176
rect 15108 16099 15160 16108
rect 15108 16065 15117 16099
rect 15117 16065 15151 16099
rect 15151 16065 15160 16099
rect 15108 16056 15160 16065
rect 16120 16056 16172 16108
rect 11520 16031 11572 16040
rect 11520 15997 11529 16031
rect 11529 15997 11563 16031
rect 11563 15997 11572 16031
rect 11520 15988 11572 15997
rect 14924 16031 14976 16040
rect 14924 15997 14933 16031
rect 14933 15997 14967 16031
rect 14967 15997 14976 16031
rect 14924 15988 14976 15997
rect 15016 16031 15068 16040
rect 15016 15997 15025 16031
rect 15025 15997 15059 16031
rect 15059 15997 15068 16031
rect 15016 15988 15068 15997
rect 15384 15988 15436 16040
rect 17132 16031 17184 16040
rect 10324 15920 10376 15972
rect 17132 15997 17141 16031
rect 17141 15997 17175 16031
rect 17175 15997 17184 16031
rect 17684 16056 17736 16108
rect 17132 15988 17184 15997
rect 18972 15988 19024 16040
rect 19064 16031 19116 16040
rect 19064 15997 19073 16031
rect 19073 15997 19107 16031
rect 19107 15997 19116 16031
rect 19064 15988 19116 15997
rect 8300 15852 8352 15904
rect 8852 15852 8904 15904
rect 9772 15852 9824 15904
rect 10876 15852 10928 15904
rect 12900 15852 12952 15904
rect 13452 15852 13504 15904
rect 16396 15852 16448 15904
rect 17592 15852 17644 15904
rect 18880 15852 18932 15904
rect 19800 16056 19852 16108
rect 20168 16235 20220 16244
rect 20168 16201 20177 16235
rect 20177 16201 20211 16235
rect 20211 16201 20220 16235
rect 20168 16192 20220 16201
rect 20996 16235 21048 16244
rect 20996 16201 21005 16235
rect 21005 16201 21039 16235
rect 21039 16201 21048 16235
rect 20996 16192 21048 16201
rect 20444 16056 20496 16108
rect 20536 16099 20588 16108
rect 20536 16065 20545 16099
rect 20545 16065 20579 16099
rect 20579 16065 20588 16099
rect 20536 16056 20588 16065
rect 20812 16099 20864 16108
rect 20812 16065 20821 16099
rect 20821 16065 20855 16099
rect 20855 16065 20864 16099
rect 20812 16056 20864 16065
rect 22100 15988 22152 16040
rect 19616 15852 19668 15904
rect 19800 15895 19852 15904
rect 19800 15861 19809 15895
rect 19809 15861 19843 15895
rect 19843 15861 19852 15895
rect 19800 15852 19852 15861
rect 20536 15852 20588 15904
rect 21456 15895 21508 15904
rect 21456 15861 21465 15895
rect 21465 15861 21499 15895
rect 21499 15861 21508 15895
rect 21456 15852 21508 15861
rect 3549 15750 3601 15802
rect 3613 15750 3665 15802
rect 3677 15750 3729 15802
rect 3741 15750 3793 15802
rect 3805 15750 3857 15802
rect 8747 15750 8799 15802
rect 8811 15750 8863 15802
rect 8875 15750 8927 15802
rect 8939 15750 8991 15802
rect 9003 15750 9055 15802
rect 13945 15750 13997 15802
rect 14009 15750 14061 15802
rect 14073 15750 14125 15802
rect 14137 15750 14189 15802
rect 14201 15750 14253 15802
rect 19143 15750 19195 15802
rect 19207 15750 19259 15802
rect 19271 15750 19323 15802
rect 19335 15750 19387 15802
rect 19399 15750 19451 15802
rect 1676 15648 1728 15700
rect 2320 15487 2372 15496
rect 1492 15351 1544 15360
rect 1492 15317 1501 15351
rect 1501 15317 1535 15351
rect 1535 15317 1544 15351
rect 1492 15308 1544 15317
rect 2320 15453 2329 15487
rect 2329 15453 2363 15487
rect 2363 15453 2372 15487
rect 2320 15444 2372 15453
rect 4160 15648 4212 15700
rect 4344 15691 4396 15700
rect 4344 15657 4353 15691
rect 4353 15657 4387 15691
rect 4387 15657 4396 15691
rect 4344 15648 4396 15657
rect 4988 15648 5040 15700
rect 6644 15648 6696 15700
rect 6828 15648 6880 15700
rect 7472 15648 7524 15700
rect 3424 15580 3476 15632
rect 2964 15555 3016 15564
rect 2964 15521 2973 15555
rect 2973 15521 3007 15555
rect 3007 15521 3016 15555
rect 2964 15512 3016 15521
rect 3884 15512 3936 15564
rect 3792 15444 3844 15496
rect 4620 15512 4672 15564
rect 5908 15580 5960 15632
rect 9312 15648 9364 15700
rect 9864 15648 9916 15700
rect 10784 15691 10836 15700
rect 10784 15657 10793 15691
rect 10793 15657 10827 15691
rect 10827 15657 10836 15691
rect 10784 15648 10836 15657
rect 11244 15648 11296 15700
rect 12900 15648 12952 15700
rect 15844 15648 15896 15700
rect 16120 15648 16172 15700
rect 19616 15648 19668 15700
rect 20812 15648 20864 15700
rect 7932 15580 7984 15632
rect 8576 15623 8628 15632
rect 8576 15589 8585 15623
rect 8585 15589 8619 15623
rect 8619 15589 8628 15623
rect 8576 15580 8628 15589
rect 6184 15555 6236 15564
rect 6184 15521 6193 15555
rect 6193 15521 6227 15555
rect 6227 15521 6236 15555
rect 6184 15512 6236 15521
rect 7288 15512 7340 15564
rect 7840 15555 7892 15564
rect 7840 15521 7849 15555
rect 7849 15521 7883 15555
rect 7883 15521 7892 15555
rect 7840 15512 7892 15521
rect 8116 15512 8168 15564
rect 9680 15512 9732 15564
rect 4252 15487 4304 15496
rect 4252 15453 4261 15487
rect 4261 15453 4295 15487
rect 4295 15453 4304 15487
rect 4252 15444 4304 15453
rect 4988 15487 5040 15496
rect 4988 15453 4997 15487
rect 4997 15453 5031 15487
rect 5031 15453 5040 15487
rect 4988 15444 5040 15453
rect 5264 15444 5316 15496
rect 2964 15308 3016 15360
rect 3148 15351 3200 15360
rect 3148 15317 3157 15351
rect 3157 15317 3191 15351
rect 3191 15317 3200 15351
rect 3148 15308 3200 15317
rect 4068 15351 4120 15360
rect 4068 15317 4077 15351
rect 4077 15317 4111 15351
rect 4111 15317 4120 15351
rect 4068 15308 4120 15317
rect 4712 15376 4764 15428
rect 11060 15580 11112 15632
rect 11980 15580 12032 15632
rect 10784 15512 10836 15564
rect 13268 15512 13320 15564
rect 8484 15444 8536 15496
rect 9404 15487 9456 15496
rect 9404 15453 9413 15487
rect 9413 15453 9447 15487
rect 9447 15453 9456 15487
rect 9404 15444 9456 15453
rect 10600 15444 10652 15496
rect 13176 15444 13228 15496
rect 13820 15444 13872 15496
rect 14924 15580 14976 15632
rect 15108 15580 15160 15632
rect 18144 15623 18196 15632
rect 16120 15512 16172 15564
rect 17132 15555 17184 15564
rect 17132 15521 17141 15555
rect 17141 15521 17175 15555
rect 17175 15521 17184 15555
rect 17132 15512 17184 15521
rect 18144 15589 18153 15623
rect 18153 15589 18187 15623
rect 18187 15589 18196 15623
rect 18144 15580 18196 15589
rect 18512 15580 18564 15632
rect 19524 15623 19576 15632
rect 19524 15589 19533 15623
rect 19533 15589 19567 15623
rect 19567 15589 19576 15623
rect 19524 15580 19576 15589
rect 20628 15580 20680 15632
rect 16304 15444 16356 15496
rect 16948 15444 17000 15496
rect 18512 15444 18564 15496
rect 18604 15444 18656 15496
rect 19708 15487 19760 15496
rect 19708 15453 19717 15487
rect 19717 15453 19751 15487
rect 19751 15453 19760 15487
rect 19708 15444 19760 15453
rect 20536 15487 20588 15496
rect 6368 15376 6420 15428
rect 5908 15308 5960 15360
rect 6644 15308 6696 15360
rect 7380 15308 7432 15360
rect 8208 15308 8260 15360
rect 8392 15376 8444 15428
rect 9772 15376 9824 15428
rect 13912 15376 13964 15428
rect 8576 15308 8628 15360
rect 9496 15351 9548 15360
rect 9496 15317 9505 15351
rect 9505 15317 9539 15351
rect 9539 15317 9548 15351
rect 9496 15308 9548 15317
rect 10968 15308 11020 15360
rect 11980 15351 12032 15360
rect 11980 15317 11989 15351
rect 11989 15317 12023 15351
rect 12023 15317 12032 15351
rect 11980 15308 12032 15317
rect 12716 15351 12768 15360
rect 12716 15317 12725 15351
rect 12725 15317 12759 15351
rect 12759 15317 12768 15351
rect 13360 15351 13412 15360
rect 12716 15308 12768 15317
rect 13360 15317 13369 15351
rect 13369 15317 13403 15351
rect 13403 15317 13412 15351
rect 13360 15308 13412 15317
rect 13728 15308 13780 15360
rect 15016 15308 15068 15360
rect 15568 15351 15620 15360
rect 15568 15317 15577 15351
rect 15577 15317 15611 15351
rect 15611 15317 15620 15351
rect 15568 15308 15620 15317
rect 15660 15351 15712 15360
rect 15660 15317 15669 15351
rect 15669 15317 15703 15351
rect 15703 15317 15712 15351
rect 15660 15308 15712 15317
rect 16396 15308 16448 15360
rect 20536 15453 20545 15487
rect 20545 15453 20579 15487
rect 20579 15453 20588 15487
rect 20536 15444 20588 15453
rect 20720 15512 20772 15564
rect 20996 15444 21048 15496
rect 17776 15351 17828 15360
rect 17776 15317 17785 15351
rect 17785 15317 17819 15351
rect 17819 15317 17828 15351
rect 18328 15351 18380 15360
rect 17776 15308 17828 15317
rect 18328 15317 18337 15351
rect 18337 15317 18371 15351
rect 18371 15317 18380 15351
rect 18328 15308 18380 15317
rect 18696 15308 18748 15360
rect 18880 15351 18932 15360
rect 18880 15317 18889 15351
rect 18889 15317 18923 15351
rect 18923 15317 18932 15351
rect 18880 15308 18932 15317
rect 19616 15308 19668 15360
rect 20168 15351 20220 15360
rect 20168 15317 20177 15351
rect 20177 15317 20211 15351
rect 20211 15317 20220 15351
rect 20168 15308 20220 15317
rect 20812 15308 20864 15360
rect 20996 15351 21048 15360
rect 20996 15317 21005 15351
rect 21005 15317 21039 15351
rect 21039 15317 21048 15351
rect 20996 15308 21048 15317
rect 21456 15351 21508 15360
rect 21456 15317 21465 15351
rect 21465 15317 21499 15351
rect 21499 15317 21508 15351
rect 21456 15308 21508 15317
rect 6148 15206 6200 15258
rect 6212 15206 6264 15258
rect 6276 15206 6328 15258
rect 6340 15206 6392 15258
rect 6404 15206 6456 15258
rect 11346 15206 11398 15258
rect 11410 15206 11462 15258
rect 11474 15206 11526 15258
rect 11538 15206 11590 15258
rect 11602 15206 11654 15258
rect 16544 15206 16596 15258
rect 16608 15206 16660 15258
rect 16672 15206 16724 15258
rect 16736 15206 16788 15258
rect 16800 15206 16852 15258
rect 21742 15206 21794 15258
rect 21806 15206 21858 15258
rect 21870 15206 21922 15258
rect 21934 15206 21986 15258
rect 21998 15206 22050 15258
rect 2412 15104 2464 15156
rect 2964 15036 3016 15088
rect 5356 15104 5408 15156
rect 6092 15147 6144 15156
rect 6092 15113 6101 15147
rect 6101 15113 6135 15147
rect 6135 15113 6144 15147
rect 6092 15104 6144 15113
rect 7564 15104 7616 15156
rect 8392 15147 8444 15156
rect 8392 15113 8401 15147
rect 8401 15113 8435 15147
rect 8435 15113 8444 15147
rect 8392 15104 8444 15113
rect 4988 15036 5040 15088
rect 1676 15011 1728 15020
rect 1676 14977 1685 15011
rect 1685 14977 1719 15011
rect 1719 14977 1728 15011
rect 1676 14968 1728 14977
rect 1860 14875 1912 14884
rect 1860 14841 1869 14875
rect 1869 14841 1903 14875
rect 1903 14841 1912 14875
rect 1860 14832 1912 14841
rect 2504 15011 2556 15020
rect 2504 14977 2513 15011
rect 2513 14977 2547 15011
rect 2547 14977 2556 15011
rect 2504 14968 2556 14977
rect 3332 14968 3384 15020
rect 4344 15011 4396 15020
rect 2412 14900 2464 14952
rect 1492 14807 1544 14816
rect 1492 14773 1501 14807
rect 1501 14773 1535 14807
rect 1535 14773 1544 14807
rect 1492 14764 1544 14773
rect 2688 14764 2740 14816
rect 3424 14764 3476 14816
rect 4344 14977 4353 15011
rect 4353 14977 4387 15011
rect 4387 14977 4396 15011
rect 4344 14968 4396 14977
rect 4896 14968 4948 15020
rect 3884 14875 3936 14884
rect 3884 14841 3893 14875
rect 3893 14841 3927 14875
rect 3927 14841 3936 14875
rect 4804 14900 4856 14952
rect 9220 15104 9272 15156
rect 9956 15104 10008 15156
rect 10784 15104 10836 15156
rect 12256 15104 12308 15156
rect 13084 15104 13136 15156
rect 13360 15104 13412 15156
rect 13912 15147 13964 15156
rect 13912 15113 13921 15147
rect 13921 15113 13955 15147
rect 13955 15113 13964 15147
rect 13912 15104 13964 15113
rect 10876 15036 10928 15088
rect 11060 15036 11112 15088
rect 15752 15104 15804 15156
rect 16120 15147 16172 15156
rect 16120 15113 16129 15147
rect 16129 15113 16163 15147
rect 16163 15113 16172 15147
rect 16120 15104 16172 15113
rect 20168 15104 20220 15156
rect 14188 15036 14240 15088
rect 5908 14968 5960 15020
rect 6000 14968 6052 15020
rect 7012 14943 7064 14952
rect 7012 14909 7021 14943
rect 7021 14909 7055 14943
rect 7055 14909 7064 14943
rect 7656 14968 7708 15020
rect 7012 14900 7064 14909
rect 3884 14832 3936 14841
rect 6000 14832 6052 14884
rect 6828 14832 6880 14884
rect 8300 14968 8352 15020
rect 9128 15011 9180 15020
rect 9128 14977 9137 15011
rect 9137 14977 9171 15011
rect 9171 14977 9180 15011
rect 9128 14968 9180 14977
rect 9220 14968 9272 15020
rect 9680 14943 9732 14952
rect 9680 14909 9689 14943
rect 9689 14909 9723 14943
rect 9723 14909 9732 14943
rect 9680 14900 9732 14909
rect 10600 14968 10652 15020
rect 13360 14968 13412 15020
rect 14280 15011 14332 15020
rect 10416 14900 10468 14952
rect 4620 14764 4672 14816
rect 6368 14807 6420 14816
rect 6368 14773 6377 14807
rect 6377 14773 6411 14807
rect 6411 14773 6420 14807
rect 6368 14764 6420 14773
rect 6644 14764 6696 14816
rect 7564 14807 7616 14816
rect 7564 14773 7573 14807
rect 7573 14773 7607 14807
rect 7607 14773 7616 14807
rect 7564 14764 7616 14773
rect 8392 14832 8444 14884
rect 9036 14832 9088 14884
rect 9496 14832 9548 14884
rect 9128 14764 9180 14816
rect 9404 14764 9456 14816
rect 11060 14900 11112 14952
rect 12256 14900 12308 14952
rect 12808 14943 12860 14952
rect 12808 14909 12817 14943
rect 12817 14909 12851 14943
rect 12851 14909 12860 14943
rect 14280 14977 14289 15011
rect 14289 14977 14323 15011
rect 14323 14977 14332 15011
rect 14280 14968 14332 14977
rect 14832 14968 14884 15020
rect 18512 15036 18564 15088
rect 19524 15036 19576 15088
rect 17132 14968 17184 15020
rect 18328 14968 18380 15020
rect 19064 14968 19116 15020
rect 12808 14900 12860 14909
rect 12624 14832 12676 14884
rect 16856 14943 16908 14952
rect 12256 14807 12308 14816
rect 12256 14773 12265 14807
rect 12265 14773 12299 14807
rect 12299 14773 12308 14807
rect 12256 14764 12308 14773
rect 12532 14764 12584 14816
rect 13820 14764 13872 14816
rect 14464 14764 14516 14816
rect 16856 14909 16865 14943
rect 16865 14909 16899 14943
rect 16899 14909 16908 14943
rect 16856 14900 16908 14909
rect 18512 14943 18564 14952
rect 18512 14909 18521 14943
rect 18521 14909 18555 14943
rect 18555 14909 18564 14943
rect 18512 14900 18564 14909
rect 15752 14764 15804 14816
rect 17776 14764 17828 14816
rect 18328 14764 18380 14816
rect 19524 14764 19576 14816
rect 20812 14968 20864 15020
rect 20996 14968 21048 15020
rect 21364 14900 21416 14952
rect 21088 14875 21140 14884
rect 21088 14841 21097 14875
rect 21097 14841 21131 14875
rect 21131 14841 21140 14875
rect 21088 14832 21140 14841
rect 20444 14764 20496 14816
rect 21456 14807 21508 14816
rect 21456 14773 21465 14807
rect 21465 14773 21499 14807
rect 21499 14773 21508 14807
rect 21456 14764 21508 14773
rect 3549 14662 3601 14714
rect 3613 14662 3665 14714
rect 3677 14662 3729 14714
rect 3741 14662 3793 14714
rect 3805 14662 3857 14714
rect 8747 14662 8799 14714
rect 8811 14662 8863 14714
rect 8875 14662 8927 14714
rect 8939 14662 8991 14714
rect 9003 14662 9055 14714
rect 13945 14662 13997 14714
rect 14009 14662 14061 14714
rect 14073 14662 14125 14714
rect 14137 14662 14189 14714
rect 14201 14662 14253 14714
rect 19143 14662 19195 14714
rect 19207 14662 19259 14714
rect 19271 14662 19323 14714
rect 19335 14662 19387 14714
rect 19399 14662 19451 14714
rect 1768 14603 1820 14612
rect 1768 14569 1777 14603
rect 1777 14569 1811 14603
rect 1811 14569 1820 14603
rect 1768 14560 1820 14569
rect 2320 14560 2372 14612
rect 3056 14603 3108 14612
rect 1676 14492 1728 14544
rect 1768 14424 1820 14476
rect 3056 14569 3065 14603
rect 3065 14569 3099 14603
rect 3099 14569 3108 14603
rect 3056 14560 3108 14569
rect 5540 14560 5592 14612
rect 3976 14492 4028 14544
rect 7656 14560 7708 14612
rect 9128 14560 9180 14612
rect 10508 14560 10560 14612
rect 11888 14603 11940 14612
rect 11888 14569 11897 14603
rect 11897 14569 11931 14603
rect 11931 14569 11940 14603
rect 11888 14560 11940 14569
rect 12624 14560 12676 14612
rect 13268 14560 13320 14612
rect 9956 14492 10008 14544
rect 10324 14492 10376 14544
rect 2320 14356 2372 14408
rect 2596 14356 2648 14408
rect 2780 14356 2832 14408
rect 2964 14356 3016 14408
rect 3240 14356 3292 14408
rect 9220 14424 9272 14476
rect 10048 14467 10100 14476
rect 4160 14356 4212 14408
rect 1492 14263 1544 14272
rect 1492 14229 1501 14263
rect 1501 14229 1535 14263
rect 1535 14229 1544 14263
rect 1492 14220 1544 14229
rect 4068 14288 4120 14340
rect 6368 14356 6420 14408
rect 8300 14399 8352 14408
rect 8300 14365 8329 14399
rect 8329 14365 8352 14399
rect 10048 14433 10057 14467
rect 10057 14433 10091 14467
rect 10091 14433 10100 14467
rect 10048 14424 10100 14433
rect 11796 14424 11848 14476
rect 11980 14467 12032 14476
rect 11980 14433 11989 14467
rect 11989 14433 12023 14467
rect 12023 14433 12032 14467
rect 11980 14424 12032 14433
rect 16396 14560 16448 14612
rect 18512 14603 18564 14612
rect 18512 14569 18521 14603
rect 18521 14569 18555 14603
rect 18555 14569 18564 14603
rect 18512 14560 18564 14569
rect 17132 14535 17184 14544
rect 17132 14501 17141 14535
rect 17141 14501 17175 14535
rect 17175 14501 17184 14535
rect 17132 14492 17184 14501
rect 19892 14560 19944 14612
rect 8300 14356 8352 14365
rect 5356 14288 5408 14340
rect 2872 14220 2924 14272
rect 3424 14220 3476 14272
rect 5172 14220 5224 14272
rect 6552 14288 6604 14340
rect 8576 14288 8628 14340
rect 7012 14263 7064 14272
rect 7012 14229 7021 14263
rect 7021 14229 7055 14263
rect 7055 14229 7064 14263
rect 7012 14220 7064 14229
rect 7748 14220 7800 14272
rect 8024 14220 8076 14272
rect 9588 14288 9640 14340
rect 10324 14399 10376 14408
rect 10324 14365 10333 14399
rect 10333 14365 10367 14399
rect 10367 14365 10376 14399
rect 10324 14356 10376 14365
rect 12624 14356 12676 14408
rect 13820 14356 13872 14408
rect 15752 14399 15804 14408
rect 15752 14365 15761 14399
rect 15761 14365 15795 14399
rect 15795 14365 15804 14399
rect 15752 14356 15804 14365
rect 17224 14424 17276 14476
rect 10600 14288 10652 14340
rect 12808 14288 12860 14340
rect 16120 14288 16172 14340
rect 16856 14356 16908 14408
rect 18788 14492 18840 14544
rect 19800 14492 19852 14544
rect 20352 14492 20404 14544
rect 19524 14424 19576 14476
rect 20628 14467 20680 14476
rect 20628 14433 20637 14467
rect 20637 14433 20671 14467
rect 20671 14433 20680 14467
rect 20628 14424 20680 14433
rect 18420 14356 18472 14408
rect 19800 14356 19852 14408
rect 20444 14399 20496 14408
rect 20444 14365 20453 14399
rect 20453 14365 20487 14399
rect 20487 14365 20496 14399
rect 20444 14356 20496 14365
rect 21272 14399 21324 14408
rect 21272 14365 21281 14399
rect 21281 14365 21315 14399
rect 21315 14365 21324 14399
rect 21272 14356 21324 14365
rect 17408 14288 17460 14340
rect 19616 14331 19668 14340
rect 19616 14297 19625 14331
rect 19625 14297 19659 14331
rect 19659 14297 19668 14331
rect 19616 14288 19668 14297
rect 8760 14263 8812 14272
rect 8760 14229 8769 14263
rect 8769 14229 8803 14263
rect 8803 14229 8812 14263
rect 8944 14263 8996 14272
rect 8760 14220 8812 14229
rect 8944 14229 8953 14263
rect 8953 14229 8987 14263
rect 8987 14229 8996 14263
rect 8944 14220 8996 14229
rect 9220 14220 9272 14272
rect 9496 14220 9548 14272
rect 9956 14220 10008 14272
rect 10140 14263 10192 14272
rect 10140 14229 10149 14263
rect 10149 14229 10183 14263
rect 10183 14229 10192 14263
rect 10140 14220 10192 14229
rect 13452 14263 13504 14272
rect 13452 14229 13461 14263
rect 13461 14229 13495 14263
rect 13495 14229 13504 14263
rect 13452 14220 13504 14229
rect 14096 14220 14148 14272
rect 14556 14220 14608 14272
rect 18420 14220 18472 14272
rect 18788 14220 18840 14272
rect 20076 14263 20128 14272
rect 20076 14229 20085 14263
rect 20085 14229 20119 14263
rect 20119 14229 20128 14263
rect 20076 14220 20128 14229
rect 20812 14220 20864 14272
rect 21456 14263 21508 14272
rect 21456 14229 21465 14263
rect 21465 14229 21499 14263
rect 21499 14229 21508 14263
rect 21456 14220 21508 14229
rect 6148 14118 6200 14170
rect 6212 14118 6264 14170
rect 6276 14118 6328 14170
rect 6340 14118 6392 14170
rect 6404 14118 6456 14170
rect 11346 14118 11398 14170
rect 11410 14118 11462 14170
rect 11474 14118 11526 14170
rect 11538 14118 11590 14170
rect 11602 14118 11654 14170
rect 16544 14118 16596 14170
rect 16608 14118 16660 14170
rect 16672 14118 16724 14170
rect 16736 14118 16788 14170
rect 16800 14118 16852 14170
rect 21742 14118 21794 14170
rect 21806 14118 21858 14170
rect 21870 14118 21922 14170
rect 21934 14118 21986 14170
rect 21998 14118 22050 14170
rect 2320 14016 2372 14068
rect 3148 14016 3200 14068
rect 4528 14016 4580 14068
rect 5908 14059 5960 14068
rect 2412 13948 2464 14000
rect 2136 13880 2188 13932
rect 2964 13923 3016 13932
rect 1584 13812 1636 13864
rect 2964 13889 2973 13923
rect 2973 13889 3007 13923
rect 3007 13889 3016 13923
rect 2964 13880 3016 13889
rect 3884 13948 3936 14000
rect 5264 13948 5316 14000
rect 5908 14025 5917 14059
rect 5917 14025 5951 14059
rect 5951 14025 5960 14059
rect 5908 14016 5960 14025
rect 6000 14016 6052 14068
rect 8944 14016 8996 14068
rect 9036 14016 9088 14068
rect 9588 14016 9640 14068
rect 6552 13948 6604 14000
rect 6920 13948 6972 14000
rect 7012 13948 7064 14000
rect 8392 13948 8444 14000
rect 8576 13948 8628 14000
rect 10784 14016 10836 14068
rect 11060 14059 11112 14068
rect 11060 14025 11069 14059
rect 11069 14025 11103 14059
rect 11103 14025 11112 14059
rect 11060 14016 11112 14025
rect 11428 14016 11480 14068
rect 12532 14016 12584 14068
rect 12716 14059 12768 14068
rect 12716 14025 12725 14059
rect 12725 14025 12759 14059
rect 12759 14025 12768 14059
rect 12716 14016 12768 14025
rect 14280 14016 14332 14068
rect 14556 14016 14608 14068
rect 14924 14016 14976 14068
rect 16948 14016 17000 14068
rect 2412 13855 2464 13864
rect 2412 13821 2421 13855
rect 2421 13821 2455 13855
rect 2455 13821 2464 13855
rect 3056 13855 3108 13864
rect 2412 13812 2464 13821
rect 3056 13821 3065 13855
rect 3065 13821 3099 13855
rect 3099 13821 3108 13855
rect 3056 13812 3108 13821
rect 2504 13744 2556 13796
rect 1492 13719 1544 13728
rect 1492 13685 1501 13719
rect 1501 13685 1535 13719
rect 1535 13685 1544 13719
rect 1492 13676 1544 13685
rect 1860 13719 1912 13728
rect 1860 13685 1869 13719
rect 1869 13685 1903 13719
rect 1903 13685 1912 13719
rect 1860 13676 1912 13685
rect 2412 13676 2464 13728
rect 4252 13812 4304 13864
rect 4620 13812 4672 13864
rect 4896 13855 4948 13864
rect 4896 13821 4905 13855
rect 4905 13821 4939 13855
rect 4939 13821 4948 13855
rect 4896 13812 4948 13821
rect 5172 13812 5224 13864
rect 5448 13855 5500 13864
rect 5448 13821 5457 13855
rect 5457 13821 5491 13855
rect 5491 13821 5500 13855
rect 5448 13812 5500 13821
rect 6000 13855 6052 13864
rect 6000 13821 6009 13855
rect 6009 13821 6043 13855
rect 6043 13821 6052 13855
rect 6000 13812 6052 13821
rect 10508 13880 10560 13932
rect 12532 13880 12584 13932
rect 13544 13880 13596 13932
rect 14096 13923 14148 13932
rect 14096 13889 14105 13923
rect 14105 13889 14139 13923
rect 14139 13889 14148 13923
rect 14096 13880 14148 13889
rect 16212 13948 16264 14000
rect 16304 13948 16356 14000
rect 17960 14016 18012 14068
rect 20168 14016 20220 14068
rect 19524 13948 19576 14000
rect 15844 13923 15896 13932
rect 15844 13889 15853 13923
rect 15853 13889 15887 13923
rect 15887 13889 15896 13923
rect 15844 13880 15896 13889
rect 17132 13923 17184 13932
rect 17132 13889 17141 13923
rect 17141 13889 17175 13923
rect 17175 13889 17184 13923
rect 17132 13880 17184 13889
rect 17316 13880 17368 13932
rect 18236 13880 18288 13932
rect 20628 13948 20680 14000
rect 7656 13855 7708 13864
rect 7656 13821 7665 13855
rect 7665 13821 7699 13855
rect 7699 13821 7708 13855
rect 7656 13812 7708 13821
rect 7748 13855 7800 13864
rect 7748 13821 7757 13855
rect 7757 13821 7791 13855
rect 7791 13821 7800 13855
rect 7748 13812 7800 13821
rect 5908 13744 5960 13796
rect 3424 13719 3476 13728
rect 3424 13685 3433 13719
rect 3433 13685 3467 13719
rect 3467 13685 3476 13719
rect 3424 13676 3476 13685
rect 8208 13676 8260 13728
rect 9404 13812 9456 13864
rect 9496 13812 9548 13864
rect 9588 13744 9640 13796
rect 10232 13812 10284 13864
rect 10600 13855 10652 13864
rect 10600 13821 10609 13855
rect 10609 13821 10643 13855
rect 10643 13821 10652 13855
rect 10600 13812 10652 13821
rect 11520 13855 11572 13864
rect 11520 13821 11529 13855
rect 11529 13821 11563 13855
rect 11563 13821 11572 13855
rect 11520 13812 11572 13821
rect 11704 13855 11756 13864
rect 11704 13821 11713 13855
rect 11713 13821 11747 13855
rect 11747 13821 11756 13855
rect 11704 13812 11756 13821
rect 11888 13812 11940 13864
rect 12256 13855 12308 13864
rect 12256 13821 12265 13855
rect 12265 13821 12299 13855
rect 12299 13821 12308 13855
rect 12256 13812 12308 13821
rect 12808 13812 12860 13864
rect 13268 13812 13320 13864
rect 14004 13812 14056 13864
rect 14740 13812 14792 13864
rect 10968 13744 11020 13796
rect 15568 13812 15620 13864
rect 17224 13855 17276 13864
rect 9128 13676 9180 13728
rect 9772 13676 9824 13728
rect 10600 13676 10652 13728
rect 11244 13676 11296 13728
rect 11980 13676 12032 13728
rect 12716 13676 12768 13728
rect 13360 13676 13412 13728
rect 13544 13676 13596 13728
rect 17224 13821 17233 13855
rect 17233 13821 17267 13855
rect 17267 13821 17276 13855
rect 17224 13812 17276 13821
rect 16120 13744 16172 13796
rect 18052 13812 18104 13864
rect 19800 13923 19852 13932
rect 19800 13889 19809 13923
rect 19809 13889 19843 13923
rect 19843 13889 19852 13923
rect 19800 13880 19852 13889
rect 20352 13880 20404 13932
rect 21548 13880 21600 13932
rect 22652 13880 22704 13932
rect 17132 13676 17184 13728
rect 21180 13719 21232 13728
rect 21180 13685 21189 13719
rect 21189 13685 21223 13719
rect 21223 13685 21232 13719
rect 21180 13676 21232 13685
rect 21456 13719 21508 13728
rect 21456 13685 21465 13719
rect 21465 13685 21499 13719
rect 21499 13685 21508 13719
rect 21456 13676 21508 13685
rect 3549 13574 3601 13626
rect 3613 13574 3665 13626
rect 3677 13574 3729 13626
rect 3741 13574 3793 13626
rect 3805 13574 3857 13626
rect 8747 13574 8799 13626
rect 8811 13574 8863 13626
rect 8875 13574 8927 13626
rect 8939 13574 8991 13626
rect 9003 13574 9055 13626
rect 13945 13574 13997 13626
rect 14009 13574 14061 13626
rect 14073 13574 14125 13626
rect 14137 13574 14189 13626
rect 14201 13574 14253 13626
rect 19143 13574 19195 13626
rect 19207 13574 19259 13626
rect 19271 13574 19323 13626
rect 19335 13574 19387 13626
rect 19399 13574 19451 13626
rect 2504 13472 2556 13524
rect 4160 13515 4212 13524
rect 4160 13481 4169 13515
rect 4169 13481 4203 13515
rect 4203 13481 4212 13515
rect 4160 13472 4212 13481
rect 5264 13515 5316 13524
rect 5264 13481 5273 13515
rect 5273 13481 5307 13515
rect 5307 13481 5316 13515
rect 5264 13472 5316 13481
rect 5448 13472 5500 13524
rect 6552 13472 6604 13524
rect 6920 13515 6972 13524
rect 6920 13481 6929 13515
rect 6929 13481 6963 13515
rect 6963 13481 6972 13515
rect 6920 13472 6972 13481
rect 7656 13472 7708 13524
rect 8392 13472 8444 13524
rect 8576 13472 8628 13524
rect 10508 13515 10560 13524
rect 204 13200 256 13252
rect 1768 13200 1820 13252
rect 1492 13175 1544 13184
rect 1492 13141 1501 13175
rect 1501 13141 1535 13175
rect 1535 13141 1544 13175
rect 1492 13132 1544 13141
rect 2596 13268 2648 13320
rect 4528 13404 4580 13456
rect 5632 13404 5684 13456
rect 7288 13404 7340 13456
rect 3332 13336 3384 13388
rect 3884 13336 3936 13388
rect 4620 13336 4672 13388
rect 5356 13336 5408 13388
rect 7748 13336 7800 13388
rect 3976 13200 4028 13252
rect 6000 13268 6052 13320
rect 5264 13200 5316 13252
rect 6552 13268 6604 13320
rect 8300 13379 8352 13388
rect 8300 13345 8309 13379
rect 8309 13345 8343 13379
rect 8343 13345 8352 13379
rect 8300 13336 8352 13345
rect 10508 13481 10517 13515
rect 10517 13481 10551 13515
rect 10551 13481 10560 13515
rect 10508 13472 10560 13481
rect 11336 13515 11388 13524
rect 11336 13481 11345 13515
rect 11345 13481 11379 13515
rect 11379 13481 11388 13515
rect 11336 13472 11388 13481
rect 11612 13515 11664 13524
rect 11612 13481 11621 13515
rect 11621 13481 11655 13515
rect 11655 13481 11664 13515
rect 11612 13472 11664 13481
rect 11980 13515 12032 13524
rect 11980 13481 11989 13515
rect 11989 13481 12023 13515
rect 12023 13481 12032 13515
rect 11980 13472 12032 13481
rect 13728 13472 13780 13524
rect 14372 13472 14424 13524
rect 15844 13472 15896 13524
rect 18236 13515 18288 13524
rect 18236 13481 18245 13515
rect 18245 13481 18279 13515
rect 18279 13481 18288 13515
rect 18236 13472 18288 13481
rect 19708 13515 19760 13524
rect 19708 13481 19717 13515
rect 19717 13481 19751 13515
rect 19751 13481 19760 13515
rect 19708 13472 19760 13481
rect 21272 13472 21324 13524
rect 16304 13447 16356 13456
rect 8944 13268 8996 13320
rect 9128 13268 9180 13320
rect 10508 13336 10560 13388
rect 11612 13268 11664 13320
rect 11888 13268 11940 13320
rect 6828 13132 6880 13184
rect 7840 13132 7892 13184
rect 8024 13132 8076 13184
rect 8576 13243 8628 13252
rect 8576 13209 8585 13243
rect 8585 13209 8619 13243
rect 8619 13209 8628 13243
rect 12624 13379 12676 13388
rect 12624 13345 12633 13379
rect 12633 13345 12667 13379
rect 12667 13345 12676 13379
rect 12624 13336 12676 13345
rect 14464 13379 14516 13388
rect 14464 13345 14473 13379
rect 14473 13345 14507 13379
rect 14507 13345 14516 13379
rect 14464 13336 14516 13345
rect 13084 13268 13136 13320
rect 14740 13311 14792 13320
rect 8576 13200 8628 13209
rect 12440 13200 12492 13252
rect 12624 13200 12676 13252
rect 13636 13200 13688 13252
rect 8852 13132 8904 13184
rect 9036 13132 9088 13184
rect 9588 13132 9640 13184
rect 11336 13132 11388 13184
rect 12072 13132 12124 13184
rect 12256 13132 12308 13184
rect 12808 13175 12860 13184
rect 12808 13141 12817 13175
rect 12817 13141 12851 13175
rect 12851 13141 12860 13175
rect 12808 13132 12860 13141
rect 13360 13175 13412 13184
rect 13360 13141 13369 13175
rect 13369 13141 13403 13175
rect 13403 13141 13412 13175
rect 13360 13132 13412 13141
rect 13544 13175 13596 13184
rect 13544 13141 13553 13175
rect 13553 13141 13587 13175
rect 13587 13141 13596 13175
rect 13544 13132 13596 13141
rect 14188 13175 14240 13184
rect 14188 13141 14197 13175
rect 14197 13141 14231 13175
rect 14231 13141 14240 13175
rect 14188 13132 14240 13141
rect 14740 13277 14774 13311
rect 14774 13277 14792 13311
rect 14740 13268 14792 13277
rect 15292 13268 15344 13320
rect 15936 13311 15988 13320
rect 15936 13277 15945 13311
rect 15945 13277 15979 13311
rect 15979 13277 15988 13311
rect 15936 13268 15988 13277
rect 16304 13413 16313 13447
rect 16313 13413 16347 13447
rect 16347 13413 16356 13447
rect 16304 13404 16356 13413
rect 20352 13404 20404 13456
rect 16948 13336 17000 13388
rect 18236 13336 18288 13388
rect 18788 13379 18840 13388
rect 18788 13345 18797 13379
rect 18797 13345 18831 13379
rect 18831 13345 18840 13379
rect 18788 13336 18840 13345
rect 19524 13336 19576 13388
rect 20168 13379 20220 13388
rect 20168 13345 20177 13379
rect 20177 13345 20211 13379
rect 20211 13345 20220 13379
rect 20168 13336 20220 13345
rect 21180 13336 21232 13388
rect 17500 13268 17552 13320
rect 19892 13268 19944 13320
rect 20076 13311 20128 13320
rect 20076 13277 20085 13311
rect 20085 13277 20119 13311
rect 20119 13277 20128 13311
rect 20076 13268 20128 13277
rect 20536 13268 20588 13320
rect 20720 13268 20772 13320
rect 21272 13311 21324 13320
rect 14648 13200 14700 13252
rect 15476 13200 15528 13252
rect 14556 13132 14608 13184
rect 14832 13132 14884 13184
rect 15200 13132 15252 13184
rect 16120 13132 16172 13184
rect 17224 13200 17276 13252
rect 17316 13200 17368 13252
rect 19064 13200 19116 13252
rect 21272 13277 21281 13311
rect 21281 13277 21315 13311
rect 21315 13277 21324 13311
rect 21272 13268 21324 13277
rect 17040 13132 17092 13184
rect 17592 13132 17644 13184
rect 18328 13132 18380 13184
rect 18696 13175 18748 13184
rect 18696 13141 18705 13175
rect 18705 13141 18739 13175
rect 18739 13141 18748 13175
rect 21088 13175 21140 13184
rect 18696 13132 18748 13141
rect 21088 13141 21097 13175
rect 21097 13141 21131 13175
rect 21131 13141 21140 13175
rect 21088 13132 21140 13141
rect 21456 13175 21508 13184
rect 21456 13141 21465 13175
rect 21465 13141 21499 13175
rect 21499 13141 21508 13175
rect 21456 13132 21508 13141
rect 22008 13132 22060 13184
rect 22836 13132 22888 13184
rect 6148 13030 6200 13082
rect 6212 13030 6264 13082
rect 6276 13030 6328 13082
rect 6340 13030 6392 13082
rect 6404 13030 6456 13082
rect 11346 13030 11398 13082
rect 11410 13030 11462 13082
rect 11474 13030 11526 13082
rect 11538 13030 11590 13082
rect 11602 13030 11654 13082
rect 16544 13030 16596 13082
rect 16608 13030 16660 13082
rect 16672 13030 16724 13082
rect 16736 13030 16788 13082
rect 16800 13030 16852 13082
rect 21742 13030 21794 13082
rect 21806 13030 21858 13082
rect 21870 13030 21922 13082
rect 21934 13030 21986 13082
rect 21998 13030 22050 13082
rect 1492 12971 1544 12980
rect 1492 12937 1501 12971
rect 1501 12937 1535 12971
rect 1535 12937 1544 12971
rect 1492 12928 1544 12937
rect 3056 12928 3108 12980
rect 2504 12903 2556 12912
rect 2504 12869 2513 12903
rect 2513 12869 2547 12903
rect 2547 12869 2556 12903
rect 2504 12860 2556 12869
rect 4068 12860 4120 12912
rect 6920 12928 6972 12980
rect 7840 12971 7892 12980
rect 7840 12937 7849 12971
rect 7849 12937 7883 12971
rect 7883 12937 7892 12971
rect 7840 12928 7892 12937
rect 8208 12971 8260 12980
rect 8208 12937 8217 12971
rect 8217 12937 8251 12971
rect 8251 12937 8260 12971
rect 8208 12928 8260 12937
rect 8760 12860 8812 12912
rect 8852 12860 8904 12912
rect 9404 12928 9456 12980
rect 10600 12928 10652 12980
rect 10784 12971 10836 12980
rect 10784 12937 10793 12971
rect 10793 12937 10827 12971
rect 10827 12937 10836 12971
rect 10784 12928 10836 12937
rect 11060 12971 11112 12980
rect 11060 12937 11069 12971
rect 11069 12937 11103 12971
rect 11103 12937 11112 12971
rect 11060 12928 11112 12937
rect 12072 12928 12124 12980
rect 14096 12971 14148 12980
rect 14096 12937 14105 12971
rect 14105 12937 14139 12971
rect 14139 12937 14148 12971
rect 14096 12928 14148 12937
rect 15660 12928 15712 12980
rect 1676 12835 1728 12844
rect 1676 12801 1685 12835
rect 1685 12801 1719 12835
rect 1719 12801 1728 12835
rect 1676 12792 1728 12801
rect 1952 12835 2004 12844
rect 1952 12801 1961 12835
rect 1961 12801 1995 12835
rect 1995 12801 2004 12835
rect 1952 12792 2004 12801
rect 2596 12792 2648 12844
rect 4252 12792 4304 12844
rect 1768 12724 1820 12776
rect 388 12656 440 12708
rect 1492 12656 1544 12708
rect 3976 12656 4028 12708
rect 5172 12767 5224 12776
rect 5172 12733 5181 12767
rect 5181 12733 5215 12767
rect 5215 12733 5224 12767
rect 6460 12792 6512 12844
rect 6920 12792 6972 12844
rect 5908 12767 5960 12776
rect 5172 12724 5224 12733
rect 5908 12733 5917 12767
rect 5917 12733 5951 12767
rect 5951 12733 5960 12767
rect 5908 12724 5960 12733
rect 6184 12656 6236 12708
rect 7472 12792 7524 12844
rect 8668 12792 8720 12844
rect 9772 12860 9824 12912
rect 10232 12860 10284 12912
rect 13268 12903 13320 12912
rect 8392 12767 8444 12776
rect 8392 12733 8401 12767
rect 8401 12733 8435 12767
rect 8435 12733 8444 12767
rect 8392 12724 8444 12733
rect 8576 12724 8628 12776
rect 10048 12792 10100 12844
rect 8944 12767 8996 12776
rect 8944 12733 8953 12767
rect 8953 12733 8987 12767
rect 8987 12733 8996 12767
rect 8944 12724 8996 12733
rect 2504 12588 2556 12640
rect 6368 12588 6420 12640
rect 7564 12588 7616 12640
rect 8484 12656 8536 12708
rect 9772 12656 9824 12708
rect 9404 12588 9456 12640
rect 10508 12724 10560 12776
rect 10600 12699 10652 12708
rect 10600 12665 10609 12699
rect 10609 12665 10643 12699
rect 10643 12665 10652 12699
rect 10600 12656 10652 12665
rect 11244 12792 11296 12844
rect 11796 12835 11848 12844
rect 11796 12801 11830 12835
rect 11830 12801 11848 12835
rect 13268 12869 13277 12903
rect 13277 12869 13311 12903
rect 13311 12869 13320 12903
rect 13268 12860 13320 12869
rect 13452 12860 13504 12912
rect 11796 12792 11848 12801
rect 13176 12792 13228 12844
rect 13084 12767 13136 12776
rect 13084 12733 13093 12767
rect 13093 12733 13127 12767
rect 13127 12733 13136 12767
rect 13084 12724 13136 12733
rect 13728 12724 13780 12776
rect 15292 12860 15344 12912
rect 16948 12928 17000 12980
rect 18052 12928 18104 12980
rect 19892 12971 19944 12980
rect 19892 12937 19901 12971
rect 19901 12937 19935 12971
rect 19935 12937 19944 12971
rect 19892 12928 19944 12937
rect 21272 12928 21324 12980
rect 16488 12860 16540 12912
rect 14372 12835 14424 12844
rect 14372 12801 14381 12835
rect 14381 12801 14415 12835
rect 14415 12801 14424 12835
rect 14372 12792 14424 12801
rect 14280 12724 14332 12776
rect 15200 12792 15252 12844
rect 15476 12792 15528 12844
rect 15660 12835 15712 12844
rect 15660 12801 15669 12835
rect 15669 12801 15703 12835
rect 15703 12801 15712 12835
rect 15660 12792 15712 12801
rect 10508 12631 10560 12640
rect 10508 12597 10517 12631
rect 10517 12597 10551 12631
rect 10551 12597 10560 12631
rect 10508 12588 10560 12597
rect 11060 12588 11112 12640
rect 14924 12767 14976 12776
rect 14924 12733 14933 12767
rect 14933 12733 14967 12767
rect 14967 12733 14976 12767
rect 14924 12724 14976 12733
rect 15568 12724 15620 12776
rect 16856 12792 16908 12844
rect 18328 12860 18380 12912
rect 20260 12860 20312 12912
rect 21180 12860 21232 12912
rect 21272 12835 21324 12844
rect 15660 12656 15712 12708
rect 13544 12588 13596 12640
rect 13728 12631 13780 12640
rect 13728 12597 13737 12631
rect 13737 12597 13771 12631
rect 13771 12597 13780 12631
rect 13728 12588 13780 12597
rect 13820 12588 13872 12640
rect 14004 12588 14056 12640
rect 14832 12588 14884 12640
rect 15936 12588 15988 12640
rect 16948 12588 17000 12640
rect 18420 12724 18472 12776
rect 18788 12767 18840 12776
rect 18788 12733 18797 12767
rect 18797 12733 18831 12767
rect 18831 12733 18840 12767
rect 18788 12724 18840 12733
rect 19432 12767 19484 12776
rect 19432 12733 19441 12767
rect 19441 12733 19475 12767
rect 19475 12733 19484 12767
rect 19432 12724 19484 12733
rect 18236 12656 18288 12708
rect 19616 12724 19668 12776
rect 21272 12801 21281 12835
rect 21281 12801 21315 12835
rect 21315 12801 21324 12835
rect 21272 12792 21324 12801
rect 18328 12588 18380 12640
rect 19432 12588 19484 12640
rect 20352 12588 20404 12640
rect 20720 12588 20772 12640
rect 20904 12588 20956 12640
rect 21456 12631 21508 12640
rect 21456 12597 21465 12631
rect 21465 12597 21499 12631
rect 21499 12597 21508 12631
rect 21456 12588 21508 12597
rect 3549 12486 3601 12538
rect 3613 12486 3665 12538
rect 3677 12486 3729 12538
rect 3741 12486 3793 12538
rect 3805 12486 3857 12538
rect 8747 12486 8799 12538
rect 8811 12486 8863 12538
rect 8875 12486 8927 12538
rect 8939 12486 8991 12538
rect 9003 12486 9055 12538
rect 13945 12486 13997 12538
rect 14009 12486 14061 12538
rect 14073 12486 14125 12538
rect 14137 12486 14189 12538
rect 14201 12486 14253 12538
rect 19143 12486 19195 12538
rect 19207 12486 19259 12538
rect 19271 12486 19323 12538
rect 19335 12486 19387 12538
rect 19399 12486 19451 12538
rect 1584 12427 1636 12436
rect 1584 12393 1593 12427
rect 1593 12393 1627 12427
rect 1627 12393 1636 12427
rect 1584 12384 1636 12393
rect 1676 12384 1728 12436
rect 3240 12384 3292 12436
rect 5172 12384 5224 12436
rect 2872 12316 2924 12368
rect 3976 12316 4028 12368
rect 9220 12384 9272 12436
rect 9496 12384 9548 12436
rect 10048 12427 10100 12436
rect 10048 12393 10057 12427
rect 10057 12393 10091 12427
rect 10091 12393 10100 12427
rect 10048 12384 10100 12393
rect 12808 12384 12860 12436
rect 4252 12248 4304 12300
rect 7196 12316 7248 12368
rect 7564 12316 7616 12368
rect 7840 12316 7892 12368
rect 13820 12384 13872 12436
rect 14832 12384 14884 12436
rect 14924 12384 14976 12436
rect 16856 12427 16908 12436
rect 16856 12393 16865 12427
rect 16865 12393 16899 12427
rect 16899 12393 16908 12427
rect 16856 12384 16908 12393
rect 16948 12384 17000 12436
rect 17592 12384 17644 12436
rect 18328 12384 18380 12436
rect 18696 12427 18748 12436
rect 18696 12393 18705 12427
rect 18705 12393 18739 12427
rect 18739 12393 18748 12427
rect 18696 12384 18748 12393
rect 1768 12180 1820 12232
rect 1952 12223 2004 12232
rect 1952 12189 1986 12223
rect 1986 12189 2004 12223
rect 1952 12180 2004 12189
rect 3332 12223 3384 12232
rect 3332 12189 3341 12223
rect 3341 12189 3375 12223
rect 3375 12189 3384 12223
rect 3332 12180 3384 12189
rect 3792 12180 3844 12232
rect 4804 12180 4856 12232
rect 5540 12180 5592 12232
rect 6368 12248 6420 12300
rect 6460 12248 6512 12300
rect 7288 12248 7340 12300
rect 7748 12248 7800 12300
rect 7932 12248 7984 12300
rect 8392 12291 8444 12300
rect 8392 12257 8401 12291
rect 8401 12257 8435 12291
rect 8435 12257 8444 12291
rect 8392 12248 8444 12257
rect 9404 12291 9456 12300
rect 9404 12257 9413 12291
rect 9413 12257 9447 12291
rect 9447 12257 9456 12291
rect 9404 12248 9456 12257
rect 9496 12291 9548 12300
rect 9496 12257 9505 12291
rect 9505 12257 9539 12291
rect 9539 12257 9548 12291
rect 9496 12248 9548 12257
rect 6552 12180 6604 12232
rect 8668 12223 8720 12232
rect 3056 12087 3108 12096
rect 3056 12053 3065 12087
rect 3065 12053 3099 12087
rect 3099 12053 3108 12087
rect 3056 12044 3108 12053
rect 3976 12087 4028 12096
rect 3976 12053 3985 12087
rect 3985 12053 4019 12087
rect 4019 12053 4028 12087
rect 3976 12044 4028 12053
rect 5632 12112 5684 12164
rect 6184 12112 6236 12164
rect 8668 12189 8677 12223
rect 8677 12189 8711 12223
rect 8711 12189 8720 12223
rect 8668 12180 8720 12189
rect 9956 12223 10008 12232
rect 9956 12189 9965 12223
rect 9965 12189 9999 12223
rect 9999 12189 10008 12223
rect 11060 12223 11112 12232
rect 9956 12180 10008 12189
rect 11060 12189 11069 12223
rect 11069 12189 11103 12223
rect 11103 12189 11112 12223
rect 11060 12180 11112 12189
rect 11796 12180 11848 12232
rect 13084 12248 13136 12300
rect 17776 12316 17828 12368
rect 21272 12316 21324 12368
rect 12808 12180 12860 12232
rect 13360 12180 13412 12232
rect 13636 12180 13688 12232
rect 6644 12087 6696 12096
rect 6644 12053 6653 12087
rect 6653 12053 6687 12087
rect 6687 12053 6696 12087
rect 6644 12044 6696 12053
rect 6736 12087 6788 12096
rect 6736 12053 6745 12087
rect 6745 12053 6779 12087
rect 6779 12053 6788 12087
rect 6736 12044 6788 12053
rect 7012 12044 7064 12096
rect 7380 12087 7432 12096
rect 7380 12053 7389 12087
rect 7389 12053 7423 12087
rect 7423 12053 7432 12087
rect 7380 12044 7432 12053
rect 7472 12044 7524 12096
rect 7840 12044 7892 12096
rect 8024 12044 8076 12096
rect 8208 12044 8260 12096
rect 8392 12044 8444 12096
rect 10600 12112 10652 12164
rect 11612 12112 11664 12164
rect 14740 12291 14792 12300
rect 14740 12257 14749 12291
rect 14749 12257 14783 12291
rect 14783 12257 14792 12291
rect 14740 12248 14792 12257
rect 15200 12248 15252 12300
rect 15476 12291 15528 12300
rect 15476 12257 15485 12291
rect 15485 12257 15519 12291
rect 15519 12257 15528 12291
rect 15476 12248 15528 12257
rect 18236 12248 18288 12300
rect 13820 12180 13872 12232
rect 9312 12087 9364 12096
rect 9312 12053 9321 12087
rect 9321 12053 9355 12087
rect 9355 12053 9364 12087
rect 9312 12044 9364 12053
rect 9404 12044 9456 12096
rect 10140 12044 10192 12096
rect 10692 12087 10744 12096
rect 10692 12053 10701 12087
rect 10701 12053 10735 12087
rect 10735 12053 10744 12087
rect 10692 12044 10744 12053
rect 12348 12044 12400 12096
rect 13452 12087 13504 12096
rect 13452 12053 13461 12087
rect 13461 12053 13495 12087
rect 13495 12053 13504 12087
rect 13452 12044 13504 12053
rect 13912 12087 13964 12096
rect 13912 12053 13921 12087
rect 13921 12053 13955 12087
rect 13955 12053 13964 12087
rect 13912 12044 13964 12053
rect 14556 12044 14608 12096
rect 15016 12087 15068 12096
rect 15016 12053 15025 12087
rect 15025 12053 15059 12087
rect 15059 12053 15068 12087
rect 16212 12112 16264 12164
rect 17316 12112 17368 12164
rect 17592 12180 17644 12232
rect 18604 12180 18656 12232
rect 20904 12248 20956 12300
rect 19800 12180 19852 12232
rect 20996 12180 21048 12232
rect 18052 12112 18104 12164
rect 18972 12112 19024 12164
rect 20720 12112 20772 12164
rect 21088 12155 21140 12164
rect 21088 12121 21097 12155
rect 21097 12121 21131 12155
rect 21131 12121 21140 12155
rect 21088 12112 21140 12121
rect 15016 12044 15068 12053
rect 15844 12044 15896 12096
rect 18144 12044 18196 12096
rect 18880 12044 18932 12096
rect 19340 12044 19392 12096
rect 21456 12087 21508 12096
rect 21456 12053 21465 12087
rect 21465 12053 21499 12087
rect 21499 12053 21508 12087
rect 21456 12044 21508 12053
rect 21732 12044 21784 12096
rect 22744 12044 22796 12096
rect 6148 11942 6200 11994
rect 6212 11942 6264 11994
rect 6276 11942 6328 11994
rect 6340 11942 6392 11994
rect 6404 11942 6456 11994
rect 11346 11942 11398 11994
rect 11410 11942 11462 11994
rect 11474 11942 11526 11994
rect 11538 11942 11590 11994
rect 11602 11942 11654 11994
rect 16544 11942 16596 11994
rect 16608 11942 16660 11994
rect 16672 11942 16724 11994
rect 16736 11942 16788 11994
rect 16800 11942 16852 11994
rect 21742 11942 21794 11994
rect 21806 11942 21858 11994
rect 21870 11942 21922 11994
rect 21934 11942 21986 11994
rect 21998 11942 22050 11994
rect 1860 11840 1912 11892
rect 2504 11840 2556 11892
rect 2964 11840 3016 11892
rect 3424 11840 3476 11892
rect 3976 11840 4028 11892
rect 4344 11883 4396 11892
rect 4344 11849 4353 11883
rect 4353 11849 4387 11883
rect 4387 11849 4396 11883
rect 4344 11840 4396 11849
rect 7380 11840 7432 11892
rect 7840 11840 7892 11892
rect 8024 11840 8076 11892
rect 1952 11747 2004 11756
rect 1952 11713 1961 11747
rect 1961 11713 1995 11747
rect 1995 11713 2004 11747
rect 1952 11704 2004 11713
rect 2228 11747 2280 11756
rect 2228 11713 2237 11747
rect 2237 11713 2271 11747
rect 2271 11713 2280 11747
rect 2228 11704 2280 11713
rect 2688 11747 2740 11756
rect 2688 11713 2697 11747
rect 2697 11713 2731 11747
rect 2731 11713 2740 11747
rect 2688 11704 2740 11713
rect 2780 11704 2832 11756
rect 2504 11679 2556 11688
rect 2504 11645 2513 11679
rect 2513 11645 2547 11679
rect 2547 11645 2556 11679
rect 2504 11636 2556 11645
rect 2596 11679 2648 11688
rect 2596 11645 2605 11679
rect 2605 11645 2639 11679
rect 2639 11645 2648 11679
rect 3884 11679 3936 11688
rect 2596 11636 2648 11645
rect 3884 11645 3893 11679
rect 3893 11645 3927 11679
rect 3927 11645 3936 11679
rect 3884 11636 3936 11645
rect 3976 11636 4028 11688
rect 6552 11772 6604 11824
rect 8300 11840 8352 11892
rect 8668 11840 8720 11892
rect 11612 11840 11664 11892
rect 11796 11840 11848 11892
rect 12256 11840 12308 11892
rect 12716 11883 12768 11892
rect 12716 11849 12725 11883
rect 12725 11849 12759 11883
rect 12759 11849 12768 11883
rect 12716 11840 12768 11849
rect 13268 11840 13320 11892
rect 13452 11840 13504 11892
rect 14096 11840 14148 11892
rect 15108 11840 15160 11892
rect 15200 11840 15252 11892
rect 15936 11840 15988 11892
rect 16396 11840 16448 11892
rect 16948 11883 17000 11892
rect 16948 11849 16957 11883
rect 16957 11849 16991 11883
rect 16991 11849 17000 11883
rect 16948 11840 17000 11849
rect 18052 11883 18104 11892
rect 18052 11849 18061 11883
rect 18061 11849 18095 11883
rect 18095 11849 18104 11883
rect 18052 11840 18104 11849
rect 18328 11840 18380 11892
rect 18696 11840 18748 11892
rect 21272 11840 21324 11892
rect 5816 11747 5868 11756
rect 5816 11713 5825 11747
rect 5825 11713 5859 11747
rect 5859 11713 5868 11747
rect 5816 11704 5868 11713
rect 7012 11704 7064 11756
rect 8852 11704 8904 11756
rect 9128 11704 9180 11756
rect 11704 11772 11756 11824
rect 12348 11772 12400 11824
rect 12716 11704 12768 11756
rect 5632 11679 5684 11688
rect 5632 11645 5641 11679
rect 5641 11645 5675 11679
rect 5675 11645 5684 11679
rect 5632 11636 5684 11645
rect 5724 11636 5776 11688
rect 3424 11568 3476 11620
rect 6736 11568 6788 11620
rect 7196 11636 7248 11688
rect 8024 11636 8076 11688
rect 9956 11679 10008 11688
rect 7840 11568 7892 11620
rect 9956 11645 9965 11679
rect 9965 11645 9999 11679
rect 9999 11645 10008 11679
rect 9956 11636 10008 11645
rect 11704 11679 11756 11688
rect 11704 11645 11713 11679
rect 11713 11645 11747 11679
rect 11747 11645 11756 11679
rect 11704 11636 11756 11645
rect 11796 11679 11848 11688
rect 11796 11645 11805 11679
rect 11805 11645 11839 11679
rect 11839 11645 11848 11679
rect 11796 11636 11848 11645
rect 12072 11636 12124 11688
rect 13728 11772 13780 11824
rect 13912 11772 13964 11824
rect 17776 11772 17828 11824
rect 13176 11704 13228 11756
rect 15568 11704 15620 11756
rect 16120 11704 16172 11756
rect 17224 11704 17276 11756
rect 17500 11704 17552 11756
rect 18328 11747 18380 11756
rect 18328 11713 18337 11747
rect 18337 11713 18371 11747
rect 18371 11713 18380 11747
rect 18788 11747 18840 11756
rect 18328 11704 18380 11713
rect 18788 11713 18797 11747
rect 18797 11713 18831 11747
rect 18831 11713 18840 11747
rect 18788 11704 18840 11713
rect 19248 11772 19300 11824
rect 19524 11772 19576 11824
rect 19800 11772 19852 11824
rect 21088 11772 21140 11824
rect 20444 11704 20496 11756
rect 20720 11747 20772 11756
rect 20720 11713 20729 11747
rect 20729 11713 20763 11747
rect 20763 11713 20772 11747
rect 20720 11704 20772 11713
rect 20812 11704 20864 11756
rect 22468 11704 22520 11756
rect 3148 11500 3200 11552
rect 3792 11500 3844 11552
rect 3884 11500 3936 11552
rect 4528 11500 4580 11552
rect 4804 11543 4856 11552
rect 4804 11509 4813 11543
rect 4813 11509 4847 11543
rect 4847 11509 4856 11543
rect 4804 11500 4856 11509
rect 5080 11543 5132 11552
rect 5080 11509 5089 11543
rect 5089 11509 5123 11543
rect 5123 11509 5132 11543
rect 5080 11500 5132 11509
rect 7012 11500 7064 11552
rect 8208 11500 8260 11552
rect 8852 11500 8904 11552
rect 9220 11500 9272 11552
rect 14556 11636 14608 11688
rect 15660 11679 15712 11688
rect 15660 11645 15669 11679
rect 15669 11645 15703 11679
rect 15703 11645 15712 11679
rect 15660 11636 15712 11645
rect 11796 11500 11848 11552
rect 12348 11543 12400 11552
rect 12348 11509 12357 11543
rect 12357 11509 12391 11543
rect 12391 11509 12400 11543
rect 12348 11500 12400 11509
rect 14372 11568 14424 11620
rect 12808 11500 12860 11552
rect 13360 11500 13412 11552
rect 13728 11500 13780 11552
rect 14832 11500 14884 11552
rect 15200 11543 15252 11552
rect 15200 11509 15209 11543
rect 15209 11509 15243 11543
rect 15243 11509 15252 11543
rect 15200 11500 15252 11509
rect 15476 11500 15528 11552
rect 16948 11568 17000 11620
rect 18052 11568 18104 11620
rect 19156 11636 19208 11688
rect 20904 11568 20956 11620
rect 16396 11543 16448 11552
rect 16396 11509 16405 11543
rect 16405 11509 16439 11543
rect 16439 11509 16448 11543
rect 16396 11500 16448 11509
rect 17040 11543 17092 11552
rect 17040 11509 17049 11543
rect 17049 11509 17083 11543
rect 17083 11509 17092 11543
rect 17040 11500 17092 11509
rect 17316 11543 17368 11552
rect 17316 11509 17325 11543
rect 17325 11509 17359 11543
rect 17359 11509 17368 11543
rect 17316 11500 17368 11509
rect 17776 11500 17828 11552
rect 18236 11500 18288 11552
rect 19524 11500 19576 11552
rect 20076 11500 20128 11552
rect 20536 11500 20588 11552
rect 3549 11398 3601 11450
rect 3613 11398 3665 11450
rect 3677 11398 3729 11450
rect 3741 11398 3793 11450
rect 3805 11398 3857 11450
rect 8747 11398 8799 11450
rect 8811 11398 8863 11450
rect 8875 11398 8927 11450
rect 8939 11398 8991 11450
rect 9003 11398 9055 11450
rect 13945 11398 13997 11450
rect 14009 11398 14061 11450
rect 14073 11398 14125 11450
rect 14137 11398 14189 11450
rect 14201 11398 14253 11450
rect 19143 11398 19195 11450
rect 19207 11398 19259 11450
rect 19271 11398 19323 11450
rect 19335 11398 19387 11450
rect 19399 11398 19451 11450
rect 1492 11339 1544 11348
rect 1492 11305 1501 11339
rect 1501 11305 1535 11339
rect 1535 11305 1544 11339
rect 1492 11296 1544 11305
rect 2320 11296 2372 11348
rect 5632 11339 5684 11348
rect 2044 11271 2096 11280
rect 2044 11237 2053 11271
rect 2053 11237 2087 11271
rect 2087 11237 2096 11271
rect 2044 11228 2096 11237
rect 3148 11228 3200 11280
rect 2504 11203 2556 11212
rect 2504 11169 2513 11203
rect 2513 11169 2547 11203
rect 2547 11169 2556 11203
rect 2504 11160 2556 11169
rect 1676 11135 1728 11144
rect 1676 11101 1685 11135
rect 1685 11101 1719 11135
rect 1719 11101 1728 11135
rect 1676 11092 1728 11101
rect 1860 11135 1912 11144
rect 1860 11101 1869 11135
rect 1869 11101 1903 11135
rect 1903 11101 1912 11135
rect 1860 11092 1912 11101
rect 2964 11135 3016 11144
rect 2964 11101 2973 11135
rect 2973 11101 3007 11135
rect 3007 11101 3016 11135
rect 2964 11092 3016 11101
rect 3332 11271 3384 11280
rect 3332 11237 3341 11271
rect 3341 11237 3375 11271
rect 3375 11237 3384 11271
rect 5632 11305 5641 11339
rect 5641 11305 5675 11339
rect 5675 11305 5684 11339
rect 5632 11296 5684 11305
rect 6644 11296 6696 11348
rect 6736 11296 6788 11348
rect 10600 11296 10652 11348
rect 12072 11296 12124 11348
rect 3332 11228 3384 11237
rect 4252 11228 4304 11280
rect 5540 11160 5592 11212
rect 8392 11228 8444 11280
rect 8668 11271 8720 11280
rect 8668 11237 8677 11271
rect 8677 11237 8711 11271
rect 8711 11237 8720 11271
rect 8668 11228 8720 11237
rect 8944 11228 8996 11280
rect 9128 11228 9180 11280
rect 10876 11228 10928 11280
rect 11980 11228 12032 11280
rect 7196 11203 7248 11212
rect 7196 11169 7205 11203
rect 7205 11169 7239 11203
rect 7239 11169 7248 11203
rect 8024 11203 8076 11212
rect 7196 11160 7248 11169
rect 8024 11169 8033 11203
rect 8033 11169 8067 11203
rect 8067 11169 8076 11203
rect 8024 11160 8076 11169
rect 9404 11160 9456 11212
rect 11060 11160 11112 11212
rect 11612 11160 11664 11212
rect 13268 11296 13320 11348
rect 15568 11296 15620 11348
rect 13360 11203 13412 11212
rect 13360 11169 13369 11203
rect 13369 11169 13403 11203
rect 13403 11169 13412 11203
rect 13360 11160 13412 11169
rect 13544 11203 13596 11212
rect 13544 11169 13553 11203
rect 13553 11169 13587 11203
rect 13587 11169 13596 11203
rect 13544 11160 13596 11169
rect 14280 11203 14332 11212
rect 14280 11169 14289 11203
rect 14289 11169 14323 11203
rect 14323 11169 14332 11203
rect 14280 11160 14332 11169
rect 16856 11228 16908 11280
rect 19892 11296 19944 11348
rect 19248 11228 19300 11280
rect 2872 11024 2924 11076
rect 5356 11092 5408 11144
rect 6552 11092 6604 11144
rect 7932 11135 7984 11144
rect 7932 11101 7941 11135
rect 7941 11101 7975 11135
rect 7975 11101 7984 11135
rect 7932 11092 7984 11101
rect 5540 11024 5592 11076
rect 5816 11024 5868 11076
rect 7840 11067 7892 11076
rect 3332 10956 3384 11008
rect 3700 10956 3752 11008
rect 3976 10999 4028 11008
rect 3976 10965 3985 10999
rect 3985 10965 4019 10999
rect 4019 10965 4028 10999
rect 3976 10956 4028 10965
rect 6000 10999 6052 11008
rect 6000 10965 6009 10999
rect 6009 10965 6043 10999
rect 6043 10965 6052 10999
rect 6000 10956 6052 10965
rect 7840 11033 7849 11067
rect 7849 11033 7883 11067
rect 7883 11033 7892 11067
rect 7840 11024 7892 11033
rect 10140 11135 10192 11144
rect 10140 11101 10158 11135
rect 10158 11101 10192 11135
rect 10140 11092 10192 11101
rect 10508 11092 10560 11144
rect 11520 11135 11572 11144
rect 11520 11101 11529 11135
rect 11529 11101 11563 11135
rect 11563 11101 11572 11135
rect 11520 11092 11572 11101
rect 11796 11092 11848 11144
rect 8208 11024 8260 11076
rect 6920 10956 6972 11008
rect 7932 10956 7984 11008
rect 8300 10956 8352 11008
rect 8668 10956 8720 11008
rect 9588 11024 9640 11076
rect 10692 11024 10744 11076
rect 12164 11024 12216 11076
rect 12808 11092 12860 11144
rect 13452 11092 13504 11144
rect 13820 11024 13872 11076
rect 15844 11092 15896 11144
rect 16948 11160 17000 11212
rect 17224 11203 17276 11212
rect 17224 11169 17233 11203
rect 17233 11169 17267 11203
rect 17267 11169 17276 11203
rect 17224 11160 17276 11169
rect 21272 11203 21324 11212
rect 9680 10956 9732 11008
rect 11980 10999 12032 11008
rect 11980 10965 11989 10999
rect 11989 10965 12023 10999
rect 12023 10965 12032 10999
rect 11980 10956 12032 10965
rect 12348 10999 12400 11008
rect 12348 10965 12357 10999
rect 12357 10965 12391 10999
rect 12391 10965 12400 10999
rect 12348 10956 12400 10965
rect 12808 10999 12860 11008
rect 12808 10965 12817 10999
rect 12817 10965 12851 10999
rect 12851 10965 12860 10999
rect 12808 10956 12860 10965
rect 12900 10999 12952 11008
rect 12900 10965 12909 10999
rect 12909 10965 12943 10999
rect 12943 10965 12952 10999
rect 13268 10999 13320 11008
rect 12900 10956 12952 10965
rect 13268 10965 13277 10999
rect 13277 10965 13311 10999
rect 13311 10965 13320 10999
rect 13268 10956 13320 10965
rect 13360 10956 13412 11008
rect 14648 11024 14700 11076
rect 15292 11024 15344 11076
rect 16212 11024 16264 11076
rect 21272 11169 21281 11203
rect 21281 11169 21315 11203
rect 21315 11169 21324 11203
rect 21272 11160 21324 11169
rect 15844 10956 15896 11008
rect 16948 10999 17000 11008
rect 16948 10965 16957 10999
rect 16957 10965 16991 10999
rect 16991 10965 17000 10999
rect 16948 10956 17000 10965
rect 19156 11092 19208 11144
rect 20904 11092 20956 11144
rect 18696 11024 18748 11076
rect 19892 11024 19944 11076
rect 21088 11067 21140 11076
rect 21088 11033 21097 11067
rect 21097 11033 21131 11067
rect 21131 11033 21140 11067
rect 21088 11024 21140 11033
rect 21364 11024 21416 11076
rect 18052 10956 18104 11008
rect 18604 10956 18656 11008
rect 19800 10956 19852 11008
rect 20812 10956 20864 11008
rect 6148 10854 6200 10906
rect 6212 10854 6264 10906
rect 6276 10854 6328 10906
rect 6340 10854 6392 10906
rect 6404 10854 6456 10906
rect 11346 10854 11398 10906
rect 11410 10854 11462 10906
rect 11474 10854 11526 10906
rect 11538 10854 11590 10906
rect 11602 10854 11654 10906
rect 16544 10854 16596 10906
rect 16608 10854 16660 10906
rect 16672 10854 16724 10906
rect 16736 10854 16788 10906
rect 16800 10854 16852 10906
rect 21742 10854 21794 10906
rect 21806 10854 21858 10906
rect 21870 10854 21922 10906
rect 21934 10854 21986 10906
rect 21998 10854 22050 10906
rect 2964 10752 3016 10804
rect 1492 10659 1544 10668
rect 1492 10625 1501 10659
rect 1501 10625 1535 10659
rect 1535 10625 1544 10659
rect 1492 10616 1544 10625
rect 1860 10616 1912 10668
rect 2044 10659 2096 10668
rect 2044 10625 2078 10659
rect 2078 10625 2096 10659
rect 2044 10616 2096 10625
rect 3976 10616 4028 10668
rect 1768 10591 1820 10600
rect 1768 10557 1777 10591
rect 1777 10557 1811 10591
rect 1811 10557 1820 10591
rect 1768 10548 1820 10557
rect 4804 10591 4856 10600
rect 4804 10557 4813 10591
rect 4813 10557 4847 10591
rect 4847 10557 4856 10591
rect 4804 10548 4856 10557
rect 5724 10684 5776 10736
rect 6000 10752 6052 10804
rect 6552 10752 6604 10804
rect 7104 10752 7156 10804
rect 9680 10795 9732 10804
rect 7840 10684 7892 10736
rect 5816 10659 5868 10668
rect 5816 10625 5825 10659
rect 5825 10625 5859 10659
rect 5859 10625 5868 10659
rect 5816 10616 5868 10625
rect 5540 10591 5592 10600
rect 5540 10557 5549 10591
rect 5549 10557 5583 10591
rect 5583 10557 5592 10591
rect 5540 10548 5592 10557
rect 6368 10548 6420 10600
rect 8024 10616 8076 10668
rect 8300 10684 8352 10736
rect 9680 10761 9689 10795
rect 9689 10761 9723 10795
rect 9723 10761 9732 10795
rect 9680 10752 9732 10761
rect 10692 10752 10744 10804
rect 11980 10752 12032 10804
rect 13268 10752 13320 10804
rect 13728 10752 13780 10804
rect 14464 10752 14516 10804
rect 7840 10548 7892 10600
rect 13544 10727 13596 10736
rect 13544 10693 13562 10727
rect 13562 10693 13596 10727
rect 13544 10684 13596 10693
rect 10876 10616 10928 10668
rect 11244 10659 11296 10668
rect 11244 10625 11253 10659
rect 11253 10625 11287 10659
rect 11287 10625 11296 10659
rect 11244 10616 11296 10625
rect 11980 10659 12032 10668
rect 11980 10625 11989 10659
rect 11989 10625 12023 10659
rect 12023 10625 12032 10659
rect 11980 10616 12032 10625
rect 14280 10684 14332 10736
rect 15292 10795 15344 10804
rect 15292 10761 15301 10795
rect 15301 10761 15335 10795
rect 15335 10761 15344 10795
rect 15292 10752 15344 10761
rect 16120 10795 16172 10804
rect 16120 10761 16129 10795
rect 16129 10761 16163 10795
rect 16163 10761 16172 10795
rect 16120 10752 16172 10761
rect 14188 10616 14240 10668
rect 14648 10684 14700 10736
rect 15108 10684 15160 10736
rect 16948 10752 17000 10804
rect 16764 10684 16816 10736
rect 17132 10727 17184 10736
rect 17132 10693 17141 10727
rect 17141 10693 17175 10727
rect 17175 10693 17184 10727
rect 17132 10684 17184 10693
rect 9680 10548 9732 10600
rect 9956 10548 10008 10600
rect 10140 10548 10192 10600
rect 10600 10591 10652 10600
rect 10600 10557 10609 10591
rect 10609 10557 10643 10591
rect 10643 10557 10652 10591
rect 10600 10548 10652 10557
rect 11704 10591 11756 10600
rect 11704 10557 11713 10591
rect 11713 10557 11747 10591
rect 11747 10557 11756 10591
rect 11704 10548 11756 10557
rect 14648 10591 14700 10600
rect 14648 10557 14657 10591
rect 14657 10557 14691 10591
rect 14691 10557 14700 10591
rect 14648 10548 14700 10557
rect 14832 10591 14884 10600
rect 14832 10557 14841 10591
rect 14841 10557 14875 10591
rect 14875 10557 14884 10591
rect 14832 10548 14884 10557
rect 15844 10616 15896 10668
rect 15660 10591 15712 10600
rect 15660 10557 15669 10591
rect 15669 10557 15703 10591
rect 15703 10557 15712 10591
rect 15660 10548 15712 10557
rect 17224 10591 17276 10600
rect 17224 10557 17233 10591
rect 17233 10557 17267 10591
rect 17267 10557 17276 10591
rect 17224 10548 17276 10557
rect 17868 10752 17920 10804
rect 18788 10752 18840 10804
rect 19616 10752 19668 10804
rect 17776 10684 17828 10736
rect 20720 10684 20772 10736
rect 21180 10684 21232 10736
rect 18328 10616 18380 10668
rect 18788 10616 18840 10668
rect 19524 10659 19576 10668
rect 19524 10625 19533 10659
rect 19533 10625 19567 10659
rect 19567 10625 19576 10659
rect 19524 10616 19576 10625
rect 20904 10616 20956 10668
rect 17776 10548 17828 10600
rect 18236 10548 18288 10600
rect 18512 10591 18564 10600
rect 18512 10557 18521 10591
rect 18521 10557 18555 10591
rect 18555 10557 18564 10591
rect 18512 10548 18564 10557
rect 19616 10591 19668 10600
rect 5172 10455 5224 10464
rect 5172 10421 5181 10455
rect 5181 10421 5215 10455
rect 5215 10421 5224 10455
rect 5172 10412 5224 10421
rect 5540 10412 5592 10464
rect 6552 10412 6604 10464
rect 7840 10455 7892 10464
rect 7840 10421 7849 10455
rect 7849 10421 7883 10455
rect 7883 10421 7892 10455
rect 13820 10480 13872 10532
rect 19616 10557 19625 10591
rect 19625 10557 19659 10591
rect 19659 10557 19668 10591
rect 19616 10548 19668 10557
rect 19800 10591 19852 10600
rect 19800 10557 19809 10591
rect 19809 10557 19843 10591
rect 19843 10557 19852 10591
rect 19800 10548 19852 10557
rect 7840 10412 7892 10421
rect 9496 10412 9548 10464
rect 12440 10455 12492 10464
rect 12440 10421 12449 10455
rect 12449 10421 12483 10455
rect 12483 10421 12492 10455
rect 12440 10412 12492 10421
rect 18144 10412 18196 10464
rect 18604 10412 18656 10464
rect 19708 10412 19760 10464
rect 3549 10310 3601 10362
rect 3613 10310 3665 10362
rect 3677 10310 3729 10362
rect 3741 10310 3793 10362
rect 3805 10310 3857 10362
rect 8747 10310 8799 10362
rect 8811 10310 8863 10362
rect 8875 10310 8927 10362
rect 8939 10310 8991 10362
rect 9003 10310 9055 10362
rect 13945 10310 13997 10362
rect 14009 10310 14061 10362
rect 14073 10310 14125 10362
rect 14137 10310 14189 10362
rect 14201 10310 14253 10362
rect 19143 10310 19195 10362
rect 19207 10310 19259 10362
rect 19271 10310 19323 10362
rect 19335 10310 19387 10362
rect 19399 10310 19451 10362
rect 756 10208 808 10260
rect 940 10208 992 10260
rect 2136 10208 2188 10260
rect 3608 10208 3660 10260
rect 4620 10208 4672 10260
rect 5356 10208 5408 10260
rect 6368 10251 6420 10260
rect 6368 10217 6377 10251
rect 6377 10217 6411 10251
rect 6411 10217 6420 10251
rect 6368 10208 6420 10217
rect 8208 10208 8260 10260
rect 10600 10208 10652 10260
rect 13820 10208 13872 10260
rect 1860 10140 1912 10192
rect 1768 10072 1820 10124
rect 572 10004 624 10056
rect 1032 10004 1084 10056
rect 1492 10047 1544 10056
rect 1492 10013 1501 10047
rect 1501 10013 1535 10047
rect 1535 10013 1544 10047
rect 1492 10004 1544 10013
rect 3240 10004 3292 10056
rect 2228 9979 2280 9988
rect 2228 9945 2262 9979
rect 2262 9945 2280 9979
rect 2228 9936 2280 9945
rect 2780 9936 2832 9988
rect 3056 9936 3108 9988
rect 1860 9911 1912 9920
rect 1860 9877 1869 9911
rect 1869 9877 1903 9911
rect 1903 9877 1912 9911
rect 1860 9868 1912 9877
rect 1952 9868 2004 9920
rect 4344 10140 4396 10192
rect 3516 10072 3568 10124
rect 3608 10047 3660 10056
rect 3608 10013 3617 10047
rect 3617 10013 3651 10047
rect 3651 10013 3660 10047
rect 3608 10004 3660 10013
rect 3884 10072 3936 10124
rect 5724 10140 5776 10192
rect 7104 10140 7156 10192
rect 7288 10140 7340 10192
rect 9956 10183 10008 10192
rect 5632 10072 5684 10124
rect 4804 10047 4856 10056
rect 4804 10013 4813 10047
rect 4813 10013 4847 10047
rect 4847 10013 4856 10047
rect 4804 10004 4856 10013
rect 5356 10004 5408 10056
rect 5908 10072 5960 10124
rect 6552 10115 6604 10124
rect 6552 10081 6561 10115
rect 6561 10081 6595 10115
rect 6595 10081 6604 10115
rect 6552 10072 6604 10081
rect 6920 10072 6972 10124
rect 7840 10072 7892 10124
rect 8300 10072 8352 10124
rect 8852 10072 8904 10124
rect 3608 9868 3660 9920
rect 4160 9868 4212 9920
rect 5540 9936 5592 9988
rect 5816 9936 5868 9988
rect 4712 9911 4764 9920
rect 4712 9877 4721 9911
rect 4721 9877 4755 9911
rect 4755 9877 4764 9911
rect 5632 9911 5684 9920
rect 4712 9868 4764 9877
rect 5632 9877 5641 9911
rect 5641 9877 5675 9911
rect 5675 9877 5684 9911
rect 5632 9868 5684 9877
rect 6460 10004 6512 10056
rect 6000 9936 6052 9988
rect 7840 9936 7892 9988
rect 6460 9868 6512 9920
rect 6644 9911 6696 9920
rect 6644 9877 6653 9911
rect 6653 9877 6687 9911
rect 6687 9877 6696 9911
rect 6644 9868 6696 9877
rect 6920 9911 6972 9920
rect 6920 9877 6929 9911
rect 6929 9877 6963 9911
rect 6963 9877 6972 9911
rect 6920 9868 6972 9877
rect 7472 9911 7524 9920
rect 7472 9877 7481 9911
rect 7481 9877 7515 9911
rect 7515 9877 7524 9911
rect 7472 9868 7524 9877
rect 7564 9911 7616 9920
rect 7564 9877 7573 9911
rect 7573 9877 7607 9911
rect 7607 9877 7616 9911
rect 8852 9936 8904 9988
rect 7564 9868 7616 9877
rect 8208 9868 8260 9920
rect 8668 9868 8720 9920
rect 8944 9911 8996 9920
rect 8944 9877 8953 9911
rect 8953 9877 8987 9911
rect 8987 9877 8996 9911
rect 8944 9868 8996 9877
rect 9128 9911 9180 9920
rect 9128 9877 9137 9911
rect 9137 9877 9171 9911
rect 9171 9877 9180 9911
rect 9128 9868 9180 9877
rect 9588 10072 9640 10124
rect 9496 10047 9548 10056
rect 9496 10013 9505 10047
rect 9505 10013 9539 10047
rect 9539 10013 9548 10047
rect 9496 10004 9548 10013
rect 9956 10149 9965 10183
rect 9965 10149 9999 10183
rect 9999 10149 10008 10183
rect 9956 10140 10008 10149
rect 14004 10140 14056 10192
rect 11704 10072 11756 10124
rect 12072 10115 12124 10124
rect 12072 10081 12081 10115
rect 12081 10081 12115 10115
rect 12115 10081 12124 10115
rect 12072 10072 12124 10081
rect 12440 10072 12492 10124
rect 12900 10072 12952 10124
rect 13268 10115 13320 10124
rect 13268 10081 13277 10115
rect 13277 10081 13311 10115
rect 13311 10081 13320 10115
rect 13268 10072 13320 10081
rect 14280 10208 14332 10260
rect 15660 10251 15712 10260
rect 15660 10217 15669 10251
rect 15669 10217 15703 10251
rect 15703 10217 15712 10251
rect 15660 10208 15712 10217
rect 15108 10140 15160 10192
rect 17224 10208 17276 10260
rect 18512 10208 18564 10260
rect 19616 10208 19668 10260
rect 16764 10183 16816 10192
rect 15660 10072 15712 10124
rect 16028 10072 16080 10124
rect 16764 10149 16773 10183
rect 16773 10149 16807 10183
rect 16807 10149 16816 10183
rect 16764 10140 16816 10149
rect 20904 10140 20956 10192
rect 12808 10047 12860 10056
rect 12808 10013 12817 10047
rect 12817 10013 12851 10047
rect 12851 10013 12860 10047
rect 12808 10004 12860 10013
rect 10784 9936 10836 9988
rect 11244 9936 11296 9988
rect 11520 9979 11572 9988
rect 11520 9945 11529 9979
rect 11529 9945 11563 9979
rect 11563 9945 11572 9979
rect 11520 9936 11572 9945
rect 11704 9936 11756 9988
rect 9772 9868 9824 9920
rect 9956 9868 10008 9920
rect 12072 9868 12124 9920
rect 13636 9936 13688 9988
rect 14556 9936 14608 9988
rect 16304 9936 16356 9988
rect 16948 10004 17000 10056
rect 19708 10115 19760 10124
rect 19708 10081 19717 10115
rect 19717 10081 19751 10115
rect 19751 10081 19760 10115
rect 19708 10072 19760 10081
rect 19800 10115 19852 10124
rect 19800 10081 19809 10115
rect 19809 10081 19843 10115
rect 19843 10081 19852 10115
rect 19800 10072 19852 10081
rect 18696 10047 18748 10056
rect 18696 10013 18705 10047
rect 18705 10013 18739 10047
rect 18739 10013 18748 10047
rect 18696 10004 18748 10013
rect 20812 10072 20864 10124
rect 21548 10072 21600 10124
rect 20720 10047 20772 10056
rect 20720 10013 20729 10047
rect 20729 10013 20763 10047
rect 20763 10013 20772 10047
rect 20720 10004 20772 10013
rect 20536 9936 20588 9988
rect 13728 9868 13780 9920
rect 16028 9911 16080 9920
rect 16028 9877 16037 9911
rect 16037 9877 16071 9911
rect 16071 9877 16080 9911
rect 16028 9868 16080 9877
rect 16120 9911 16172 9920
rect 16120 9877 16129 9911
rect 16129 9877 16163 9911
rect 16163 9877 16172 9911
rect 16120 9868 16172 9877
rect 16948 9868 17000 9920
rect 18052 9868 18104 9920
rect 18512 9868 18564 9920
rect 18696 9868 18748 9920
rect 18788 9868 18840 9920
rect 19892 9868 19944 9920
rect 20812 9868 20864 9920
rect 6148 9766 6200 9818
rect 6212 9766 6264 9818
rect 6276 9766 6328 9818
rect 6340 9766 6392 9818
rect 6404 9766 6456 9818
rect 11346 9766 11398 9818
rect 11410 9766 11462 9818
rect 11474 9766 11526 9818
rect 11538 9766 11590 9818
rect 11602 9766 11654 9818
rect 16544 9766 16596 9818
rect 16608 9766 16660 9818
rect 16672 9766 16724 9818
rect 16736 9766 16788 9818
rect 16800 9766 16852 9818
rect 21742 9766 21794 9818
rect 21806 9766 21858 9818
rect 21870 9766 21922 9818
rect 21934 9766 21986 9818
rect 21998 9766 22050 9818
rect 1860 9664 1912 9716
rect 3056 9664 3108 9716
rect 3240 9664 3292 9716
rect 7288 9664 7340 9716
rect 7472 9664 7524 9716
rect 8300 9664 8352 9716
rect 1492 9639 1544 9648
rect 1492 9605 1501 9639
rect 1501 9605 1535 9639
rect 1535 9605 1544 9639
rect 1492 9596 1544 9605
rect 3424 9596 3476 9648
rect 2320 9528 2372 9580
rect 2504 9528 2556 9580
rect 1952 9503 2004 9512
rect 1952 9469 1961 9503
rect 1961 9469 1995 9503
rect 1995 9469 2004 9503
rect 1952 9460 2004 9469
rect 2136 9503 2188 9512
rect 2136 9469 2145 9503
rect 2145 9469 2179 9503
rect 2179 9469 2188 9503
rect 2136 9460 2188 9469
rect 3608 9528 3660 9580
rect 3700 9528 3752 9580
rect 4160 9528 4212 9580
rect 4528 9528 4580 9580
rect 4712 9571 4764 9580
rect 4712 9537 4721 9571
rect 4721 9537 4755 9571
rect 4755 9537 4764 9571
rect 4712 9528 4764 9537
rect 5264 9528 5316 9580
rect 6184 9571 6236 9580
rect 6184 9537 6193 9571
rect 6193 9537 6227 9571
rect 6227 9537 6236 9571
rect 6184 9528 6236 9537
rect 1860 9392 1912 9444
rect 3056 9460 3108 9512
rect 4804 9503 4856 9512
rect 1492 9324 1544 9376
rect 2688 9392 2740 9444
rect 4068 9435 4120 9444
rect 2228 9324 2280 9376
rect 4068 9401 4077 9435
rect 4077 9401 4111 9435
rect 4111 9401 4120 9435
rect 4068 9392 4120 9401
rect 4804 9469 4813 9503
rect 4813 9469 4847 9503
rect 4847 9469 4856 9503
rect 4804 9460 4856 9469
rect 5632 9503 5684 9512
rect 5632 9469 5641 9503
rect 5641 9469 5675 9503
rect 5675 9469 5684 9503
rect 5632 9460 5684 9469
rect 7840 9596 7892 9648
rect 8208 9596 8260 9648
rect 6644 9571 6696 9580
rect 6644 9537 6653 9571
rect 6653 9537 6687 9571
rect 6687 9537 6696 9571
rect 6644 9528 6696 9537
rect 8392 9571 8444 9580
rect 7012 9503 7064 9512
rect 7012 9469 7021 9503
rect 7021 9469 7055 9503
rect 7055 9469 7064 9503
rect 7012 9460 7064 9469
rect 8024 9503 8076 9512
rect 8024 9469 8033 9503
rect 8033 9469 8067 9503
rect 8067 9469 8076 9503
rect 8024 9460 8076 9469
rect 8392 9537 8401 9571
rect 8401 9537 8435 9571
rect 8435 9537 8444 9571
rect 8392 9528 8444 9537
rect 8300 9460 8352 9512
rect 8659 9571 8711 9580
rect 8659 9537 8668 9571
rect 8668 9537 8702 9571
rect 8702 9537 8711 9571
rect 9128 9596 9180 9648
rect 10692 9664 10744 9716
rect 12532 9664 12584 9716
rect 13268 9664 13320 9716
rect 10232 9639 10284 9648
rect 10232 9605 10241 9639
rect 10241 9605 10275 9639
rect 10275 9605 10284 9639
rect 10876 9639 10928 9648
rect 10232 9596 10284 9605
rect 10876 9605 10885 9639
rect 10885 9605 10919 9639
rect 10919 9605 10928 9639
rect 10876 9596 10928 9605
rect 12992 9596 13044 9648
rect 13636 9596 13688 9648
rect 15384 9664 15436 9716
rect 15568 9596 15620 9648
rect 16304 9664 16356 9716
rect 18236 9664 18288 9716
rect 18328 9664 18380 9716
rect 16028 9596 16080 9648
rect 16212 9596 16264 9648
rect 8659 9528 8711 9537
rect 7564 9392 7616 9444
rect 7656 9392 7708 9444
rect 10140 9528 10192 9580
rect 10692 9571 10744 9580
rect 10692 9537 10701 9571
rect 10701 9537 10735 9571
rect 10735 9537 10744 9571
rect 10692 9528 10744 9537
rect 10416 9503 10468 9512
rect 10416 9469 10425 9503
rect 10425 9469 10459 9503
rect 10459 9469 10468 9503
rect 10416 9460 10468 9469
rect 10508 9460 10560 9512
rect 11336 9528 11388 9580
rect 11612 9528 11664 9580
rect 12440 9528 12492 9580
rect 13728 9528 13780 9580
rect 11060 9460 11112 9512
rect 11520 9460 11572 9512
rect 11704 9503 11756 9512
rect 11704 9469 11713 9503
rect 11713 9469 11747 9503
rect 11747 9469 11756 9503
rect 11704 9460 11756 9469
rect 12624 9503 12676 9512
rect 12624 9469 12633 9503
rect 12633 9469 12667 9503
rect 12667 9469 12676 9503
rect 12624 9460 12676 9469
rect 15476 9528 15528 9580
rect 15752 9571 15804 9580
rect 15752 9537 15761 9571
rect 15761 9537 15795 9571
rect 15795 9537 15804 9571
rect 15752 9528 15804 9537
rect 14924 9460 14976 9512
rect 16304 9528 16356 9580
rect 17132 9571 17184 9580
rect 17132 9537 17141 9571
rect 17141 9537 17175 9571
rect 17175 9537 17184 9571
rect 17132 9528 17184 9537
rect 17960 9571 18012 9580
rect 17960 9537 17969 9571
rect 17969 9537 18003 9571
rect 18003 9537 18012 9571
rect 17960 9528 18012 9537
rect 18788 9571 18840 9580
rect 18788 9537 18797 9571
rect 18797 9537 18831 9571
rect 18831 9537 18840 9571
rect 18788 9528 18840 9537
rect 19524 9664 19576 9716
rect 19800 9664 19852 9716
rect 20628 9664 20680 9716
rect 20996 9664 21048 9716
rect 21180 9664 21232 9716
rect 20720 9596 20772 9648
rect 20904 9596 20956 9648
rect 15292 9435 15344 9444
rect 15292 9401 15301 9435
rect 15301 9401 15335 9435
rect 15335 9401 15344 9435
rect 15292 9392 15344 9401
rect 16948 9503 17000 9512
rect 16948 9469 16957 9503
rect 16957 9469 16991 9503
rect 16991 9469 17000 9503
rect 16948 9460 17000 9469
rect 17408 9392 17460 9444
rect 17776 9460 17828 9512
rect 18052 9503 18104 9512
rect 18052 9469 18061 9503
rect 18061 9469 18095 9503
rect 18095 9469 18104 9503
rect 18052 9460 18104 9469
rect 18144 9503 18196 9512
rect 18144 9469 18153 9503
rect 18153 9469 18187 9503
rect 18187 9469 18196 9503
rect 18144 9460 18196 9469
rect 19616 9528 19668 9580
rect 20996 9571 21048 9580
rect 3792 9324 3844 9376
rect 4252 9324 4304 9376
rect 4436 9324 4488 9376
rect 5448 9324 5500 9376
rect 6460 9367 6512 9376
rect 6460 9333 6469 9367
rect 6469 9333 6503 9367
rect 6503 9333 6512 9367
rect 6460 9324 6512 9333
rect 6552 9324 6604 9376
rect 12808 9324 12860 9376
rect 12900 9324 12952 9376
rect 14280 9367 14332 9376
rect 14280 9333 14289 9367
rect 14289 9333 14323 9367
rect 14323 9333 14332 9367
rect 14280 9324 14332 9333
rect 14648 9367 14700 9376
rect 14648 9333 14657 9367
rect 14657 9333 14691 9367
rect 14691 9333 14700 9367
rect 14648 9324 14700 9333
rect 15108 9324 15160 9376
rect 15568 9324 15620 9376
rect 17684 9324 17736 9376
rect 17776 9324 17828 9376
rect 18328 9324 18380 9376
rect 18696 9324 18748 9376
rect 20536 9460 20588 9512
rect 19616 9392 19668 9444
rect 20996 9537 21005 9571
rect 21005 9537 21039 9571
rect 21039 9537 21048 9571
rect 20996 9528 21048 9537
rect 21548 9528 21600 9580
rect 22928 9528 22980 9580
rect 21272 9503 21324 9512
rect 21272 9469 21281 9503
rect 21281 9469 21315 9503
rect 21315 9469 21324 9503
rect 21272 9460 21324 9469
rect 22928 9392 22980 9444
rect 19708 9324 19760 9376
rect 19892 9324 19944 9376
rect 20444 9324 20496 9376
rect 3549 9222 3601 9274
rect 3613 9222 3665 9274
rect 3677 9222 3729 9274
rect 3741 9222 3793 9274
rect 3805 9222 3857 9274
rect 8747 9222 8799 9274
rect 8811 9222 8863 9274
rect 8875 9222 8927 9274
rect 8939 9222 8991 9274
rect 9003 9222 9055 9274
rect 13945 9222 13997 9274
rect 14009 9222 14061 9274
rect 14073 9222 14125 9274
rect 14137 9222 14189 9274
rect 14201 9222 14253 9274
rect 19143 9222 19195 9274
rect 19207 9222 19259 9274
rect 19271 9222 19323 9274
rect 19335 9222 19387 9274
rect 19399 9222 19451 9274
rect 2136 9163 2188 9172
rect 2136 9129 2145 9163
rect 2145 9129 2179 9163
rect 2179 9129 2188 9163
rect 2136 9120 2188 9129
rect 2228 9163 2280 9172
rect 2228 9129 2237 9163
rect 2237 9129 2271 9163
rect 2271 9129 2280 9163
rect 2228 9120 2280 9129
rect 2596 9120 2648 9172
rect 4620 9163 4672 9172
rect 4620 9129 4629 9163
rect 4629 9129 4663 9163
rect 4663 9129 4672 9163
rect 4620 9120 4672 9129
rect 5264 9163 5316 9172
rect 5264 9129 5273 9163
rect 5273 9129 5307 9163
rect 5307 9129 5316 9163
rect 5264 9120 5316 9129
rect 5632 9120 5684 9172
rect 7012 9120 7064 9172
rect 8668 9120 8720 9172
rect 10416 9120 10468 9172
rect 1584 9027 1636 9036
rect 1584 8993 1593 9027
rect 1593 8993 1627 9027
rect 1627 8993 1636 9027
rect 3700 9052 3752 9104
rect 4160 9052 4212 9104
rect 4804 9052 4856 9104
rect 7840 9095 7892 9104
rect 7840 9061 7849 9095
rect 7849 9061 7883 9095
rect 7883 9061 7892 9095
rect 7840 9052 7892 9061
rect 1584 8984 1636 8993
rect 3976 8984 4028 9036
rect 4252 9027 4304 9036
rect 4252 8993 4261 9027
rect 4261 8993 4295 9027
rect 4295 8993 4304 9027
rect 4252 8984 4304 8993
rect 4344 9027 4396 9036
rect 4344 8993 4353 9027
rect 4353 8993 4387 9027
rect 4387 8993 4396 9027
rect 4344 8984 4396 8993
rect 5908 9027 5960 9036
rect 5908 8993 5917 9027
rect 5917 8993 5951 9027
rect 5951 8993 5960 9027
rect 5908 8984 5960 8993
rect 6460 8984 6512 9036
rect 6644 8984 6696 9036
rect 7564 9027 7616 9036
rect 7564 8993 7573 9027
rect 7573 8993 7607 9027
rect 7607 8993 7616 9027
rect 7564 8984 7616 8993
rect 1400 8916 1452 8968
rect 2964 8916 3016 8968
rect 3332 8959 3384 8968
rect 3332 8925 3350 8959
rect 3350 8925 3384 8959
rect 3332 8916 3384 8925
rect 4436 8916 4488 8968
rect 2412 8848 2464 8900
rect 1768 8823 1820 8832
rect 1768 8789 1777 8823
rect 1777 8789 1811 8823
rect 1811 8789 1820 8823
rect 1768 8780 1820 8789
rect 4160 8780 4212 8832
rect 5080 8916 5132 8968
rect 5264 8780 5316 8832
rect 5540 8780 5592 8832
rect 5816 8848 5868 8900
rect 7012 8916 7064 8968
rect 8576 9052 8628 9104
rect 8668 9027 8720 9036
rect 8668 8993 8677 9027
rect 8677 8993 8711 9027
rect 8711 8993 8720 9027
rect 8668 8984 8720 8993
rect 8392 8916 8444 8968
rect 10968 9120 11020 9172
rect 11336 9120 11388 9172
rect 13636 9120 13688 9172
rect 14096 9120 14148 9172
rect 14464 9120 14516 9172
rect 13360 8984 13412 9036
rect 13820 8984 13872 9036
rect 16856 9120 16908 9172
rect 17132 9163 17184 9172
rect 17132 9129 17141 9163
rect 17141 9129 17175 9163
rect 17175 9129 17184 9163
rect 17132 9120 17184 9129
rect 17316 9120 17368 9172
rect 18696 9120 18748 9172
rect 18788 9120 18840 9172
rect 20260 9120 20312 9172
rect 20720 9163 20772 9172
rect 20720 9129 20729 9163
rect 20729 9129 20763 9163
rect 20763 9129 20772 9163
rect 20720 9120 20772 9129
rect 17408 9052 17460 9104
rect 17132 8984 17184 9036
rect 18144 8984 18196 9036
rect 18788 9027 18840 9036
rect 6644 8848 6696 8900
rect 9036 8848 9088 8900
rect 6920 8780 6972 8832
rect 7380 8823 7432 8832
rect 7380 8789 7389 8823
rect 7389 8789 7423 8823
rect 7423 8789 7432 8823
rect 7380 8780 7432 8789
rect 7656 8780 7708 8832
rect 8576 8780 8628 8832
rect 10784 8823 10836 8832
rect 10784 8789 10793 8823
rect 10793 8789 10827 8823
rect 10827 8789 10836 8823
rect 10784 8780 10836 8789
rect 11060 8823 11112 8832
rect 11060 8789 11069 8823
rect 11069 8789 11103 8823
rect 11103 8789 11112 8823
rect 11060 8780 11112 8789
rect 11704 8848 11756 8900
rect 12900 8959 12952 8968
rect 12900 8925 12909 8959
rect 12909 8925 12943 8959
rect 12943 8925 12952 8959
rect 12900 8916 12952 8925
rect 14096 8959 14148 8968
rect 12808 8848 12860 8900
rect 14096 8925 14105 8959
rect 14105 8925 14139 8959
rect 14139 8925 14148 8959
rect 14096 8916 14148 8925
rect 13360 8848 13412 8900
rect 13728 8848 13780 8900
rect 12532 8823 12584 8832
rect 12532 8789 12541 8823
rect 12541 8789 12575 8823
rect 12575 8789 12584 8823
rect 12532 8780 12584 8789
rect 12900 8780 12952 8832
rect 13544 8823 13596 8832
rect 13544 8789 13553 8823
rect 13553 8789 13587 8823
rect 13587 8789 13596 8823
rect 13544 8780 13596 8789
rect 15476 8916 15528 8968
rect 15200 8848 15252 8900
rect 18788 8993 18797 9027
rect 18797 8993 18831 9027
rect 18831 8993 18840 9027
rect 18788 8984 18840 8993
rect 21272 9027 21324 9036
rect 18604 8916 18656 8968
rect 19064 8916 19116 8968
rect 21272 8993 21281 9027
rect 21281 8993 21315 9027
rect 21315 8993 21324 9027
rect 21272 8984 21324 8993
rect 16028 8848 16080 8900
rect 18144 8848 18196 8900
rect 18972 8891 19024 8900
rect 18972 8857 18981 8891
rect 18981 8857 19015 8891
rect 19015 8857 19024 8891
rect 18972 8848 19024 8857
rect 15292 8780 15344 8832
rect 15752 8780 15804 8832
rect 16120 8780 16172 8832
rect 18328 8823 18380 8832
rect 18328 8789 18337 8823
rect 18337 8789 18371 8823
rect 18371 8789 18380 8823
rect 18328 8780 18380 8789
rect 18788 8780 18840 8832
rect 19892 8848 19944 8900
rect 21548 8848 21600 8900
rect 19248 8780 19300 8832
rect 19800 8780 19852 8832
rect 20628 8823 20680 8832
rect 20628 8789 20637 8823
rect 20637 8789 20671 8823
rect 20671 8789 20680 8823
rect 20628 8780 20680 8789
rect 21180 8823 21232 8832
rect 21180 8789 21189 8823
rect 21189 8789 21223 8823
rect 21223 8789 21232 8823
rect 21180 8780 21232 8789
rect 6148 8678 6200 8730
rect 6212 8678 6264 8730
rect 6276 8678 6328 8730
rect 6340 8678 6392 8730
rect 6404 8678 6456 8730
rect 11346 8678 11398 8730
rect 11410 8678 11462 8730
rect 11474 8678 11526 8730
rect 11538 8678 11590 8730
rect 11602 8678 11654 8730
rect 16544 8678 16596 8730
rect 16608 8678 16660 8730
rect 16672 8678 16724 8730
rect 16736 8678 16788 8730
rect 16800 8678 16852 8730
rect 21742 8678 21794 8730
rect 21806 8678 21858 8730
rect 21870 8678 21922 8730
rect 21934 8678 21986 8730
rect 21998 8678 22050 8730
rect 2136 8576 2188 8628
rect 2320 8619 2372 8628
rect 2320 8585 2329 8619
rect 2329 8585 2363 8619
rect 2363 8585 2372 8619
rect 2320 8576 2372 8585
rect 2412 8619 2464 8628
rect 2412 8585 2421 8619
rect 2421 8585 2455 8619
rect 2455 8585 2464 8619
rect 2412 8576 2464 8585
rect 3148 8576 3200 8628
rect 3332 8576 3384 8628
rect 3884 8619 3936 8628
rect 3884 8585 3893 8619
rect 3893 8585 3927 8619
rect 3927 8585 3936 8619
rect 3884 8576 3936 8585
rect 4712 8576 4764 8628
rect 5632 8619 5684 8628
rect 5632 8585 5641 8619
rect 5641 8585 5675 8619
rect 5675 8585 5684 8619
rect 5632 8576 5684 8585
rect 6092 8576 6144 8628
rect 7012 8576 7064 8628
rect 7564 8576 7616 8628
rect 8024 8576 8076 8628
rect 9588 8619 9640 8628
rect 9588 8585 9597 8619
rect 9597 8585 9631 8619
rect 9631 8585 9640 8619
rect 9588 8576 9640 8585
rect 10140 8619 10192 8628
rect 10140 8585 10149 8619
rect 10149 8585 10183 8619
rect 10183 8585 10192 8619
rect 10140 8576 10192 8585
rect 10508 8619 10560 8628
rect 10508 8585 10517 8619
rect 10517 8585 10551 8619
rect 10551 8585 10560 8619
rect 10508 8576 10560 8585
rect 10600 8576 10652 8628
rect 12900 8576 12952 8628
rect 13268 8576 13320 8628
rect 13820 8576 13872 8628
rect 18052 8576 18104 8628
rect 18328 8619 18380 8628
rect 18328 8585 18337 8619
rect 18337 8585 18371 8619
rect 18371 8585 18380 8619
rect 18328 8576 18380 8585
rect 18420 8576 18472 8628
rect 18788 8576 18840 8628
rect 18880 8576 18932 8628
rect 6828 8508 6880 8560
rect 7472 8508 7524 8560
rect 1952 8483 2004 8492
rect 1952 8449 1961 8483
rect 1961 8449 1995 8483
rect 1995 8449 2004 8483
rect 1952 8440 2004 8449
rect 3148 8440 3200 8492
rect 3884 8440 3936 8492
rect 4528 8440 4580 8492
rect 4804 8483 4856 8492
rect 4804 8449 4813 8483
rect 4813 8449 4847 8483
rect 4847 8449 4856 8483
rect 4804 8440 4856 8449
rect 6092 8440 6144 8492
rect 7564 8440 7616 8492
rect 1584 8372 1636 8424
rect 1860 8415 1912 8424
rect 1860 8381 1869 8415
rect 1869 8381 1903 8415
rect 1903 8381 1912 8415
rect 1860 8372 1912 8381
rect 3056 8415 3108 8424
rect 3056 8381 3065 8415
rect 3065 8381 3099 8415
rect 3099 8381 3108 8415
rect 3056 8372 3108 8381
rect 3516 8372 3568 8424
rect 4620 8372 4672 8424
rect 5264 8372 5316 8424
rect 5908 8415 5960 8424
rect 5908 8381 5917 8415
rect 5917 8381 5951 8415
rect 5951 8381 5960 8415
rect 5908 8372 5960 8381
rect 2320 8304 2372 8356
rect 5080 8304 5132 8356
rect 5632 8304 5684 8356
rect 6184 8304 6236 8356
rect 4252 8236 4304 8288
rect 4804 8236 4856 8288
rect 5172 8236 5224 8288
rect 7748 8440 7800 8492
rect 9036 8483 9088 8492
rect 9036 8449 9045 8483
rect 9045 8449 9079 8483
rect 9079 8449 9088 8483
rect 9036 8440 9088 8449
rect 9220 8440 9272 8492
rect 10508 8440 10560 8492
rect 12624 8483 12676 8492
rect 9680 8415 9732 8424
rect 9680 8381 9689 8415
rect 9689 8381 9723 8415
rect 9723 8381 9732 8415
rect 9680 8372 9732 8381
rect 10416 8372 10468 8424
rect 12624 8449 12642 8483
rect 12642 8449 12676 8483
rect 12624 8440 12676 8449
rect 12808 8440 12860 8492
rect 13636 8508 13688 8560
rect 14004 8508 14056 8560
rect 15844 8551 15896 8560
rect 15844 8517 15853 8551
rect 15853 8517 15887 8551
rect 15887 8517 15896 8551
rect 15844 8508 15896 8517
rect 16212 8508 16264 8560
rect 17132 8508 17184 8560
rect 14096 8483 14148 8492
rect 14096 8449 14105 8483
rect 14105 8449 14139 8483
rect 14139 8449 14148 8483
rect 14096 8440 14148 8449
rect 14924 8440 14976 8492
rect 11612 8372 11664 8424
rect 11796 8372 11848 8424
rect 12992 8372 13044 8424
rect 13636 8372 13688 8424
rect 14740 8372 14792 8424
rect 15200 8415 15252 8424
rect 15200 8381 15209 8415
rect 15209 8381 15243 8415
rect 15243 8381 15252 8415
rect 15200 8372 15252 8381
rect 8024 8304 8076 8356
rect 8300 8304 8352 8356
rect 9128 8304 9180 8356
rect 10232 8304 10284 8356
rect 7012 8236 7064 8288
rect 9772 8236 9824 8288
rect 11060 8236 11112 8288
rect 11336 8236 11388 8288
rect 11704 8236 11756 8288
rect 12900 8304 12952 8356
rect 14004 8304 14056 8356
rect 14188 8304 14240 8356
rect 15016 8304 15068 8356
rect 13820 8236 13872 8288
rect 14832 8236 14884 8288
rect 15568 8372 15620 8424
rect 15752 8372 15804 8424
rect 18972 8508 19024 8560
rect 19340 8576 19392 8628
rect 19892 8576 19944 8628
rect 20260 8619 20312 8628
rect 20260 8585 20269 8619
rect 20269 8585 20303 8619
rect 20303 8585 20312 8619
rect 20260 8576 20312 8585
rect 20444 8619 20496 8628
rect 20444 8585 20453 8619
rect 20453 8585 20487 8619
rect 20487 8585 20496 8619
rect 20444 8576 20496 8585
rect 18420 8483 18472 8492
rect 18420 8449 18429 8483
rect 18429 8449 18463 8483
rect 18463 8449 18472 8483
rect 18420 8440 18472 8449
rect 18880 8440 18932 8492
rect 19248 8440 19300 8492
rect 19800 8483 19852 8492
rect 19800 8449 19818 8483
rect 19818 8449 19852 8483
rect 19800 8440 19852 8449
rect 20720 8483 20772 8492
rect 20720 8449 20729 8483
rect 20729 8449 20763 8483
rect 20763 8449 20772 8483
rect 20720 8440 20772 8449
rect 16580 8372 16632 8424
rect 18512 8372 18564 8424
rect 15660 8304 15712 8356
rect 16304 8347 16356 8356
rect 16304 8313 16313 8347
rect 16313 8313 16347 8347
rect 16347 8313 16356 8347
rect 16304 8304 16356 8313
rect 16948 8304 17000 8356
rect 18236 8304 18288 8356
rect 15844 8236 15896 8288
rect 16212 8236 16264 8288
rect 18144 8236 18196 8288
rect 18696 8236 18748 8288
rect 19064 8236 19116 8288
rect 20720 8304 20772 8356
rect 21732 8304 21784 8356
rect 22928 8304 22980 8356
rect 3549 8134 3601 8186
rect 3613 8134 3665 8186
rect 3677 8134 3729 8186
rect 3741 8134 3793 8186
rect 3805 8134 3857 8186
rect 8747 8134 8799 8186
rect 8811 8134 8863 8186
rect 8875 8134 8927 8186
rect 8939 8134 8991 8186
rect 9003 8134 9055 8186
rect 13945 8134 13997 8186
rect 14009 8134 14061 8186
rect 14073 8134 14125 8186
rect 14137 8134 14189 8186
rect 14201 8134 14253 8186
rect 19143 8134 19195 8186
rect 19207 8134 19259 8186
rect 19271 8134 19323 8186
rect 19335 8134 19387 8186
rect 19399 8134 19451 8186
rect 1768 8032 1820 8084
rect 1860 8032 1912 8084
rect 2964 8032 3016 8084
rect 4988 8032 5040 8084
rect 5356 8032 5408 8084
rect 5724 8032 5776 8084
rect 7380 8032 7432 8084
rect 7748 8032 7800 8084
rect 9312 8032 9364 8084
rect 9772 8032 9824 8084
rect 11796 8032 11848 8084
rect 12440 8032 12492 8084
rect 13268 8032 13320 8084
rect 13912 8032 13964 8084
rect 15108 8032 15160 8084
rect 16028 8032 16080 8084
rect 16120 8032 16172 8084
rect 17316 8032 17368 8084
rect 17960 8032 18012 8084
rect 18420 8032 18472 8084
rect 20996 8032 21048 8084
rect 21088 8032 21140 8084
rect 3240 7964 3292 8016
rect 5448 7964 5500 8016
rect 2688 7896 2740 7948
rect 3056 7896 3108 7948
rect 3516 7896 3568 7948
rect 3976 7896 4028 7948
rect 4252 7939 4304 7948
rect 4252 7905 4261 7939
rect 4261 7905 4295 7939
rect 4295 7905 4304 7939
rect 4252 7896 4304 7905
rect 4344 7939 4396 7948
rect 4344 7905 4353 7939
rect 4353 7905 4387 7939
rect 4387 7905 4396 7939
rect 4344 7896 4396 7905
rect 4896 7896 4948 7948
rect 5172 7896 5224 7948
rect 2044 7828 2096 7880
rect 2228 7828 2280 7880
rect 4804 7828 4856 7880
rect 5448 7828 5500 7880
rect 6276 7964 6328 8016
rect 6000 7896 6052 7948
rect 5816 7828 5868 7880
rect 6184 7871 6236 7880
rect 6184 7837 6193 7871
rect 6193 7837 6227 7871
rect 6227 7837 6236 7871
rect 6828 7896 6880 7948
rect 7840 7896 7892 7948
rect 8116 7896 8168 7948
rect 8760 7896 8812 7948
rect 8852 7896 8904 7948
rect 6184 7828 6236 7837
rect 2596 7760 2648 7812
rect 2504 7692 2556 7744
rect 3792 7760 3844 7812
rect 3516 7692 3568 7744
rect 3976 7692 4028 7744
rect 4528 7760 4580 7812
rect 5356 7760 5408 7812
rect 6552 7760 6604 7812
rect 7748 7828 7800 7880
rect 9312 7871 9364 7880
rect 9312 7837 9321 7871
rect 9321 7837 9355 7871
rect 9355 7837 9364 7871
rect 11244 7964 11296 8016
rect 12624 7964 12676 8016
rect 16580 8007 16632 8016
rect 11336 7896 11388 7948
rect 13728 7896 13780 7948
rect 14740 7896 14792 7948
rect 15200 7896 15252 7948
rect 15292 7896 15344 7948
rect 16580 7973 16589 8007
rect 16589 7973 16623 8007
rect 16623 7973 16632 8007
rect 16580 7964 16632 7973
rect 20444 7964 20496 8016
rect 20536 7964 20588 8016
rect 21456 7964 21508 8016
rect 17224 7896 17276 7948
rect 9312 7828 9364 7837
rect 10600 7828 10652 7880
rect 10784 7828 10836 7880
rect 6920 7760 6972 7812
rect 8300 7760 8352 7812
rect 10876 7760 10928 7812
rect 12532 7828 12584 7880
rect 12992 7828 13044 7880
rect 13360 7871 13412 7880
rect 13360 7837 13369 7871
rect 13369 7837 13403 7871
rect 13403 7837 13412 7871
rect 13360 7828 13412 7837
rect 14464 7828 14516 7880
rect 14648 7828 14700 7880
rect 12624 7760 12676 7812
rect 12808 7760 12860 7812
rect 14372 7803 14424 7812
rect 14372 7769 14381 7803
rect 14381 7769 14415 7803
rect 14415 7769 14424 7803
rect 14372 7760 14424 7769
rect 16212 7760 16264 7812
rect 17408 7871 17460 7880
rect 17408 7837 17417 7871
rect 17417 7837 17451 7871
rect 17451 7837 17460 7871
rect 17408 7828 17460 7837
rect 18604 7896 18656 7948
rect 20628 7896 20680 7948
rect 20812 7896 20864 7948
rect 18972 7828 19024 7880
rect 19064 7828 19116 7880
rect 19892 7871 19944 7880
rect 19892 7837 19901 7871
rect 19901 7837 19935 7871
rect 19935 7837 19944 7871
rect 19892 7828 19944 7837
rect 21088 7896 21140 7948
rect 4712 7692 4764 7744
rect 4896 7735 4948 7744
rect 4896 7701 4905 7735
rect 4905 7701 4939 7735
rect 4939 7701 4948 7735
rect 4896 7692 4948 7701
rect 5816 7692 5868 7744
rect 5908 7692 5960 7744
rect 6644 7692 6696 7744
rect 7748 7735 7800 7744
rect 7748 7701 7757 7735
rect 7757 7701 7791 7735
rect 7791 7701 7800 7735
rect 7748 7692 7800 7701
rect 8116 7735 8168 7744
rect 8116 7701 8125 7735
rect 8125 7701 8159 7735
rect 8159 7701 8168 7735
rect 8576 7735 8628 7744
rect 8116 7692 8168 7701
rect 8576 7701 8585 7735
rect 8585 7701 8619 7735
rect 8619 7701 8628 7735
rect 8576 7692 8628 7701
rect 8668 7692 8720 7744
rect 9772 7735 9824 7744
rect 9772 7701 9781 7735
rect 9781 7701 9815 7735
rect 9815 7701 9824 7735
rect 9772 7692 9824 7701
rect 10232 7692 10284 7744
rect 11244 7692 11296 7744
rect 12256 7692 12308 7744
rect 12992 7735 13044 7744
rect 12992 7701 13001 7735
rect 13001 7701 13035 7735
rect 13035 7701 13044 7735
rect 12992 7692 13044 7701
rect 13636 7692 13688 7744
rect 15292 7692 15344 7744
rect 15936 7692 15988 7744
rect 17592 7692 17644 7744
rect 17960 7692 18012 7744
rect 19340 7692 19392 7744
rect 20720 7692 20772 7744
rect 21088 7692 21140 7744
rect 6148 7590 6200 7642
rect 6212 7590 6264 7642
rect 6276 7590 6328 7642
rect 6340 7590 6392 7642
rect 6404 7590 6456 7642
rect 11346 7590 11398 7642
rect 11410 7590 11462 7642
rect 11474 7590 11526 7642
rect 11538 7590 11590 7642
rect 11602 7590 11654 7642
rect 16544 7590 16596 7642
rect 16608 7590 16660 7642
rect 16672 7590 16724 7642
rect 16736 7590 16788 7642
rect 16800 7590 16852 7642
rect 21742 7590 21794 7642
rect 21806 7590 21858 7642
rect 21870 7590 21922 7642
rect 21934 7590 21986 7642
rect 21998 7590 22050 7642
rect 1584 7531 1636 7540
rect 1584 7497 1593 7531
rect 1593 7497 1627 7531
rect 1627 7497 1636 7531
rect 1584 7488 1636 7497
rect 2412 7488 2464 7540
rect 2596 7488 2648 7540
rect 4528 7488 4580 7540
rect 5172 7488 5224 7540
rect 6000 7488 6052 7540
rect 6828 7488 6880 7540
rect 6920 7488 6972 7540
rect 8760 7488 8812 7540
rect 10140 7531 10192 7540
rect 2780 7420 2832 7472
rect 1400 7395 1452 7404
rect 1400 7361 1409 7395
rect 1409 7361 1443 7395
rect 1443 7361 1452 7395
rect 1400 7352 1452 7361
rect 4896 7420 4948 7472
rect 5448 7420 5500 7472
rect 8392 7420 8444 7472
rect 3424 7352 3476 7404
rect 4528 7352 4580 7404
rect 4620 7352 4672 7404
rect 4804 7327 4856 7336
rect 4804 7293 4813 7327
rect 4813 7293 4847 7327
rect 4847 7293 4856 7327
rect 4804 7284 4856 7293
rect 4252 7148 4304 7200
rect 5172 7148 5224 7200
rect 6920 7352 6972 7404
rect 8300 7352 8352 7404
rect 8852 7352 8904 7404
rect 10140 7497 10149 7531
rect 10149 7497 10183 7531
rect 10183 7497 10192 7531
rect 10140 7488 10192 7497
rect 11244 7488 11296 7540
rect 12992 7488 13044 7540
rect 13636 7531 13688 7540
rect 13636 7497 13645 7531
rect 13645 7497 13679 7531
rect 13679 7497 13688 7531
rect 13636 7488 13688 7497
rect 9680 7420 9732 7472
rect 10324 7420 10376 7472
rect 10876 7420 10928 7472
rect 9496 7352 9548 7404
rect 9864 7352 9916 7404
rect 10968 7352 11020 7404
rect 11152 7395 11204 7404
rect 11152 7361 11161 7395
rect 11161 7361 11195 7395
rect 11195 7361 11204 7395
rect 11152 7352 11204 7361
rect 14556 7488 14608 7540
rect 14832 7488 14884 7540
rect 15016 7488 15068 7540
rect 15292 7488 15344 7540
rect 18144 7488 18196 7540
rect 7104 7284 7156 7336
rect 7380 7284 7432 7336
rect 9312 7327 9364 7336
rect 9312 7293 9321 7327
rect 9321 7293 9355 7327
rect 9355 7293 9364 7327
rect 9312 7284 9364 7293
rect 6644 7148 6696 7200
rect 7104 7191 7156 7200
rect 7104 7157 7113 7191
rect 7113 7157 7147 7191
rect 7147 7157 7156 7191
rect 7104 7148 7156 7157
rect 7656 7148 7708 7200
rect 9220 7216 9272 7268
rect 11980 7352 12032 7404
rect 12072 7352 12124 7404
rect 12256 7352 12308 7404
rect 12716 7395 12768 7404
rect 12716 7361 12725 7395
rect 12725 7361 12759 7395
rect 12759 7361 12768 7395
rect 12716 7352 12768 7361
rect 13544 7352 13596 7404
rect 14556 7352 14608 7404
rect 11704 7284 11756 7336
rect 12624 7284 12676 7336
rect 9680 7216 9732 7268
rect 10876 7216 10928 7268
rect 11244 7216 11296 7268
rect 13360 7284 13412 7336
rect 13268 7216 13320 7268
rect 13544 7216 13596 7268
rect 13728 7216 13780 7268
rect 14924 7284 14976 7336
rect 15200 7327 15252 7336
rect 15200 7293 15209 7327
rect 15209 7293 15243 7327
rect 15243 7293 15252 7327
rect 15200 7284 15252 7293
rect 15476 7395 15528 7404
rect 15476 7361 15485 7395
rect 15485 7361 15519 7395
rect 15519 7361 15528 7395
rect 15476 7352 15528 7361
rect 16212 7352 16264 7404
rect 16396 7352 16448 7404
rect 15844 7284 15896 7336
rect 16028 7327 16080 7336
rect 16028 7293 16037 7327
rect 16037 7293 16071 7327
rect 16071 7293 16080 7327
rect 16028 7284 16080 7293
rect 16488 7284 16540 7336
rect 17316 7284 17368 7336
rect 18144 7327 18196 7336
rect 18144 7293 18153 7327
rect 18153 7293 18187 7327
rect 18187 7293 18196 7327
rect 18144 7284 18196 7293
rect 18696 7488 18748 7540
rect 19800 7488 19852 7540
rect 19984 7488 20036 7540
rect 21180 7531 21232 7540
rect 21180 7497 21189 7531
rect 21189 7497 21223 7531
rect 21223 7497 21232 7531
rect 21180 7488 21232 7497
rect 18604 7463 18656 7472
rect 18604 7429 18638 7463
rect 18638 7429 18656 7463
rect 18604 7420 18656 7429
rect 20260 7463 20312 7472
rect 20260 7429 20269 7463
rect 20269 7429 20303 7463
rect 20303 7429 20312 7463
rect 20260 7420 20312 7429
rect 21456 7463 21508 7472
rect 21456 7429 21465 7463
rect 21465 7429 21499 7463
rect 21499 7429 21508 7463
rect 21456 7420 21508 7429
rect 19984 7395 20036 7404
rect 19984 7361 19993 7395
rect 19993 7361 20027 7395
rect 20027 7361 20036 7395
rect 19984 7352 20036 7361
rect 19340 7284 19392 7336
rect 21088 7352 21140 7404
rect 15292 7216 15344 7268
rect 9864 7148 9916 7200
rect 10968 7148 11020 7200
rect 11612 7148 11664 7200
rect 12256 7148 12308 7200
rect 12992 7148 13044 7200
rect 14832 7148 14884 7200
rect 15384 7148 15436 7200
rect 16212 7191 16264 7200
rect 16212 7157 16221 7191
rect 16221 7157 16255 7191
rect 16255 7157 16264 7191
rect 16212 7148 16264 7157
rect 17776 7216 17828 7268
rect 20904 7284 20956 7336
rect 21180 7284 21232 7336
rect 20812 7216 20864 7268
rect 17500 7191 17552 7200
rect 17500 7157 17509 7191
rect 17509 7157 17543 7191
rect 17543 7157 17552 7191
rect 17500 7148 17552 7157
rect 17684 7148 17736 7200
rect 20260 7148 20312 7200
rect 3549 7046 3601 7098
rect 3613 7046 3665 7098
rect 3677 7046 3729 7098
rect 3741 7046 3793 7098
rect 3805 7046 3857 7098
rect 8747 7046 8799 7098
rect 8811 7046 8863 7098
rect 8875 7046 8927 7098
rect 8939 7046 8991 7098
rect 9003 7046 9055 7098
rect 13945 7046 13997 7098
rect 14009 7046 14061 7098
rect 14073 7046 14125 7098
rect 14137 7046 14189 7098
rect 14201 7046 14253 7098
rect 19143 7046 19195 7098
rect 19207 7046 19259 7098
rect 19271 7046 19323 7098
rect 19335 7046 19387 7098
rect 19399 7046 19451 7098
rect 3608 6987 3660 6996
rect 3608 6953 3617 6987
rect 3617 6953 3651 6987
rect 3651 6953 3660 6987
rect 3608 6944 3660 6953
rect 3976 6944 4028 6996
rect 5080 6944 5132 6996
rect 10232 6944 10284 6996
rect 10876 6944 10928 6996
rect 12808 6944 12860 6996
rect 13360 6944 13412 6996
rect 572 6808 624 6860
rect 1492 6808 1544 6860
rect 2504 6808 2556 6860
rect 2780 6808 2832 6860
rect 3608 6808 3660 6860
rect 4528 6876 4580 6928
rect 2136 6740 2188 6792
rect 2872 6740 2924 6792
rect 3148 6783 3200 6792
rect 3148 6749 3157 6783
rect 3157 6749 3191 6783
rect 3191 6749 3200 6783
rect 3148 6740 3200 6749
rect 3240 6783 3292 6792
rect 3240 6749 3249 6783
rect 3249 6749 3283 6783
rect 3283 6749 3292 6783
rect 3240 6740 3292 6749
rect 3424 6740 3476 6792
rect 20 6672 72 6724
rect 940 6672 992 6724
rect 2596 6715 2648 6724
rect 2596 6681 2605 6715
rect 2605 6681 2639 6715
rect 2639 6681 2648 6715
rect 2596 6672 2648 6681
rect 3884 6672 3936 6724
rect 4068 6672 4120 6724
rect 5264 6851 5316 6860
rect 5264 6817 5273 6851
rect 5273 6817 5307 6851
rect 5307 6817 5316 6851
rect 5264 6808 5316 6817
rect 5080 6740 5132 6792
rect 5908 6876 5960 6928
rect 8300 6876 8352 6928
rect 5632 6808 5684 6860
rect 7012 6808 7064 6860
rect 8392 6808 8444 6860
rect 6460 6783 6512 6792
rect 6460 6749 6469 6783
rect 6469 6749 6503 6783
rect 6503 6749 6512 6783
rect 6460 6740 6512 6749
rect 8852 6808 8904 6860
rect 9496 6851 9548 6860
rect 9496 6817 9505 6851
rect 9505 6817 9539 6851
rect 9539 6817 9548 6851
rect 9496 6808 9548 6817
rect 2136 6604 2188 6656
rect 4988 6647 5040 6656
rect 4988 6613 4997 6647
rect 4997 6613 5031 6647
rect 5031 6613 5040 6647
rect 4988 6604 5040 6613
rect 5080 6647 5132 6656
rect 5080 6613 5089 6647
rect 5089 6613 5123 6647
rect 5123 6613 5132 6647
rect 5080 6604 5132 6613
rect 5264 6604 5316 6656
rect 5816 6647 5868 6656
rect 5816 6613 5825 6647
rect 5825 6613 5859 6647
rect 5859 6613 5868 6647
rect 5816 6604 5868 6613
rect 6552 6604 6604 6656
rect 6644 6604 6696 6656
rect 8576 6783 8628 6792
rect 8576 6749 8585 6783
rect 8585 6749 8619 6783
rect 8619 6749 8628 6783
rect 8576 6740 8628 6749
rect 10140 6876 10192 6928
rect 11612 6876 11664 6928
rect 10048 6740 10100 6792
rect 10600 6740 10652 6792
rect 7288 6604 7340 6656
rect 7564 6604 7616 6656
rect 8116 6672 8168 6724
rect 8392 6672 8444 6724
rect 10692 6672 10744 6724
rect 11980 6876 12032 6928
rect 14464 6944 14516 6996
rect 15108 6944 15160 6996
rect 12164 6808 12216 6860
rect 8944 6647 8996 6656
rect 8944 6613 8953 6647
rect 8953 6613 8987 6647
rect 8987 6613 8996 6647
rect 8944 6604 8996 6613
rect 9588 6604 9640 6656
rect 9864 6647 9916 6656
rect 9864 6613 9873 6647
rect 9873 6613 9907 6647
rect 9907 6613 9916 6647
rect 9864 6604 9916 6613
rect 10416 6604 10468 6656
rect 11796 6672 11848 6724
rect 12348 6672 12400 6724
rect 12624 6851 12676 6860
rect 12624 6817 12633 6851
rect 12633 6817 12667 6851
rect 12667 6817 12676 6851
rect 12624 6808 12676 6817
rect 13084 6808 13136 6860
rect 15568 6808 15620 6860
rect 16488 6808 16540 6860
rect 14096 6783 14148 6792
rect 13544 6672 13596 6724
rect 14096 6749 14105 6783
rect 14105 6749 14139 6783
rect 14139 6749 14148 6783
rect 14096 6740 14148 6749
rect 15108 6740 15160 6792
rect 13820 6672 13872 6724
rect 15200 6672 15252 6724
rect 15936 6715 15988 6724
rect 15936 6681 15945 6715
rect 15945 6681 15979 6715
rect 15979 6681 15988 6715
rect 15936 6672 15988 6681
rect 18328 6944 18380 6996
rect 19984 6987 20036 6996
rect 18328 6808 18380 6860
rect 18788 6808 18840 6860
rect 19984 6953 19993 6987
rect 19993 6953 20027 6987
rect 20027 6953 20036 6987
rect 19984 6944 20036 6953
rect 18972 6876 19024 6928
rect 19156 6808 19208 6860
rect 19800 6808 19852 6860
rect 16948 6740 17000 6792
rect 11336 6647 11388 6656
rect 11336 6613 11345 6647
rect 11345 6613 11379 6647
rect 11379 6613 11388 6647
rect 11336 6604 11388 6613
rect 13084 6604 13136 6656
rect 13360 6647 13412 6656
rect 13360 6613 13369 6647
rect 13369 6613 13403 6647
rect 13403 6613 13412 6647
rect 13360 6604 13412 6613
rect 13636 6604 13688 6656
rect 14188 6604 14240 6656
rect 15476 6647 15528 6656
rect 15476 6613 15485 6647
rect 15485 6613 15519 6647
rect 15519 6613 15528 6647
rect 15476 6604 15528 6613
rect 15568 6647 15620 6656
rect 15568 6613 15577 6647
rect 15577 6613 15611 6647
rect 15611 6613 15620 6647
rect 16028 6647 16080 6656
rect 15568 6604 15620 6613
rect 16028 6613 16037 6647
rect 16037 6613 16071 6647
rect 16071 6613 16080 6647
rect 16028 6604 16080 6613
rect 16856 6604 16908 6656
rect 18696 6740 18748 6792
rect 20904 6808 20956 6860
rect 18144 6672 18196 6724
rect 20628 6740 20680 6792
rect 19800 6672 19852 6724
rect 20260 6672 20312 6724
rect 17960 6604 18012 6656
rect 18328 6604 18380 6656
rect 18972 6604 19024 6656
rect 19248 6604 19300 6656
rect 19708 6604 19760 6656
rect 19892 6604 19944 6656
rect 6148 6502 6200 6554
rect 6212 6502 6264 6554
rect 6276 6502 6328 6554
rect 6340 6502 6392 6554
rect 6404 6502 6456 6554
rect 11346 6502 11398 6554
rect 11410 6502 11462 6554
rect 11474 6502 11526 6554
rect 11538 6502 11590 6554
rect 11602 6502 11654 6554
rect 16544 6502 16596 6554
rect 16608 6502 16660 6554
rect 16672 6502 16724 6554
rect 16736 6502 16788 6554
rect 16800 6502 16852 6554
rect 21742 6502 21794 6554
rect 21806 6502 21858 6554
rect 21870 6502 21922 6554
rect 21934 6502 21986 6554
rect 21998 6502 22050 6554
rect 1952 6400 2004 6452
rect 2228 6443 2280 6452
rect 2228 6409 2237 6443
rect 2237 6409 2271 6443
rect 2271 6409 2280 6443
rect 2228 6400 2280 6409
rect 2872 6400 2924 6452
rect 7288 6400 7340 6452
rect 8300 6400 8352 6452
rect 8668 6400 8720 6452
rect 1492 6375 1544 6384
rect 1492 6341 1501 6375
rect 1501 6341 1535 6375
rect 1535 6341 1544 6375
rect 1492 6332 1544 6341
rect 1768 6332 1820 6384
rect 3148 6375 3200 6384
rect 3148 6341 3157 6375
rect 3157 6341 3191 6375
rect 3191 6341 3200 6375
rect 3148 6332 3200 6341
rect 2780 6307 2832 6316
rect 2780 6273 2789 6307
rect 2789 6273 2823 6307
rect 2823 6273 2832 6307
rect 6552 6332 6604 6384
rect 2780 6264 2832 6273
rect 2688 6196 2740 6248
rect 4252 6264 4304 6316
rect 4528 6264 4580 6316
rect 4896 6307 4948 6316
rect 4896 6273 4905 6307
rect 4905 6273 4939 6307
rect 4939 6273 4948 6307
rect 4896 6264 4948 6273
rect 5356 6264 5408 6316
rect 6184 6264 6236 6316
rect 6368 6264 6420 6316
rect 7012 6264 7064 6316
rect 4344 6196 4396 6248
rect 3148 6128 3200 6180
rect 3240 6128 3292 6180
rect 5080 6128 5132 6180
rect 5632 6196 5684 6248
rect 6644 6196 6696 6248
rect 7380 6239 7432 6248
rect 7380 6205 7389 6239
rect 7389 6205 7423 6239
rect 7423 6205 7432 6239
rect 7380 6196 7432 6205
rect 8208 6332 8260 6384
rect 9588 6332 9640 6384
rect 9128 6264 9180 6316
rect 9772 6264 9824 6316
rect 10048 6332 10100 6384
rect 10324 6307 10376 6316
rect 10324 6273 10342 6307
rect 10342 6273 10376 6307
rect 10324 6264 10376 6273
rect 9496 6196 9548 6248
rect 10600 6332 10652 6384
rect 11888 6400 11940 6452
rect 12440 6400 12492 6452
rect 16028 6400 16080 6452
rect 13820 6332 13872 6384
rect 16580 6400 16632 6452
rect 17040 6400 17092 6452
rect 14004 6307 14056 6316
rect 11980 6239 12032 6248
rect 11980 6205 11989 6239
rect 11989 6205 12023 6239
rect 12023 6205 12032 6239
rect 11980 6196 12032 6205
rect 14004 6273 14013 6307
rect 14013 6273 14047 6307
rect 14047 6273 14056 6307
rect 14004 6264 14056 6273
rect 14096 6264 14148 6316
rect 15476 6264 15528 6316
rect 15844 6264 15896 6316
rect 16028 6264 16080 6316
rect 16304 6332 16356 6384
rect 16764 6332 16816 6384
rect 17040 6307 17092 6316
rect 12900 6239 12952 6248
rect 5724 6128 5776 6180
rect 4620 6103 4672 6112
rect 4620 6069 4629 6103
rect 4629 6069 4663 6103
rect 4663 6069 4672 6103
rect 4620 6060 4672 6069
rect 4896 6060 4948 6112
rect 5356 6103 5408 6112
rect 5356 6069 5365 6103
rect 5365 6069 5399 6103
rect 5399 6069 5408 6103
rect 5356 6060 5408 6069
rect 5448 6060 5500 6112
rect 7840 6128 7892 6180
rect 8208 6128 8260 6180
rect 8944 6128 8996 6180
rect 9404 6128 9456 6180
rect 10784 6128 10836 6180
rect 11612 6128 11664 6180
rect 12900 6205 12909 6239
rect 12909 6205 12943 6239
rect 12943 6205 12952 6239
rect 12900 6196 12952 6205
rect 13820 6196 13872 6248
rect 15752 6196 15804 6248
rect 17040 6273 17049 6307
rect 17049 6273 17083 6307
rect 17083 6273 17092 6307
rect 17040 6264 17092 6273
rect 18420 6332 18472 6384
rect 18604 6400 18656 6452
rect 19248 6443 19300 6452
rect 19248 6409 19257 6443
rect 19257 6409 19291 6443
rect 19291 6409 19300 6443
rect 19248 6400 19300 6409
rect 19708 6443 19760 6452
rect 19708 6409 19717 6443
rect 19717 6409 19751 6443
rect 19751 6409 19760 6443
rect 19708 6400 19760 6409
rect 19800 6443 19852 6452
rect 19800 6409 19809 6443
rect 19809 6409 19843 6443
rect 19843 6409 19852 6443
rect 19800 6400 19852 6409
rect 20720 6400 20772 6452
rect 21364 6443 21416 6452
rect 21364 6409 21373 6443
rect 21373 6409 21407 6443
rect 21407 6409 21416 6443
rect 21364 6400 21416 6409
rect 21456 6400 21508 6452
rect 21732 6400 21784 6452
rect 17592 6307 17644 6316
rect 17592 6273 17626 6307
rect 17626 6273 17644 6307
rect 17592 6264 17644 6273
rect 18788 6264 18840 6316
rect 19524 6264 19576 6316
rect 20168 6307 20220 6316
rect 20168 6273 20177 6307
rect 20177 6273 20211 6307
rect 20211 6273 20220 6307
rect 20168 6264 20220 6273
rect 20720 6264 20772 6316
rect 14464 6128 14516 6180
rect 16212 6128 16264 6180
rect 17040 6128 17092 6180
rect 17132 6128 17184 6180
rect 5908 6060 5960 6112
rect 6276 6060 6328 6112
rect 8300 6060 8352 6112
rect 9680 6060 9732 6112
rect 10692 6060 10744 6112
rect 10876 6103 10928 6112
rect 10876 6069 10885 6103
rect 10885 6069 10919 6103
rect 10919 6069 10928 6103
rect 10876 6060 10928 6069
rect 11244 6060 11296 6112
rect 12992 6060 13044 6112
rect 13544 6103 13596 6112
rect 13544 6069 13553 6103
rect 13553 6069 13587 6103
rect 13587 6069 13596 6103
rect 13544 6060 13596 6069
rect 14004 6060 14056 6112
rect 14372 6103 14424 6112
rect 14372 6069 14381 6103
rect 14381 6069 14415 6103
rect 14415 6069 14424 6103
rect 14372 6060 14424 6069
rect 14832 6060 14884 6112
rect 16120 6060 16172 6112
rect 18604 6196 18656 6248
rect 20260 6239 20312 6248
rect 20260 6205 20269 6239
rect 20269 6205 20303 6239
rect 20303 6205 20312 6239
rect 20260 6196 20312 6205
rect 20812 6239 20864 6248
rect 20812 6205 20821 6239
rect 20821 6205 20855 6239
rect 20855 6205 20864 6239
rect 20812 6196 20864 6205
rect 18972 6060 19024 6112
rect 21548 6103 21600 6112
rect 21548 6069 21557 6103
rect 21557 6069 21591 6103
rect 21591 6069 21600 6103
rect 21548 6060 21600 6069
rect 3549 5958 3601 6010
rect 3613 5958 3665 6010
rect 3677 5958 3729 6010
rect 3741 5958 3793 6010
rect 3805 5958 3857 6010
rect 8747 5958 8799 6010
rect 8811 5958 8863 6010
rect 8875 5958 8927 6010
rect 8939 5958 8991 6010
rect 9003 5958 9055 6010
rect 13945 5958 13997 6010
rect 14009 5958 14061 6010
rect 14073 5958 14125 6010
rect 14137 5958 14189 6010
rect 14201 5958 14253 6010
rect 19143 5958 19195 6010
rect 19207 5958 19259 6010
rect 19271 5958 19323 6010
rect 19335 5958 19387 6010
rect 19399 5958 19451 6010
rect 3884 5856 3936 5908
rect 2872 5720 2924 5772
rect 3884 5720 3936 5772
rect 2596 5584 2648 5636
rect 2688 5584 2740 5636
rect 2136 5516 2188 5568
rect 3148 5559 3200 5568
rect 3148 5525 3157 5559
rect 3157 5525 3191 5559
rect 3191 5525 3200 5559
rect 3148 5516 3200 5525
rect 4988 5856 5040 5908
rect 5908 5899 5960 5908
rect 5908 5865 5917 5899
rect 5917 5865 5951 5899
rect 5951 5865 5960 5899
rect 5908 5856 5960 5865
rect 6184 5899 6236 5908
rect 6184 5865 6193 5899
rect 6193 5865 6227 5899
rect 6227 5865 6236 5899
rect 6184 5856 6236 5865
rect 6552 5856 6604 5908
rect 10600 5856 10652 5908
rect 10876 5856 10928 5908
rect 4252 5788 4304 5840
rect 6276 5788 6328 5840
rect 6368 5788 6420 5840
rect 7288 5788 7340 5840
rect 7932 5788 7984 5840
rect 8116 5788 8168 5840
rect 9588 5788 9640 5840
rect 10968 5788 11020 5840
rect 14648 5856 14700 5908
rect 18328 5856 18380 5908
rect 18420 5856 18472 5908
rect 19524 5899 19576 5908
rect 15476 5788 15528 5840
rect 17316 5831 17368 5840
rect 6644 5720 6696 5772
rect 7380 5763 7432 5772
rect 7380 5729 7389 5763
rect 7389 5729 7423 5763
rect 7423 5729 7432 5763
rect 7380 5720 7432 5729
rect 8760 5720 8812 5772
rect 9680 5720 9732 5772
rect 9864 5763 9916 5772
rect 9864 5729 9873 5763
rect 9873 5729 9907 5763
rect 9907 5729 9916 5763
rect 9864 5720 9916 5729
rect 10876 5720 10928 5772
rect 13176 5763 13228 5772
rect 5724 5695 5776 5704
rect 5724 5661 5733 5695
rect 5733 5661 5767 5695
rect 5767 5661 5776 5695
rect 5724 5652 5776 5661
rect 7472 5652 7524 5704
rect 7748 5652 7800 5704
rect 10600 5652 10652 5704
rect 4160 5627 4212 5636
rect 4160 5593 4169 5627
rect 4169 5593 4203 5627
rect 4203 5593 4212 5627
rect 4160 5584 4212 5593
rect 4252 5516 4304 5568
rect 4988 5584 5040 5636
rect 5632 5559 5684 5568
rect 5632 5525 5641 5559
rect 5641 5525 5675 5559
rect 5675 5525 5684 5559
rect 5632 5516 5684 5525
rect 5724 5516 5776 5568
rect 6368 5516 6420 5568
rect 6460 5516 6512 5568
rect 6828 5584 6880 5636
rect 8208 5584 8260 5636
rect 8668 5584 8720 5636
rect 6920 5516 6972 5568
rect 7472 5559 7524 5568
rect 7472 5525 7481 5559
rect 7481 5525 7515 5559
rect 7515 5525 7524 5559
rect 7472 5516 7524 5525
rect 7932 5559 7984 5568
rect 7932 5525 7941 5559
rect 7941 5525 7975 5559
rect 7975 5525 7984 5559
rect 7932 5516 7984 5525
rect 8576 5516 8628 5568
rect 9404 5584 9456 5636
rect 9864 5584 9916 5636
rect 11336 5584 11388 5636
rect 10140 5559 10192 5568
rect 10140 5525 10149 5559
rect 10149 5525 10183 5559
rect 10183 5525 10192 5559
rect 10508 5559 10560 5568
rect 10140 5516 10192 5525
rect 10508 5525 10517 5559
rect 10517 5525 10551 5559
rect 10551 5525 10560 5559
rect 10508 5516 10560 5525
rect 11244 5516 11296 5568
rect 11612 5516 11664 5568
rect 12164 5652 12216 5704
rect 13176 5729 13185 5763
rect 13185 5729 13219 5763
rect 13219 5729 13228 5763
rect 13176 5720 13228 5729
rect 13636 5720 13688 5772
rect 13084 5695 13136 5704
rect 13084 5661 13093 5695
rect 13093 5661 13127 5695
rect 13127 5661 13136 5695
rect 13084 5652 13136 5661
rect 14280 5720 14332 5772
rect 14464 5763 14516 5772
rect 14464 5729 14473 5763
rect 14473 5729 14507 5763
rect 14507 5729 14516 5763
rect 16580 5763 16632 5772
rect 14464 5720 14516 5729
rect 14924 5652 14976 5704
rect 11980 5584 12032 5636
rect 13912 5584 13964 5636
rect 12164 5559 12216 5568
rect 12164 5525 12173 5559
rect 12173 5525 12207 5559
rect 12207 5525 12216 5559
rect 12164 5516 12216 5525
rect 12716 5559 12768 5568
rect 12716 5525 12725 5559
rect 12725 5525 12759 5559
rect 12759 5525 12768 5559
rect 12716 5516 12768 5525
rect 13544 5559 13596 5568
rect 13544 5525 13553 5559
rect 13553 5525 13587 5559
rect 13587 5525 13596 5559
rect 13544 5516 13596 5525
rect 13820 5516 13872 5568
rect 14188 5516 14240 5568
rect 14464 5516 14516 5568
rect 15384 5652 15436 5704
rect 16580 5729 16589 5763
rect 16589 5729 16623 5763
rect 16623 5729 16632 5763
rect 16580 5720 16632 5729
rect 17316 5797 17325 5831
rect 17325 5797 17359 5831
rect 17359 5797 17368 5831
rect 17316 5788 17368 5797
rect 17592 5788 17644 5840
rect 19524 5865 19533 5899
rect 19533 5865 19567 5899
rect 19567 5865 19576 5899
rect 19524 5856 19576 5865
rect 20168 5856 20220 5908
rect 20996 5856 21048 5908
rect 21272 5788 21324 5840
rect 16764 5695 16816 5704
rect 16304 5627 16356 5636
rect 16304 5593 16322 5627
rect 16322 5593 16356 5627
rect 16764 5661 16773 5695
rect 16773 5661 16807 5695
rect 16807 5661 16816 5695
rect 16764 5652 16816 5661
rect 17040 5695 17092 5704
rect 17040 5661 17049 5695
rect 17049 5661 17083 5695
rect 17083 5661 17092 5695
rect 17040 5652 17092 5661
rect 18788 5720 18840 5772
rect 17868 5652 17920 5704
rect 18880 5652 18932 5704
rect 19064 5652 19116 5704
rect 19892 5695 19944 5704
rect 19892 5661 19901 5695
rect 19901 5661 19935 5695
rect 19935 5661 19944 5695
rect 19892 5652 19944 5661
rect 20444 5720 20496 5772
rect 21272 5652 21324 5704
rect 22560 5652 22612 5704
rect 16304 5584 16356 5593
rect 18144 5584 18196 5636
rect 18788 5627 18840 5636
rect 18788 5593 18797 5627
rect 18797 5593 18831 5627
rect 18831 5593 18840 5627
rect 18788 5584 18840 5593
rect 19708 5584 19760 5636
rect 21732 5584 21784 5636
rect 15384 5516 15436 5568
rect 16764 5516 16816 5568
rect 17132 5516 17184 5568
rect 17868 5516 17920 5568
rect 20720 5559 20772 5568
rect 20720 5525 20729 5559
rect 20729 5525 20763 5559
rect 20763 5525 20772 5559
rect 20720 5516 20772 5525
rect 388 5448 440 5500
rect 940 5448 992 5500
rect 6148 5414 6200 5466
rect 6212 5414 6264 5466
rect 6276 5414 6328 5466
rect 6340 5414 6392 5466
rect 6404 5414 6456 5466
rect 11346 5414 11398 5466
rect 11410 5414 11462 5466
rect 11474 5414 11526 5466
rect 11538 5414 11590 5466
rect 11602 5414 11654 5466
rect 16544 5414 16596 5466
rect 16608 5414 16660 5466
rect 16672 5414 16724 5466
rect 16736 5414 16788 5466
rect 16800 5414 16852 5466
rect 21742 5414 21794 5466
rect 21806 5414 21858 5466
rect 21870 5414 21922 5466
rect 21934 5414 21986 5466
rect 21998 5414 22050 5466
rect 3332 5355 3384 5364
rect 3332 5321 3341 5355
rect 3341 5321 3375 5355
rect 3375 5321 3384 5355
rect 3332 5312 3384 5321
rect 4068 5355 4120 5364
rect 4068 5321 4077 5355
rect 4077 5321 4111 5355
rect 4111 5321 4120 5355
rect 4068 5312 4120 5321
rect 4436 5312 4488 5364
rect 204 5244 256 5296
rect 1032 5244 1084 5296
rect 3516 5244 3568 5296
rect 2044 5176 2096 5228
rect 3332 5176 3384 5228
rect 3884 5176 3936 5228
rect 4160 5176 4212 5228
rect 1768 5108 1820 5160
rect 3056 5108 3108 5160
rect 5540 5244 5592 5296
rect 4160 5040 4212 5092
rect 4988 5176 5040 5228
rect 5724 5312 5776 5364
rect 5908 5312 5960 5364
rect 7472 5312 7524 5364
rect 8024 5312 8076 5364
rect 8760 5312 8812 5364
rect 10140 5312 10192 5364
rect 10784 5355 10836 5364
rect 10784 5321 10793 5355
rect 10793 5321 10827 5355
rect 10827 5321 10836 5355
rect 10784 5312 10836 5321
rect 11612 5312 11664 5364
rect 11888 5312 11940 5364
rect 12164 5312 12216 5364
rect 12256 5312 12308 5364
rect 12624 5312 12676 5364
rect 14372 5312 14424 5364
rect 17500 5312 17552 5364
rect 19432 5312 19484 5364
rect 7288 5244 7340 5296
rect 6276 5176 6328 5228
rect 7012 5176 7064 5228
rect 6644 5108 6696 5160
rect 7012 5040 7064 5092
rect 8024 5176 8076 5228
rect 9680 5244 9732 5296
rect 13728 5244 13780 5296
rect 16948 5244 17000 5296
rect 17224 5244 17276 5296
rect 7840 5108 7892 5160
rect 9312 5176 9364 5228
rect 10048 5219 10100 5228
rect 10048 5185 10057 5219
rect 10057 5185 10091 5219
rect 10091 5185 10100 5219
rect 10048 5176 10100 5185
rect 10508 5176 10560 5228
rect 11612 5176 11664 5228
rect 11888 5219 11940 5228
rect 11888 5185 11897 5219
rect 11897 5185 11931 5219
rect 11931 5185 11940 5219
rect 11888 5176 11940 5185
rect 11980 5176 12032 5228
rect 12256 5176 12308 5228
rect 12716 5176 12768 5228
rect 13084 5176 13136 5228
rect 14832 5176 14884 5228
rect 15108 5176 15160 5228
rect 15660 5219 15712 5228
rect 15660 5185 15669 5219
rect 15669 5185 15703 5219
rect 15703 5185 15712 5219
rect 15660 5176 15712 5185
rect 17592 5219 17644 5228
rect 17592 5185 17601 5219
rect 17601 5185 17635 5219
rect 17635 5185 17644 5219
rect 17592 5176 17644 5185
rect 10692 5108 10744 5160
rect 11152 5108 11204 5160
rect 2504 5015 2556 5024
rect 2504 4981 2513 5015
rect 2513 4981 2547 5015
rect 2547 4981 2556 5015
rect 2504 4972 2556 4981
rect 2872 5015 2924 5024
rect 2872 4981 2881 5015
rect 2881 4981 2915 5015
rect 2915 4981 2924 5015
rect 2872 4972 2924 4981
rect 3332 4972 3384 5024
rect 4252 4972 4304 5024
rect 4436 4972 4488 5024
rect 5724 4972 5776 5024
rect 6368 5015 6420 5024
rect 6368 4981 6377 5015
rect 6377 4981 6411 5015
rect 6411 4981 6420 5015
rect 6368 4972 6420 4981
rect 7288 5015 7340 5024
rect 7288 4981 7297 5015
rect 7297 4981 7331 5015
rect 7331 4981 7340 5015
rect 7288 4972 7340 4981
rect 7748 5040 7800 5092
rect 15200 5108 15252 5160
rect 16488 5108 16540 5160
rect 17316 5108 17368 5160
rect 18236 5176 18288 5228
rect 18420 5219 18472 5228
rect 18420 5185 18454 5219
rect 18454 5185 18472 5219
rect 19616 5244 19668 5296
rect 20904 5312 20956 5364
rect 21364 5355 21416 5364
rect 21364 5321 21373 5355
rect 21373 5321 21407 5355
rect 21407 5321 21416 5355
rect 21364 5312 21416 5321
rect 21732 5312 21784 5364
rect 22468 5312 22520 5364
rect 21456 5287 21508 5296
rect 21456 5253 21465 5287
rect 21465 5253 21499 5287
rect 21499 5253 21508 5287
rect 21456 5244 21508 5253
rect 18420 5176 18472 5185
rect 20260 5176 20312 5228
rect 21364 5176 21416 5228
rect 22744 5176 22796 5228
rect 16396 5040 16448 5092
rect 8944 4972 8996 5024
rect 10140 4972 10192 5024
rect 10324 5015 10376 5024
rect 10324 4981 10333 5015
rect 10333 4981 10367 5015
rect 10367 4981 10376 5015
rect 10324 4972 10376 4981
rect 11888 4972 11940 5024
rect 12348 4972 12400 5024
rect 13268 4972 13320 5024
rect 13452 4972 13504 5024
rect 13544 5015 13596 5024
rect 13544 4981 13553 5015
rect 13553 4981 13587 5015
rect 13587 4981 13596 5015
rect 15200 5015 15252 5024
rect 13544 4972 13596 4981
rect 15200 4981 15209 5015
rect 15209 4981 15243 5015
rect 15243 4981 15252 5015
rect 15200 4972 15252 4981
rect 18512 4972 18564 5024
rect 18880 4972 18932 5024
rect 20812 5108 20864 5160
rect 21456 5108 21508 5160
rect 3549 4870 3601 4922
rect 3613 4870 3665 4922
rect 3677 4870 3729 4922
rect 3741 4870 3793 4922
rect 3805 4870 3857 4922
rect 8747 4870 8799 4922
rect 8811 4870 8863 4922
rect 8875 4870 8927 4922
rect 8939 4870 8991 4922
rect 9003 4870 9055 4922
rect 13945 4870 13997 4922
rect 14009 4870 14061 4922
rect 14073 4870 14125 4922
rect 14137 4870 14189 4922
rect 14201 4870 14253 4922
rect 19143 4870 19195 4922
rect 19207 4870 19259 4922
rect 19271 4870 19323 4922
rect 19335 4870 19387 4922
rect 19399 4870 19451 4922
rect 2136 4768 2188 4820
rect 1952 4675 2004 4684
rect 1952 4641 1961 4675
rect 1961 4641 1995 4675
rect 1995 4641 2004 4675
rect 1952 4632 2004 4641
rect 2872 4700 2924 4752
rect 3148 4768 3200 4820
rect 5632 4768 5684 4820
rect 5816 4768 5868 4820
rect 6276 4811 6328 4820
rect 6276 4777 6285 4811
rect 6285 4777 6319 4811
rect 6319 4777 6328 4811
rect 6276 4768 6328 4777
rect 7564 4768 7616 4820
rect 8668 4768 8720 4820
rect 9036 4768 9088 4820
rect 3240 4700 3292 4752
rect 2596 4675 2648 4684
rect 2596 4641 2605 4675
rect 2605 4641 2639 4675
rect 2639 4641 2648 4675
rect 3332 4675 3384 4684
rect 2596 4632 2648 4641
rect 3332 4641 3341 4675
rect 3341 4641 3375 4675
rect 3375 4641 3384 4675
rect 3332 4632 3384 4641
rect 4068 4632 4120 4684
rect 4804 4700 4856 4752
rect 5356 4700 5408 4752
rect 5724 4675 5776 4684
rect 940 4564 992 4616
rect 2412 4607 2464 4616
rect 2412 4573 2421 4607
rect 2421 4573 2455 4607
rect 2455 4573 2464 4607
rect 2412 4564 2464 4573
rect 5724 4641 5733 4675
rect 5733 4641 5767 4675
rect 5767 4641 5776 4675
rect 5724 4632 5776 4641
rect 5816 4675 5868 4684
rect 5816 4641 5825 4675
rect 5825 4641 5859 4675
rect 5859 4641 5868 4675
rect 5816 4632 5868 4641
rect 6828 4632 6880 4684
rect 7472 4632 7524 4684
rect 8208 4632 8260 4684
rect 8484 4700 8536 4752
rect 9956 4768 10008 4820
rect 10600 4811 10652 4820
rect 10600 4777 10609 4811
rect 10609 4777 10643 4811
rect 10643 4777 10652 4811
rect 10600 4768 10652 4777
rect 10784 4768 10836 4820
rect 12440 4768 12492 4820
rect 12992 4768 13044 4820
rect 5080 4564 5132 4616
rect 6368 4564 6420 4616
rect 6644 4564 6696 4616
rect 1768 4496 1820 4548
rect 2228 4496 2280 4548
rect 2596 4496 2648 4548
rect 4436 4496 4488 4548
rect 1032 4428 1084 4480
rect 1400 4428 1452 4480
rect 2044 4471 2096 4480
rect 2044 4437 2053 4471
rect 2053 4437 2087 4471
rect 2087 4437 2096 4471
rect 2044 4428 2096 4437
rect 2412 4428 2464 4480
rect 4804 4428 4856 4480
rect 5080 4428 5132 4480
rect 5908 4496 5960 4548
rect 6184 4539 6236 4548
rect 6184 4505 6193 4539
rect 6193 4505 6227 4539
rect 6227 4505 6236 4539
rect 6184 4496 6236 4505
rect 5632 4428 5684 4480
rect 8668 4564 8720 4616
rect 9680 4632 9732 4684
rect 9772 4632 9824 4684
rect 11152 4675 11204 4684
rect 11152 4641 11161 4675
rect 11161 4641 11195 4675
rect 11195 4641 11204 4675
rect 11152 4632 11204 4641
rect 10232 4607 10284 4616
rect 10232 4573 10241 4607
rect 10241 4573 10275 4607
rect 10275 4573 10284 4607
rect 10968 4607 11020 4616
rect 10232 4564 10284 4573
rect 10968 4573 10977 4607
rect 10977 4573 11011 4607
rect 11011 4573 11020 4607
rect 10968 4564 11020 4573
rect 7656 4496 7708 4548
rect 7840 4471 7892 4480
rect 7840 4437 7849 4471
rect 7849 4437 7883 4471
rect 7883 4437 7892 4471
rect 7840 4428 7892 4437
rect 7932 4471 7984 4480
rect 7932 4437 7941 4471
rect 7941 4437 7975 4471
rect 7975 4437 7984 4471
rect 7932 4428 7984 4437
rect 8944 4428 8996 4480
rect 9220 4428 9272 4480
rect 13084 4743 13136 4752
rect 13084 4709 13093 4743
rect 13093 4709 13127 4743
rect 13127 4709 13136 4743
rect 13084 4700 13136 4709
rect 11980 4675 12032 4684
rect 11980 4641 11989 4675
rect 11989 4641 12023 4675
rect 12023 4641 12032 4675
rect 11980 4632 12032 4641
rect 12716 4632 12768 4684
rect 12992 4632 13044 4684
rect 13360 4632 13412 4684
rect 13728 4675 13780 4684
rect 13728 4641 13737 4675
rect 13737 4641 13771 4675
rect 13771 4641 13780 4675
rect 17684 4768 17736 4820
rect 18236 4768 18288 4820
rect 18880 4768 18932 4820
rect 13728 4632 13780 4641
rect 14464 4675 14516 4684
rect 14464 4641 14473 4675
rect 14473 4641 14507 4675
rect 14507 4641 14516 4675
rect 14464 4632 14516 4641
rect 16304 4632 16356 4684
rect 16948 4632 17000 4684
rect 17684 4675 17736 4684
rect 17684 4641 17693 4675
rect 17693 4641 17727 4675
rect 17727 4641 17736 4675
rect 17684 4632 17736 4641
rect 18052 4632 18104 4684
rect 22008 4700 22060 4752
rect 22652 4700 22704 4752
rect 18880 4675 18932 4684
rect 18880 4641 18889 4675
rect 18889 4641 18923 4675
rect 18923 4641 18932 4675
rect 18880 4632 18932 4641
rect 19616 4632 19668 4684
rect 21916 4632 21968 4684
rect 12900 4564 12952 4616
rect 13084 4564 13136 4616
rect 14556 4564 14608 4616
rect 15292 4607 15344 4616
rect 15292 4573 15301 4607
rect 15301 4573 15335 4607
rect 15335 4573 15344 4607
rect 15292 4564 15344 4573
rect 15568 4564 15620 4616
rect 16396 4564 16448 4616
rect 16580 4564 16632 4616
rect 20996 4607 21048 4616
rect 20996 4573 21005 4607
rect 21005 4573 21039 4607
rect 21039 4573 21048 4607
rect 20996 4564 21048 4573
rect 12532 4496 12584 4548
rect 12716 4539 12768 4548
rect 12716 4505 12725 4539
rect 12725 4505 12759 4539
rect 12759 4505 12768 4539
rect 12716 4496 12768 4505
rect 15108 4496 15160 4548
rect 11980 4428 12032 4480
rect 13176 4471 13228 4480
rect 13176 4437 13185 4471
rect 13185 4437 13219 4471
rect 13219 4437 13228 4471
rect 13176 4428 13228 4437
rect 14556 4471 14608 4480
rect 14556 4437 14565 4471
rect 14565 4437 14599 4471
rect 14599 4437 14608 4471
rect 14556 4428 14608 4437
rect 15752 4471 15804 4480
rect 15752 4437 15761 4471
rect 15761 4437 15795 4471
rect 15795 4437 15804 4471
rect 15752 4428 15804 4437
rect 16120 4496 16172 4548
rect 16948 4496 17000 4548
rect 17224 4496 17276 4548
rect 17776 4496 17828 4548
rect 16396 4428 16448 4480
rect 16764 4428 16816 4480
rect 17960 4428 18012 4480
rect 18328 4471 18380 4480
rect 18328 4437 18337 4471
rect 18337 4437 18371 4471
rect 18371 4437 18380 4471
rect 18328 4428 18380 4437
rect 18604 4428 18656 4480
rect 19524 4471 19576 4480
rect 19524 4437 19533 4471
rect 19533 4437 19567 4471
rect 19567 4437 19576 4471
rect 19524 4428 19576 4437
rect 19616 4471 19668 4480
rect 19616 4437 19625 4471
rect 19625 4437 19659 4471
rect 19659 4437 19668 4471
rect 19984 4471 20036 4480
rect 19616 4428 19668 4437
rect 19984 4437 19993 4471
rect 19993 4437 20027 4471
rect 20027 4437 20036 4471
rect 19984 4428 20036 4437
rect 20076 4471 20128 4480
rect 20076 4437 20085 4471
rect 20085 4437 20119 4471
rect 20119 4437 20128 4471
rect 20076 4428 20128 4437
rect 6148 4326 6200 4378
rect 6212 4326 6264 4378
rect 6276 4326 6328 4378
rect 6340 4326 6392 4378
rect 6404 4326 6456 4378
rect 11346 4326 11398 4378
rect 11410 4326 11462 4378
rect 11474 4326 11526 4378
rect 11538 4326 11590 4378
rect 11602 4326 11654 4378
rect 16544 4326 16596 4378
rect 16608 4326 16660 4378
rect 16672 4326 16724 4378
rect 16736 4326 16788 4378
rect 16800 4326 16852 4378
rect 21742 4326 21794 4378
rect 21806 4326 21858 4378
rect 21870 4326 21922 4378
rect 21934 4326 21986 4378
rect 21998 4326 22050 4378
rect 2044 4224 2096 4276
rect 4160 4267 4212 4276
rect 4160 4233 4169 4267
rect 4169 4233 4203 4267
rect 4203 4233 4212 4267
rect 4160 4224 4212 4233
rect 4436 4224 4488 4276
rect 5816 4267 5868 4276
rect 5816 4233 5825 4267
rect 5825 4233 5859 4267
rect 5859 4233 5868 4267
rect 5816 4224 5868 4233
rect 6092 4224 6144 4276
rect 5264 4156 5316 4208
rect 5356 4156 5408 4208
rect 6920 4224 6972 4276
rect 7104 4224 7156 4276
rect 11980 4224 12032 4276
rect 12532 4267 12584 4276
rect 1492 4088 1544 4140
rect 1676 3995 1728 4004
rect 1676 3961 1685 3995
rect 1685 3961 1719 3995
rect 1719 3961 1728 3995
rect 1676 3952 1728 3961
rect 2780 4131 2832 4140
rect 2780 4097 2789 4131
rect 2789 4097 2823 4131
rect 2823 4097 2832 4131
rect 2780 4088 2832 4097
rect 3332 4088 3384 4140
rect 4252 4131 4304 4140
rect 4252 4097 4261 4131
rect 4261 4097 4295 4131
rect 4295 4097 4304 4131
rect 4252 4088 4304 4097
rect 4988 4131 5040 4140
rect 4988 4097 4997 4131
rect 4997 4097 5031 4131
rect 5031 4097 5040 4131
rect 4988 4088 5040 4097
rect 6368 4131 6420 4140
rect 2136 4063 2188 4072
rect 2136 4029 2145 4063
rect 2145 4029 2179 4063
rect 2179 4029 2188 4063
rect 2136 4020 2188 4029
rect 5080 4063 5132 4072
rect 5080 4029 5089 4063
rect 5089 4029 5123 4063
rect 5123 4029 5132 4063
rect 5080 4020 5132 4029
rect 2688 3995 2740 4004
rect 2688 3961 2697 3995
rect 2697 3961 2731 3995
rect 2731 3961 2740 3995
rect 2688 3952 2740 3961
rect 4252 3952 4304 4004
rect 4896 3952 4948 4004
rect 6000 4063 6052 4072
rect 6000 4029 6009 4063
rect 6009 4029 6043 4063
rect 6043 4029 6052 4063
rect 6000 4020 6052 4029
rect 6368 4097 6377 4131
rect 6377 4097 6411 4131
rect 6411 4097 6420 4131
rect 6368 4088 6420 4097
rect 6736 4088 6788 4140
rect 7196 4156 7248 4208
rect 7380 4156 7432 4208
rect 7472 4156 7524 4208
rect 7932 4156 7984 4208
rect 8116 4156 8168 4208
rect 9036 4199 9088 4208
rect 9036 4165 9045 4199
rect 9045 4165 9079 4199
rect 9079 4165 9088 4199
rect 9036 4156 9088 4165
rect 11244 4156 11296 4208
rect 12532 4233 12541 4267
rect 12541 4233 12575 4267
rect 12575 4233 12584 4267
rect 12532 4224 12584 4233
rect 13176 4224 13228 4276
rect 13452 4224 13504 4276
rect 12440 4156 12492 4208
rect 7564 4088 7616 4140
rect 8392 4088 8444 4140
rect 9588 4131 9640 4140
rect 9588 4097 9597 4131
rect 9597 4097 9631 4131
rect 9631 4097 9640 4131
rect 9588 4088 9640 4097
rect 10324 4088 10376 4140
rect 11612 4131 11664 4140
rect 7012 4063 7064 4072
rect 7012 4029 7021 4063
rect 7021 4029 7055 4063
rect 7055 4029 7064 4063
rect 7012 4020 7064 4029
rect 9680 4020 9732 4072
rect 10232 4063 10284 4072
rect 10232 4029 10241 4063
rect 10241 4029 10275 4063
rect 10275 4029 10284 4063
rect 10232 4020 10284 4029
rect 5540 3952 5592 4004
rect 6644 3952 6696 4004
rect 8208 3952 8260 4004
rect 8576 3995 8628 4004
rect 8576 3961 8585 3995
rect 8585 3961 8619 3995
rect 8619 3961 8628 3995
rect 8576 3952 8628 3961
rect 11612 4097 11621 4131
rect 11621 4097 11655 4131
rect 11655 4097 11664 4131
rect 11612 4088 11664 4097
rect 12072 4088 12124 4140
rect 13268 4088 13320 4140
rect 15108 4224 15160 4276
rect 15936 4267 15988 4276
rect 15936 4233 15945 4267
rect 15945 4233 15979 4267
rect 15979 4233 15988 4267
rect 15936 4224 15988 4233
rect 16396 4156 16448 4208
rect 17684 4224 17736 4276
rect 18420 4224 18472 4276
rect 20076 4224 20128 4276
rect 17040 4156 17092 4208
rect 18236 4156 18288 4208
rect 19800 4156 19852 4208
rect 4620 3927 4672 3936
rect 4620 3893 4629 3927
rect 4629 3893 4663 3927
rect 4663 3893 4672 3927
rect 6552 3927 6604 3936
rect 4620 3884 4672 3893
rect 6552 3893 6561 3927
rect 6561 3893 6595 3927
rect 6595 3893 6604 3927
rect 6552 3884 6604 3893
rect 6736 3884 6788 3936
rect 10508 3952 10560 4004
rect 12992 4020 13044 4072
rect 13176 4063 13228 4072
rect 13176 4029 13185 4063
rect 13185 4029 13219 4063
rect 13219 4029 13228 4063
rect 13176 4020 13228 4029
rect 13544 4020 13596 4072
rect 8944 3884 8996 3936
rect 9220 3884 9272 3936
rect 9496 3927 9548 3936
rect 9496 3893 9505 3927
rect 9505 3893 9539 3927
rect 9539 3893 9548 3927
rect 9496 3884 9548 3893
rect 9680 3884 9732 3936
rect 10692 3884 10744 3936
rect 13728 3952 13780 4004
rect 14280 4020 14332 4072
rect 15292 4063 15344 4072
rect 15292 4029 15301 4063
rect 15301 4029 15335 4063
rect 15335 4029 15344 4063
rect 15292 4020 15344 4029
rect 17224 4131 17276 4140
rect 17224 4097 17258 4131
rect 17258 4097 17276 4131
rect 17224 4088 17276 4097
rect 18880 4088 18932 4140
rect 15844 4063 15896 4072
rect 15844 4029 15853 4063
rect 15853 4029 15887 4063
rect 15887 4029 15896 4063
rect 16396 4063 16448 4072
rect 15844 4020 15896 4029
rect 16396 4029 16405 4063
rect 16405 4029 16439 4063
rect 16439 4029 16448 4063
rect 16396 4020 16448 4029
rect 18420 4020 18472 4072
rect 18696 4063 18748 4072
rect 18696 4029 18705 4063
rect 18705 4029 18739 4063
rect 18739 4029 18748 4063
rect 18696 4020 18748 4029
rect 19064 4020 19116 4072
rect 19984 4088 20036 4140
rect 20352 4088 20404 4140
rect 15016 3952 15068 4004
rect 12072 3927 12124 3936
rect 12072 3893 12081 3927
rect 12081 3893 12115 3927
rect 12115 3893 12124 3927
rect 12072 3884 12124 3893
rect 12348 3927 12400 3936
rect 12348 3893 12357 3927
rect 12357 3893 12391 3927
rect 12391 3893 12400 3927
rect 12348 3884 12400 3893
rect 12992 3927 13044 3936
rect 12992 3893 13001 3927
rect 13001 3893 13035 3927
rect 13035 3893 13044 3927
rect 12992 3884 13044 3893
rect 14464 3884 14516 3936
rect 14556 3884 14608 3936
rect 16304 3927 16356 3936
rect 16304 3893 16313 3927
rect 16313 3893 16347 3927
rect 16347 3893 16356 3927
rect 16304 3884 16356 3893
rect 16856 3927 16908 3936
rect 16856 3893 16865 3927
rect 16865 3893 16899 3927
rect 16899 3893 16908 3927
rect 16856 3884 16908 3893
rect 19616 3952 19668 4004
rect 20812 4020 20864 4072
rect 19984 3952 20036 4004
rect 20444 3884 20496 3936
rect 3549 3782 3601 3834
rect 3613 3782 3665 3834
rect 3677 3782 3729 3834
rect 3741 3782 3793 3834
rect 3805 3782 3857 3834
rect 8747 3782 8799 3834
rect 8811 3782 8863 3834
rect 8875 3782 8927 3834
rect 8939 3782 8991 3834
rect 9003 3782 9055 3834
rect 13945 3782 13997 3834
rect 14009 3782 14061 3834
rect 14073 3782 14125 3834
rect 14137 3782 14189 3834
rect 14201 3782 14253 3834
rect 19143 3782 19195 3834
rect 19207 3782 19259 3834
rect 19271 3782 19323 3834
rect 19335 3782 19387 3834
rect 19399 3782 19451 3834
rect 756 3612 808 3664
rect 1952 3612 2004 3664
rect 3332 3655 3384 3664
rect 3332 3621 3341 3655
rect 3341 3621 3375 3655
rect 3375 3621 3384 3655
rect 3332 3612 3384 3621
rect 3516 3680 3568 3732
rect 5172 3723 5224 3732
rect 5172 3689 5181 3723
rect 5181 3689 5215 3723
rect 5215 3689 5224 3723
rect 5172 3680 5224 3689
rect 5908 3680 5960 3732
rect 3792 3612 3844 3664
rect 6000 3612 6052 3664
rect 7840 3680 7892 3732
rect 7932 3680 7984 3732
rect 10324 3680 10376 3732
rect 11612 3680 11664 3732
rect 12164 3680 12216 3732
rect 13268 3680 13320 3732
rect 16120 3680 16172 3732
rect 16304 3680 16356 3732
rect 6828 3612 6880 3664
rect 1400 3519 1452 3528
rect 1400 3485 1409 3519
rect 1409 3485 1443 3519
rect 1443 3485 1452 3519
rect 1400 3476 1452 3485
rect 1216 3408 1268 3460
rect 2780 3476 2832 3528
rect 3424 3519 3476 3528
rect 3424 3485 3433 3519
rect 3433 3485 3467 3519
rect 3467 3485 3476 3519
rect 3424 3476 3476 3485
rect 6276 3544 6328 3596
rect 8208 3612 8260 3664
rect 8300 3587 8352 3596
rect 8300 3553 8309 3587
rect 8309 3553 8343 3587
rect 8343 3553 8352 3587
rect 8300 3544 8352 3553
rect 10876 3612 10928 3664
rect 12440 3612 12492 3664
rect 13544 3612 13596 3664
rect 7840 3519 7892 3528
rect 1584 3383 1636 3392
rect 1584 3349 1593 3383
rect 1593 3349 1627 3383
rect 1627 3349 1636 3383
rect 1584 3340 1636 3349
rect 2504 3408 2556 3460
rect 4160 3408 4212 3460
rect 4712 3408 4764 3460
rect 5356 3451 5408 3460
rect 5356 3417 5365 3451
rect 5365 3417 5399 3451
rect 5399 3417 5408 3451
rect 5356 3408 5408 3417
rect 5448 3408 5500 3460
rect 6644 3408 6696 3460
rect 7840 3485 7849 3519
rect 7849 3485 7883 3519
rect 7883 3485 7892 3519
rect 7840 3476 7892 3485
rect 8024 3476 8076 3528
rect 8944 3519 8996 3528
rect 8944 3485 8953 3519
rect 8953 3485 8987 3519
rect 8987 3485 8996 3519
rect 8944 3476 8996 3485
rect 14556 3587 14608 3596
rect 10508 3476 10560 3528
rect 10876 3476 10928 3528
rect 14556 3553 14565 3587
rect 14565 3553 14599 3587
rect 14599 3553 14608 3587
rect 14556 3544 14608 3553
rect 15292 3612 15344 3664
rect 13268 3476 13320 3528
rect 13636 3476 13688 3528
rect 3056 3340 3108 3392
rect 3884 3340 3936 3392
rect 4252 3340 4304 3392
rect 5264 3340 5316 3392
rect 5908 3383 5960 3392
rect 5908 3349 5917 3383
rect 5917 3349 5951 3383
rect 5951 3349 5960 3383
rect 5908 3340 5960 3349
rect 6000 3383 6052 3392
rect 6000 3349 6009 3383
rect 6009 3349 6043 3383
rect 6043 3349 6052 3383
rect 6000 3340 6052 3349
rect 6276 3340 6328 3392
rect 7380 3340 7432 3392
rect 10140 3408 10192 3460
rect 10692 3408 10744 3460
rect 7748 3340 7800 3392
rect 8024 3340 8076 3392
rect 8392 3383 8444 3392
rect 8392 3349 8401 3383
rect 8401 3349 8435 3383
rect 8435 3349 8444 3383
rect 8392 3340 8444 3349
rect 9404 3340 9456 3392
rect 10232 3340 10284 3392
rect 13176 3408 13228 3460
rect 14740 3476 14792 3528
rect 17224 3544 17276 3596
rect 18696 3680 18748 3732
rect 20720 3680 20772 3732
rect 18420 3612 18472 3664
rect 18788 3612 18840 3664
rect 18328 3587 18380 3596
rect 15016 3408 15068 3460
rect 13544 3340 13596 3392
rect 13912 3383 13964 3392
rect 13912 3349 13921 3383
rect 13921 3349 13955 3383
rect 13955 3349 13964 3383
rect 13912 3340 13964 3349
rect 14188 3340 14240 3392
rect 14280 3340 14332 3392
rect 15200 3383 15252 3392
rect 15200 3349 15209 3383
rect 15209 3349 15243 3383
rect 15243 3349 15252 3383
rect 17040 3519 17092 3528
rect 17040 3485 17049 3519
rect 17049 3485 17083 3519
rect 17083 3485 17092 3519
rect 18328 3553 18337 3587
rect 18337 3553 18371 3587
rect 18371 3553 18380 3587
rect 18328 3544 18380 3553
rect 17040 3476 17092 3485
rect 16028 3408 16080 3460
rect 16396 3408 16448 3460
rect 16856 3408 16908 3460
rect 17868 3408 17920 3460
rect 18236 3476 18288 3528
rect 18880 3476 18932 3528
rect 19064 3519 19116 3528
rect 19064 3485 19073 3519
rect 19073 3485 19107 3519
rect 19107 3485 19116 3519
rect 19064 3476 19116 3485
rect 18696 3408 18748 3460
rect 15200 3340 15252 3349
rect 15752 3340 15804 3392
rect 16304 3340 16356 3392
rect 17132 3340 17184 3392
rect 17500 3340 17552 3392
rect 17684 3340 17736 3392
rect 18144 3340 18196 3392
rect 19432 3408 19484 3460
rect 19892 3476 19944 3528
rect 20260 3612 20312 3664
rect 21364 3612 21416 3664
rect 20904 3544 20956 3596
rect 20352 3519 20404 3528
rect 20352 3485 20361 3519
rect 20361 3485 20395 3519
rect 20395 3485 20404 3519
rect 20352 3476 20404 3485
rect 22100 3476 22152 3528
rect 20812 3451 20864 3460
rect 18880 3383 18932 3392
rect 18880 3349 18889 3383
rect 18889 3349 18923 3383
rect 18923 3349 18932 3383
rect 19892 3383 19944 3392
rect 18880 3340 18932 3349
rect 19892 3349 19901 3383
rect 19901 3349 19935 3383
rect 19935 3349 19944 3383
rect 19892 3340 19944 3349
rect 20812 3417 20821 3451
rect 20821 3417 20855 3451
rect 20855 3417 20864 3451
rect 20812 3408 20864 3417
rect 21088 3408 21140 3460
rect 20720 3340 20772 3392
rect 6148 3238 6200 3290
rect 6212 3238 6264 3290
rect 6276 3238 6328 3290
rect 6340 3238 6392 3290
rect 6404 3238 6456 3290
rect 11346 3238 11398 3290
rect 11410 3238 11462 3290
rect 11474 3238 11526 3290
rect 11538 3238 11590 3290
rect 11602 3238 11654 3290
rect 16544 3238 16596 3290
rect 16608 3238 16660 3290
rect 16672 3238 16724 3290
rect 16736 3238 16788 3290
rect 16800 3238 16852 3290
rect 21742 3238 21794 3290
rect 21806 3238 21858 3290
rect 21870 3238 21922 3290
rect 21934 3238 21986 3290
rect 21998 3238 22050 3290
rect 2412 3179 2464 3188
rect 2412 3145 2421 3179
rect 2421 3145 2455 3179
rect 2455 3145 2464 3179
rect 2412 3136 2464 3145
rect 4620 3136 4672 3188
rect 4712 3136 4764 3188
rect 5816 3136 5868 3188
rect 5908 3136 5960 3188
rect 6552 3136 6604 3188
rect 6828 3136 6880 3188
rect 7012 3136 7064 3188
rect 7840 3136 7892 3188
rect 7932 3136 7984 3188
rect 9404 3179 9456 3188
rect 1124 3068 1176 3120
rect 4068 3068 4120 3120
rect 2688 3000 2740 3052
rect 3332 3043 3384 3052
rect 3332 3009 3341 3043
rect 3341 3009 3375 3043
rect 3375 3009 3384 3043
rect 3332 3000 3384 3009
rect 2504 2932 2556 2984
rect 3516 2932 3568 2984
rect 4160 2932 4212 2984
rect 1860 2864 1912 2916
rect 1768 2839 1820 2848
rect 1768 2805 1777 2839
rect 1777 2805 1811 2839
rect 1811 2805 1820 2839
rect 1768 2796 1820 2805
rect 2044 2839 2096 2848
rect 2044 2805 2053 2839
rect 2053 2805 2087 2839
rect 2087 2805 2096 2839
rect 2044 2796 2096 2805
rect 2136 2796 2188 2848
rect 4252 2796 4304 2848
rect 4896 3000 4948 3052
rect 5448 3068 5500 3120
rect 6736 3000 6788 3052
rect 6920 3000 6972 3052
rect 7288 2932 7340 2984
rect 7656 3043 7708 3052
rect 7656 3009 7665 3043
rect 7665 3009 7699 3043
rect 7699 3009 7708 3043
rect 7656 3000 7708 3009
rect 7472 2932 7524 2984
rect 8300 2932 8352 2984
rect 8576 2975 8628 2984
rect 8576 2941 8585 2975
rect 8585 2941 8619 2975
rect 8619 2941 8628 2975
rect 9404 3145 9413 3179
rect 9413 3145 9447 3179
rect 9447 3145 9456 3179
rect 9404 3136 9456 3145
rect 10324 3136 10376 3188
rect 9220 3068 9272 3120
rect 9772 3068 9824 3120
rect 12348 3136 12400 3188
rect 13544 3136 13596 3188
rect 14280 3179 14332 3188
rect 14280 3145 14289 3179
rect 14289 3145 14323 3179
rect 14323 3145 14332 3179
rect 14280 3136 14332 3145
rect 14464 3136 14516 3188
rect 16396 3136 16448 3188
rect 10232 3043 10284 3052
rect 8576 2932 8628 2941
rect 8944 2932 8996 2984
rect 10232 3009 10255 3043
rect 10255 3009 10284 3043
rect 10232 3000 10284 3009
rect 11888 3009 11897 3036
rect 11897 3009 11931 3036
rect 11931 3009 11940 3036
rect 11888 2984 11940 3009
rect 4620 2864 4672 2916
rect 5816 2864 5868 2916
rect 7932 2864 7984 2916
rect 8208 2864 8260 2916
rect 9864 2932 9916 2984
rect 11060 2932 11112 2984
rect 5540 2796 5592 2848
rect 7196 2796 7248 2848
rect 7840 2796 7892 2848
rect 8116 2839 8168 2848
rect 8116 2805 8125 2839
rect 8125 2805 8159 2839
rect 8159 2805 8168 2839
rect 8116 2796 8168 2805
rect 8300 2796 8352 2848
rect 10968 2864 11020 2916
rect 12532 3068 12584 3120
rect 12348 3043 12400 3052
rect 12348 3009 12357 3043
rect 12357 3009 12391 3043
rect 12391 3009 12400 3043
rect 12348 3000 12400 3009
rect 11244 2796 11296 2848
rect 12808 2932 12860 2984
rect 12532 2839 12584 2848
rect 12532 2805 12541 2839
rect 12541 2805 12575 2839
rect 12575 2805 12584 2839
rect 12532 2796 12584 2805
rect 13912 3043 13964 3052
rect 13912 3009 13941 3043
rect 13941 3009 13964 3043
rect 13912 3000 13964 3009
rect 14832 3068 14884 3120
rect 14648 3043 14700 3052
rect 14648 3009 14657 3043
rect 14657 3009 14691 3043
rect 14691 3009 14700 3043
rect 14648 3000 14700 3009
rect 15660 3068 15712 3120
rect 15476 3000 15528 3052
rect 16120 3043 16172 3052
rect 16120 3009 16129 3043
rect 16129 3009 16163 3043
rect 16163 3009 16172 3043
rect 16120 3000 16172 3009
rect 14280 2932 14332 2984
rect 15016 2932 15068 2984
rect 16488 3000 16540 3052
rect 16948 3043 17000 3052
rect 16948 3009 16957 3043
rect 16957 3009 16991 3043
rect 16991 3009 17000 3043
rect 16948 3000 17000 3009
rect 17316 3000 17368 3052
rect 17592 3136 17644 3188
rect 18144 3179 18196 3188
rect 18144 3145 18153 3179
rect 18153 3145 18187 3179
rect 18187 3145 18196 3179
rect 18144 3136 18196 3145
rect 17960 3068 18012 3120
rect 18880 3068 18932 3120
rect 19524 3068 19576 3120
rect 16764 2932 16816 2984
rect 17868 3000 17920 3052
rect 18604 2975 18656 2984
rect 18604 2941 18613 2975
rect 18613 2941 18647 2975
rect 18647 2941 18656 2975
rect 18604 2932 18656 2941
rect 18696 2975 18748 2984
rect 18696 2941 18705 2975
rect 18705 2941 18739 2975
rect 18739 2941 18748 2975
rect 18696 2932 18748 2941
rect 19800 2932 19852 2984
rect 20076 3043 20128 3052
rect 20076 3009 20085 3043
rect 20085 3009 20119 3043
rect 20119 3009 20128 3043
rect 20076 3000 20128 3009
rect 20444 3043 20496 3052
rect 20444 3009 20453 3043
rect 20453 3009 20487 3043
rect 20487 3009 20496 3043
rect 20444 3000 20496 3009
rect 22192 3136 22244 3188
rect 22284 3068 22336 3120
rect 22376 3000 22428 3052
rect 21180 2932 21232 2984
rect 15384 2864 15436 2916
rect 15660 2864 15712 2916
rect 14372 2796 14424 2848
rect 15476 2796 15528 2848
rect 15936 2839 15988 2848
rect 15936 2805 15945 2839
rect 15945 2805 15979 2839
rect 15979 2805 15988 2839
rect 15936 2796 15988 2805
rect 19616 2864 19668 2916
rect 20628 2864 20680 2916
rect 16672 2839 16724 2848
rect 16672 2805 16681 2839
rect 16681 2805 16715 2839
rect 16715 2805 16724 2839
rect 16672 2796 16724 2805
rect 17224 2839 17276 2848
rect 17224 2805 17233 2839
rect 17233 2805 17267 2839
rect 17267 2805 17276 2839
rect 17224 2796 17276 2805
rect 18052 2796 18104 2848
rect 18696 2796 18748 2848
rect 18880 2796 18932 2848
rect 18972 2796 19024 2848
rect 19064 2796 19116 2848
rect 20352 2796 20404 2848
rect 21364 2796 21416 2848
rect 3549 2694 3601 2746
rect 3613 2694 3665 2746
rect 3677 2694 3729 2746
rect 3741 2694 3793 2746
rect 3805 2694 3857 2746
rect 8747 2694 8799 2746
rect 8811 2694 8863 2746
rect 8875 2694 8927 2746
rect 8939 2694 8991 2746
rect 9003 2694 9055 2746
rect 13945 2694 13997 2746
rect 14009 2694 14061 2746
rect 14073 2694 14125 2746
rect 14137 2694 14189 2746
rect 14201 2694 14253 2746
rect 19143 2694 19195 2746
rect 19207 2694 19259 2746
rect 19271 2694 19323 2746
rect 19335 2694 19387 2746
rect 19399 2694 19451 2746
rect 2780 2592 2832 2644
rect 4252 2592 4304 2644
rect 5632 2635 5684 2644
rect 5632 2601 5641 2635
rect 5641 2601 5675 2635
rect 5675 2601 5684 2635
rect 5632 2592 5684 2601
rect 6828 2592 6880 2644
rect 7472 2635 7524 2644
rect 7472 2601 7481 2635
rect 7481 2601 7515 2635
rect 7515 2601 7524 2635
rect 7472 2592 7524 2601
rect 7656 2635 7708 2644
rect 7656 2601 7665 2635
rect 7665 2601 7699 2635
rect 7699 2601 7708 2635
rect 7656 2592 7708 2601
rect 8024 2592 8076 2644
rect 3240 2524 3292 2576
rect 3608 2567 3660 2576
rect 3608 2533 3617 2567
rect 3617 2533 3651 2567
rect 3651 2533 3660 2567
rect 3608 2524 3660 2533
rect 3700 2524 3752 2576
rect 3976 2524 4028 2576
rect 4160 2567 4212 2576
rect 4160 2533 4169 2567
rect 4169 2533 4203 2567
rect 4203 2533 4212 2567
rect 4160 2524 4212 2533
rect 5540 2524 5592 2576
rect 5908 2524 5960 2576
rect 2044 2456 2096 2508
rect 2780 2388 2832 2440
rect 2688 2320 2740 2372
rect 3608 2320 3660 2372
rect 3976 2363 4028 2372
rect 3976 2329 3985 2363
rect 3985 2329 4019 2363
rect 4019 2329 4028 2363
rect 3976 2320 4028 2329
rect 5264 2456 5316 2508
rect 4896 2388 4948 2440
rect 6000 2388 6052 2440
rect 7104 2456 7156 2508
rect 8300 2524 8352 2576
rect 7380 2456 7432 2508
rect 8208 2499 8260 2508
rect 8208 2465 8217 2499
rect 8217 2465 8251 2499
rect 8251 2465 8260 2499
rect 8208 2456 8260 2465
rect 9864 2592 9916 2644
rect 10876 2592 10928 2644
rect 11152 2592 11204 2644
rect 14648 2592 14700 2644
rect 15844 2592 15896 2644
rect 17684 2592 17736 2644
rect 20076 2592 20128 2644
rect 8668 2567 8720 2576
rect 8668 2533 8677 2567
rect 8677 2533 8711 2567
rect 8711 2533 8720 2567
rect 8668 2524 8720 2533
rect 9772 2524 9824 2576
rect 12348 2567 12400 2576
rect 12348 2533 12357 2567
rect 12357 2533 12391 2567
rect 12391 2533 12400 2567
rect 12348 2524 12400 2533
rect 13636 2524 13688 2576
rect 15108 2524 15160 2576
rect 16212 2524 16264 2576
rect 17316 2524 17368 2576
rect 18420 2524 18472 2576
rect 18604 2524 18656 2576
rect 4620 2320 4672 2372
rect 5816 2252 5868 2304
rect 6644 2320 6696 2372
rect 6736 2320 6788 2372
rect 7656 2320 7708 2372
rect 8116 2388 8168 2440
rect 8392 2388 8444 2440
rect 8668 2388 8720 2440
rect 9404 2431 9456 2440
rect 9404 2397 9413 2431
rect 9413 2397 9447 2431
rect 9447 2397 9456 2431
rect 9404 2388 9456 2397
rect 12072 2456 12124 2508
rect 9956 2388 10008 2440
rect 11704 2388 11756 2440
rect 11888 2431 11940 2440
rect 11888 2397 11897 2431
rect 11897 2397 11931 2431
rect 11931 2397 11940 2431
rect 11888 2388 11940 2397
rect 12348 2388 12400 2440
rect 13176 2456 13228 2508
rect 13360 2431 13412 2440
rect 9312 2295 9364 2304
rect 9312 2261 9321 2295
rect 9321 2261 9355 2295
rect 9355 2261 9364 2295
rect 9312 2252 9364 2261
rect 9496 2252 9548 2304
rect 10232 2252 10284 2304
rect 13360 2397 13369 2431
rect 13369 2397 13403 2431
rect 13403 2397 13412 2431
rect 13360 2388 13412 2397
rect 13728 2388 13780 2440
rect 15016 2388 15068 2440
rect 15936 2456 15988 2508
rect 15292 2431 15344 2440
rect 15292 2397 15301 2431
rect 15301 2397 15335 2431
rect 15335 2397 15344 2431
rect 15660 2431 15712 2440
rect 15292 2388 15344 2397
rect 15660 2397 15669 2431
rect 15669 2397 15703 2431
rect 15703 2397 15712 2431
rect 15660 2388 15712 2397
rect 16672 2388 16724 2440
rect 17224 2388 17276 2440
rect 18144 2456 18196 2508
rect 19800 2499 19852 2508
rect 19800 2465 19809 2499
rect 19809 2465 19843 2499
rect 19843 2465 19852 2499
rect 19800 2456 19852 2465
rect 22928 2456 22980 2508
rect 17960 2388 18012 2440
rect 10600 2295 10652 2304
rect 10600 2261 10609 2295
rect 10609 2261 10643 2295
rect 10643 2261 10652 2295
rect 12072 2295 12124 2304
rect 10600 2252 10652 2261
rect 12072 2261 12081 2295
rect 12081 2261 12115 2295
rect 12115 2261 12124 2295
rect 12072 2252 12124 2261
rect 12532 2252 12584 2304
rect 12900 2252 12952 2304
rect 13268 2252 13320 2304
rect 14004 2320 14056 2372
rect 13820 2252 13872 2304
rect 14464 2252 14516 2304
rect 14740 2320 14792 2372
rect 17040 2320 17092 2372
rect 18328 2388 18380 2440
rect 18512 2431 18564 2440
rect 18512 2397 18521 2431
rect 18521 2397 18555 2431
rect 18555 2397 18564 2431
rect 18512 2388 18564 2397
rect 18972 2388 19024 2440
rect 19708 2388 19760 2440
rect 20536 2388 20588 2440
rect 20720 2431 20772 2440
rect 20720 2397 20729 2431
rect 20729 2397 20763 2431
rect 20763 2397 20772 2431
rect 20720 2388 20772 2397
rect 21548 2388 21600 2440
rect 16396 2295 16448 2304
rect 16396 2261 16405 2295
rect 16405 2261 16439 2295
rect 16439 2261 16448 2295
rect 16396 2252 16448 2261
rect 16948 2252 17000 2304
rect 20168 2320 20220 2372
rect 21272 2252 21324 2304
rect 6148 2150 6200 2202
rect 6212 2150 6264 2202
rect 6276 2150 6328 2202
rect 6340 2150 6392 2202
rect 6404 2150 6456 2202
rect 11346 2150 11398 2202
rect 11410 2150 11462 2202
rect 11474 2150 11526 2202
rect 11538 2150 11590 2202
rect 11602 2150 11654 2202
rect 16544 2150 16596 2202
rect 16608 2150 16660 2202
rect 16672 2150 16724 2202
rect 16736 2150 16788 2202
rect 16800 2150 16852 2202
rect 21742 2150 21794 2202
rect 21806 2150 21858 2202
rect 21870 2150 21922 2202
rect 21934 2150 21986 2202
rect 21998 2150 22050 2202
rect 3976 2048 4028 2100
rect 1308 1980 1360 2032
rect 5264 1980 5316 2032
rect 5540 2048 5592 2100
rect 10232 2048 10284 2100
rect 11060 2048 11112 2100
rect 12348 2048 12400 2100
rect 16396 2048 16448 2100
rect 18328 2048 18380 2100
rect 19892 2048 19944 2100
rect 7380 1980 7432 2032
rect 7472 1980 7524 2032
rect 12256 1980 12308 2032
rect 12624 1980 12676 2032
rect 15660 1980 15712 2032
rect 17500 1980 17552 2032
rect 19800 1980 19852 2032
rect 1860 1912 1912 1964
rect 5448 1912 5500 1964
rect 5816 1912 5868 1964
rect 8576 1912 8628 1964
rect 14556 1912 14608 1964
rect 19248 1912 19300 1964
rect 6644 1844 6696 1896
rect 8852 1844 8904 1896
rect 10784 1844 10836 1896
rect 14924 1844 14976 1896
rect 19156 1844 19208 1896
rect 3792 1776 3844 1828
rect 7564 1776 7616 1828
rect 14464 1776 14516 1828
rect 19984 1776 20036 1828
rect 3608 1708 3660 1760
rect 6736 1708 6788 1760
rect 1492 1640 1544 1692
rect 9680 1640 9732 1692
rect 8116 1300 8168 1352
rect 10600 1300 10652 1352
rect 5080 1164 5132 1216
rect 17132 1300 17184 1352
rect 5724 1096 5776 1148
rect 16120 1232 16172 1284
rect 7472 76 7524 128
rect 22836 76 22888 128
rect 3976 8 4028 60
rect 20444 8 20496 60
<< metal2 >>
rect 124 22222 520 22250
rect 20 19440 72 19446
rect 20 19382 72 19388
rect 32 16318 60 19382
rect 20 16312 72 16318
rect 20 16254 72 16260
rect 124 15978 152 22222
rect 492 22114 520 22222
rect 570 22200 626 23000
rect 938 22200 994 23000
rect 1306 22200 1362 23000
rect 1674 22200 1730 23000
rect 2042 22200 2098 23000
rect 2318 22264 2374 22273
rect 584 22114 612 22200
rect 492 22086 612 22114
rect 952 19446 980 22200
rect 1122 21312 1178 21321
rect 1032 21276 1084 21282
rect 1122 21247 1178 21256
rect 1032 21218 1084 21224
rect 940 19440 992 19446
rect 940 19382 992 19388
rect 1044 16574 1072 21218
rect 1136 16726 1164 21247
rect 1216 21208 1268 21214
rect 1216 21150 1268 21156
rect 1124 16720 1176 16726
rect 1124 16662 1176 16668
rect 1044 16546 1164 16574
rect 940 16312 992 16318
rect 938 16280 940 16289
rect 992 16280 994 16289
rect 938 16215 994 16224
rect 112 15972 164 15978
rect 112 15914 164 15920
rect 938 14240 994 14249
rect 32 14198 938 14226
rect 32 6730 60 14198
rect 938 14175 994 14184
rect 938 13968 994 13977
rect 860 13926 938 13954
rect 204 13252 256 13258
rect 204 13194 256 13200
rect 20 6724 72 6730
rect 20 6666 72 6672
rect 216 5302 244 13194
rect 388 12708 440 12714
rect 388 12650 440 12656
rect 400 5506 428 12650
rect 756 10260 808 10266
rect 756 10202 808 10208
rect 572 10056 624 10062
rect 572 9998 624 10004
rect 584 6866 612 9998
rect 572 6860 624 6866
rect 572 6802 624 6808
rect 388 5500 440 5506
rect 388 5442 440 5448
rect 204 5296 256 5302
rect 204 5238 256 5244
rect 768 3670 796 10202
rect 756 3664 808 3670
rect 756 3606 808 3612
rect 860 3346 888 13926
rect 938 13903 994 13912
rect 1030 13424 1086 13433
rect 1030 13359 1086 13368
rect 938 13152 994 13161
rect 938 13087 994 13096
rect 952 10266 980 13087
rect 940 10260 992 10266
rect 940 10202 992 10208
rect 1044 10062 1072 13359
rect 1032 10056 1084 10062
rect 1032 9998 1084 10004
rect 940 6724 992 6730
rect 940 6666 992 6672
rect 952 6361 980 6666
rect 938 6352 994 6361
rect 938 6287 994 6296
rect 938 5536 994 5545
rect 938 5471 940 5480
rect 992 5471 994 5480
rect 940 5442 992 5448
rect 952 4622 980 5442
rect 1032 5296 1084 5302
rect 1032 5238 1084 5244
rect 1044 4729 1072 5238
rect 1030 4720 1086 4729
rect 1030 4655 1086 4664
rect 940 4616 992 4622
rect 940 4558 992 4564
rect 1032 4480 1084 4486
rect 1032 4422 1084 4428
rect 938 3360 994 3369
rect 860 3318 938 3346
rect 938 3295 994 3304
rect 1044 649 1072 4422
rect 1136 3126 1164 16546
rect 1228 3466 1256 21150
rect 1320 17513 1348 22200
rect 1584 21140 1636 21146
rect 1584 21082 1636 21088
rect 1492 20256 1544 20262
rect 1490 20224 1492 20233
rect 1544 20224 1546 20233
rect 1490 20159 1546 20168
rect 1492 19712 1544 19718
rect 1492 19654 1544 19660
rect 1504 19417 1532 19654
rect 1490 19408 1546 19417
rect 1400 19372 1452 19378
rect 1490 19343 1546 19352
rect 1400 19314 1452 19320
rect 1306 17504 1362 17513
rect 1306 17439 1362 17448
rect 1412 17338 1440 19314
rect 1492 19168 1544 19174
rect 1492 19110 1544 19116
rect 1504 19009 1532 19110
rect 1490 19000 1546 19009
rect 1490 18935 1546 18944
rect 1492 18624 1544 18630
rect 1490 18592 1492 18601
rect 1544 18592 1546 18601
rect 1490 18527 1546 18536
rect 1492 18080 1544 18086
rect 1492 18022 1544 18028
rect 1504 17785 1532 18022
rect 1596 17882 1624 21082
rect 1688 19394 1716 22200
rect 1766 21448 1822 21457
rect 1766 21383 1822 21392
rect 1780 19514 1808 21383
rect 2056 21146 2084 22200
rect 2318 22199 2374 22208
rect 2410 22200 2466 23000
rect 2778 22200 2834 23000
rect 3146 22200 3202 23000
rect 3514 22200 3570 23000
rect 3882 22200 3938 23000
rect 4250 22200 4306 23000
rect 4356 22222 4568 22250
rect 2044 21140 2096 21146
rect 2044 21082 2096 21088
rect 2226 21040 2282 21049
rect 2044 21004 2096 21010
rect 2226 20975 2282 20984
rect 2044 20946 2096 20952
rect 1952 20800 2004 20806
rect 1952 20742 2004 20748
rect 1858 20632 1914 20641
rect 1858 20567 1860 20576
rect 1912 20567 1914 20576
rect 1860 20538 1912 20544
rect 1964 20466 1992 20742
rect 2056 20466 2084 20946
rect 2134 20904 2190 20913
rect 2134 20839 2190 20848
rect 1952 20460 2004 20466
rect 1952 20402 2004 20408
rect 2044 20460 2096 20466
rect 2044 20402 2096 20408
rect 2148 20262 2176 20839
rect 2136 20256 2188 20262
rect 2134 20224 2136 20233
rect 2188 20224 2190 20233
rect 2134 20159 2190 20168
rect 2240 20058 2268 20975
rect 2332 20058 2360 22199
rect 2424 21298 2452 22200
rect 2424 21270 2544 21298
rect 2412 21140 2464 21146
rect 2412 21082 2464 21088
rect 2228 20052 2280 20058
rect 2228 19994 2280 20000
rect 2320 20052 2372 20058
rect 2320 19994 2372 20000
rect 2424 19854 2452 21082
rect 1952 19848 2004 19854
rect 1858 19816 1914 19825
rect 2320 19848 2372 19854
rect 1952 19790 2004 19796
rect 2042 19816 2098 19825
rect 1858 19751 1914 19760
rect 1872 19718 1900 19751
rect 1860 19712 1912 19718
rect 1860 19654 1912 19660
rect 1768 19508 1820 19514
rect 1768 19450 1820 19456
rect 1688 19366 1808 19394
rect 1584 17876 1636 17882
rect 1584 17818 1636 17824
rect 1490 17776 1546 17785
rect 1490 17711 1546 17720
rect 1584 17740 1636 17746
rect 1584 17682 1636 17688
rect 1492 17536 1544 17542
rect 1492 17478 1544 17484
rect 1400 17332 1452 17338
rect 1400 17274 1452 17280
rect 1400 16992 1452 16998
rect 1504 16969 1532 17478
rect 1400 16934 1452 16940
rect 1490 16960 1546 16969
rect 1308 16652 1360 16658
rect 1308 16594 1360 16600
rect 1216 3460 1268 3466
rect 1216 3402 1268 3408
rect 1124 3120 1176 3126
rect 1124 3062 1176 3068
rect 1320 2038 1348 16594
rect 1412 16590 1440 16934
rect 1490 16895 1546 16904
rect 1400 16584 1452 16590
rect 1596 16574 1624 17682
rect 1676 17672 1728 17678
rect 1676 17614 1728 17620
rect 1400 16526 1452 16532
rect 1504 16546 1624 16574
rect 1504 15994 1532 16546
rect 1584 16448 1636 16454
rect 1584 16390 1636 16396
rect 1596 16153 1624 16390
rect 1582 16144 1638 16153
rect 1582 16079 1638 16088
rect 1412 15966 1532 15994
rect 1412 8974 1440 15966
rect 1492 15904 1544 15910
rect 1492 15846 1544 15852
rect 1504 15745 1532 15846
rect 1490 15736 1546 15745
rect 1688 15706 1716 17614
rect 1490 15671 1546 15680
rect 1676 15700 1728 15706
rect 1676 15642 1728 15648
rect 1492 15360 1544 15366
rect 1490 15328 1492 15337
rect 1544 15328 1546 15337
rect 1490 15263 1546 15272
rect 1676 15020 1728 15026
rect 1676 14962 1728 14968
rect 1492 14816 1544 14822
rect 1492 14758 1544 14764
rect 1504 14521 1532 14758
rect 1688 14550 1716 14962
rect 1780 14618 1808 19366
rect 1858 18184 1914 18193
rect 1858 18119 1860 18128
rect 1912 18119 1914 18128
rect 1860 18090 1912 18096
rect 1860 17536 1912 17542
rect 1860 17478 1912 17484
rect 1872 17377 1900 17478
rect 1858 17368 1914 17377
rect 1858 17303 1914 17312
rect 1858 16552 1914 16561
rect 1858 16487 1914 16496
rect 1872 16454 1900 16487
rect 1860 16448 1912 16454
rect 1860 16390 1912 16396
rect 1964 16017 1992 19790
rect 2320 19790 2372 19796
rect 2412 19848 2464 19854
rect 2412 19790 2464 19796
rect 2042 19751 2098 19760
rect 2056 19378 2084 19751
rect 2044 19372 2096 19378
rect 2044 19314 2096 19320
rect 2136 19372 2188 19378
rect 2136 19314 2188 19320
rect 2044 18624 2096 18630
rect 2044 18566 2096 18572
rect 2056 18290 2084 18566
rect 2044 18284 2096 18290
rect 2044 18226 2096 18232
rect 2148 17082 2176 19314
rect 2228 19168 2280 19174
rect 2228 19110 2280 19116
rect 2240 18902 2268 19110
rect 2228 18896 2280 18902
rect 2228 18838 2280 18844
rect 2228 18760 2280 18766
rect 2228 18702 2280 18708
rect 2240 17882 2268 18702
rect 2228 17876 2280 17882
rect 2228 17818 2280 17824
rect 2228 17672 2280 17678
rect 2228 17614 2280 17620
rect 2240 17105 2268 17614
rect 2056 17054 2176 17082
rect 2226 17096 2282 17105
rect 2056 16697 2084 17054
rect 2226 17031 2282 17040
rect 2136 16992 2188 16998
rect 2188 16952 2268 16980
rect 2136 16934 2188 16940
rect 2042 16688 2098 16697
rect 2042 16623 2098 16632
rect 2044 16584 2096 16590
rect 2044 16526 2096 16532
rect 2056 16250 2084 16526
rect 2240 16522 2268 16952
rect 2228 16516 2280 16522
rect 2228 16458 2280 16464
rect 2044 16244 2096 16250
rect 2044 16186 2096 16192
rect 2136 16108 2188 16114
rect 2136 16050 2188 16056
rect 1950 16008 2006 16017
rect 1950 15943 2006 15952
rect 1858 14920 1914 14929
rect 1858 14855 1860 14864
rect 1912 14855 1914 14864
rect 1860 14826 1912 14832
rect 1768 14612 1820 14618
rect 1768 14554 1820 14560
rect 1676 14544 1728 14550
rect 1490 14512 1546 14521
rect 1676 14486 1728 14492
rect 1780 14482 1808 14554
rect 1490 14447 1546 14456
rect 1768 14476 1820 14482
rect 1768 14418 1820 14424
rect 1492 14272 1544 14278
rect 1492 14214 1544 14220
rect 1504 14113 1532 14214
rect 1490 14104 1546 14113
rect 2148 14090 2176 16050
rect 2240 16046 2268 16458
rect 2228 16040 2280 16046
rect 2228 15982 2280 15988
rect 2332 15609 2360 19790
rect 2516 19145 2544 21270
rect 2596 20460 2648 20466
rect 2596 20402 2648 20408
rect 2688 20460 2740 20466
rect 2688 20402 2740 20408
rect 2502 19136 2558 19145
rect 2502 19071 2558 19080
rect 2608 18873 2636 20402
rect 2594 18864 2650 18873
rect 2594 18799 2650 18808
rect 2596 18760 2648 18766
rect 2700 18737 2728 20402
rect 2596 18702 2648 18708
rect 2686 18728 2742 18737
rect 2504 18624 2556 18630
rect 2424 18584 2504 18612
rect 2424 18290 2452 18584
rect 2504 18566 2556 18572
rect 2412 18284 2464 18290
rect 2412 18226 2464 18232
rect 2504 18284 2556 18290
rect 2504 18226 2556 18232
rect 2412 18080 2464 18086
rect 2412 18022 2464 18028
rect 2424 16130 2452 18022
rect 2516 16574 2544 18226
rect 2608 17785 2636 18702
rect 2686 18663 2742 18672
rect 2688 18624 2740 18630
rect 2688 18566 2740 18572
rect 2594 17776 2650 17785
rect 2594 17711 2650 17720
rect 2700 16998 2728 18566
rect 2688 16992 2740 16998
rect 2688 16934 2740 16940
rect 2596 16788 2648 16794
rect 2700 16776 2728 16934
rect 2648 16748 2728 16776
rect 2596 16730 2648 16736
rect 2686 16688 2742 16697
rect 2686 16623 2742 16632
rect 2516 16546 2636 16574
rect 2608 16153 2636 16546
rect 2594 16144 2650 16153
rect 2424 16102 2544 16130
rect 2412 16040 2464 16046
rect 2412 15982 2464 15988
rect 2318 15600 2374 15609
rect 2318 15535 2374 15544
rect 2320 15496 2372 15502
rect 2320 15438 2372 15444
rect 2332 14618 2360 15438
rect 2424 15162 2452 15982
rect 2412 15156 2464 15162
rect 2412 15098 2464 15104
rect 2516 15026 2544 16102
rect 2594 16079 2650 16088
rect 2504 15020 2556 15026
rect 2504 14962 2556 14968
rect 2412 14952 2464 14958
rect 2412 14894 2464 14900
rect 2320 14612 2372 14618
rect 2320 14554 2372 14560
rect 2320 14408 2372 14414
rect 2320 14350 2372 14356
rect 2148 14062 2268 14090
rect 2332 14074 2360 14350
rect 1490 14039 1546 14048
rect 2136 13932 2188 13938
rect 2136 13874 2188 13880
rect 1584 13864 1636 13870
rect 1584 13806 1636 13812
rect 1492 13728 1544 13734
rect 1490 13696 1492 13705
rect 1544 13696 1546 13705
rect 1490 13631 1546 13640
rect 1490 13288 1546 13297
rect 1490 13223 1546 13232
rect 1504 13190 1532 13223
rect 1492 13184 1544 13190
rect 1492 13126 1544 13132
rect 1492 12980 1544 12986
rect 1492 12922 1544 12928
rect 1504 12889 1532 12922
rect 1490 12880 1546 12889
rect 1490 12815 1546 12824
rect 1490 12744 1546 12753
rect 1490 12679 1492 12688
rect 1544 12679 1546 12688
rect 1492 12650 1544 12656
rect 1596 12442 1624 13806
rect 1860 13728 1912 13734
rect 1860 13670 1912 13676
rect 1766 13288 1822 13297
rect 1766 13223 1768 13232
rect 1820 13223 1822 13232
rect 1768 13194 1820 13200
rect 1676 12844 1728 12850
rect 1676 12786 1728 12792
rect 1688 12442 1716 12786
rect 1768 12776 1820 12782
rect 1768 12718 1820 12724
rect 1584 12436 1636 12442
rect 1584 12378 1636 12384
rect 1676 12436 1728 12442
rect 1676 12378 1728 12384
rect 1780 12238 1808 12718
rect 1872 12481 1900 13670
rect 1952 12844 2004 12850
rect 1952 12786 2004 12792
rect 1858 12472 1914 12481
rect 1858 12407 1914 12416
rect 1964 12238 1992 12786
rect 1768 12232 1820 12238
rect 1768 12174 1820 12180
rect 1952 12232 2004 12238
rect 1952 12174 2004 12180
rect 2042 12200 2098 12209
rect 2042 12135 2098 12144
rect 1490 12064 1546 12073
rect 1490 11999 1546 12008
rect 1504 11354 1532 11999
rect 1860 11892 1912 11898
rect 1860 11834 1912 11840
rect 1492 11348 1544 11354
rect 1492 11290 1544 11296
rect 1872 11257 1900 11834
rect 1950 11792 2006 11801
rect 1950 11727 1952 11736
rect 2004 11727 2006 11736
rect 1952 11698 2004 11704
rect 2056 11286 2084 12135
rect 2044 11280 2096 11286
rect 1858 11248 1914 11257
rect 2044 11222 2096 11228
rect 1858 11183 1914 11192
rect 1872 11150 1900 11183
rect 1676 11144 1728 11150
rect 1676 11086 1728 11092
rect 1860 11144 1912 11150
rect 1860 11086 1912 11092
rect 1490 10840 1546 10849
rect 1490 10775 1546 10784
rect 1504 10674 1532 10775
rect 1492 10668 1544 10674
rect 1492 10610 1544 10616
rect 1490 10432 1546 10441
rect 1490 10367 1546 10376
rect 1504 10062 1532 10367
rect 1492 10056 1544 10062
rect 1492 9998 1544 10004
rect 1492 9648 1544 9654
rect 1490 9616 1492 9625
rect 1544 9616 1546 9625
rect 1490 9551 1546 9560
rect 1492 9376 1544 9382
rect 1492 9318 1544 9324
rect 1400 8968 1452 8974
rect 1400 8910 1452 8916
rect 1398 8800 1454 8809
rect 1398 8735 1454 8744
rect 1412 7410 1440 8735
rect 1400 7404 1452 7410
rect 1400 7346 1452 7352
rect 1504 7256 1532 9318
rect 1584 9036 1636 9042
rect 1584 8978 1636 8984
rect 1596 8430 1624 8978
rect 1584 8424 1636 8430
rect 1584 8366 1636 8372
rect 1582 8256 1638 8265
rect 1582 8191 1638 8200
rect 1596 7546 1624 8191
rect 1584 7540 1636 7546
rect 1584 7482 1636 7488
rect 1412 7228 1532 7256
rect 1412 4486 1440 7228
rect 1490 7168 1546 7177
rect 1490 7103 1546 7112
rect 1504 6866 1532 7103
rect 1492 6860 1544 6866
rect 1492 6802 1544 6808
rect 1504 6390 1532 6802
rect 1492 6384 1544 6390
rect 1492 6326 1544 6332
rect 1400 4480 1452 4486
rect 1400 4422 1452 4428
rect 1398 4312 1454 4321
rect 1398 4247 1454 4256
rect 1412 3534 1440 4247
rect 1492 4140 1544 4146
rect 1492 4082 1544 4088
rect 1400 3528 1452 3534
rect 1400 3470 1452 3476
rect 1308 2032 1360 2038
rect 1308 1974 1360 1980
rect 1504 1698 1532 4082
rect 1688 4010 1716 11086
rect 1860 10668 1912 10674
rect 1860 10610 1912 10616
rect 2044 10668 2096 10674
rect 2044 10610 2096 10616
rect 1768 10600 1820 10606
rect 1872 10577 1900 10610
rect 1768 10542 1820 10548
rect 1858 10568 1914 10577
rect 1780 10130 1808 10542
rect 1858 10503 1914 10512
rect 1860 10192 1912 10198
rect 1858 10160 1860 10169
rect 1912 10160 1914 10169
rect 1768 10124 1820 10130
rect 1858 10095 1914 10104
rect 1768 10066 1820 10072
rect 1860 9920 1912 9926
rect 1860 9862 1912 9868
rect 1952 9920 2004 9926
rect 2056 9908 2084 10610
rect 2148 10266 2176 13874
rect 2240 11914 2268 14062
rect 2320 14068 2372 14074
rect 2320 14010 2372 14016
rect 2424 14006 2452 14894
rect 2412 14000 2464 14006
rect 2412 13942 2464 13948
rect 2516 13954 2544 14962
rect 2700 14822 2728 16623
rect 2688 14816 2740 14822
rect 2688 14758 2740 14764
rect 2792 14414 2820 22200
rect 2872 20528 2924 20534
rect 2870 20496 2872 20505
rect 2924 20496 2926 20505
rect 2870 20431 2926 20440
rect 2964 20460 3016 20466
rect 2964 20402 3016 20408
rect 2870 19136 2926 19145
rect 2870 19071 2926 19080
rect 2596 14408 2648 14414
rect 2780 14408 2832 14414
rect 2648 14368 2728 14396
rect 2596 14350 2648 14356
rect 2516 13926 2636 13954
rect 2412 13864 2464 13870
rect 2410 13832 2412 13841
rect 2464 13832 2466 13841
rect 2410 13767 2466 13776
rect 2504 13796 2556 13802
rect 2504 13738 2556 13744
rect 2412 13728 2464 13734
rect 2412 13670 2464 13676
rect 2240 11886 2360 11914
rect 2228 11756 2280 11762
rect 2228 11698 2280 11704
rect 2240 11665 2268 11698
rect 2226 11656 2282 11665
rect 2226 11591 2282 11600
rect 2332 11354 2360 11886
rect 2320 11348 2372 11354
rect 2320 11290 2372 11296
rect 2136 10260 2188 10266
rect 2136 10202 2188 10208
rect 2228 9988 2280 9994
rect 2228 9930 2280 9936
rect 2004 9880 2084 9908
rect 1952 9862 2004 9868
rect 1872 9722 1900 9862
rect 1860 9716 1912 9722
rect 1860 9658 1912 9664
rect 1964 9518 1992 9862
rect 2042 9752 2098 9761
rect 2042 9687 2098 9696
rect 1952 9512 2004 9518
rect 1952 9454 2004 9460
rect 1860 9444 1912 9450
rect 1860 9386 1912 9392
rect 1872 8945 1900 9386
rect 1858 8936 1914 8945
rect 1858 8871 1914 8880
rect 1768 8832 1820 8838
rect 1768 8774 1820 8780
rect 1780 8090 1808 8774
rect 1952 8492 2004 8498
rect 1952 8434 2004 8440
rect 1860 8424 1912 8430
rect 1860 8366 1912 8372
rect 1872 8090 1900 8366
rect 1768 8084 1820 8090
rect 1768 8026 1820 8032
rect 1860 8084 1912 8090
rect 1860 8026 1912 8032
rect 1766 7712 1822 7721
rect 1766 7647 1822 7656
rect 1780 6390 1808 7647
rect 1964 6458 1992 8434
rect 2056 7886 2084 9687
rect 2136 9512 2188 9518
rect 2136 9454 2188 9460
rect 2148 9178 2176 9454
rect 2240 9382 2268 9930
rect 2320 9580 2372 9586
rect 2320 9522 2372 9528
rect 2228 9376 2280 9382
rect 2228 9318 2280 9324
rect 2240 9178 2268 9318
rect 2136 9172 2188 9178
rect 2136 9114 2188 9120
rect 2228 9172 2280 9178
rect 2228 9114 2280 9120
rect 2134 8664 2190 8673
rect 2332 8634 2360 9522
rect 2424 9058 2452 13670
rect 2516 13530 2544 13738
rect 2504 13524 2556 13530
rect 2504 13466 2556 13472
rect 2516 12918 2544 13466
rect 2608 13326 2636 13926
rect 2596 13320 2648 13326
rect 2596 13262 2648 13268
rect 2504 12912 2556 12918
rect 2504 12854 2556 12860
rect 2608 12850 2636 13262
rect 2596 12844 2648 12850
rect 2596 12786 2648 12792
rect 2504 12640 2556 12646
rect 2504 12582 2556 12588
rect 2516 11898 2544 12582
rect 2700 11937 2728 14368
rect 2884 14396 2912 19071
rect 2976 18737 3004 20402
rect 3160 20040 3188 22200
rect 3332 20460 3384 20466
rect 3332 20402 3384 20408
rect 3160 20012 3280 20040
rect 3146 19952 3202 19961
rect 3146 19887 3202 19896
rect 3160 19854 3188 19887
rect 3148 19848 3200 19854
rect 3148 19790 3200 19796
rect 3056 19780 3108 19786
rect 3056 19722 3108 19728
rect 3068 19446 3096 19722
rect 3148 19712 3200 19718
rect 3148 19654 3200 19660
rect 3056 19440 3108 19446
rect 3056 19382 3108 19388
rect 3056 19168 3108 19174
rect 3056 19110 3108 19116
rect 2962 18728 3018 18737
rect 2962 18663 3018 18672
rect 3068 18426 3096 19110
rect 3160 18970 3188 19654
rect 3148 18964 3200 18970
rect 3148 18906 3200 18912
rect 3148 18624 3200 18630
rect 3148 18566 3200 18572
rect 3160 18426 3188 18566
rect 3056 18420 3108 18426
rect 3056 18362 3108 18368
rect 3148 18420 3200 18426
rect 3148 18362 3200 18368
rect 3056 18284 3108 18290
rect 3056 18226 3108 18232
rect 2964 18216 3016 18222
rect 2964 18158 3016 18164
rect 2976 17202 3004 18158
rect 2964 17196 3016 17202
rect 2964 17138 3016 17144
rect 2976 15570 3004 17138
rect 2964 15564 3016 15570
rect 2964 15506 3016 15512
rect 2964 15360 3016 15366
rect 2964 15302 3016 15308
rect 2976 15094 3004 15302
rect 2964 15088 3016 15094
rect 2964 15030 3016 15036
rect 3068 14618 3096 18226
rect 3252 17746 3280 20012
rect 3344 19281 3372 20402
rect 3528 20369 3556 22200
rect 3896 21026 3924 22200
rect 4066 21856 4122 21865
rect 4066 21791 4122 21800
rect 3896 20998 4016 21026
rect 3884 20936 3936 20942
rect 3884 20878 3936 20884
rect 3896 20602 3924 20878
rect 3884 20596 3936 20602
rect 3884 20538 3936 20544
rect 3988 20482 4016 20998
rect 4080 20806 4108 21791
rect 4068 20800 4120 20806
rect 4068 20742 4120 20748
rect 4160 20528 4212 20534
rect 3988 20454 4108 20482
rect 4160 20470 4212 20476
rect 3976 20392 4028 20398
rect 3514 20360 3570 20369
rect 3424 20324 3476 20330
rect 3976 20334 4028 20340
rect 3514 20295 3570 20304
rect 3424 20266 3476 20272
rect 3436 19417 3464 20266
rect 3884 20256 3936 20262
rect 3884 20198 3936 20204
rect 3549 20156 3857 20165
rect 3549 20154 3555 20156
rect 3611 20154 3635 20156
rect 3691 20154 3715 20156
rect 3771 20154 3795 20156
rect 3851 20154 3857 20156
rect 3611 20102 3613 20154
rect 3793 20102 3795 20154
rect 3549 20100 3555 20102
rect 3611 20100 3635 20102
rect 3691 20100 3715 20102
rect 3771 20100 3795 20102
rect 3851 20100 3857 20102
rect 3549 20091 3857 20100
rect 3896 19854 3924 20198
rect 3884 19848 3936 19854
rect 3884 19790 3936 19796
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 3608 19372 3660 19378
rect 3608 19314 3660 19320
rect 3330 19272 3386 19281
rect 3330 19207 3386 19216
rect 3424 19236 3476 19242
rect 3424 19178 3476 19184
rect 3332 19168 3384 19174
rect 3332 19110 3384 19116
rect 3344 18834 3372 19110
rect 3436 18834 3464 19178
rect 3620 19174 3648 19314
rect 3608 19168 3660 19174
rect 3608 19110 3660 19116
rect 3884 19168 3936 19174
rect 3884 19110 3936 19116
rect 3549 19068 3857 19077
rect 3549 19066 3555 19068
rect 3611 19066 3635 19068
rect 3691 19066 3715 19068
rect 3771 19066 3795 19068
rect 3851 19066 3857 19068
rect 3611 19014 3613 19066
rect 3793 19014 3795 19066
rect 3549 19012 3555 19014
rect 3611 19012 3635 19014
rect 3691 19012 3715 19014
rect 3771 19012 3795 19014
rect 3851 19012 3857 19014
rect 3549 19003 3857 19012
rect 3896 18834 3924 19110
rect 3332 18828 3384 18834
rect 3332 18770 3384 18776
rect 3424 18828 3476 18834
rect 3424 18770 3476 18776
rect 3884 18828 3936 18834
rect 3884 18770 3936 18776
rect 3332 18624 3384 18630
rect 3332 18566 3384 18572
rect 3344 18358 3372 18566
rect 3332 18352 3384 18358
rect 3332 18294 3384 18300
rect 3332 17808 3384 17814
rect 3332 17750 3384 17756
rect 3240 17740 3292 17746
rect 3240 17682 3292 17688
rect 3344 17610 3372 17750
rect 3332 17604 3384 17610
rect 3332 17546 3384 17552
rect 3148 17536 3200 17542
rect 3148 17478 3200 17484
rect 3240 17536 3292 17542
rect 3240 17478 3292 17484
rect 3160 16794 3188 17478
rect 3148 16788 3200 16794
rect 3148 16730 3200 16736
rect 3252 16130 3280 17478
rect 3436 17354 3464 18770
rect 3988 18766 4016 20334
rect 4080 19802 4108 20454
rect 4172 20097 4200 20470
rect 4158 20088 4214 20097
rect 4158 20023 4214 20032
rect 4264 19922 4292 22200
rect 4252 19916 4304 19922
rect 4252 19858 4304 19864
rect 4080 19774 4200 19802
rect 4068 19712 4120 19718
rect 4068 19654 4120 19660
rect 4080 18766 4108 19654
rect 3976 18760 4028 18766
rect 3976 18702 4028 18708
rect 4068 18760 4120 18766
rect 4068 18702 4120 18708
rect 3988 18306 4016 18702
rect 4066 18456 4122 18465
rect 4066 18391 4068 18400
rect 4120 18391 4122 18400
rect 4068 18362 4120 18368
rect 3988 18278 4108 18306
rect 3976 18148 4028 18154
rect 3976 18090 4028 18096
rect 3549 17980 3857 17989
rect 3549 17978 3555 17980
rect 3611 17978 3635 17980
rect 3691 17978 3715 17980
rect 3771 17978 3795 17980
rect 3851 17978 3857 17980
rect 3611 17926 3613 17978
rect 3793 17926 3795 17978
rect 3549 17924 3555 17926
rect 3611 17924 3635 17926
rect 3691 17924 3715 17926
rect 3771 17924 3795 17926
rect 3851 17924 3857 17926
rect 3549 17915 3857 17924
rect 3700 17740 3752 17746
rect 3700 17682 3752 17688
rect 3712 17610 3740 17682
rect 3884 17672 3936 17678
rect 3884 17614 3936 17620
rect 3608 17604 3660 17610
rect 3608 17546 3660 17552
rect 3700 17604 3752 17610
rect 3700 17546 3752 17552
rect 3160 16102 3280 16130
rect 3344 17326 3464 17354
rect 3160 15978 3188 16102
rect 3240 16040 3292 16046
rect 3240 15982 3292 15988
rect 3148 15972 3200 15978
rect 3148 15914 3200 15920
rect 3148 15360 3200 15366
rect 3148 15302 3200 15308
rect 3056 14612 3108 14618
rect 3056 14554 3108 14560
rect 2964 14408 3016 14414
rect 2884 14368 2964 14396
rect 2780 14350 2832 14356
rect 2964 14350 3016 14356
rect 2686 11928 2742 11937
rect 2504 11892 2556 11898
rect 2686 11863 2742 11872
rect 2504 11834 2556 11840
rect 2792 11762 2820 14350
rect 2872 14272 2924 14278
rect 2872 14214 2924 14220
rect 2884 12374 2912 14214
rect 3160 14074 3188 15302
rect 3252 15065 3280 15982
rect 3238 15056 3294 15065
rect 3344 15026 3372 17326
rect 3620 17270 3648 17546
rect 3792 17536 3844 17542
rect 3792 17478 3844 17484
rect 3424 17264 3476 17270
rect 3424 17206 3476 17212
rect 3608 17264 3660 17270
rect 3804 17241 3832 17478
rect 3608 17206 3660 17212
rect 3790 17232 3846 17241
rect 3436 16726 3464 17206
rect 3790 17167 3846 17176
rect 3549 16892 3857 16901
rect 3549 16890 3555 16892
rect 3611 16890 3635 16892
rect 3691 16890 3715 16892
rect 3771 16890 3795 16892
rect 3851 16890 3857 16892
rect 3611 16838 3613 16890
rect 3793 16838 3795 16890
rect 3549 16836 3555 16838
rect 3611 16836 3635 16838
rect 3691 16836 3715 16838
rect 3771 16836 3795 16838
rect 3851 16836 3857 16838
rect 3549 16827 3857 16836
rect 3896 16726 3924 17614
rect 3424 16720 3476 16726
rect 3424 16662 3476 16668
rect 3884 16720 3936 16726
rect 3884 16662 3936 16668
rect 3988 16590 4016 18090
rect 4080 18086 4108 18278
rect 4068 18080 4120 18086
rect 4068 18022 4120 18028
rect 4068 17536 4120 17542
rect 4068 17478 4120 17484
rect 4080 17270 4108 17478
rect 4068 17264 4120 17270
rect 4068 17206 4120 17212
rect 4066 16960 4122 16969
rect 4066 16895 4122 16904
rect 3976 16584 4028 16590
rect 3976 16526 4028 16532
rect 4080 16436 4108 16895
rect 4172 16538 4200 19774
rect 4252 19780 4304 19786
rect 4252 19722 4304 19728
rect 4264 18630 4292 19722
rect 4252 18624 4304 18630
rect 4252 18566 4304 18572
rect 4264 17134 4292 18566
rect 4356 17678 4384 22222
rect 4540 22114 4568 22222
rect 4618 22200 4674 23000
rect 4986 22200 5042 23000
rect 5354 22200 5410 23000
rect 5722 22200 5778 23000
rect 6090 22200 6146 23000
rect 6458 22200 6514 23000
rect 6826 22200 6882 23000
rect 7194 22200 7250 23000
rect 7562 22200 7618 23000
rect 7930 22200 7986 23000
rect 8298 22200 8354 23000
rect 8666 22200 8722 23000
rect 9034 22200 9090 23000
rect 9402 22200 9458 23000
rect 9770 22200 9826 23000
rect 10138 22200 10194 23000
rect 10506 22200 10562 23000
rect 10874 22200 10930 23000
rect 11242 22200 11298 23000
rect 11610 22200 11666 23000
rect 11978 22200 12034 23000
rect 12346 22200 12402 23000
rect 12714 22200 12770 23000
rect 13082 22200 13138 23000
rect 13450 22200 13506 23000
rect 13818 22200 13874 23000
rect 14186 22200 14242 23000
rect 14554 22200 14610 23000
rect 14922 22200 14978 23000
rect 15290 22200 15346 23000
rect 15658 22200 15714 23000
rect 16026 22200 16082 23000
rect 16394 22200 16450 23000
rect 16762 22200 16818 23000
rect 17130 22200 17186 23000
rect 17498 22200 17554 23000
rect 17866 22200 17922 23000
rect 18234 22200 18290 23000
rect 18602 22200 18658 23000
rect 18970 22200 19026 23000
rect 19338 22200 19394 23000
rect 19706 22200 19762 23000
rect 20074 22200 20130 23000
rect 20442 22200 20498 23000
rect 20810 22200 20866 23000
rect 21178 22200 21234 23000
rect 21546 22200 21602 23000
rect 21652 22222 21864 22250
rect 4632 22114 4660 22200
rect 4540 22086 4660 22114
rect 4712 20460 4764 20466
rect 4712 20402 4764 20408
rect 4618 20360 4674 20369
rect 4618 20295 4674 20304
rect 4632 19854 4660 20295
rect 4620 19848 4672 19854
rect 4620 19790 4672 19796
rect 4436 19780 4488 19786
rect 4436 19722 4488 19728
rect 4448 18834 4476 19722
rect 4528 19712 4580 19718
rect 4528 19654 4580 19660
rect 4540 19553 4568 19654
rect 4526 19544 4582 19553
rect 4526 19479 4582 19488
rect 4528 19304 4580 19310
rect 4528 19246 4580 19252
rect 4436 18828 4488 18834
rect 4436 18770 4488 18776
rect 4434 18320 4490 18329
rect 4434 18255 4490 18264
rect 4344 17672 4396 17678
rect 4344 17614 4396 17620
rect 4252 17128 4304 17134
rect 4252 17070 4304 17076
rect 4356 16697 4384 17614
rect 4448 17542 4476 18255
rect 4436 17536 4488 17542
rect 4436 17478 4488 17484
rect 4342 16688 4398 16697
rect 4342 16623 4398 16632
rect 4172 16522 4384 16538
rect 4172 16516 4396 16522
rect 4172 16510 4344 16516
rect 4344 16458 4396 16464
rect 3988 16408 4108 16436
rect 4160 16448 4212 16454
rect 3884 16040 3936 16046
rect 3422 16008 3478 16017
rect 3884 15982 3936 15988
rect 3422 15943 3478 15952
rect 3436 15638 3464 15943
rect 3549 15804 3857 15813
rect 3549 15802 3555 15804
rect 3611 15802 3635 15804
rect 3691 15802 3715 15804
rect 3771 15802 3795 15804
rect 3851 15802 3857 15804
rect 3611 15750 3613 15802
rect 3793 15750 3795 15802
rect 3549 15748 3555 15750
rect 3611 15748 3635 15750
rect 3691 15748 3715 15750
rect 3771 15748 3795 15750
rect 3851 15748 3857 15750
rect 3549 15739 3857 15748
rect 3424 15632 3476 15638
rect 3424 15574 3476 15580
rect 3896 15570 3924 15982
rect 3884 15564 3936 15570
rect 3884 15506 3936 15512
rect 3792 15496 3844 15502
rect 3790 15464 3792 15473
rect 3844 15464 3846 15473
rect 3790 15399 3846 15408
rect 3238 14991 3294 15000
rect 3332 15020 3384 15026
rect 3252 14498 3280 14991
rect 3332 14962 3384 14968
rect 3896 14890 3924 15506
rect 3884 14884 3936 14890
rect 3884 14826 3936 14832
rect 3424 14816 3476 14822
rect 3424 14758 3476 14764
rect 3252 14470 3372 14498
rect 3240 14408 3292 14414
rect 3240 14350 3292 14356
rect 3148 14068 3200 14074
rect 3148 14010 3200 14016
rect 2964 13932 3016 13938
rect 2964 13874 3016 13880
rect 2872 12368 2924 12374
rect 2872 12310 2924 12316
rect 2976 11898 3004 13874
rect 3056 13864 3108 13870
rect 3056 13806 3108 13812
rect 3068 12986 3096 13806
rect 3056 12980 3108 12986
rect 3056 12922 3108 12928
rect 3252 12442 3280 14350
rect 3344 13705 3372 14470
rect 3436 14278 3464 14758
rect 3549 14716 3857 14725
rect 3549 14714 3555 14716
rect 3611 14714 3635 14716
rect 3691 14714 3715 14716
rect 3771 14714 3795 14716
rect 3851 14714 3857 14716
rect 3611 14662 3613 14714
rect 3793 14662 3795 14714
rect 3549 14660 3555 14662
rect 3611 14660 3635 14662
rect 3691 14660 3715 14662
rect 3771 14660 3795 14662
rect 3851 14660 3857 14662
rect 3549 14651 3857 14660
rect 3988 14550 4016 16408
rect 4160 16390 4212 16396
rect 4172 15706 4200 16390
rect 4342 16280 4398 16289
rect 4342 16215 4398 16224
rect 4252 15904 4304 15910
rect 4252 15846 4304 15852
rect 4160 15700 4212 15706
rect 4160 15642 4212 15648
rect 4066 15600 4122 15609
rect 4264 15586 4292 15846
rect 4356 15706 4384 16215
rect 4448 16114 4476 17478
rect 4540 16697 4568 19246
rect 4632 17649 4660 19790
rect 4724 18834 4752 20402
rect 4896 19916 4948 19922
rect 4896 19858 4948 19864
rect 4804 19848 4856 19854
rect 4804 19790 4856 19796
rect 4816 19378 4844 19790
rect 4804 19372 4856 19378
rect 4804 19314 4856 19320
rect 4712 18828 4764 18834
rect 4712 18770 4764 18776
rect 4724 18465 4752 18770
rect 4710 18456 4766 18465
rect 4710 18391 4766 18400
rect 4712 18284 4764 18290
rect 4712 18226 4764 18232
rect 4618 17640 4674 17649
rect 4618 17575 4674 17584
rect 4724 17542 4752 18226
rect 4816 17678 4844 19314
rect 4908 19145 4936 19858
rect 5000 19802 5028 22200
rect 5368 20505 5396 22200
rect 5354 20496 5410 20505
rect 5354 20431 5410 20440
rect 5356 20256 5408 20262
rect 5540 20256 5592 20262
rect 5356 20198 5408 20204
rect 5460 20204 5540 20210
rect 5460 20198 5592 20204
rect 5000 19774 5212 19802
rect 5080 19712 5132 19718
rect 5080 19654 5132 19660
rect 5092 19174 5120 19654
rect 4988 19168 5040 19174
rect 4894 19136 4950 19145
rect 4988 19110 5040 19116
rect 5080 19168 5132 19174
rect 5080 19110 5132 19116
rect 4894 19071 4950 19080
rect 5000 18714 5028 19110
rect 5000 18686 5120 18714
rect 4896 18624 4948 18630
rect 4896 18566 4948 18572
rect 4988 18624 5040 18630
rect 4988 18566 5040 18572
rect 4804 17672 4856 17678
rect 4804 17614 4856 17620
rect 4712 17536 4764 17542
rect 4712 17478 4764 17484
rect 4804 17196 4856 17202
rect 4804 17138 4856 17144
rect 4620 16992 4672 16998
rect 4620 16934 4672 16940
rect 4526 16688 4582 16697
rect 4526 16623 4582 16632
rect 4632 16182 4660 16934
rect 4816 16833 4844 17138
rect 4802 16824 4858 16833
rect 4802 16759 4858 16768
rect 4712 16584 4764 16590
rect 4764 16544 4844 16572
rect 4712 16526 4764 16532
rect 4620 16176 4672 16182
rect 4620 16118 4672 16124
rect 4436 16108 4488 16114
rect 4436 16050 4488 16056
rect 4344 15700 4396 15706
rect 4344 15642 4396 15648
rect 4356 15609 4384 15642
rect 4066 15535 4122 15544
rect 4172 15558 4292 15586
rect 4342 15600 4398 15609
rect 4080 15366 4108 15535
rect 4068 15360 4120 15366
rect 4068 15302 4120 15308
rect 3976 14544 4028 14550
rect 3976 14486 4028 14492
rect 4172 14414 4200 15558
rect 4342 15535 4398 15544
rect 4620 15564 4672 15570
rect 4620 15506 4672 15512
rect 4252 15496 4304 15502
rect 4250 15464 4252 15473
rect 4304 15464 4306 15473
rect 4250 15399 4306 15408
rect 4264 14657 4292 15399
rect 4344 15020 4396 15026
rect 4344 14962 4396 14968
rect 4250 14648 4306 14657
rect 4250 14583 4306 14592
rect 4160 14408 4212 14414
rect 4160 14350 4212 14356
rect 4068 14340 4120 14346
rect 4068 14282 4120 14288
rect 3424 14272 3476 14278
rect 3424 14214 3476 14220
rect 3884 14000 3936 14006
rect 3884 13942 3936 13948
rect 3424 13728 3476 13734
rect 3330 13696 3386 13705
rect 3424 13670 3476 13676
rect 3330 13631 3386 13640
rect 3332 13388 3384 13394
rect 3332 13330 3384 13336
rect 3240 12436 3292 12442
rect 3240 12378 3292 12384
rect 3344 12322 3372 13330
rect 3252 12294 3372 12322
rect 3056 12096 3108 12102
rect 3056 12038 3108 12044
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 2688 11756 2740 11762
rect 2688 11698 2740 11704
rect 2780 11756 2832 11762
rect 2780 11698 2832 11704
rect 2504 11688 2556 11694
rect 2504 11630 2556 11636
rect 2596 11688 2648 11694
rect 2596 11630 2648 11636
rect 2516 11218 2544 11630
rect 2504 11212 2556 11218
rect 2504 11154 2556 11160
rect 2502 10704 2558 10713
rect 2502 10639 2558 10648
rect 2516 10033 2544 10639
rect 2502 10024 2558 10033
rect 2502 9959 2558 9968
rect 2516 9586 2544 9959
rect 2504 9580 2556 9586
rect 2504 9522 2556 9528
rect 2608 9178 2636 11630
rect 2700 9450 2728 11698
rect 2964 11144 3016 11150
rect 2964 11086 3016 11092
rect 2872 11076 2924 11082
rect 2872 11018 2924 11024
rect 2780 9988 2832 9994
rect 2780 9930 2832 9936
rect 2688 9444 2740 9450
rect 2688 9386 2740 9392
rect 2596 9172 2648 9178
rect 2596 9114 2648 9120
rect 2424 9030 2544 9058
rect 2412 8900 2464 8906
rect 2412 8842 2464 8848
rect 2424 8634 2452 8842
rect 2134 8599 2136 8608
rect 2188 8599 2190 8608
rect 2320 8628 2372 8634
rect 2136 8570 2188 8576
rect 2320 8570 2372 8576
rect 2412 8628 2464 8634
rect 2412 8570 2464 8576
rect 2320 8356 2372 8362
rect 2320 8298 2372 8304
rect 2044 7880 2096 7886
rect 2044 7822 2096 7828
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 2042 7440 2098 7449
rect 2042 7375 2098 7384
rect 1952 6452 2004 6458
rect 1952 6394 2004 6400
rect 1768 6384 1820 6390
rect 1768 6326 1820 6332
rect 2056 5234 2084 7375
rect 2136 6792 2188 6798
rect 2134 6760 2136 6769
rect 2188 6760 2190 6769
rect 2134 6695 2190 6704
rect 2136 6656 2188 6662
rect 2136 6598 2188 6604
rect 2148 6338 2176 6598
rect 2240 6458 2268 7822
rect 2228 6452 2280 6458
rect 2228 6394 2280 6400
rect 2148 6310 2268 6338
rect 2136 5568 2188 5574
rect 2136 5510 2188 5516
rect 2044 5228 2096 5234
rect 2044 5170 2096 5176
rect 1768 5160 1820 5166
rect 1766 5128 1768 5137
rect 1820 5128 1822 5137
rect 1766 5063 1822 5072
rect 1950 5128 2006 5137
rect 1950 5063 2006 5072
rect 1964 4690 1992 5063
rect 2148 4826 2176 5510
rect 2136 4820 2188 4826
rect 2136 4762 2188 4768
rect 1952 4684 2004 4690
rect 1952 4626 2004 4632
rect 1768 4548 1820 4554
rect 1768 4490 1820 4496
rect 1780 4321 1808 4490
rect 2044 4480 2096 4486
rect 2044 4422 2096 4428
rect 1766 4312 1822 4321
rect 2056 4282 2084 4422
rect 1766 4247 1822 4256
rect 2044 4276 2096 4282
rect 2044 4218 2096 4224
rect 2148 4078 2176 4762
rect 2240 4554 2268 6310
rect 2228 4548 2280 4554
rect 2228 4490 2280 4496
rect 2136 4072 2188 4078
rect 2136 4014 2188 4020
rect 1676 4004 1728 4010
rect 1676 3946 1728 3952
rect 1952 3664 2004 3670
rect 1950 3632 1952 3641
rect 2004 3632 2006 3641
rect 1950 3567 2006 3576
rect 1584 3392 1636 3398
rect 1584 3334 1636 3340
rect 1492 1692 1544 1698
rect 1492 1634 1544 1640
rect 1596 1329 1624 3334
rect 2332 2938 2360 8298
rect 2516 7750 2544 9030
rect 2792 8537 2820 9930
rect 2778 8528 2834 8537
rect 2778 8463 2834 8472
rect 2688 7948 2740 7954
rect 2688 7890 2740 7896
rect 2596 7812 2648 7818
rect 2596 7754 2648 7760
rect 2504 7744 2556 7750
rect 2504 7686 2556 7692
rect 2412 7540 2464 7546
rect 2412 7482 2464 7488
rect 2424 4622 2452 7482
rect 2516 7313 2544 7686
rect 2608 7546 2636 7754
rect 2596 7540 2648 7546
rect 2596 7482 2648 7488
rect 2502 7304 2558 7313
rect 2502 7239 2558 7248
rect 2504 6860 2556 6866
rect 2504 6802 2556 6808
rect 2516 5681 2544 6802
rect 2594 6760 2650 6769
rect 2594 6695 2596 6704
rect 2648 6695 2650 6704
rect 2596 6666 2648 6672
rect 2700 6254 2728 7890
rect 2792 7478 2820 8463
rect 2884 7970 2912 11018
rect 2976 10810 3004 11086
rect 2964 10804 3016 10810
rect 2964 10746 3016 10752
rect 3068 9994 3096 12038
rect 3148 11552 3200 11558
rect 3148 11494 3200 11500
rect 3160 11286 3188 11494
rect 3148 11280 3200 11286
rect 3148 11222 3200 11228
rect 3252 10146 3280 12294
rect 3332 12232 3384 12238
rect 3332 12174 3384 12180
rect 3344 11286 3372 12174
rect 3436 11898 3464 13670
rect 3549 13628 3857 13637
rect 3549 13626 3555 13628
rect 3611 13626 3635 13628
rect 3691 13626 3715 13628
rect 3771 13626 3795 13628
rect 3851 13626 3857 13628
rect 3611 13574 3613 13626
rect 3793 13574 3795 13626
rect 3549 13572 3555 13574
rect 3611 13572 3635 13574
rect 3691 13572 3715 13574
rect 3771 13572 3795 13574
rect 3851 13572 3857 13574
rect 3549 13563 3857 13572
rect 3896 13394 3924 13942
rect 3884 13388 3936 13394
rect 3884 13330 3936 13336
rect 3976 13252 4028 13258
rect 3976 13194 4028 13200
rect 3988 12714 4016 13194
rect 4080 13025 4108 14282
rect 4172 13530 4200 14350
rect 4252 13864 4304 13870
rect 4356 13841 4384 14962
rect 4632 14822 4660 15506
rect 4712 15428 4764 15434
rect 4712 15370 4764 15376
rect 4620 14816 4672 14822
rect 4620 14758 4672 14764
rect 4528 14068 4580 14074
rect 4528 14010 4580 14016
rect 4252 13806 4304 13812
rect 4342 13832 4398 13841
rect 4160 13524 4212 13530
rect 4160 13466 4212 13472
rect 4066 13016 4122 13025
rect 4066 12951 4122 12960
rect 4068 12912 4120 12918
rect 4068 12854 4120 12860
rect 3976 12708 4028 12714
rect 3976 12650 4028 12656
rect 3549 12540 3857 12549
rect 3549 12538 3555 12540
rect 3611 12538 3635 12540
rect 3691 12538 3715 12540
rect 3771 12538 3795 12540
rect 3851 12538 3857 12540
rect 3611 12486 3613 12538
rect 3793 12486 3795 12538
rect 3549 12484 3555 12486
rect 3611 12484 3635 12486
rect 3691 12484 3715 12486
rect 3771 12484 3795 12486
rect 3851 12484 3857 12486
rect 3549 12475 3857 12484
rect 3988 12434 4016 12650
rect 3896 12406 4016 12434
rect 3792 12232 3844 12238
rect 3792 12174 3844 12180
rect 3424 11892 3476 11898
rect 3424 11834 3476 11840
rect 3424 11620 3476 11626
rect 3424 11562 3476 11568
rect 3332 11280 3384 11286
rect 3332 11222 3384 11228
rect 3332 11008 3384 11014
rect 3332 10950 3384 10956
rect 3160 10118 3280 10146
rect 3056 9988 3108 9994
rect 3056 9930 3108 9936
rect 3054 9752 3110 9761
rect 3054 9687 3056 9696
rect 3108 9687 3110 9696
rect 3056 9658 3108 9664
rect 3056 9512 3108 9518
rect 3056 9454 3108 9460
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 2976 8090 3004 8910
rect 3068 8430 3096 9454
rect 3160 8634 3188 10118
rect 3240 10056 3292 10062
rect 3240 9998 3292 10004
rect 3252 9722 3280 9998
rect 3240 9716 3292 9722
rect 3240 9658 3292 9664
rect 3344 9602 3372 10950
rect 3436 10112 3464 11562
rect 3804 11558 3832 12174
rect 3896 11694 3924 12406
rect 3976 12368 4028 12374
rect 3974 12336 3976 12345
rect 4028 12336 4030 12345
rect 3974 12271 4030 12280
rect 3976 12096 4028 12102
rect 3976 12038 4028 12044
rect 3988 11898 4016 12038
rect 3976 11892 4028 11898
rect 3976 11834 4028 11840
rect 3884 11688 3936 11694
rect 3884 11630 3936 11636
rect 3976 11688 4028 11694
rect 3976 11630 4028 11636
rect 3792 11552 3844 11558
rect 3792 11494 3844 11500
rect 3884 11552 3936 11558
rect 3884 11494 3936 11500
rect 3549 11452 3857 11461
rect 3549 11450 3555 11452
rect 3611 11450 3635 11452
rect 3691 11450 3715 11452
rect 3771 11450 3795 11452
rect 3851 11450 3857 11452
rect 3611 11398 3613 11450
rect 3793 11398 3795 11450
rect 3549 11396 3555 11398
rect 3611 11396 3635 11398
rect 3691 11396 3715 11398
rect 3771 11396 3795 11398
rect 3851 11396 3857 11398
rect 3549 11387 3857 11396
rect 3896 11336 3924 11494
rect 3712 11308 3924 11336
rect 3712 11014 3740 11308
rect 3988 11098 4016 11630
rect 3896 11070 4016 11098
rect 3700 11008 3752 11014
rect 3700 10950 3752 10956
rect 3896 10713 3924 11070
rect 3976 11008 4028 11014
rect 3976 10950 4028 10956
rect 3882 10704 3938 10713
rect 3988 10674 4016 10950
rect 3882 10639 3938 10648
rect 3976 10668 4028 10674
rect 3976 10610 4028 10616
rect 3549 10364 3857 10373
rect 3549 10362 3555 10364
rect 3611 10362 3635 10364
rect 3691 10362 3715 10364
rect 3771 10362 3795 10364
rect 3851 10362 3857 10364
rect 3611 10310 3613 10362
rect 3793 10310 3795 10362
rect 3549 10308 3555 10310
rect 3611 10308 3635 10310
rect 3691 10308 3715 10310
rect 3771 10308 3795 10310
rect 3851 10308 3857 10310
rect 3549 10299 3857 10308
rect 3608 10260 3660 10266
rect 3608 10202 3660 10208
rect 3516 10124 3568 10130
rect 3436 10084 3516 10112
rect 3516 10066 3568 10072
rect 3424 9648 3476 9654
rect 3252 9574 3372 9602
rect 3422 9616 3424 9625
rect 3476 9616 3478 9625
rect 3148 8628 3200 8634
rect 3148 8570 3200 8576
rect 3148 8492 3200 8498
rect 3252 8480 3280 9574
rect 3422 9551 3478 9560
rect 3528 9500 3556 10066
rect 3620 10062 3648 10202
rect 3884 10124 3936 10130
rect 3884 10066 3936 10072
rect 3608 10056 3660 10062
rect 3608 9998 3660 10004
rect 3608 9920 3660 9926
rect 3608 9862 3660 9868
rect 3620 9761 3648 9862
rect 3606 9752 3662 9761
rect 3606 9687 3662 9696
rect 3790 9752 3846 9761
rect 3790 9687 3846 9696
rect 3620 9586 3648 9687
rect 3608 9580 3660 9586
rect 3608 9522 3660 9528
rect 3700 9580 3752 9586
rect 3700 9522 3752 9528
rect 3330 9480 3386 9489
rect 3330 9415 3386 9424
rect 3436 9472 3556 9500
rect 3712 9489 3740 9522
rect 3698 9480 3754 9489
rect 3344 8974 3372 9415
rect 3332 8968 3384 8974
rect 3332 8910 3384 8916
rect 3332 8628 3384 8634
rect 3332 8570 3384 8576
rect 3200 8452 3280 8480
rect 3148 8434 3200 8440
rect 3056 8424 3108 8430
rect 3056 8366 3108 8372
rect 2964 8084 3016 8090
rect 2964 8026 3016 8032
rect 2884 7942 3004 7970
rect 3068 7954 3096 8366
rect 2780 7472 2832 7478
rect 2780 7414 2832 7420
rect 2792 6866 2820 7414
rect 2870 6896 2926 6905
rect 2780 6860 2832 6866
rect 2870 6831 2926 6840
rect 2780 6802 2832 6808
rect 2884 6798 2912 6831
rect 2872 6792 2924 6798
rect 2872 6734 2924 6740
rect 2872 6452 2924 6458
rect 2872 6394 2924 6400
rect 2780 6316 2832 6322
rect 2780 6258 2832 6264
rect 2688 6248 2740 6254
rect 2688 6190 2740 6196
rect 2792 5953 2820 6258
rect 2778 5944 2834 5953
rect 2778 5879 2834 5888
rect 2884 5778 2912 6394
rect 2872 5772 2924 5778
rect 2872 5714 2924 5720
rect 2502 5672 2558 5681
rect 2502 5607 2558 5616
rect 2596 5636 2648 5642
rect 2596 5578 2648 5584
rect 2688 5636 2740 5642
rect 2688 5578 2740 5584
rect 2504 5024 2556 5030
rect 2504 4966 2556 4972
rect 2516 4729 2544 4966
rect 2502 4720 2558 4729
rect 2608 4690 2636 5578
rect 2502 4655 2558 4664
rect 2596 4684 2648 4690
rect 2596 4626 2648 4632
rect 2412 4616 2464 4622
rect 2412 4558 2464 4564
rect 2596 4548 2648 4554
rect 2596 4490 2648 4496
rect 2412 4480 2464 4486
rect 2412 4422 2464 4428
rect 2424 3194 2452 4422
rect 2504 3460 2556 3466
rect 2504 3402 2556 3408
rect 2412 3188 2464 3194
rect 2412 3130 2464 3136
rect 2516 2990 2544 3402
rect 1860 2916 1912 2922
rect 1860 2858 1912 2864
rect 1964 2910 2360 2938
rect 2504 2984 2556 2990
rect 2504 2926 2556 2932
rect 1768 2848 1820 2854
rect 1768 2790 1820 2796
rect 1780 2417 1808 2790
rect 1766 2408 1822 2417
rect 1766 2343 1822 2352
rect 1872 1970 1900 2858
rect 1860 1964 1912 1970
rect 1860 1906 1912 1912
rect 1582 1320 1638 1329
rect 1582 1255 1638 1264
rect 1964 1034 1992 2910
rect 2044 2848 2096 2854
rect 2044 2790 2096 2796
rect 2136 2848 2188 2854
rect 2136 2790 2188 2796
rect 2056 2514 2084 2790
rect 2044 2508 2096 2514
rect 2044 2450 2096 2456
rect 1780 1006 1992 1034
rect 1504 870 1624 898
rect 1504 800 1532 870
rect 1030 640 1086 649
rect 1030 575 1086 584
rect 1490 0 1546 800
rect 1596 762 1624 870
rect 1780 762 1808 1006
rect 1872 870 1992 898
rect 1872 800 1900 870
rect 1596 734 1808 762
rect 1858 0 1914 800
rect 1964 762 1992 870
rect 2148 762 2176 2790
rect 2226 2544 2282 2553
rect 2226 2479 2282 2488
rect 2240 800 2268 2479
rect 2608 800 2636 4490
rect 2700 4010 2728 5578
rect 2884 5114 2912 5714
rect 2792 5086 2912 5114
rect 2792 4146 2820 5086
rect 2872 5024 2924 5030
rect 2872 4966 2924 4972
rect 2884 4758 2912 4966
rect 2872 4752 2924 4758
rect 2872 4694 2924 4700
rect 2870 4448 2926 4457
rect 2870 4383 2926 4392
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 2688 4004 2740 4010
rect 2688 3946 2740 3952
rect 2792 3534 2820 4082
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 2688 3052 2740 3058
rect 2688 2994 2740 3000
rect 2700 2961 2728 2994
rect 2686 2952 2742 2961
rect 2686 2887 2742 2896
rect 2778 2680 2834 2689
rect 2778 2615 2780 2624
rect 2832 2615 2834 2624
rect 2780 2586 2832 2592
rect 2686 2544 2742 2553
rect 2686 2479 2742 2488
rect 2700 2378 2728 2479
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 2688 2372 2740 2378
rect 2688 2314 2740 2320
rect 2792 1057 2820 2382
rect 2884 1442 2912 4383
rect 2976 1601 3004 7942
rect 3056 7948 3108 7954
rect 3056 7890 3108 7896
rect 3160 7834 3188 8434
rect 3240 8016 3292 8022
rect 3240 7958 3292 7964
rect 3068 7806 3188 7834
rect 3068 5273 3096 7806
rect 3252 6798 3280 7958
rect 3148 6792 3200 6798
rect 3146 6760 3148 6769
rect 3240 6792 3292 6798
rect 3200 6760 3202 6769
rect 3240 6734 3292 6740
rect 3146 6695 3202 6704
rect 3146 6488 3202 6497
rect 3146 6423 3202 6432
rect 3160 6390 3188 6423
rect 3148 6384 3200 6390
rect 3148 6326 3200 6332
rect 3146 6216 3202 6225
rect 3146 6151 3148 6160
rect 3200 6151 3202 6160
rect 3240 6180 3292 6186
rect 3148 6122 3200 6128
rect 3240 6122 3292 6128
rect 3148 5568 3200 5574
rect 3148 5510 3200 5516
rect 3054 5264 3110 5273
rect 3054 5199 3110 5208
rect 3056 5160 3108 5166
rect 3056 5102 3108 5108
rect 3068 4706 3096 5102
rect 3160 4826 3188 5510
rect 3148 4820 3200 4826
rect 3148 4762 3200 4768
rect 3252 4758 3280 6122
rect 3344 5370 3372 8570
rect 3436 8401 3464 9472
rect 3698 9415 3754 9424
rect 3804 9382 3832 9687
rect 3792 9376 3844 9382
rect 3792 9318 3844 9324
rect 3549 9276 3857 9285
rect 3549 9274 3555 9276
rect 3611 9274 3635 9276
rect 3691 9274 3715 9276
rect 3771 9274 3795 9276
rect 3851 9274 3857 9276
rect 3611 9222 3613 9274
rect 3793 9222 3795 9274
rect 3549 9220 3555 9222
rect 3611 9220 3635 9222
rect 3691 9220 3715 9222
rect 3771 9220 3795 9222
rect 3851 9220 3857 9222
rect 3549 9211 3857 9220
rect 3700 9104 3752 9110
rect 3606 9072 3662 9081
rect 3662 9052 3700 9058
rect 3662 9046 3752 9052
rect 3662 9030 3740 9046
rect 3606 9007 3662 9016
rect 3896 8634 3924 10066
rect 3988 9042 4016 10610
rect 4080 9625 4108 12854
rect 4264 12850 4292 13806
rect 4342 13767 4398 13776
rect 4540 13462 4568 14010
rect 4620 13864 4672 13870
rect 4620 13806 4672 13812
rect 4528 13456 4580 13462
rect 4528 13398 4580 13404
rect 4632 13394 4660 13806
rect 4620 13388 4672 13394
rect 4620 13330 4672 13336
rect 4252 12844 4304 12850
rect 4252 12786 4304 12792
rect 4264 12306 4292 12786
rect 4252 12300 4304 12306
rect 4252 12242 4304 12248
rect 4342 11928 4398 11937
rect 4342 11863 4344 11872
rect 4396 11863 4398 11872
rect 4344 11834 4396 11840
rect 4528 11552 4580 11558
rect 4528 11494 4580 11500
rect 4434 11384 4490 11393
rect 4434 11319 4490 11328
rect 4252 11280 4304 11286
rect 4252 11222 4304 11228
rect 4158 10024 4214 10033
rect 4158 9959 4214 9968
rect 4172 9926 4200 9959
rect 4160 9920 4212 9926
rect 4160 9862 4212 9868
rect 4066 9616 4122 9625
rect 4066 9551 4122 9560
rect 4160 9580 4212 9586
rect 4160 9522 4212 9528
rect 4066 9480 4122 9489
rect 4066 9415 4068 9424
rect 4120 9415 4122 9424
rect 4068 9386 4120 9392
rect 4066 9344 4122 9353
rect 4066 9279 4122 9288
rect 3976 9036 4028 9042
rect 3976 8978 4028 8984
rect 3884 8628 3936 8634
rect 3884 8570 3936 8576
rect 3884 8492 3936 8498
rect 3884 8434 3936 8440
rect 3516 8424 3568 8430
rect 3422 8392 3478 8401
rect 3516 8366 3568 8372
rect 3422 8327 3478 8336
rect 3528 8276 3556 8366
rect 3436 8248 3556 8276
rect 3436 7410 3464 8248
rect 3549 8188 3857 8197
rect 3549 8186 3555 8188
rect 3611 8186 3635 8188
rect 3691 8186 3715 8188
rect 3771 8186 3795 8188
rect 3851 8186 3857 8188
rect 3611 8134 3613 8186
rect 3793 8134 3795 8186
rect 3549 8132 3555 8134
rect 3611 8132 3635 8134
rect 3691 8132 3715 8134
rect 3771 8132 3795 8134
rect 3851 8132 3857 8134
rect 3549 8123 3857 8132
rect 3896 7993 3924 8434
rect 3974 8120 4030 8129
rect 3974 8055 4030 8064
rect 3882 7984 3938 7993
rect 3516 7948 3568 7954
rect 3988 7954 4016 8055
rect 3882 7919 3938 7928
rect 3976 7948 4028 7954
rect 3516 7890 3568 7896
rect 3976 7890 4028 7896
rect 3528 7750 3556 7890
rect 3790 7848 3846 7857
rect 3790 7783 3792 7792
rect 3844 7783 3846 7792
rect 3792 7754 3844 7760
rect 3516 7744 3568 7750
rect 3516 7686 3568 7692
rect 3976 7744 4028 7750
rect 3976 7686 4028 7692
rect 3528 7585 3556 7686
rect 3514 7576 3570 7585
rect 3514 7511 3570 7520
rect 3424 7404 3476 7410
rect 3424 7346 3476 7352
rect 3549 7100 3857 7109
rect 3549 7098 3555 7100
rect 3611 7098 3635 7100
rect 3691 7098 3715 7100
rect 3771 7098 3795 7100
rect 3851 7098 3857 7100
rect 3611 7046 3613 7098
rect 3793 7046 3795 7098
rect 3549 7044 3555 7046
rect 3611 7044 3635 7046
rect 3691 7044 3715 7046
rect 3771 7044 3795 7046
rect 3851 7044 3857 7046
rect 3549 7035 3857 7044
rect 3988 7002 4016 7686
rect 3608 6996 3660 7002
rect 3608 6938 3660 6944
rect 3976 6996 4028 7002
rect 3976 6938 4028 6944
rect 3620 6866 3648 6938
rect 4080 6882 4108 9279
rect 4172 9110 4200 9522
rect 4264 9489 4292 11222
rect 4344 10192 4396 10198
rect 4344 10134 4396 10140
rect 4250 9480 4306 9489
rect 4250 9415 4306 9424
rect 4252 9376 4304 9382
rect 4252 9318 4304 9324
rect 4160 9104 4212 9110
rect 4160 9046 4212 9052
rect 4264 9042 4292 9318
rect 4356 9042 4384 10134
rect 4448 9466 4476 11319
rect 4540 9586 4568 11494
rect 4632 11257 4660 13330
rect 4724 11665 4752 15370
rect 4816 14958 4844 16544
rect 4908 16454 4936 18566
rect 5000 17338 5028 18566
rect 5092 18426 5120 18686
rect 5080 18420 5132 18426
rect 5080 18362 5132 18368
rect 5184 18193 5212 19774
rect 5368 19446 5396 20198
rect 5460 20182 5580 20198
rect 5460 19786 5488 20182
rect 5630 20088 5686 20097
rect 5630 20023 5686 20032
rect 5448 19780 5500 19786
rect 5448 19722 5500 19728
rect 5460 19530 5488 19722
rect 5460 19514 5580 19530
rect 5460 19508 5592 19514
rect 5460 19502 5540 19508
rect 5540 19450 5592 19456
rect 5356 19440 5408 19446
rect 5356 19382 5408 19388
rect 5644 19334 5672 20023
rect 5736 19938 5764 22200
rect 6104 20890 6132 22200
rect 6012 20862 6132 20890
rect 6472 20890 6500 22200
rect 6472 20862 6592 20890
rect 5908 20392 5960 20398
rect 5908 20334 5960 20340
rect 5736 19910 5856 19938
rect 5724 19780 5776 19786
rect 5724 19722 5776 19728
rect 5552 19306 5672 19334
rect 5354 19000 5410 19009
rect 5354 18935 5410 18944
rect 5368 18902 5396 18935
rect 5356 18896 5408 18902
rect 5356 18838 5408 18844
rect 5356 18624 5408 18630
rect 5356 18566 5408 18572
rect 5262 18320 5318 18329
rect 5262 18255 5264 18264
rect 5316 18255 5318 18264
rect 5264 18226 5316 18232
rect 5170 18184 5226 18193
rect 5170 18119 5226 18128
rect 5264 18080 5316 18086
rect 5264 18022 5316 18028
rect 5276 17882 5304 18022
rect 5264 17876 5316 17882
rect 5264 17818 5316 17824
rect 5264 17604 5316 17610
rect 5264 17546 5316 17552
rect 4988 17332 5040 17338
rect 4988 17274 5040 17280
rect 4988 17196 5040 17202
rect 4988 17138 5040 17144
rect 4896 16448 4948 16454
rect 4896 16390 4948 16396
rect 5000 15706 5028 17138
rect 5078 17096 5134 17105
rect 5078 17031 5134 17040
rect 5172 17060 5224 17066
rect 4988 15700 5040 15706
rect 4988 15642 5040 15648
rect 4988 15496 5040 15502
rect 5092 15484 5120 17031
rect 5172 17002 5224 17008
rect 5184 16017 5212 17002
rect 5276 16182 5304 17546
rect 5368 16658 5396 18566
rect 5552 18465 5580 19306
rect 5632 18828 5684 18834
rect 5632 18770 5684 18776
rect 5538 18456 5594 18465
rect 5538 18391 5594 18400
rect 5448 18284 5500 18290
rect 5448 18226 5500 18232
rect 5460 17921 5488 18226
rect 5540 18216 5592 18222
rect 5540 18158 5592 18164
rect 5446 17912 5502 17921
rect 5552 17882 5580 18158
rect 5446 17847 5502 17856
rect 5540 17876 5592 17882
rect 5540 17818 5592 17824
rect 5644 17610 5672 18770
rect 5632 17604 5684 17610
rect 5632 17546 5684 17552
rect 5448 17536 5500 17542
rect 5448 17478 5500 17484
rect 5460 17134 5488 17478
rect 5538 17368 5594 17377
rect 5538 17303 5540 17312
rect 5592 17303 5594 17312
rect 5540 17274 5592 17280
rect 5538 17232 5594 17241
rect 5538 17167 5594 17176
rect 5448 17128 5500 17134
rect 5448 17070 5500 17076
rect 5460 16658 5488 17070
rect 5356 16652 5408 16658
rect 5356 16594 5408 16600
rect 5448 16652 5500 16658
rect 5448 16594 5500 16600
rect 5264 16176 5316 16182
rect 5264 16118 5316 16124
rect 5170 16008 5226 16017
rect 5170 15943 5226 15952
rect 5448 15904 5500 15910
rect 5448 15846 5500 15852
rect 5460 15609 5488 15846
rect 5262 15600 5318 15609
rect 5262 15535 5318 15544
rect 5446 15600 5502 15609
rect 5446 15535 5502 15544
rect 5276 15502 5304 15535
rect 5040 15456 5120 15484
rect 4988 15438 5040 15444
rect 5092 15314 5120 15456
rect 5264 15496 5316 15502
rect 5264 15438 5316 15444
rect 5092 15286 5396 15314
rect 5368 15162 5396 15286
rect 5356 15156 5408 15162
rect 5356 15098 5408 15104
rect 4988 15088 5040 15094
rect 4988 15030 5040 15036
rect 4896 15020 4948 15026
rect 4896 14962 4948 14968
rect 4804 14952 4856 14958
rect 4804 14894 4856 14900
rect 4908 13870 4936 14962
rect 4896 13864 4948 13870
rect 4896 13806 4948 13812
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 4710 11656 4766 11665
rect 4710 11591 4766 11600
rect 4816 11558 4844 12174
rect 4804 11552 4856 11558
rect 4802 11520 4804 11529
rect 4856 11520 4858 11529
rect 4802 11455 4858 11464
rect 4618 11248 4674 11257
rect 4618 11183 4674 11192
rect 4710 10704 4766 10713
rect 4710 10639 4766 10648
rect 4620 10260 4672 10266
rect 4620 10202 4672 10208
rect 4528 9580 4580 9586
rect 4528 9522 4580 9528
rect 4448 9438 4568 9466
rect 4436 9376 4488 9382
rect 4436 9318 4488 9324
rect 4252 9036 4304 9042
rect 4252 8978 4304 8984
rect 4344 9036 4396 9042
rect 4344 8978 4396 8984
rect 4448 8974 4476 9318
rect 4436 8968 4488 8974
rect 4436 8910 4488 8916
rect 4160 8832 4212 8838
rect 4160 8774 4212 8780
rect 3608 6860 3660 6866
rect 3608 6802 3660 6808
rect 3988 6854 4108 6882
rect 3424 6792 3476 6798
rect 3424 6734 3476 6740
rect 3436 5522 3464 6734
rect 3884 6724 3936 6730
rect 3884 6666 3936 6672
rect 3549 6012 3857 6021
rect 3549 6010 3555 6012
rect 3611 6010 3635 6012
rect 3691 6010 3715 6012
rect 3771 6010 3795 6012
rect 3851 6010 3857 6012
rect 3611 5958 3613 6010
rect 3793 5958 3795 6010
rect 3549 5956 3555 5958
rect 3611 5956 3635 5958
rect 3691 5956 3715 5958
rect 3771 5956 3795 5958
rect 3851 5956 3857 5958
rect 3549 5947 3857 5956
rect 3896 5914 3924 6666
rect 3884 5908 3936 5914
rect 3884 5850 3936 5856
rect 3884 5772 3936 5778
rect 3884 5714 3936 5720
rect 3896 5681 3924 5714
rect 3882 5672 3938 5681
rect 3882 5607 3938 5616
rect 3436 5494 3556 5522
rect 3332 5364 3384 5370
rect 3384 5324 3464 5352
rect 3332 5306 3384 5312
rect 3330 5264 3386 5273
rect 3330 5199 3332 5208
rect 3384 5199 3386 5208
rect 3332 5170 3384 5176
rect 3332 5024 3384 5030
rect 3332 4966 3384 4972
rect 3240 4752 3292 4758
rect 3068 4678 3188 4706
rect 3240 4694 3292 4700
rect 3344 4690 3372 4966
rect 3056 3392 3108 3398
rect 3056 3334 3108 3340
rect 2962 1592 3018 1601
rect 2962 1527 3018 1536
rect 2884 1414 3004 1442
rect 2778 1048 2834 1057
rect 2778 983 2834 992
rect 2976 800 3004 1414
rect 1964 734 2176 762
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3068 762 3096 3334
rect 3160 1193 3188 4678
rect 3332 4684 3384 4690
rect 3332 4626 3384 4632
rect 3436 4570 3464 5324
rect 3528 5302 3556 5494
rect 3516 5296 3568 5302
rect 3516 5238 3568 5244
rect 3884 5228 3936 5234
rect 3884 5170 3936 5176
rect 3549 4924 3857 4933
rect 3549 4922 3555 4924
rect 3611 4922 3635 4924
rect 3691 4922 3715 4924
rect 3771 4922 3795 4924
rect 3851 4922 3857 4924
rect 3611 4870 3613 4922
rect 3793 4870 3795 4922
rect 3549 4868 3555 4870
rect 3611 4868 3635 4870
rect 3691 4868 3715 4870
rect 3771 4868 3795 4870
rect 3851 4868 3857 4870
rect 3549 4859 3857 4868
rect 3896 4593 3924 5170
rect 3252 4542 3464 4570
rect 3882 4584 3938 4593
rect 3252 2582 3280 4542
rect 3882 4519 3938 4528
rect 3332 4140 3384 4146
rect 3332 4082 3384 4088
rect 3344 3670 3372 4082
rect 3549 3836 3857 3845
rect 3549 3834 3555 3836
rect 3611 3834 3635 3836
rect 3691 3834 3715 3836
rect 3771 3834 3795 3836
rect 3851 3834 3857 3836
rect 3611 3782 3613 3834
rect 3793 3782 3795 3834
rect 3549 3780 3555 3782
rect 3611 3780 3635 3782
rect 3691 3780 3715 3782
rect 3771 3780 3795 3782
rect 3851 3780 3857 3782
rect 3549 3771 3857 3780
rect 3516 3732 3568 3738
rect 3516 3674 3568 3680
rect 3332 3664 3384 3670
rect 3332 3606 3384 3612
rect 3422 3632 3478 3641
rect 3422 3567 3478 3576
rect 3436 3534 3464 3567
rect 3424 3528 3476 3534
rect 3424 3470 3476 3476
rect 3436 3097 3464 3470
rect 3422 3088 3478 3097
rect 3332 3052 3384 3058
rect 3422 3023 3478 3032
rect 3332 2994 3384 3000
rect 3240 2576 3292 2582
rect 3240 2518 3292 2524
rect 3344 2009 3372 2994
rect 3528 2990 3556 3674
rect 3792 3664 3844 3670
rect 3790 3632 3792 3641
rect 3844 3632 3846 3641
rect 3790 3567 3846 3576
rect 3884 3392 3936 3398
rect 3884 3334 3936 3340
rect 3516 2984 3568 2990
rect 3516 2926 3568 2932
rect 3549 2748 3857 2757
rect 3549 2746 3555 2748
rect 3611 2746 3635 2748
rect 3691 2746 3715 2748
rect 3771 2746 3795 2748
rect 3851 2746 3857 2748
rect 3611 2694 3613 2746
rect 3793 2694 3795 2746
rect 3549 2692 3555 2694
rect 3611 2692 3635 2694
rect 3691 2692 3715 2694
rect 3771 2692 3795 2694
rect 3851 2692 3857 2694
rect 3549 2683 3857 2692
rect 3608 2576 3660 2582
rect 3606 2544 3608 2553
rect 3700 2576 3752 2582
rect 3660 2544 3662 2553
rect 3700 2518 3752 2524
rect 3606 2479 3662 2488
rect 3608 2372 3660 2378
rect 3608 2314 3660 2320
rect 3330 2000 3386 2009
rect 3330 1935 3386 1944
rect 3620 1766 3648 2314
rect 3608 1760 3660 1766
rect 3608 1702 3660 1708
rect 3146 1184 3202 1193
rect 3146 1119 3202 1128
rect 3422 1184 3478 1193
rect 3422 1119 3478 1128
rect 3436 921 3464 1119
rect 3422 912 3478 921
rect 3252 870 3372 898
rect 3252 762 3280 870
rect 3344 800 3372 870
rect 3422 847 3478 856
rect 3712 898 3740 2518
rect 3790 2272 3846 2281
rect 3790 2207 3846 2216
rect 3804 1834 3832 2207
rect 3792 1828 3844 1834
rect 3792 1770 3844 1776
rect 3896 1193 3924 3334
rect 3988 3233 4016 6854
rect 4068 6724 4120 6730
rect 4172 6712 4200 8774
rect 4540 8498 4568 9438
rect 4632 9178 4660 10202
rect 4724 9926 4752 10639
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 4816 10062 4844 10542
rect 4804 10056 4856 10062
rect 4804 9998 4856 10004
rect 4712 9920 4764 9926
rect 4710 9888 4712 9897
rect 4764 9888 4766 9897
rect 4710 9823 4766 9832
rect 4712 9580 4764 9586
rect 4712 9522 4764 9528
rect 4620 9172 4672 9178
rect 4620 9114 4672 9120
rect 4618 9072 4674 9081
rect 4618 9007 4674 9016
rect 4528 8492 4580 8498
rect 4528 8434 4580 8440
rect 4632 8430 4660 9007
rect 4724 8634 4752 9522
rect 4804 9512 4856 9518
rect 4804 9454 4856 9460
rect 4816 9110 4844 9454
rect 4804 9104 4856 9110
rect 4804 9046 4856 9052
rect 4802 8664 4858 8673
rect 4712 8628 4764 8634
rect 4802 8599 4858 8608
rect 4712 8570 4764 8576
rect 4816 8498 4844 8599
rect 4804 8492 4856 8498
rect 4724 8452 4804 8480
rect 4620 8424 4672 8430
rect 4618 8392 4620 8401
rect 4672 8392 4674 8401
rect 4618 8327 4674 8336
rect 4252 8288 4304 8294
rect 4252 8230 4304 8236
rect 4264 7954 4292 8230
rect 4724 8072 4752 8452
rect 4804 8434 4856 8440
rect 4804 8288 4856 8294
rect 4804 8230 4856 8236
rect 4632 8044 4752 8072
rect 4252 7948 4304 7954
rect 4252 7890 4304 7896
rect 4344 7948 4396 7954
rect 4344 7890 4396 7896
rect 4252 7200 4304 7206
rect 4356 7188 4384 7890
rect 4528 7812 4580 7818
rect 4528 7754 4580 7760
rect 4540 7546 4568 7754
rect 4632 7562 4660 8044
rect 4710 7984 4766 7993
rect 4710 7919 4766 7928
rect 4724 7750 4752 7919
rect 4816 7886 4844 8230
rect 4908 7954 4936 13806
rect 5000 8090 5028 15030
rect 5552 14618 5580 17167
rect 5644 16658 5672 17546
rect 5632 16652 5684 16658
rect 5632 16594 5684 16600
rect 5644 16250 5672 16594
rect 5632 16244 5684 16250
rect 5632 16186 5684 16192
rect 5540 14612 5592 14618
rect 5540 14554 5592 14560
rect 5356 14340 5408 14346
rect 5356 14282 5408 14288
rect 5172 14272 5224 14278
rect 5172 14214 5224 14220
rect 5184 13870 5212 14214
rect 5264 14000 5316 14006
rect 5264 13942 5316 13948
rect 5172 13864 5224 13870
rect 5172 13806 5224 13812
rect 5276 13530 5304 13942
rect 5264 13524 5316 13530
rect 5264 13466 5316 13472
rect 5368 13394 5396 14282
rect 5630 14104 5686 14113
rect 5630 14039 5686 14048
rect 5448 13864 5500 13870
rect 5448 13806 5500 13812
rect 5460 13530 5488 13806
rect 5448 13524 5500 13530
rect 5448 13466 5500 13472
rect 5644 13462 5672 14039
rect 5632 13456 5684 13462
rect 5632 13398 5684 13404
rect 5356 13388 5408 13394
rect 5356 13330 5408 13336
rect 5264 13252 5316 13258
rect 5264 13194 5316 13200
rect 5172 12776 5224 12782
rect 5172 12718 5224 12724
rect 5184 12442 5212 12718
rect 5172 12436 5224 12442
rect 5276 12434 5304 13194
rect 5276 12406 5488 12434
rect 5172 12378 5224 12384
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 5092 8974 5120 11494
rect 5356 11144 5408 11150
rect 5356 11086 5408 11092
rect 5172 10464 5224 10470
rect 5172 10406 5224 10412
rect 5080 8968 5132 8974
rect 5080 8910 5132 8916
rect 5092 8362 5120 8910
rect 5080 8356 5132 8362
rect 5080 8298 5132 8304
rect 5184 8294 5212 10406
rect 5368 10266 5396 11086
rect 5356 10260 5408 10266
rect 5356 10202 5408 10208
rect 5356 10056 5408 10062
rect 5356 9998 5408 10004
rect 5264 9580 5316 9586
rect 5264 9522 5316 9528
rect 5276 9178 5304 9522
rect 5264 9172 5316 9178
rect 5264 9114 5316 9120
rect 5264 8832 5316 8838
rect 5264 8774 5316 8780
rect 5276 8673 5304 8774
rect 5262 8664 5318 8673
rect 5262 8599 5318 8608
rect 5262 8528 5318 8537
rect 5368 8514 5396 9998
rect 5460 9602 5488 12406
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5552 11218 5580 12174
rect 5632 12164 5684 12170
rect 5632 12106 5684 12112
rect 5644 11694 5672 12106
rect 5736 11801 5764 19722
rect 5828 18737 5856 19910
rect 5920 18873 5948 20334
rect 5906 18864 5962 18873
rect 5906 18799 5962 18808
rect 5814 18728 5870 18737
rect 5814 18663 5870 18672
rect 5816 18624 5868 18630
rect 5816 18566 5868 18572
rect 5908 18624 5960 18630
rect 5908 18566 5960 18572
rect 5828 18426 5856 18566
rect 5920 18426 5948 18566
rect 5816 18420 5868 18426
rect 5816 18362 5868 18368
rect 5908 18420 5960 18426
rect 5908 18362 5960 18368
rect 5814 18320 5870 18329
rect 5814 18255 5816 18264
rect 5868 18255 5870 18264
rect 5816 18226 5868 18232
rect 5828 16969 5856 18226
rect 6012 18086 6040 20862
rect 6148 20700 6456 20709
rect 6148 20698 6154 20700
rect 6210 20698 6234 20700
rect 6290 20698 6314 20700
rect 6370 20698 6394 20700
rect 6450 20698 6456 20700
rect 6210 20646 6212 20698
rect 6392 20646 6394 20698
rect 6148 20644 6154 20646
rect 6210 20644 6234 20646
rect 6290 20644 6314 20646
rect 6370 20644 6394 20646
rect 6450 20644 6456 20646
rect 6148 20635 6456 20644
rect 6148 19612 6456 19621
rect 6148 19610 6154 19612
rect 6210 19610 6234 19612
rect 6290 19610 6314 19612
rect 6370 19610 6394 19612
rect 6450 19610 6456 19612
rect 6210 19558 6212 19610
rect 6392 19558 6394 19610
rect 6148 19556 6154 19558
rect 6210 19556 6234 19558
rect 6290 19556 6314 19558
rect 6370 19556 6394 19558
rect 6450 19556 6456 19558
rect 6148 19547 6456 19556
rect 6564 19394 6592 20862
rect 6840 20346 6868 22200
rect 7102 21448 7158 21457
rect 7102 21383 7158 21392
rect 7116 21185 7144 21383
rect 7102 21176 7158 21185
rect 7102 21111 7158 21120
rect 7104 20460 7156 20466
rect 7104 20402 7156 20408
rect 6472 19366 6592 19394
rect 6656 20318 6868 20346
rect 6276 19304 6328 19310
rect 6472 19281 6500 19366
rect 6276 19246 6328 19252
rect 6458 19272 6514 19281
rect 6288 18970 6316 19246
rect 6458 19207 6514 19216
rect 6276 18964 6328 18970
rect 6276 18906 6328 18912
rect 6288 18766 6316 18906
rect 6276 18760 6328 18766
rect 6472 18737 6500 19207
rect 6552 19168 6604 19174
rect 6552 19110 6604 19116
rect 6276 18702 6328 18708
rect 6458 18728 6514 18737
rect 6458 18663 6514 18672
rect 6564 18578 6592 19110
rect 6656 18698 6684 20318
rect 6828 20256 6880 20262
rect 6828 20198 6880 20204
rect 6736 20052 6788 20058
rect 6736 19994 6788 20000
rect 6748 19446 6776 19994
rect 6840 19854 6868 20198
rect 6828 19848 6880 19854
rect 6828 19790 6880 19796
rect 6736 19440 6788 19446
rect 6736 19382 6788 19388
rect 7116 19378 7144 20402
rect 7104 19372 7156 19378
rect 7104 19314 7156 19320
rect 7012 19304 7064 19310
rect 7012 19246 7064 19252
rect 7024 19174 7052 19246
rect 6736 19168 6788 19174
rect 6920 19168 6972 19174
rect 6788 19128 6868 19156
rect 6736 19110 6788 19116
rect 6736 18964 6788 18970
rect 6736 18906 6788 18912
rect 6644 18692 6696 18698
rect 6644 18634 6696 18640
rect 6564 18550 6684 18578
rect 6148 18524 6456 18533
rect 6148 18522 6154 18524
rect 6210 18522 6234 18524
rect 6290 18522 6314 18524
rect 6370 18522 6394 18524
rect 6450 18522 6456 18524
rect 6210 18470 6212 18522
rect 6392 18470 6394 18522
rect 6148 18468 6154 18470
rect 6210 18468 6234 18470
rect 6290 18468 6314 18470
rect 6370 18468 6394 18470
rect 6450 18468 6456 18470
rect 6148 18459 6456 18468
rect 6552 18284 6604 18290
rect 6552 18226 6604 18232
rect 6184 18216 6236 18222
rect 6184 18158 6236 18164
rect 6368 18216 6420 18222
rect 6368 18158 6420 18164
rect 6000 18080 6052 18086
rect 6000 18022 6052 18028
rect 5906 17912 5962 17921
rect 5906 17847 5962 17856
rect 5920 17746 5948 17847
rect 6012 17814 6040 18022
rect 6000 17808 6052 17814
rect 6000 17750 6052 17756
rect 5908 17740 5960 17746
rect 5908 17682 5960 17688
rect 6092 17672 6144 17678
rect 6012 17632 6092 17660
rect 5906 17504 5962 17513
rect 5906 17439 5962 17448
rect 5920 17202 5948 17439
rect 5908 17196 5960 17202
rect 5908 17138 5960 17144
rect 6012 16998 6040 17632
rect 6092 17614 6144 17620
rect 6196 17542 6224 18158
rect 6276 18080 6328 18086
rect 6276 18022 6328 18028
rect 6288 17610 6316 18022
rect 6380 17678 6408 18158
rect 6368 17672 6420 17678
rect 6368 17614 6420 17620
rect 6276 17604 6328 17610
rect 6276 17546 6328 17552
rect 6184 17536 6236 17542
rect 6184 17478 6236 17484
rect 6148 17436 6456 17445
rect 6148 17434 6154 17436
rect 6210 17434 6234 17436
rect 6290 17434 6314 17436
rect 6370 17434 6394 17436
rect 6450 17434 6456 17436
rect 6210 17382 6212 17434
rect 6392 17382 6394 17434
rect 6148 17380 6154 17382
rect 6210 17380 6234 17382
rect 6290 17380 6314 17382
rect 6370 17380 6394 17382
rect 6450 17380 6456 17382
rect 6148 17371 6456 17380
rect 6276 17332 6328 17338
rect 6276 17274 6328 17280
rect 6184 17128 6236 17134
rect 6184 17070 6236 17076
rect 6000 16992 6052 16998
rect 5814 16960 5870 16969
rect 6000 16934 6052 16940
rect 5814 16895 5870 16904
rect 5816 16788 5868 16794
rect 5816 16730 5868 16736
rect 5828 11880 5856 16730
rect 6000 16720 6052 16726
rect 6000 16662 6052 16668
rect 5908 16516 5960 16522
rect 5908 16458 5960 16464
rect 5920 15638 5948 16458
rect 6012 16250 6040 16662
rect 6196 16658 6224 17070
rect 6288 16794 6316 17274
rect 6276 16788 6328 16794
rect 6276 16730 6328 16736
rect 6184 16652 6236 16658
rect 6184 16594 6236 16600
rect 6148 16348 6456 16357
rect 6148 16346 6154 16348
rect 6210 16346 6234 16348
rect 6290 16346 6314 16348
rect 6370 16346 6394 16348
rect 6450 16346 6456 16348
rect 6210 16294 6212 16346
rect 6392 16294 6394 16346
rect 6148 16292 6154 16294
rect 6210 16292 6234 16294
rect 6290 16292 6314 16294
rect 6370 16292 6394 16294
rect 6450 16292 6456 16294
rect 6148 16283 6456 16292
rect 6000 16244 6052 16250
rect 6000 16186 6052 16192
rect 6184 16176 6236 16182
rect 6184 16118 6236 16124
rect 6000 16108 6052 16114
rect 6000 16050 6052 16056
rect 5908 15632 5960 15638
rect 5908 15574 5960 15580
rect 5908 15360 5960 15366
rect 5906 15328 5908 15337
rect 5960 15328 5962 15337
rect 5906 15263 5962 15272
rect 6012 15026 6040 16050
rect 6196 15570 6224 16118
rect 6368 16040 6420 16046
rect 6368 15982 6420 15988
rect 6184 15564 6236 15570
rect 6184 15506 6236 15512
rect 6380 15434 6408 15982
rect 6564 15910 6592 18226
rect 6656 17270 6684 18550
rect 6644 17264 6696 17270
rect 6644 17206 6696 17212
rect 6644 17128 6696 17134
rect 6642 17096 6644 17105
rect 6696 17096 6698 17105
rect 6642 17031 6698 17040
rect 6644 16992 6696 16998
rect 6644 16934 6696 16940
rect 6656 16590 6684 16934
rect 6644 16584 6696 16590
rect 6644 16526 6696 16532
rect 6642 16144 6698 16153
rect 6642 16079 6698 16088
rect 6552 15904 6604 15910
rect 6552 15846 6604 15852
rect 6656 15706 6684 16079
rect 6644 15700 6696 15706
rect 6644 15642 6696 15648
rect 6368 15428 6420 15434
rect 6368 15370 6420 15376
rect 6644 15360 6696 15366
rect 6642 15328 6644 15337
rect 6696 15328 6698 15337
rect 6148 15260 6456 15269
rect 6642 15263 6698 15272
rect 6148 15258 6154 15260
rect 6210 15258 6234 15260
rect 6290 15258 6314 15260
rect 6370 15258 6394 15260
rect 6450 15258 6456 15260
rect 6210 15206 6212 15258
rect 6392 15206 6394 15258
rect 6148 15204 6154 15206
rect 6210 15204 6234 15206
rect 6290 15204 6314 15206
rect 6370 15204 6394 15206
rect 6450 15204 6456 15206
rect 6148 15195 6456 15204
rect 6092 15156 6144 15162
rect 6092 15098 6144 15104
rect 5908 15020 5960 15026
rect 5908 14962 5960 14968
rect 6000 15020 6052 15026
rect 6000 14962 6052 14968
rect 5920 14074 5948 14962
rect 6104 14929 6132 15098
rect 6090 14920 6146 14929
rect 6000 14884 6052 14890
rect 6090 14855 6146 14864
rect 6000 14826 6052 14832
rect 6012 14074 6040 14826
rect 6368 14816 6420 14822
rect 6368 14758 6420 14764
rect 6644 14816 6696 14822
rect 6644 14758 6696 14764
rect 6380 14414 6408 14758
rect 6368 14408 6420 14414
rect 6368 14350 6420 14356
rect 6552 14340 6604 14346
rect 6552 14282 6604 14288
rect 6148 14172 6456 14181
rect 6148 14170 6154 14172
rect 6210 14170 6234 14172
rect 6290 14170 6314 14172
rect 6370 14170 6394 14172
rect 6450 14170 6456 14172
rect 6210 14118 6212 14170
rect 6392 14118 6394 14170
rect 6148 14116 6154 14118
rect 6210 14116 6234 14118
rect 6290 14116 6314 14118
rect 6370 14116 6394 14118
rect 6450 14116 6456 14118
rect 6148 14107 6456 14116
rect 5908 14068 5960 14074
rect 5908 14010 5960 14016
rect 6000 14068 6052 14074
rect 6000 14010 6052 14016
rect 6564 14006 6592 14282
rect 6552 14000 6604 14006
rect 6552 13942 6604 13948
rect 6000 13864 6052 13870
rect 6000 13806 6052 13812
rect 5908 13796 5960 13802
rect 5908 13738 5960 13744
rect 5920 12782 5948 13738
rect 6012 13326 6040 13806
rect 6564 13530 6592 13942
rect 6552 13524 6604 13530
rect 6552 13466 6604 13472
rect 6000 13320 6052 13326
rect 6000 13262 6052 13268
rect 6552 13320 6604 13326
rect 6656 13308 6684 14758
rect 6748 13410 6776 18906
rect 6840 18873 6868 19128
rect 6920 19110 6972 19116
rect 7012 19168 7064 19174
rect 7012 19110 7064 19116
rect 6826 18864 6882 18873
rect 6826 18799 6882 18808
rect 6932 18698 6960 19110
rect 7116 18986 7144 19314
rect 7024 18958 7144 18986
rect 6920 18692 6972 18698
rect 6920 18634 6972 18640
rect 6918 18592 6974 18601
rect 6918 18527 6974 18536
rect 6826 18456 6882 18465
rect 6826 18391 6882 18400
rect 6840 18154 6868 18391
rect 6932 18358 6960 18527
rect 6920 18352 6972 18358
rect 6920 18294 6972 18300
rect 6828 18148 6880 18154
rect 6828 18090 6880 18096
rect 6932 17610 6960 18294
rect 6920 17604 6972 17610
rect 6920 17546 6972 17552
rect 6932 17377 6960 17546
rect 6918 17368 6974 17377
rect 6918 17303 6974 17312
rect 6920 17264 6972 17270
rect 6920 17206 6972 17212
rect 6828 17196 6880 17202
rect 6828 17138 6880 17144
rect 6840 16538 6868 17138
rect 6932 16726 6960 17206
rect 7024 17066 7052 18958
rect 7208 18358 7236 22200
rect 7380 20800 7432 20806
rect 7380 20742 7432 20748
rect 7286 20496 7342 20505
rect 7286 20431 7288 20440
rect 7340 20431 7342 20440
rect 7288 20402 7340 20408
rect 7288 19372 7340 19378
rect 7288 19314 7340 19320
rect 7300 18426 7328 19314
rect 7288 18420 7340 18426
rect 7288 18362 7340 18368
rect 7196 18352 7248 18358
rect 7196 18294 7248 18300
rect 7104 18148 7156 18154
rect 7104 18090 7156 18096
rect 7012 17060 7064 17066
rect 7012 17002 7064 17008
rect 6920 16720 6972 16726
rect 6920 16662 6972 16668
rect 7010 16688 7066 16697
rect 7010 16623 7066 16632
rect 6918 16552 6974 16561
rect 6840 16510 6918 16538
rect 6918 16487 6974 16496
rect 6828 16448 6880 16454
rect 6828 16390 6880 16396
rect 6920 16448 6972 16454
rect 6920 16390 6972 16396
rect 6840 15706 6868 16390
rect 6828 15700 6880 15706
rect 6828 15642 6880 15648
rect 6932 15484 6960 16390
rect 7024 16182 7052 16623
rect 7012 16176 7064 16182
rect 7012 16118 7064 16124
rect 6840 15456 6960 15484
rect 6840 14890 6868 15456
rect 7012 14952 7064 14958
rect 7012 14894 7064 14900
rect 6828 14884 6880 14890
rect 6828 14826 6880 14832
rect 7024 14278 7052 14894
rect 7012 14272 7064 14278
rect 7012 14214 7064 14220
rect 6826 14104 6882 14113
rect 6826 14039 6882 14048
rect 6840 13705 6868 14039
rect 7024 14006 7052 14214
rect 6920 14000 6972 14006
rect 6920 13942 6972 13948
rect 7012 14000 7064 14006
rect 7012 13942 7064 13948
rect 6826 13696 6882 13705
rect 6826 13631 6882 13640
rect 6932 13530 6960 13942
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 6748 13382 7052 13410
rect 6604 13280 6684 13308
rect 6552 13262 6604 13268
rect 6828 13184 6880 13190
rect 6828 13126 6880 13132
rect 6148 13084 6456 13093
rect 6148 13082 6154 13084
rect 6210 13082 6234 13084
rect 6290 13082 6314 13084
rect 6370 13082 6394 13084
rect 6450 13082 6456 13084
rect 6210 13030 6212 13082
rect 6392 13030 6394 13082
rect 6148 13028 6154 13030
rect 6210 13028 6234 13030
rect 6290 13028 6314 13030
rect 6370 13028 6394 13030
rect 6450 13028 6456 13030
rect 6148 13019 6456 13028
rect 6460 12844 6512 12850
rect 6460 12786 6512 12792
rect 5908 12776 5960 12782
rect 5908 12718 5960 12724
rect 5920 12481 5948 12718
rect 6184 12708 6236 12714
rect 6184 12650 6236 12656
rect 5906 12472 5962 12481
rect 5906 12407 5962 12416
rect 6196 12170 6224 12650
rect 6368 12640 6420 12646
rect 6368 12582 6420 12588
rect 6380 12306 6408 12582
rect 6472 12306 6500 12786
rect 6368 12300 6420 12306
rect 6368 12242 6420 12248
rect 6460 12300 6512 12306
rect 6460 12242 6512 12248
rect 6552 12232 6604 12238
rect 6552 12174 6604 12180
rect 6184 12164 6236 12170
rect 6184 12106 6236 12112
rect 6148 11996 6456 12005
rect 6148 11994 6154 11996
rect 6210 11994 6234 11996
rect 6290 11994 6314 11996
rect 6370 11994 6394 11996
rect 6450 11994 6456 11996
rect 6210 11942 6212 11994
rect 6392 11942 6394 11994
rect 6148 11940 6154 11942
rect 6210 11940 6234 11942
rect 6290 11940 6314 11942
rect 6370 11940 6394 11942
rect 6450 11940 6456 11942
rect 6148 11931 6456 11940
rect 5828 11852 5948 11880
rect 5722 11792 5778 11801
rect 5722 11727 5778 11736
rect 5816 11756 5868 11762
rect 5816 11698 5868 11704
rect 5632 11688 5684 11694
rect 5632 11630 5684 11636
rect 5724 11688 5776 11694
rect 5724 11630 5776 11636
rect 5644 11354 5672 11630
rect 5632 11348 5684 11354
rect 5632 11290 5684 11296
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5540 11076 5592 11082
rect 5540 11018 5592 11024
rect 5552 10606 5580 11018
rect 5736 10742 5764 11630
rect 5828 11082 5856 11698
rect 5816 11076 5868 11082
rect 5816 11018 5868 11024
rect 5724 10736 5776 10742
rect 5724 10678 5776 10684
rect 5816 10668 5868 10674
rect 5816 10610 5868 10616
rect 5540 10600 5592 10606
rect 5540 10542 5592 10548
rect 5552 10470 5580 10542
rect 5540 10464 5592 10470
rect 5592 10424 5672 10452
rect 5540 10406 5592 10412
rect 5644 10130 5672 10424
rect 5724 10192 5776 10198
rect 5724 10134 5776 10140
rect 5632 10124 5684 10130
rect 5632 10066 5684 10072
rect 5540 9988 5592 9994
rect 5540 9930 5592 9936
rect 5552 9674 5580 9930
rect 5632 9920 5684 9926
rect 5736 9908 5764 10134
rect 5828 9994 5856 10610
rect 5920 10130 5948 11852
rect 6564 11830 6592 12174
rect 6644 12096 6696 12102
rect 6644 12038 6696 12044
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 6552 11824 6604 11830
rect 6552 11766 6604 11772
rect 6656 11354 6684 12038
rect 6748 11626 6776 12038
rect 6736 11620 6788 11626
rect 6736 11562 6788 11568
rect 6644 11348 6696 11354
rect 6644 11290 6696 11296
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 6552 11144 6604 11150
rect 6552 11086 6604 11092
rect 6000 11008 6052 11014
rect 6000 10950 6052 10956
rect 6012 10810 6040 10950
rect 6148 10908 6456 10917
rect 6148 10906 6154 10908
rect 6210 10906 6234 10908
rect 6290 10906 6314 10908
rect 6370 10906 6394 10908
rect 6450 10906 6456 10908
rect 6210 10854 6212 10906
rect 6392 10854 6394 10906
rect 6148 10852 6154 10854
rect 6210 10852 6234 10854
rect 6290 10852 6314 10854
rect 6370 10852 6394 10854
rect 6450 10852 6456 10854
rect 6148 10843 6456 10852
rect 6564 10810 6592 11086
rect 6000 10804 6052 10810
rect 6000 10746 6052 10752
rect 6552 10804 6604 10810
rect 6552 10746 6604 10752
rect 6368 10600 6420 10606
rect 6368 10542 6420 10548
rect 6380 10266 6408 10542
rect 6564 10470 6592 10746
rect 6552 10464 6604 10470
rect 6552 10406 6604 10412
rect 6550 10296 6606 10305
rect 6368 10260 6420 10266
rect 6550 10231 6606 10240
rect 6368 10202 6420 10208
rect 6564 10130 6592 10231
rect 5908 10124 5960 10130
rect 5908 10066 5960 10072
rect 6552 10124 6604 10130
rect 6552 10066 6604 10072
rect 6460 10056 6512 10062
rect 6460 9998 6512 10004
rect 5816 9988 5868 9994
rect 6000 9988 6052 9994
rect 5816 9930 5868 9936
rect 5929 9948 6000 9976
rect 5929 9908 5957 9948
rect 6000 9930 6052 9936
rect 6472 9926 6500 9998
rect 5684 9880 5764 9908
rect 5889 9880 5957 9908
rect 6460 9920 6512 9926
rect 5632 9862 5684 9868
rect 5889 9674 5917 9880
rect 6460 9862 6512 9868
rect 6644 9920 6696 9926
rect 6644 9862 6696 9868
rect 6148 9820 6456 9829
rect 6148 9818 6154 9820
rect 6210 9818 6234 9820
rect 6290 9818 6314 9820
rect 6370 9818 6394 9820
rect 6450 9818 6456 9820
rect 6210 9766 6212 9818
rect 6392 9766 6394 9818
rect 6148 9764 6154 9766
rect 6210 9764 6234 9766
rect 6290 9764 6314 9766
rect 6370 9764 6394 9766
rect 6450 9764 6456 9766
rect 6148 9755 6456 9764
rect 6656 9674 6684 9862
rect 5552 9646 5856 9674
rect 5889 9646 6040 9674
rect 5460 9574 5764 9602
rect 5632 9512 5684 9518
rect 5632 9454 5684 9460
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 5318 8486 5396 8514
rect 5262 8463 5318 8472
rect 5276 8430 5304 8463
rect 5264 8424 5316 8430
rect 5264 8366 5316 8372
rect 5172 8288 5224 8294
rect 5078 8256 5134 8265
rect 5172 8230 5224 8236
rect 5078 8191 5134 8200
rect 4988 8084 5040 8090
rect 4988 8026 5040 8032
rect 4896 7948 4948 7954
rect 4896 7890 4948 7896
rect 4804 7880 4856 7886
rect 4804 7822 4856 7828
rect 4712 7744 4764 7750
rect 4712 7686 4764 7692
rect 4528 7540 4580 7546
rect 4632 7534 4752 7562
rect 4528 7482 4580 7488
rect 4724 7449 4752 7534
rect 4710 7440 4766 7449
rect 4528 7404 4580 7410
rect 4528 7346 4580 7352
rect 4620 7404 4672 7410
rect 4710 7375 4766 7384
rect 4620 7346 4672 7352
rect 4304 7160 4384 7188
rect 4252 7142 4304 7148
rect 4120 6684 4200 6712
rect 4068 6666 4120 6672
rect 4264 6322 4292 7142
rect 4434 7032 4490 7041
rect 4434 6967 4490 6976
rect 4252 6316 4304 6322
rect 4252 6258 4304 6264
rect 4344 6248 4396 6254
rect 4344 6190 4396 6196
rect 4158 5944 4214 5953
rect 4158 5879 4214 5888
rect 4172 5828 4200 5879
rect 4252 5840 4304 5846
rect 4172 5800 4252 5828
rect 4252 5782 4304 5788
rect 4160 5636 4212 5642
rect 4160 5578 4212 5584
rect 4066 5400 4122 5409
rect 4066 5335 4068 5344
rect 4120 5335 4122 5344
rect 4068 5306 4120 5312
rect 4172 5234 4200 5578
rect 4252 5568 4304 5574
rect 4252 5510 4304 5516
rect 4264 5409 4292 5510
rect 4250 5400 4306 5409
rect 4250 5335 4306 5344
rect 4160 5228 4212 5234
rect 4160 5170 4212 5176
rect 4160 5092 4212 5098
rect 4160 5034 4212 5040
rect 4068 4684 4120 4690
rect 4068 4626 4120 4632
rect 4080 3448 4108 4626
rect 4172 4282 4200 5034
rect 4252 5024 4304 5030
rect 4252 4966 4304 4972
rect 4160 4276 4212 4282
rect 4160 4218 4212 4224
rect 4264 4146 4292 4966
rect 4252 4140 4304 4146
rect 4252 4082 4304 4088
rect 4252 4004 4304 4010
rect 4252 3946 4304 3952
rect 4264 3641 4292 3946
rect 4250 3632 4306 3641
rect 4250 3567 4306 3576
rect 4160 3460 4212 3466
rect 4080 3420 4160 3448
rect 4160 3402 4212 3408
rect 3974 3224 4030 3233
rect 3974 3159 4030 3168
rect 4068 3120 4120 3126
rect 4068 3062 4120 3068
rect 3974 2816 4030 2825
rect 3974 2751 4030 2760
rect 3988 2582 4016 2751
rect 3976 2576 4028 2582
rect 3976 2518 4028 2524
rect 3976 2372 4028 2378
rect 3976 2314 4028 2320
rect 3988 2106 4016 2314
rect 3976 2100 4028 2106
rect 3976 2042 4028 2048
rect 3882 1184 3938 1193
rect 3882 1119 3938 1128
rect 3712 870 3832 898
rect 3712 800 3740 870
rect 3068 734 3280 762
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 3804 762 3832 870
rect 4080 800 4108 3062
rect 4172 2990 4200 3402
rect 4252 3392 4304 3398
rect 4252 3334 4304 3340
rect 4160 2984 4212 2990
rect 4160 2926 4212 2932
rect 4264 2854 4292 3334
rect 4252 2848 4304 2854
rect 4252 2790 4304 2796
rect 4158 2680 4214 2689
rect 4356 2666 4384 6190
rect 4448 5370 4476 6967
rect 4540 6934 4568 7346
rect 4528 6928 4580 6934
rect 4528 6870 4580 6876
rect 4528 6316 4580 6322
rect 4528 6258 4580 6264
rect 4436 5364 4488 5370
rect 4436 5306 4488 5312
rect 4540 5250 4568 6258
rect 4632 6118 4660 7346
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 4632 5681 4660 6054
rect 4618 5672 4674 5681
rect 4618 5607 4674 5616
rect 4448 5222 4568 5250
rect 4448 5030 4476 5222
rect 4436 5024 4488 5030
rect 4724 4978 4752 7375
rect 4816 7342 4844 7822
rect 4896 7744 4948 7750
rect 4896 7686 4948 7692
rect 4908 7478 4936 7686
rect 4896 7472 4948 7478
rect 4896 7414 4948 7420
rect 4804 7336 4856 7342
rect 4804 7278 4856 7284
rect 4816 5953 4844 7278
rect 4908 6322 4936 7414
rect 5092 7002 5120 8191
rect 5172 7948 5224 7954
rect 5172 7890 5224 7896
rect 5184 7546 5212 7890
rect 5172 7540 5224 7546
rect 5172 7482 5224 7488
rect 5172 7200 5224 7206
rect 5172 7142 5224 7148
rect 5080 6996 5132 7002
rect 5080 6938 5132 6944
rect 5080 6792 5132 6798
rect 5080 6734 5132 6740
rect 5092 6662 5120 6734
rect 4988 6656 5040 6662
rect 4988 6598 5040 6604
rect 5080 6656 5132 6662
rect 5080 6598 5132 6604
rect 4896 6316 4948 6322
rect 4896 6258 4948 6264
rect 4896 6112 4948 6118
rect 4896 6054 4948 6060
rect 4802 5944 4858 5953
rect 4802 5879 4858 5888
rect 4436 4966 4488 4972
rect 4540 4950 4752 4978
rect 4436 4548 4488 4554
rect 4436 4490 4488 4496
rect 4448 4282 4476 4490
rect 4436 4276 4488 4282
rect 4436 4218 4488 4224
rect 4434 2952 4490 2961
rect 4434 2887 4490 2896
rect 4264 2650 4384 2666
rect 4158 2615 4214 2624
rect 4252 2644 4384 2650
rect 4172 2582 4200 2615
rect 4304 2638 4384 2644
rect 4252 2586 4304 2592
rect 4160 2576 4212 2582
rect 4160 2518 4212 2524
rect 4448 898 4476 2887
rect 4540 2360 4568 4950
rect 4908 4842 4936 6054
rect 5000 5914 5028 6598
rect 5092 6186 5120 6598
rect 5080 6180 5132 6186
rect 5080 6122 5132 6128
rect 4988 5908 5040 5914
rect 4988 5850 5040 5856
rect 4988 5636 5040 5642
rect 4988 5578 5040 5584
rect 5000 5234 5028 5578
rect 4988 5228 5040 5234
rect 4988 5170 5040 5176
rect 5078 4992 5134 5001
rect 5078 4927 5134 4936
rect 4724 4814 4936 4842
rect 4986 4856 5042 4865
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 4632 3194 4660 3878
rect 4724 3777 4752 4814
rect 4986 4791 5042 4800
rect 4804 4752 4856 4758
rect 4804 4694 4856 4700
rect 4816 4486 4844 4694
rect 4804 4480 4856 4486
rect 4804 4422 4856 4428
rect 5000 4146 5028 4791
rect 5092 4622 5120 4927
rect 5080 4616 5132 4622
rect 5080 4558 5132 4564
rect 5080 4480 5132 4486
rect 5078 4448 5080 4457
rect 5132 4448 5134 4457
rect 5078 4383 5134 4392
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 5080 4072 5132 4078
rect 5080 4014 5132 4020
rect 4896 4004 4948 4010
rect 4896 3946 4948 3952
rect 4710 3768 4766 3777
rect 4710 3703 4766 3712
rect 4802 3632 4858 3641
rect 4802 3567 4858 3576
rect 4712 3460 4764 3466
rect 4712 3402 4764 3408
rect 4724 3194 4752 3402
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 4620 2916 4672 2922
rect 4620 2858 4672 2864
rect 4632 2825 4660 2858
rect 4618 2816 4674 2825
rect 4618 2751 4674 2760
rect 4620 2372 4672 2378
rect 4540 2332 4620 2360
rect 4620 2314 4672 2320
rect 4448 870 4568 898
rect 4448 800 4476 870
rect 3804 734 4016 762
rect 3988 66 4016 734
rect 3976 60 4028 66
rect 3976 2 4028 8
rect 4066 0 4122 800
rect 4434 0 4490 800
rect 4540 762 4568 870
rect 4816 800 4844 3567
rect 4908 3058 4936 3946
rect 4896 3052 4948 3058
rect 4896 2994 4948 3000
rect 4908 2446 4936 2994
rect 4896 2440 4948 2446
rect 4896 2382 4948 2388
rect 4986 2408 5042 2417
rect 4986 2343 5042 2352
rect 5000 1465 5028 2343
rect 4986 1456 5042 1465
rect 4986 1391 5042 1400
rect 5092 1222 5120 4014
rect 5184 3738 5212 7142
rect 5276 6866 5304 8366
rect 5356 8084 5408 8090
rect 5356 8026 5408 8032
rect 5368 7818 5396 8026
rect 5460 8022 5488 9318
rect 5644 9178 5672 9454
rect 5632 9172 5684 9178
rect 5632 9114 5684 9120
rect 5630 9072 5686 9081
rect 5630 9007 5686 9016
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 5448 8016 5500 8022
rect 5448 7958 5500 7964
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 5356 7812 5408 7818
rect 5356 7754 5408 7760
rect 5460 7585 5488 7822
rect 5446 7576 5502 7585
rect 5446 7511 5502 7520
rect 5448 7472 5500 7478
rect 5448 7414 5500 7420
rect 5354 6896 5410 6905
rect 5264 6860 5316 6866
rect 5354 6831 5410 6840
rect 5264 6802 5316 6808
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 5276 4214 5304 6598
rect 5368 6322 5396 6831
rect 5460 6633 5488 7414
rect 5446 6624 5502 6633
rect 5446 6559 5502 6568
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 5368 6225 5396 6258
rect 5354 6216 5410 6225
rect 5354 6151 5410 6160
rect 5356 6112 5408 6118
rect 5356 6054 5408 6060
rect 5448 6112 5500 6118
rect 5448 6054 5500 6060
rect 5368 4758 5396 6054
rect 5460 5817 5488 6054
rect 5446 5808 5502 5817
rect 5446 5743 5502 5752
rect 5552 5386 5580 8774
rect 5644 8634 5672 9007
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 5632 8356 5684 8362
rect 5632 8298 5684 8304
rect 5644 8265 5672 8298
rect 5630 8256 5686 8265
rect 5630 8191 5686 8200
rect 5736 8090 5764 9574
rect 5828 8906 5856 9646
rect 5908 9036 5960 9042
rect 5908 8978 5960 8984
rect 5816 8900 5868 8906
rect 5816 8842 5868 8848
rect 5814 8664 5870 8673
rect 5814 8599 5870 8608
rect 5828 8265 5856 8599
rect 5920 8430 5948 8978
rect 5908 8424 5960 8430
rect 5908 8366 5960 8372
rect 5814 8256 5870 8265
rect 6012 8242 6040 9646
rect 6564 9646 6684 9674
rect 6184 9580 6236 9586
rect 6564 9568 6592 9646
rect 6236 9540 6592 9568
rect 6644 9580 6696 9586
rect 6184 9522 6236 9528
rect 6644 9522 6696 9528
rect 6196 9353 6224 9522
rect 6460 9376 6512 9382
rect 6182 9344 6238 9353
rect 6460 9318 6512 9324
rect 6552 9376 6604 9382
rect 6552 9318 6604 9324
rect 6182 9279 6238 9288
rect 6472 9042 6500 9318
rect 6460 9036 6512 9042
rect 6460 8978 6512 8984
rect 6148 8732 6456 8741
rect 6148 8730 6154 8732
rect 6210 8730 6234 8732
rect 6290 8730 6314 8732
rect 6370 8730 6394 8732
rect 6450 8730 6456 8732
rect 6210 8678 6212 8730
rect 6392 8678 6394 8730
rect 6148 8676 6154 8678
rect 6210 8676 6234 8678
rect 6290 8676 6314 8678
rect 6370 8676 6394 8678
rect 6450 8676 6456 8678
rect 6148 8667 6456 8676
rect 6092 8628 6144 8634
rect 6564 8616 6592 9318
rect 6656 9042 6684 9522
rect 6644 9036 6696 9042
rect 6644 8978 6696 8984
rect 6642 8936 6698 8945
rect 6642 8871 6644 8880
rect 6696 8871 6698 8880
rect 6644 8842 6696 8848
rect 6748 8786 6776 11290
rect 6144 8588 6592 8616
rect 6656 8758 6776 8786
rect 6092 8570 6144 8576
rect 6092 8492 6144 8498
rect 6092 8434 6144 8440
rect 5814 8191 5870 8200
rect 5920 8214 6040 8242
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 5920 7970 5948 8214
rect 6104 7993 6132 8434
rect 6184 8356 6236 8362
rect 6184 8298 6236 8304
rect 5644 7942 5948 7970
rect 6090 7984 6146 7993
rect 6000 7948 6052 7954
rect 5644 7721 5672 7942
rect 6090 7919 6146 7928
rect 6000 7890 6052 7896
rect 5816 7880 5868 7886
rect 5736 7840 5816 7868
rect 5630 7712 5686 7721
rect 5630 7647 5686 7656
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 5644 6254 5672 6802
rect 5632 6248 5684 6254
rect 5632 6190 5684 6196
rect 5644 5574 5672 6190
rect 5736 6186 5764 7840
rect 5816 7822 5868 7828
rect 5816 7744 5868 7750
rect 5816 7686 5868 7692
rect 5908 7744 5960 7750
rect 5908 7686 5960 7692
rect 5828 6746 5856 7686
rect 5920 6934 5948 7686
rect 6012 7546 6040 7890
rect 6196 7886 6224 8298
rect 6656 8129 6684 8758
rect 6840 8650 6868 13126
rect 6920 12980 6972 12986
rect 6920 12922 6972 12928
rect 6932 12850 6960 12922
rect 6920 12844 6972 12850
rect 6920 12786 6972 12792
rect 7024 12102 7052 13382
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 7024 11762 7052 12038
rect 7012 11756 7064 11762
rect 7012 11698 7064 11704
rect 7012 11552 7064 11558
rect 7012 11494 7064 11500
rect 6920 11008 6972 11014
rect 6920 10950 6972 10956
rect 6932 10130 6960 10950
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 6932 9761 6960 9862
rect 6918 9752 6974 9761
rect 6918 9687 6974 9696
rect 6932 8838 6960 9687
rect 7024 9602 7052 11494
rect 7116 10810 7144 18090
rect 7288 17876 7340 17882
rect 7288 17818 7340 17824
rect 7196 17536 7248 17542
rect 7196 17478 7248 17484
rect 7208 16522 7236 17478
rect 7300 17134 7328 17818
rect 7288 17128 7340 17134
rect 7288 17070 7340 17076
rect 7300 16658 7328 17070
rect 7288 16652 7340 16658
rect 7288 16594 7340 16600
rect 7196 16516 7248 16522
rect 7196 16458 7248 16464
rect 7196 16108 7248 16114
rect 7196 16050 7248 16056
rect 7208 12374 7236 16050
rect 7300 15570 7328 16594
rect 7392 16454 7420 20742
rect 7472 19848 7524 19854
rect 7472 19790 7524 19796
rect 7484 19334 7512 19790
rect 7576 19530 7604 22200
rect 7838 20360 7894 20369
rect 7838 20295 7894 20304
rect 7748 20256 7800 20262
rect 7748 20198 7800 20204
rect 7760 20097 7788 20198
rect 7746 20088 7802 20097
rect 7746 20023 7802 20032
rect 7748 19712 7800 19718
rect 7748 19654 7800 19660
rect 7576 19502 7696 19530
rect 7484 19310 7604 19334
rect 7484 19306 7616 19310
rect 7564 19304 7616 19306
rect 7564 19246 7616 19252
rect 7576 18834 7604 19246
rect 7668 19174 7696 19502
rect 7760 19310 7788 19654
rect 7748 19304 7800 19310
rect 7748 19246 7800 19252
rect 7656 19168 7708 19174
rect 7656 19110 7708 19116
rect 7564 18828 7616 18834
rect 7564 18770 7616 18776
rect 7760 18766 7788 19246
rect 7748 18760 7800 18766
rect 7748 18702 7800 18708
rect 7656 18624 7708 18630
rect 7656 18566 7708 18572
rect 7748 18624 7800 18630
rect 7748 18566 7800 18572
rect 7852 18578 7880 20295
rect 7944 20058 7972 22200
rect 8312 20262 8340 22200
rect 8680 20466 8708 22200
rect 9048 21026 9076 22200
rect 9048 20998 9168 21026
rect 9140 20942 9168 20998
rect 9128 20936 9180 20942
rect 9128 20878 9180 20884
rect 9140 20466 9168 20878
rect 8668 20460 8720 20466
rect 8668 20402 8720 20408
rect 9128 20460 9180 20466
rect 9128 20402 9180 20408
rect 8392 20392 8444 20398
rect 8392 20334 8444 20340
rect 8300 20256 8352 20262
rect 8300 20198 8352 20204
rect 7932 20052 7984 20058
rect 7932 19994 7984 20000
rect 8312 19922 8340 20198
rect 8404 19922 8432 20334
rect 8300 19916 8352 19922
rect 8300 19858 8352 19864
rect 8392 19916 8444 19922
rect 8392 19858 8444 19864
rect 8680 19802 8708 20402
rect 9312 20256 9364 20262
rect 9312 20198 9364 20204
rect 8747 20156 9055 20165
rect 8747 20154 8753 20156
rect 8809 20154 8833 20156
rect 8889 20154 8913 20156
rect 8969 20154 8993 20156
rect 9049 20154 9055 20156
rect 8809 20102 8811 20154
rect 8991 20102 8993 20154
rect 8747 20100 8753 20102
rect 8809 20100 8833 20102
rect 8889 20100 8913 20102
rect 8969 20100 8993 20102
rect 9049 20100 9055 20102
rect 8747 20091 9055 20100
rect 8392 19780 8444 19786
rect 8680 19774 8892 19802
rect 8392 19722 8444 19728
rect 8300 19712 8352 19718
rect 8300 19654 8352 19660
rect 8206 19544 8262 19553
rect 8206 19479 8208 19488
rect 8260 19479 8262 19488
rect 8208 19450 8260 19456
rect 7932 19440 7984 19446
rect 7984 19388 8156 19394
rect 7932 19382 8156 19388
rect 7944 19366 8156 19382
rect 7932 19304 7984 19310
rect 7932 19246 7984 19252
rect 7944 18970 7972 19246
rect 7932 18964 7984 18970
rect 7932 18906 7984 18912
rect 8128 18902 8156 19366
rect 8206 19000 8262 19009
rect 8206 18935 8262 18944
rect 8116 18896 8168 18902
rect 8116 18838 8168 18844
rect 8220 18698 8248 18935
rect 8208 18692 8260 18698
rect 8208 18634 8260 18640
rect 8312 18630 8340 19654
rect 8404 19242 8432 19722
rect 8576 19712 8628 19718
rect 8576 19654 8628 19660
rect 8760 19712 8812 19718
rect 8760 19654 8812 19660
rect 8484 19372 8536 19378
rect 8484 19314 8536 19320
rect 8392 19236 8444 19242
rect 8392 19178 8444 19184
rect 8024 18624 8076 18630
rect 7668 18358 7696 18566
rect 7472 18352 7524 18358
rect 7472 18294 7524 18300
rect 7656 18352 7708 18358
rect 7656 18294 7708 18300
rect 7484 17354 7512 18294
rect 7760 18086 7788 18566
rect 7852 18550 7972 18578
rect 8024 18566 8076 18572
rect 8116 18624 8168 18630
rect 8116 18566 8168 18572
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 7840 18420 7892 18426
rect 7840 18362 7892 18368
rect 7748 18080 7800 18086
rect 7852 18057 7880 18362
rect 7748 18022 7800 18028
rect 7838 18048 7894 18057
rect 7838 17983 7894 17992
rect 7564 17536 7616 17542
rect 7562 17504 7564 17513
rect 7616 17504 7618 17513
rect 7562 17439 7618 17448
rect 7746 17504 7802 17513
rect 7746 17439 7802 17448
rect 7654 17368 7710 17377
rect 7484 17326 7604 17354
rect 7472 17196 7524 17202
rect 7472 17138 7524 17144
rect 7380 16448 7432 16454
rect 7380 16390 7432 16396
rect 7484 16153 7512 17138
rect 7470 16144 7526 16153
rect 7470 16079 7526 16088
rect 7472 15700 7524 15706
rect 7472 15642 7524 15648
rect 7288 15564 7340 15570
rect 7288 15506 7340 15512
rect 7380 15360 7432 15366
rect 7380 15302 7432 15308
rect 7288 13456 7340 13462
rect 7288 13398 7340 13404
rect 7196 12368 7248 12374
rect 7196 12310 7248 12316
rect 7300 12306 7328 13398
rect 7392 12434 7420 15302
rect 7484 12850 7512 15642
rect 7576 15162 7604 17326
rect 7654 17303 7710 17312
rect 7668 16697 7696 17303
rect 7760 17241 7788 17439
rect 7944 17320 7972 18550
rect 8036 17338 8064 18566
rect 8128 17882 8156 18566
rect 8300 18420 8352 18426
rect 8220 18380 8300 18408
rect 8116 17876 8168 17882
rect 8116 17818 8168 17824
rect 8116 17740 8168 17746
rect 8116 17682 8168 17688
rect 7852 17292 7972 17320
rect 8024 17332 8076 17338
rect 7746 17232 7802 17241
rect 7746 17167 7802 17176
rect 7746 17096 7802 17105
rect 7746 17031 7802 17040
rect 7760 16794 7788 17031
rect 7748 16788 7800 16794
rect 7748 16730 7800 16736
rect 7654 16688 7710 16697
rect 7654 16623 7710 16632
rect 7748 16584 7800 16590
rect 7746 16552 7748 16561
rect 7800 16552 7802 16561
rect 7746 16487 7802 16496
rect 7852 16114 7880 17292
rect 8024 17274 8076 17280
rect 7932 17196 7984 17202
rect 7932 17138 7984 17144
rect 7944 16697 7972 17138
rect 7930 16688 7986 16697
rect 8128 16674 8156 17682
rect 8220 17542 8248 18380
rect 8300 18362 8352 18368
rect 8404 18306 8432 19178
rect 8496 18970 8524 19314
rect 8484 18964 8536 18970
rect 8484 18906 8536 18912
rect 8484 18624 8536 18630
rect 8484 18566 8536 18572
rect 8312 18278 8432 18306
rect 8312 18222 8340 18278
rect 8300 18216 8352 18222
rect 8300 18158 8352 18164
rect 8392 18148 8444 18154
rect 8392 18090 8444 18096
rect 8404 17814 8432 18090
rect 8496 18057 8524 18566
rect 8588 18222 8616 19654
rect 8668 19440 8720 19446
rect 8668 19382 8720 19388
rect 8680 18970 8708 19382
rect 8772 19310 8800 19654
rect 8760 19304 8812 19310
rect 8760 19246 8812 19252
rect 8864 19242 8892 19774
rect 9128 19372 9180 19378
rect 9128 19314 9180 19320
rect 8852 19236 8904 19242
rect 8852 19178 8904 19184
rect 8747 19068 9055 19077
rect 8747 19066 8753 19068
rect 8809 19066 8833 19068
rect 8889 19066 8913 19068
rect 8969 19066 8993 19068
rect 9049 19066 9055 19068
rect 8809 19014 8811 19066
rect 8991 19014 8993 19066
rect 8747 19012 8753 19014
rect 8809 19012 8833 19014
rect 8889 19012 8913 19014
rect 8969 19012 8993 19014
rect 9049 19012 9055 19014
rect 8747 19003 9055 19012
rect 8668 18964 8720 18970
rect 8668 18906 8720 18912
rect 8760 18624 8812 18630
rect 8760 18566 8812 18572
rect 8772 18358 8800 18566
rect 8760 18352 8812 18358
rect 8760 18294 8812 18300
rect 8576 18216 8628 18222
rect 8760 18216 8812 18222
rect 8576 18158 8628 18164
rect 8680 18176 8760 18204
rect 8482 18048 8538 18057
rect 8482 17983 8538 17992
rect 8482 17912 8538 17921
rect 8482 17847 8538 17856
rect 8392 17808 8444 17814
rect 8392 17750 8444 17756
rect 8496 17542 8524 17847
rect 8588 17746 8616 18158
rect 8576 17740 8628 17746
rect 8576 17682 8628 17688
rect 8208 17536 8260 17542
rect 8208 17478 8260 17484
rect 8484 17536 8536 17542
rect 8484 17478 8536 17484
rect 8208 17332 8260 17338
rect 8208 17274 8260 17280
rect 8220 16969 8248 17274
rect 8680 17270 8708 18176
rect 8760 18158 8812 18164
rect 8747 17980 9055 17989
rect 8747 17978 8753 17980
rect 8809 17978 8833 17980
rect 8889 17978 8913 17980
rect 8969 17978 8993 17980
rect 9049 17978 9055 17980
rect 8809 17926 8811 17978
rect 8991 17926 8993 17978
rect 8747 17924 8753 17926
rect 8809 17924 8833 17926
rect 8889 17924 8913 17926
rect 8969 17924 8993 17926
rect 9049 17924 9055 17926
rect 8747 17915 9055 17924
rect 8850 17776 8906 17785
rect 9034 17776 9090 17785
rect 8850 17711 8906 17720
rect 8944 17740 8996 17746
rect 8864 17542 8892 17711
rect 9034 17711 9090 17720
rect 8944 17682 8996 17688
rect 8852 17536 8904 17542
rect 8852 17478 8904 17484
rect 8864 17338 8892 17478
rect 8852 17332 8904 17338
rect 8852 17274 8904 17280
rect 8484 17264 8536 17270
rect 8668 17264 8720 17270
rect 8484 17206 8536 17212
rect 8588 17224 8668 17252
rect 8300 17128 8352 17134
rect 8300 17070 8352 17076
rect 8206 16960 8262 16969
rect 8206 16895 8262 16904
rect 7930 16623 7932 16632
rect 7984 16623 7986 16632
rect 8036 16646 8156 16674
rect 7932 16594 7984 16600
rect 7840 16108 7892 16114
rect 7840 16050 7892 16056
rect 7932 15632 7984 15638
rect 7654 15600 7710 15609
rect 7654 15535 7710 15544
rect 7838 15600 7894 15609
rect 7932 15574 7984 15580
rect 7838 15535 7840 15544
rect 7668 15337 7696 15535
rect 7892 15535 7894 15544
rect 7840 15506 7892 15512
rect 7654 15328 7710 15337
rect 7654 15263 7710 15272
rect 7564 15156 7616 15162
rect 7564 15098 7616 15104
rect 7656 15020 7708 15026
rect 7656 14962 7708 14968
rect 7564 14816 7616 14822
rect 7564 14758 7616 14764
rect 7472 12844 7524 12850
rect 7472 12786 7524 12792
rect 7576 12646 7604 14758
rect 7668 14618 7696 14962
rect 7656 14612 7708 14618
rect 7656 14554 7708 14560
rect 7748 14272 7800 14278
rect 7748 14214 7800 14220
rect 7760 13870 7788 14214
rect 7656 13864 7708 13870
rect 7656 13806 7708 13812
rect 7748 13864 7800 13870
rect 7748 13806 7800 13812
rect 7668 13530 7696 13806
rect 7656 13524 7708 13530
rect 7656 13466 7708 13472
rect 7760 13394 7788 13806
rect 7748 13388 7800 13394
rect 7748 13330 7800 13336
rect 7944 13274 7972 15574
rect 8036 14278 8064 16646
rect 8116 16584 8168 16590
rect 8312 16574 8340 17070
rect 8392 17060 8444 17066
rect 8392 17002 8444 17008
rect 8404 16726 8432 17002
rect 8392 16720 8444 16726
rect 8392 16662 8444 16668
rect 8116 16526 8168 16532
rect 8220 16546 8340 16574
rect 8390 16552 8446 16561
rect 8128 16114 8156 16526
rect 8116 16108 8168 16114
rect 8116 16050 8168 16056
rect 8116 15564 8168 15570
rect 8116 15506 8168 15512
rect 8024 14272 8076 14278
rect 8024 14214 8076 14220
rect 7668 13246 7972 13274
rect 7564 12640 7616 12646
rect 7564 12582 7616 12588
rect 7392 12406 7512 12434
rect 7288 12300 7340 12306
rect 7288 12242 7340 12248
rect 7484 12186 7512 12406
rect 7564 12368 7616 12374
rect 7564 12310 7616 12316
rect 7300 12158 7512 12186
rect 7196 11688 7248 11694
rect 7196 11630 7248 11636
rect 7208 11218 7236 11630
rect 7196 11212 7248 11218
rect 7196 11154 7248 11160
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 7116 10198 7144 10746
rect 7300 10441 7328 12158
rect 7380 12096 7432 12102
rect 7378 12064 7380 12073
rect 7472 12096 7524 12102
rect 7432 12064 7434 12073
rect 7472 12038 7524 12044
rect 7378 11999 7434 12008
rect 7392 11898 7420 11999
rect 7380 11892 7432 11898
rect 7380 11834 7432 11840
rect 7392 11801 7420 11834
rect 7378 11792 7434 11801
rect 7378 11727 7434 11736
rect 7286 10432 7342 10441
rect 7286 10367 7342 10376
rect 7484 10282 7512 12038
rect 7208 10254 7512 10282
rect 7104 10192 7156 10198
rect 7104 10134 7156 10140
rect 7024 9574 7144 9602
rect 7012 9512 7064 9518
rect 7012 9454 7064 9460
rect 7024 9178 7052 9454
rect 7012 9172 7064 9178
rect 7012 9114 7064 9120
rect 7012 8968 7064 8974
rect 7012 8910 7064 8916
rect 6920 8832 6972 8838
rect 7024 8809 7052 8910
rect 6920 8774 6972 8780
rect 7010 8800 7066 8809
rect 6748 8622 6868 8650
rect 6642 8120 6698 8129
rect 6642 8055 6698 8064
rect 6276 8016 6328 8022
rect 6274 7984 6276 7993
rect 6328 7984 6330 7993
rect 6274 7919 6330 7928
rect 6184 7880 6236 7886
rect 6184 7822 6236 7828
rect 6552 7812 6604 7818
rect 6552 7754 6604 7760
rect 6148 7644 6456 7653
rect 6148 7642 6154 7644
rect 6210 7642 6234 7644
rect 6290 7642 6314 7644
rect 6370 7642 6394 7644
rect 6450 7642 6456 7644
rect 6210 7590 6212 7642
rect 6392 7590 6394 7642
rect 6148 7588 6154 7590
rect 6210 7588 6234 7590
rect 6290 7588 6314 7590
rect 6370 7588 6394 7590
rect 6450 7588 6456 7590
rect 6148 7579 6456 7588
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 5908 6928 5960 6934
rect 5908 6870 5960 6876
rect 5828 6718 5948 6746
rect 5816 6656 5868 6662
rect 5816 6598 5868 6604
rect 5724 6180 5776 6186
rect 5724 6122 5776 6128
rect 5724 5704 5776 5710
rect 5722 5672 5724 5681
rect 5776 5672 5778 5681
rect 5722 5607 5778 5616
rect 5632 5568 5684 5574
rect 5632 5510 5684 5516
rect 5724 5568 5776 5574
rect 5724 5510 5776 5516
rect 5644 5409 5672 5510
rect 5460 5358 5580 5386
rect 5630 5400 5686 5409
rect 5356 4752 5408 4758
rect 5356 4694 5408 4700
rect 5264 4208 5316 4214
rect 5264 4150 5316 4156
rect 5356 4208 5408 4214
rect 5356 4150 5408 4156
rect 5368 4026 5396 4150
rect 5276 3998 5396 4026
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 5276 3398 5304 3998
rect 5460 3890 5488 5358
rect 5736 5370 5764 5510
rect 5630 5335 5686 5344
rect 5724 5364 5776 5370
rect 5540 5296 5592 5302
rect 5540 5238 5592 5244
rect 5552 4010 5580 5238
rect 5644 4826 5672 5335
rect 5724 5306 5776 5312
rect 5828 5137 5856 6598
rect 5920 6118 5948 6718
rect 5908 6112 5960 6118
rect 5908 6054 5960 6060
rect 5906 5944 5962 5953
rect 5906 5879 5908 5888
rect 5960 5879 5962 5888
rect 5908 5850 5960 5856
rect 5906 5536 5962 5545
rect 5906 5471 5962 5480
rect 5920 5370 5948 5471
rect 5908 5364 5960 5370
rect 5908 5306 5960 5312
rect 5814 5128 5870 5137
rect 5814 5063 5870 5072
rect 5724 5024 5776 5030
rect 5724 4966 5776 4972
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 5736 4690 5764 4966
rect 5816 4820 5868 4826
rect 5816 4762 5868 4768
rect 5828 4690 5856 4762
rect 5724 4684 5776 4690
rect 5724 4626 5776 4632
rect 5816 4684 5868 4690
rect 5816 4626 5868 4632
rect 5630 4584 5686 4593
rect 5630 4519 5686 4528
rect 5814 4584 5870 4593
rect 5814 4519 5870 4528
rect 5908 4548 5960 4554
rect 5644 4486 5672 4519
rect 5632 4480 5684 4486
rect 5632 4422 5684 4428
rect 5828 4282 5856 4519
rect 5908 4490 5960 4496
rect 5920 4457 5948 4490
rect 5906 4448 5962 4457
rect 5906 4383 5962 4392
rect 5816 4276 5868 4282
rect 5816 4218 5868 4224
rect 6012 4162 6040 7482
rect 6458 6896 6514 6905
rect 6458 6831 6514 6840
rect 6472 6798 6500 6831
rect 6460 6792 6512 6798
rect 6460 6734 6512 6740
rect 6564 6662 6592 7754
rect 6644 7744 6696 7750
rect 6642 7712 6644 7721
rect 6696 7712 6698 7721
rect 6642 7647 6698 7656
rect 6656 7313 6684 7647
rect 6642 7304 6698 7313
rect 6642 7239 6698 7248
rect 6644 7200 6696 7206
rect 6644 7142 6696 7148
rect 6656 6905 6684 7142
rect 6642 6896 6698 6905
rect 6642 6831 6698 6840
rect 6552 6656 6604 6662
rect 6552 6598 6604 6604
rect 6644 6656 6696 6662
rect 6644 6598 6696 6604
rect 6148 6556 6456 6565
rect 6148 6554 6154 6556
rect 6210 6554 6234 6556
rect 6290 6554 6314 6556
rect 6370 6554 6394 6556
rect 6450 6554 6456 6556
rect 6210 6502 6212 6554
rect 6392 6502 6394 6554
rect 6148 6500 6154 6502
rect 6210 6500 6234 6502
rect 6290 6500 6314 6502
rect 6370 6500 6394 6502
rect 6450 6500 6456 6502
rect 6148 6491 6456 6500
rect 6564 6390 6592 6598
rect 6552 6384 6604 6390
rect 6656 6361 6684 6598
rect 6552 6326 6604 6332
rect 6642 6352 6698 6361
rect 6184 6316 6236 6322
rect 6184 6258 6236 6264
rect 6368 6316 6420 6322
rect 6642 6287 6698 6296
rect 6368 6258 6420 6264
rect 6196 5914 6224 6258
rect 6380 6225 6408 6258
rect 6644 6248 6696 6254
rect 6366 6216 6422 6225
rect 6644 6190 6696 6196
rect 6366 6151 6422 6160
rect 6276 6112 6328 6118
rect 6276 6054 6328 6060
rect 6184 5908 6236 5914
rect 6184 5850 6236 5856
rect 6288 5846 6316 6054
rect 6552 5908 6604 5914
rect 6552 5850 6604 5856
rect 6276 5840 6328 5846
rect 6276 5782 6328 5788
rect 6368 5840 6420 5846
rect 6368 5782 6420 5788
rect 6458 5808 6514 5817
rect 6288 5681 6316 5782
rect 6274 5672 6330 5681
rect 6274 5607 6330 5616
rect 6380 5574 6408 5782
rect 6458 5743 6514 5752
rect 6472 5574 6500 5743
rect 6368 5568 6420 5574
rect 6368 5510 6420 5516
rect 6460 5568 6512 5574
rect 6460 5510 6512 5516
rect 6148 5468 6456 5477
rect 6148 5466 6154 5468
rect 6210 5466 6234 5468
rect 6290 5466 6314 5468
rect 6370 5466 6394 5468
rect 6450 5466 6456 5468
rect 6210 5414 6212 5466
rect 6392 5414 6394 5466
rect 6148 5412 6154 5414
rect 6210 5412 6234 5414
rect 6290 5412 6314 5414
rect 6370 5412 6394 5414
rect 6450 5412 6456 5414
rect 6148 5403 6456 5412
rect 6182 5264 6238 5273
rect 6182 5199 6238 5208
rect 6276 5228 6328 5234
rect 6196 4554 6224 5199
rect 6276 5170 6328 5176
rect 6288 5001 6316 5170
rect 6368 5024 6420 5030
rect 6274 4992 6330 5001
rect 6368 4966 6420 4972
rect 6274 4927 6330 4936
rect 6274 4856 6330 4865
rect 6274 4791 6276 4800
rect 6328 4791 6330 4800
rect 6276 4762 6328 4768
rect 6380 4622 6408 4966
rect 6368 4616 6420 4622
rect 6368 4558 6420 4564
rect 6184 4548 6236 4554
rect 6184 4490 6236 4496
rect 6148 4380 6456 4389
rect 6148 4378 6154 4380
rect 6210 4378 6234 4380
rect 6290 4378 6314 4380
rect 6370 4378 6394 4380
rect 6450 4378 6456 4380
rect 6210 4326 6212 4378
rect 6392 4326 6394 4378
rect 6148 4324 6154 4326
rect 6210 4324 6234 4326
rect 6290 4324 6314 4326
rect 6370 4324 6394 4326
rect 6450 4324 6456 4326
rect 6148 4315 6456 4324
rect 6092 4276 6144 4282
rect 6092 4218 6144 4224
rect 5644 4134 6040 4162
rect 5540 4004 5592 4010
rect 5540 3946 5592 3952
rect 5460 3862 5580 3890
rect 5356 3460 5408 3466
rect 5356 3402 5408 3408
rect 5448 3460 5500 3466
rect 5448 3402 5500 3408
rect 5264 3392 5316 3398
rect 5368 3369 5396 3402
rect 5264 3334 5316 3340
rect 5354 3360 5410 3369
rect 5354 3295 5410 3304
rect 5460 3126 5488 3402
rect 5448 3120 5500 3126
rect 5552 3097 5580 3862
rect 5448 3062 5500 3068
rect 5538 3088 5594 3097
rect 5538 3023 5594 3032
rect 5540 2848 5592 2854
rect 5540 2790 5592 2796
rect 5446 2680 5502 2689
rect 5446 2615 5502 2624
rect 5264 2508 5316 2514
rect 5264 2450 5316 2456
rect 5276 2038 5304 2450
rect 5264 2032 5316 2038
rect 5264 1974 5316 1980
rect 5276 1442 5304 1974
rect 5460 1970 5488 2615
rect 5552 2582 5580 2790
rect 5644 2650 5672 4134
rect 6000 4072 6052 4078
rect 5920 4032 6000 4060
rect 5920 3738 5948 4032
rect 6000 4014 6052 4020
rect 5998 3904 6054 3913
rect 5998 3839 6054 3848
rect 5908 3732 5960 3738
rect 5908 3674 5960 3680
rect 6012 3670 6040 3839
rect 6000 3664 6052 3670
rect 6000 3606 6052 3612
rect 6104 3482 6132 4218
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 6380 4049 6408 4082
rect 6366 4040 6422 4049
rect 6366 3975 6422 3984
rect 6564 3942 6592 5850
rect 6656 5778 6684 6190
rect 6644 5772 6696 5778
rect 6644 5714 6696 5720
rect 6656 5166 6684 5714
rect 6644 5160 6696 5166
rect 6644 5102 6696 5108
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 6656 4010 6684 4558
rect 6748 4146 6776 8622
rect 6828 8560 6880 8566
rect 6932 8537 6960 8774
rect 7010 8735 7066 8744
rect 7024 8634 7052 8735
rect 7012 8628 7064 8634
rect 7012 8570 7064 8576
rect 6828 8502 6880 8508
rect 6918 8528 6974 8537
rect 6840 7954 6868 8502
rect 6918 8463 6974 8472
rect 7012 8288 7064 8294
rect 6932 8248 7012 8276
rect 6828 7948 6880 7954
rect 6828 7890 6880 7896
rect 6840 7546 6868 7890
rect 6932 7818 6960 8248
rect 7012 8230 7064 8236
rect 7010 8120 7066 8129
rect 7010 8055 7066 8064
rect 6920 7812 6972 7818
rect 6920 7754 6972 7760
rect 6932 7546 6960 7754
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6920 7540 6972 7546
rect 6920 7482 6972 7488
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 6828 5636 6880 5642
rect 6828 5578 6880 5584
rect 6840 5137 6868 5578
rect 6932 5574 6960 7346
rect 7024 6866 7052 8055
rect 7116 7342 7144 9574
rect 7104 7336 7156 7342
rect 7104 7278 7156 7284
rect 7104 7200 7156 7206
rect 7104 7142 7156 7148
rect 7012 6860 7064 6866
rect 7012 6802 7064 6808
rect 7010 6488 7066 6497
rect 7010 6423 7066 6432
rect 7024 6322 7052 6423
rect 7012 6316 7064 6322
rect 7012 6258 7064 6264
rect 6920 5568 6972 5574
rect 6920 5510 6972 5516
rect 6826 5128 6882 5137
rect 6826 5063 6882 5072
rect 6828 4684 6880 4690
rect 6828 4626 6880 4632
rect 6736 4140 6788 4146
rect 6736 4082 6788 4088
rect 6644 4004 6696 4010
rect 6644 3946 6696 3952
rect 6552 3936 6604 3942
rect 6552 3878 6604 3884
rect 6550 3768 6606 3777
rect 6550 3703 6606 3712
rect 6276 3596 6328 3602
rect 6276 3538 6328 3544
rect 5736 3454 6132 3482
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 5540 2576 5592 2582
rect 5540 2518 5592 2524
rect 5538 2408 5594 2417
rect 5538 2343 5594 2352
rect 5552 2106 5580 2343
rect 5540 2100 5592 2106
rect 5540 2042 5592 2048
rect 5448 1964 5500 1970
rect 5448 1906 5500 1912
rect 5538 1864 5594 1873
rect 5538 1799 5594 1808
rect 5184 1414 5304 1442
rect 5080 1216 5132 1222
rect 5080 1158 5132 1164
rect 5184 800 5212 1414
rect 5552 800 5580 1799
rect 5736 1154 5764 3454
rect 6288 3398 6316 3538
rect 5908 3392 5960 3398
rect 5908 3334 5960 3340
rect 6000 3392 6052 3398
rect 6000 3334 6052 3340
rect 6276 3392 6328 3398
rect 6276 3334 6328 3340
rect 5920 3194 5948 3334
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 5908 3188 5960 3194
rect 5908 3130 5960 3136
rect 5828 2922 5856 3130
rect 5816 2916 5868 2922
rect 5816 2858 5868 2864
rect 5908 2576 5960 2582
rect 5908 2518 5960 2524
rect 5920 2417 5948 2518
rect 6012 2446 6040 3334
rect 6148 3292 6456 3301
rect 6148 3290 6154 3292
rect 6210 3290 6234 3292
rect 6290 3290 6314 3292
rect 6370 3290 6394 3292
rect 6450 3290 6456 3292
rect 6210 3238 6212 3290
rect 6392 3238 6394 3290
rect 6148 3236 6154 3238
rect 6210 3236 6234 3238
rect 6290 3236 6314 3238
rect 6370 3236 6394 3238
rect 6450 3236 6456 3238
rect 6148 3227 6456 3236
rect 6564 3194 6592 3703
rect 6656 3466 6684 3946
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6644 3460 6696 3466
rect 6644 3402 6696 3408
rect 6552 3188 6604 3194
rect 6552 3130 6604 3136
rect 6656 2938 6684 3402
rect 6748 3058 6776 3878
rect 6840 3670 6868 4626
rect 6932 4282 6960 5510
rect 7010 5400 7066 5409
rect 7010 5335 7066 5344
rect 7024 5234 7052 5335
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 7012 5092 7064 5098
rect 7012 5034 7064 5040
rect 6920 4276 6972 4282
rect 6920 4218 6972 4224
rect 7024 4078 7052 5034
rect 7116 4282 7144 7142
rect 7104 4276 7156 4282
rect 7104 4218 7156 4224
rect 7208 4214 7236 10254
rect 7288 10192 7340 10198
rect 7576 10180 7604 12310
rect 7288 10134 7340 10140
rect 7392 10152 7604 10180
rect 7300 9722 7328 10134
rect 7288 9716 7340 9722
rect 7288 9658 7340 9664
rect 7392 8922 7420 10152
rect 7472 9920 7524 9926
rect 7472 9862 7524 9868
rect 7564 9920 7616 9926
rect 7564 9862 7616 9868
rect 7484 9722 7512 9862
rect 7472 9716 7524 9722
rect 7472 9658 7524 9664
rect 7576 9450 7604 9862
rect 7668 9761 7696 13246
rect 8036 13190 8064 14214
rect 7840 13184 7892 13190
rect 7840 13126 7892 13132
rect 8024 13184 8076 13190
rect 8024 13126 8076 13132
rect 7852 12986 7880 13126
rect 7840 12980 7892 12986
rect 7840 12922 7892 12928
rect 7840 12368 7892 12374
rect 7840 12310 7892 12316
rect 7748 12300 7800 12306
rect 7748 12242 7800 12248
rect 7654 9752 7710 9761
rect 7654 9687 7710 9696
rect 7668 9450 7696 9687
rect 7564 9444 7616 9450
rect 7564 9386 7616 9392
rect 7656 9444 7708 9450
rect 7656 9386 7708 9392
rect 7470 9208 7526 9217
rect 7470 9143 7526 9152
rect 7300 8894 7420 8922
rect 7300 6662 7328 8894
rect 7380 8832 7432 8838
rect 7380 8774 7432 8780
rect 7392 8090 7420 8774
rect 7484 8566 7512 9143
rect 7564 9036 7616 9042
rect 7564 8978 7616 8984
rect 7576 8634 7604 8978
rect 7656 8832 7708 8838
rect 7656 8774 7708 8780
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 7472 8560 7524 8566
rect 7472 8502 7524 8508
rect 7562 8528 7618 8537
rect 7562 8463 7564 8472
rect 7616 8463 7618 8472
rect 7564 8434 7616 8440
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7380 7336 7432 7342
rect 7380 7278 7432 7284
rect 7470 7304 7526 7313
rect 7288 6656 7340 6662
rect 7288 6598 7340 6604
rect 7300 6458 7328 6598
rect 7288 6452 7340 6458
rect 7288 6394 7340 6400
rect 7392 6338 7420 7278
rect 7470 7239 7526 7248
rect 7300 6310 7420 6338
rect 7300 5846 7328 6310
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 7288 5840 7340 5846
rect 7288 5782 7340 5788
rect 7300 5545 7328 5782
rect 7392 5778 7420 6190
rect 7380 5772 7432 5778
rect 7380 5714 7432 5720
rect 7286 5536 7342 5545
rect 7286 5471 7342 5480
rect 7286 5400 7342 5409
rect 7286 5335 7342 5344
rect 7300 5302 7328 5335
rect 7288 5296 7340 5302
rect 7288 5238 7340 5244
rect 7288 5024 7340 5030
rect 7288 4966 7340 4972
rect 7196 4208 7248 4214
rect 7196 4150 7248 4156
rect 7012 4072 7064 4078
rect 7012 4014 7064 4020
rect 6828 3664 6880 3670
rect 6828 3606 6880 3612
rect 6918 3360 6974 3369
rect 6918 3295 6974 3304
rect 6826 3224 6882 3233
rect 6826 3159 6828 3168
rect 6880 3159 6882 3168
rect 6828 3130 6880 3136
rect 6932 3058 6960 3295
rect 7024 3194 7052 4014
rect 7102 3904 7158 3913
rect 7102 3839 7158 3848
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 7010 3088 7066 3097
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 6920 3052 6972 3058
rect 7010 3023 7066 3032
rect 6920 2994 6972 3000
rect 6656 2910 6776 2938
rect 6550 2816 6606 2825
rect 6550 2751 6606 2760
rect 6000 2440 6052 2446
rect 5906 2408 5962 2417
rect 6000 2382 6052 2388
rect 5906 2343 5962 2352
rect 5816 2304 5868 2310
rect 5816 2246 5868 2252
rect 5906 2272 5962 2281
rect 5828 1970 5856 2246
rect 5906 2207 5962 2216
rect 5816 1964 5868 1970
rect 5816 1906 5868 1912
rect 5724 1148 5776 1154
rect 5724 1090 5776 1096
rect 5920 800 5948 2207
rect 6148 2204 6456 2213
rect 6148 2202 6154 2204
rect 6210 2202 6234 2204
rect 6290 2202 6314 2204
rect 6370 2202 6394 2204
rect 6450 2202 6456 2204
rect 6210 2150 6212 2202
rect 6392 2150 6394 2202
rect 6148 2148 6154 2150
rect 6210 2148 6234 2150
rect 6290 2148 6314 2150
rect 6370 2148 6394 2150
rect 6450 2148 6456 2150
rect 6148 2139 6456 2148
rect 6288 870 6408 898
rect 6288 800 6316 870
rect 4540 734 4660 762
rect 4632 105 4660 734
rect 4618 96 4674 105
rect 4618 31 4674 40
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5906 0 5962 800
rect 6274 0 6330 800
rect 6380 762 6408 870
rect 6564 762 6592 2751
rect 6748 2378 6776 2910
rect 6826 2816 6882 2825
rect 6826 2751 6882 2760
rect 6840 2650 6868 2751
rect 6828 2644 6880 2650
rect 6828 2586 6880 2592
rect 6644 2372 6696 2378
rect 6644 2314 6696 2320
rect 6736 2372 6788 2378
rect 6736 2314 6788 2320
rect 6656 1902 6684 2314
rect 6644 1896 6696 1902
rect 6644 1838 6696 1844
rect 6734 1864 6790 1873
rect 6734 1799 6790 1808
rect 6748 1766 6776 1799
rect 6736 1760 6788 1766
rect 6736 1702 6788 1708
rect 6748 1442 6776 1702
rect 6656 1414 6776 1442
rect 6656 800 6684 1414
rect 7024 800 7052 3023
rect 7116 2514 7144 3839
rect 7208 2854 7236 4150
rect 7300 2990 7328 4966
rect 7392 4214 7420 5714
rect 7484 5710 7512 7239
rect 7668 7206 7696 8774
rect 7760 8498 7788 12242
rect 7852 12102 7880 12310
rect 7932 12300 7984 12306
rect 7932 12242 7984 12248
rect 7840 12096 7892 12102
rect 7840 12038 7892 12044
rect 7840 11892 7892 11898
rect 7840 11834 7892 11840
rect 7852 11626 7880 11834
rect 7840 11620 7892 11626
rect 7840 11562 7892 11568
rect 7944 11150 7972 12242
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 8036 11898 8064 12038
rect 8024 11892 8076 11898
rect 8024 11834 8076 11840
rect 8024 11688 8076 11694
rect 8024 11630 8076 11636
rect 8036 11218 8064 11630
rect 8024 11212 8076 11218
rect 8024 11154 8076 11160
rect 7932 11144 7984 11150
rect 7838 11112 7894 11121
rect 7932 11086 7984 11092
rect 7838 11047 7840 11056
rect 7892 11047 7894 11056
rect 7840 11018 7892 11024
rect 7932 11008 7984 11014
rect 7932 10950 7984 10956
rect 7840 10736 7892 10742
rect 7944 10724 7972 10950
rect 7892 10696 7972 10724
rect 7840 10678 7892 10684
rect 7852 10606 7880 10678
rect 8036 10674 8064 11154
rect 8024 10668 8076 10674
rect 8024 10610 8076 10616
rect 7840 10600 7892 10606
rect 7840 10542 7892 10548
rect 7840 10464 7892 10470
rect 7840 10406 7892 10412
rect 8022 10432 8078 10441
rect 7852 10130 7880 10406
rect 8022 10367 8078 10376
rect 7840 10124 7892 10130
rect 7840 10066 7892 10072
rect 7840 9988 7892 9994
rect 7840 9930 7892 9936
rect 7852 9761 7880 9930
rect 8036 9874 8064 10367
rect 8128 10169 8156 15506
rect 8220 15366 8248 16546
rect 8390 16487 8446 16496
rect 8300 15904 8352 15910
rect 8300 15846 8352 15852
rect 8208 15360 8260 15366
rect 8208 15302 8260 15308
rect 8312 15026 8340 15846
rect 8404 15434 8432 16487
rect 8496 15502 8524 17206
rect 8588 15638 8616 17224
rect 8864 17241 8892 17274
rect 8668 17206 8720 17212
rect 8850 17232 8906 17241
rect 8850 17167 8906 17176
rect 8956 17134 8984 17682
rect 9048 17513 9076 17711
rect 9034 17504 9090 17513
rect 9034 17439 9090 17448
rect 9036 17264 9088 17270
rect 9036 17206 9088 17212
rect 8944 17128 8996 17134
rect 8944 17070 8996 17076
rect 9048 17066 9076 17206
rect 9036 17060 9088 17066
rect 9036 17002 9088 17008
rect 8747 16892 9055 16901
rect 8747 16890 8753 16892
rect 8809 16890 8833 16892
rect 8889 16890 8913 16892
rect 8969 16890 8993 16892
rect 9049 16890 9055 16892
rect 8809 16838 8811 16890
rect 8991 16838 8993 16890
rect 8747 16836 8753 16838
rect 8809 16836 8833 16838
rect 8889 16836 8913 16838
rect 8969 16836 8993 16838
rect 9049 16836 9055 16838
rect 8747 16827 9055 16836
rect 9140 16776 9168 19314
rect 9324 19258 9352 20198
rect 8864 16748 9168 16776
rect 9232 19230 9352 19258
rect 8668 16720 8720 16726
rect 8668 16662 8720 16668
rect 8758 16688 8814 16697
rect 8576 15632 8628 15638
rect 8576 15574 8628 15580
rect 8484 15496 8536 15502
rect 8680 15473 8708 16662
rect 8758 16623 8814 16632
rect 8772 16114 8800 16623
rect 8864 16454 8892 16748
rect 9126 16688 9182 16697
rect 9126 16623 9182 16632
rect 8852 16448 8904 16454
rect 8852 16390 8904 16396
rect 8944 16448 8996 16454
rect 8944 16390 8996 16396
rect 8760 16108 8812 16114
rect 8760 16050 8812 16056
rect 8852 15904 8904 15910
rect 8956 15892 8984 16390
rect 8904 15864 8984 15892
rect 8852 15846 8904 15852
rect 8747 15804 9055 15813
rect 8747 15802 8753 15804
rect 8809 15802 8833 15804
rect 8889 15802 8913 15804
rect 8969 15802 8993 15804
rect 9049 15802 9055 15804
rect 8809 15750 8811 15802
rect 8991 15750 8993 15802
rect 8747 15748 8753 15750
rect 8809 15748 8833 15750
rect 8889 15748 8913 15750
rect 8969 15748 8993 15750
rect 9049 15748 9055 15750
rect 8747 15739 9055 15748
rect 9140 15586 9168 16623
rect 9048 15558 9168 15586
rect 8484 15438 8536 15444
rect 8666 15464 8722 15473
rect 8392 15428 8444 15434
rect 8666 15399 8722 15408
rect 8392 15370 8444 15376
rect 8576 15360 8628 15366
rect 8390 15328 8446 15337
rect 8390 15263 8446 15272
rect 8574 15328 8576 15337
rect 8628 15328 8630 15337
rect 8574 15263 8630 15272
rect 8404 15162 8432 15263
rect 8392 15156 8444 15162
rect 8392 15098 8444 15104
rect 8300 15020 8352 15026
rect 8300 14962 8352 14968
rect 8312 14498 8340 14962
rect 9048 14890 9076 15558
rect 9232 15162 9260 19230
rect 9416 18714 9444 22200
rect 9784 20602 9812 22200
rect 9772 20596 9824 20602
rect 10152 20584 10180 22200
rect 10152 20556 10272 20584
rect 9772 20538 9824 20544
rect 9496 20392 9548 20398
rect 9496 20334 9548 20340
rect 9508 19417 9536 20334
rect 9494 19408 9550 19417
rect 9494 19343 9550 19352
rect 9588 19168 9640 19174
rect 9588 19110 9640 19116
rect 9680 19168 9732 19174
rect 9680 19110 9732 19116
rect 9600 18834 9628 19110
rect 9588 18828 9640 18834
rect 9588 18770 9640 18776
rect 9416 18686 9536 18714
rect 9312 18624 9364 18630
rect 9312 18566 9364 18572
rect 9404 18624 9456 18630
rect 9404 18566 9456 18572
rect 9324 18426 9352 18566
rect 9312 18420 9364 18426
rect 9312 18362 9364 18368
rect 9312 18080 9364 18086
rect 9312 18022 9364 18028
rect 9324 17762 9352 18022
rect 9416 17882 9444 18566
rect 9508 18290 9536 18686
rect 9692 18442 9720 19110
rect 9784 18766 9812 20538
rect 10140 20460 10192 20466
rect 10140 20402 10192 20408
rect 9772 18760 9824 18766
rect 9772 18702 9824 18708
rect 9864 18692 9916 18698
rect 9864 18634 9916 18640
rect 9772 18624 9824 18630
rect 9772 18566 9824 18572
rect 9784 18465 9812 18566
rect 9600 18414 9720 18442
rect 9770 18456 9826 18465
rect 9496 18284 9548 18290
rect 9496 18226 9548 18232
rect 9404 17876 9456 17882
rect 9404 17818 9456 17824
rect 9324 17734 9444 17762
rect 9416 16674 9444 17734
rect 9508 16794 9536 18226
rect 9600 17377 9628 18414
rect 9770 18391 9826 18400
rect 9876 18290 9904 18634
rect 10152 18426 10180 20402
rect 10244 20330 10272 20556
rect 10520 20466 10548 22200
rect 10888 20602 10916 22200
rect 10876 20596 10928 20602
rect 10876 20538 10928 20544
rect 10600 20528 10652 20534
rect 10600 20470 10652 20476
rect 10508 20460 10560 20466
rect 10508 20402 10560 20408
rect 10416 20392 10468 20398
rect 10416 20334 10468 20340
rect 10232 20324 10284 20330
rect 10232 20266 10284 20272
rect 10428 19530 10456 20334
rect 10232 19508 10284 19514
rect 10428 19502 10548 19530
rect 10232 19450 10284 19456
rect 10244 19417 10272 19450
rect 10416 19440 10468 19446
rect 10230 19408 10286 19417
rect 10416 19382 10468 19388
rect 10230 19343 10286 19352
rect 10232 18760 10284 18766
rect 10232 18702 10284 18708
rect 10244 18601 10272 18702
rect 10230 18592 10286 18601
rect 10230 18527 10286 18536
rect 10140 18420 10192 18426
rect 10140 18362 10192 18368
rect 10428 18290 10456 19382
rect 9864 18284 9916 18290
rect 9864 18226 9916 18232
rect 10416 18284 10468 18290
rect 10416 18226 10468 18232
rect 9956 18216 10008 18222
rect 10008 18176 10088 18204
rect 9956 18158 10008 18164
rect 9680 18080 9732 18086
rect 9680 18022 9732 18028
rect 9586 17368 9642 17377
rect 9586 17303 9642 17312
rect 9496 16788 9548 16794
rect 9496 16730 9548 16736
rect 9416 16646 9628 16674
rect 9600 16522 9628 16646
rect 9588 16516 9640 16522
rect 9588 16458 9640 16464
rect 9692 16289 9720 18022
rect 9772 17876 9824 17882
rect 9772 17818 9824 17824
rect 9784 17610 9812 17818
rect 9772 17604 9824 17610
rect 9772 17546 9824 17552
rect 9954 17504 10010 17513
rect 9954 17439 10010 17448
rect 9968 17270 9996 17439
rect 9956 17264 10008 17270
rect 9956 17206 10008 17212
rect 9864 17196 9916 17202
rect 9864 17138 9916 17144
rect 9876 16794 9904 17138
rect 9864 16788 9916 16794
rect 9864 16730 9916 16736
rect 9772 16652 9824 16658
rect 9772 16594 9824 16600
rect 9956 16652 10008 16658
rect 9956 16594 10008 16600
rect 9678 16280 9734 16289
rect 9678 16215 9734 16224
rect 9404 16108 9456 16114
rect 9404 16050 9456 16056
rect 9310 15872 9366 15881
rect 9310 15807 9366 15816
rect 9324 15706 9352 15807
rect 9312 15700 9364 15706
rect 9312 15642 9364 15648
rect 9416 15502 9444 16050
rect 9680 16040 9732 16046
rect 9680 15982 9732 15988
rect 9588 15972 9640 15978
rect 9588 15914 9640 15920
rect 9404 15496 9456 15502
rect 9404 15438 9456 15444
rect 9496 15360 9548 15366
rect 9496 15302 9548 15308
rect 9220 15156 9272 15162
rect 9220 15098 9272 15104
rect 9126 15056 9182 15065
rect 9126 14991 9128 15000
rect 9180 14991 9182 15000
rect 9220 15020 9272 15026
rect 9128 14962 9180 14968
rect 9220 14962 9272 14968
rect 8392 14884 8444 14890
rect 8392 14826 8444 14832
rect 9036 14884 9088 14890
rect 9036 14826 9088 14832
rect 8404 14793 8432 14826
rect 9128 14816 9180 14822
rect 8390 14784 8446 14793
rect 9128 14758 9180 14764
rect 8390 14719 8446 14728
rect 8747 14716 9055 14725
rect 8747 14714 8753 14716
rect 8809 14714 8833 14716
rect 8889 14714 8913 14716
rect 8969 14714 8993 14716
rect 9049 14714 9055 14716
rect 8809 14662 8811 14714
rect 8991 14662 8993 14714
rect 8747 14660 8753 14662
rect 8809 14660 8833 14662
rect 8889 14660 8913 14662
rect 8969 14660 8993 14662
rect 9049 14660 9055 14662
rect 8482 14648 8538 14657
rect 8747 14651 9055 14660
rect 9140 14618 9168 14758
rect 8482 14583 8538 14592
rect 9128 14612 9180 14618
rect 8312 14470 8432 14498
rect 8300 14408 8352 14414
rect 8300 14350 8352 14356
rect 8208 13728 8260 13734
rect 8208 13670 8260 13676
rect 8220 13274 8248 13670
rect 8312 13394 8340 14350
rect 8404 14006 8432 14470
rect 8392 14000 8444 14006
rect 8392 13942 8444 13948
rect 8404 13530 8432 13942
rect 8392 13524 8444 13530
rect 8392 13466 8444 13472
rect 8300 13388 8352 13394
rect 8352 13348 8432 13376
rect 8300 13330 8352 13336
rect 8220 13246 8340 13274
rect 8206 13152 8262 13161
rect 8206 13087 8262 13096
rect 8220 12986 8248 13087
rect 8208 12980 8260 12986
rect 8208 12922 8260 12928
rect 8312 12481 8340 13246
rect 8404 12782 8432 13348
rect 8392 12776 8444 12782
rect 8392 12718 8444 12724
rect 8496 12714 8524 14583
rect 9128 14554 9180 14560
rect 9232 14482 9260 14962
rect 9508 14890 9536 15302
rect 9496 14884 9548 14890
rect 9496 14826 9548 14832
rect 9404 14816 9456 14822
rect 9404 14758 9456 14764
rect 9600 14770 9628 15914
rect 9692 15570 9720 15982
rect 9784 15910 9812 16594
rect 9864 16448 9916 16454
rect 9864 16390 9916 16396
rect 9772 15904 9824 15910
rect 9772 15846 9824 15852
rect 9876 15706 9904 16390
rect 9864 15700 9916 15706
rect 9864 15642 9916 15648
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 9692 14958 9720 15506
rect 9772 15428 9824 15434
rect 9772 15370 9824 15376
rect 9680 14952 9732 14958
rect 9680 14894 9732 14900
rect 9220 14476 9272 14482
rect 9220 14418 9272 14424
rect 8576 14340 8628 14346
rect 8576 14282 8628 14288
rect 8588 14006 8616 14282
rect 9232 14278 9260 14418
rect 8760 14272 8812 14278
rect 8758 14240 8760 14249
rect 8944 14272 8996 14278
rect 8812 14240 8814 14249
rect 8944 14214 8996 14220
rect 9220 14272 9272 14278
rect 9220 14214 9272 14220
rect 8758 14175 8814 14184
rect 8956 14074 8984 14214
rect 8944 14068 8996 14074
rect 8944 14010 8996 14016
rect 9036 14068 9088 14074
rect 9036 14010 9088 14016
rect 8576 14000 8628 14006
rect 8576 13942 8628 13948
rect 9048 13716 9076 14010
rect 9416 13870 9444 14758
rect 9600 14742 9720 14770
rect 9588 14340 9640 14346
rect 9588 14282 9640 14288
rect 9496 14272 9548 14278
rect 9494 14240 9496 14249
rect 9548 14240 9550 14249
rect 9494 14175 9550 14184
rect 9600 14074 9628 14282
rect 9588 14068 9640 14074
rect 9588 14010 9640 14016
rect 9404 13864 9456 13870
rect 9404 13806 9456 13812
rect 9496 13864 9548 13870
rect 9496 13806 9548 13812
rect 8680 13688 9076 13716
rect 9128 13728 9180 13734
rect 8574 13560 8630 13569
rect 8574 13495 8576 13504
rect 8628 13495 8630 13504
rect 8576 13466 8628 13472
rect 8576 13252 8628 13258
rect 8576 13194 8628 13200
rect 8588 12782 8616 13194
rect 8680 13138 8708 13688
rect 9128 13670 9180 13676
rect 8747 13628 9055 13637
rect 8747 13626 8753 13628
rect 8809 13626 8833 13628
rect 8889 13626 8913 13628
rect 8969 13626 8993 13628
rect 9049 13626 9055 13628
rect 8809 13574 8811 13626
rect 8991 13574 8993 13626
rect 8747 13572 8753 13574
rect 8809 13572 8833 13574
rect 8889 13572 8913 13574
rect 8969 13572 8993 13574
rect 9049 13572 9055 13574
rect 8747 13563 9055 13572
rect 9140 13326 9168 13670
rect 8944 13320 8996 13326
rect 8944 13262 8996 13268
rect 9128 13320 9180 13326
rect 9128 13262 9180 13268
rect 8852 13184 8904 13190
rect 8680 13110 8800 13138
rect 8852 13126 8904 13132
rect 8772 12918 8800 13110
rect 8864 12918 8892 13126
rect 8760 12912 8812 12918
rect 8760 12854 8812 12860
rect 8852 12912 8904 12918
rect 8852 12854 8904 12860
rect 8668 12844 8720 12850
rect 8668 12786 8720 12792
rect 8576 12776 8628 12782
rect 8576 12718 8628 12724
rect 8484 12708 8536 12714
rect 8484 12650 8536 12656
rect 8588 12594 8616 12718
rect 8496 12566 8616 12594
rect 8298 12472 8354 12481
rect 8298 12407 8354 12416
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 8220 11558 8248 12038
rect 8312 11898 8340 12407
rect 8390 12336 8446 12345
rect 8390 12271 8392 12280
rect 8444 12271 8446 12280
rect 8392 12242 8444 12248
rect 8392 12096 8444 12102
rect 8392 12038 8444 12044
rect 8300 11892 8352 11898
rect 8300 11834 8352 11840
rect 8208 11552 8260 11558
rect 8208 11494 8260 11500
rect 8298 11520 8354 11529
rect 8298 11455 8354 11464
rect 8208 11076 8260 11082
rect 8208 11018 8260 11024
rect 8220 10266 8248 11018
rect 8312 11014 8340 11455
rect 8404 11393 8432 12038
rect 8390 11384 8446 11393
rect 8390 11319 8446 11328
rect 8392 11280 8444 11286
rect 8392 11222 8444 11228
rect 8300 11008 8352 11014
rect 8300 10950 8352 10956
rect 8300 10736 8352 10742
rect 8300 10678 8352 10684
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 8114 10160 8170 10169
rect 8312 10130 8340 10678
rect 8114 10095 8170 10104
rect 8300 10124 8352 10130
rect 8300 10066 8352 10072
rect 8208 9920 8260 9926
rect 8114 9888 8170 9897
rect 8036 9846 8114 9874
rect 8208 9862 8260 9868
rect 8114 9823 8170 9832
rect 7838 9752 7894 9761
rect 7838 9687 7894 9696
rect 7840 9648 7892 9654
rect 7892 9608 7972 9636
rect 7840 9590 7892 9596
rect 7838 9208 7894 9217
rect 7838 9143 7894 9152
rect 7852 9110 7880 9143
rect 7840 9104 7892 9110
rect 7840 9046 7892 9052
rect 7748 8492 7800 8498
rect 7748 8434 7800 8440
rect 7838 8256 7894 8265
rect 7838 8191 7894 8200
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 7760 7886 7788 8026
rect 7852 7954 7880 8191
rect 7840 7948 7892 7954
rect 7840 7890 7892 7896
rect 7748 7880 7800 7886
rect 7748 7822 7800 7828
rect 7748 7744 7800 7750
rect 7748 7686 7800 7692
rect 7656 7200 7708 7206
rect 7656 7142 7708 7148
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 7472 5704 7524 5710
rect 7472 5646 7524 5652
rect 7472 5568 7524 5574
rect 7472 5510 7524 5516
rect 7484 5370 7512 5510
rect 7472 5364 7524 5370
rect 7472 5306 7524 5312
rect 7576 4826 7604 6598
rect 7564 4820 7616 4826
rect 7564 4762 7616 4768
rect 7472 4684 7524 4690
rect 7472 4626 7524 4632
rect 7484 4214 7512 4626
rect 7576 4457 7604 4762
rect 7668 4554 7696 7142
rect 7760 5710 7788 7686
rect 7840 6180 7892 6186
rect 7840 6122 7892 6128
rect 7748 5704 7800 5710
rect 7748 5646 7800 5652
rect 7852 5545 7880 6122
rect 7944 5846 7972 9608
rect 8024 9512 8076 9518
rect 8024 9454 8076 9460
rect 8036 8634 8064 9454
rect 8128 9217 8156 9823
rect 8220 9761 8248 9862
rect 8206 9752 8262 9761
rect 8312 9722 8340 10066
rect 8206 9687 8262 9696
rect 8300 9716 8352 9722
rect 8300 9658 8352 9664
rect 8208 9648 8260 9654
rect 8208 9590 8260 9596
rect 8220 9364 8248 9590
rect 8312 9518 8340 9658
rect 8404 9586 8432 11222
rect 8392 9580 8444 9586
rect 8392 9522 8444 9528
rect 8300 9512 8352 9518
rect 8300 9454 8352 9460
rect 8220 9336 8340 9364
rect 8114 9208 8170 9217
rect 8114 9143 8170 9152
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 8206 8528 8262 8537
rect 8206 8463 8262 8472
rect 8024 8356 8076 8362
rect 8024 8298 8076 8304
rect 8036 8072 8064 8298
rect 8036 8044 8156 8072
rect 8128 7954 8156 8044
rect 8116 7948 8168 7954
rect 8116 7890 8168 7896
rect 8116 7744 8168 7750
rect 8116 7686 8168 7692
rect 8022 7032 8078 7041
rect 8022 6967 8078 6976
rect 8036 6089 8064 6967
rect 8128 6730 8156 7686
rect 8116 6724 8168 6730
rect 8116 6666 8168 6672
rect 8220 6474 8248 8463
rect 8312 8362 8340 9336
rect 8404 8974 8432 9522
rect 8392 8968 8444 8974
rect 8392 8910 8444 8916
rect 8300 8356 8352 8362
rect 8300 8298 8352 8304
rect 8298 8256 8354 8265
rect 8298 8191 8354 8200
rect 8312 7818 8340 8191
rect 8300 7812 8352 7818
rect 8300 7754 8352 7760
rect 8404 7478 8432 8910
rect 8392 7472 8444 7478
rect 8392 7414 8444 7420
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 8312 6934 8340 7346
rect 8300 6928 8352 6934
rect 8300 6870 8352 6876
rect 8404 6866 8432 7414
rect 8392 6860 8444 6866
rect 8392 6802 8444 6808
rect 8392 6724 8444 6730
rect 8392 6666 8444 6672
rect 8298 6624 8354 6633
rect 8298 6559 8354 6568
rect 8128 6446 8248 6474
rect 8312 6458 8340 6559
rect 8300 6452 8352 6458
rect 8022 6080 8078 6089
rect 8128 6066 8156 6446
rect 8300 6394 8352 6400
rect 8208 6384 8260 6390
rect 8208 6326 8260 6332
rect 8220 6186 8248 6326
rect 8208 6180 8260 6186
rect 8208 6122 8260 6128
rect 8300 6112 8352 6118
rect 8128 6038 8248 6066
rect 8300 6054 8352 6060
rect 8022 6015 8078 6024
rect 7932 5840 7984 5846
rect 7932 5782 7984 5788
rect 7932 5568 7984 5574
rect 7838 5536 7894 5545
rect 7932 5510 7984 5516
rect 7838 5471 7894 5480
rect 7852 5166 7880 5471
rect 7840 5160 7892 5166
rect 7840 5102 7892 5108
rect 7748 5092 7800 5098
rect 7748 5034 7800 5040
rect 7656 4548 7708 4554
rect 7656 4490 7708 4496
rect 7562 4448 7618 4457
rect 7562 4383 7618 4392
rect 7380 4208 7432 4214
rect 7380 4150 7432 4156
rect 7472 4208 7524 4214
rect 7472 4150 7524 4156
rect 7392 3398 7420 4150
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7380 3392 7432 3398
rect 7380 3334 7432 3340
rect 7288 2984 7340 2990
rect 7288 2926 7340 2932
rect 7196 2848 7248 2854
rect 7196 2790 7248 2796
rect 7392 2514 7420 3334
rect 7472 2984 7524 2990
rect 7472 2926 7524 2932
rect 7484 2825 7512 2926
rect 7470 2816 7526 2825
rect 7470 2751 7526 2760
rect 7472 2644 7524 2650
rect 7472 2586 7524 2592
rect 7104 2508 7156 2514
rect 7104 2450 7156 2456
rect 7380 2508 7432 2514
rect 7380 2450 7432 2456
rect 7484 2038 7512 2586
rect 7380 2032 7432 2038
rect 7380 1974 7432 1980
rect 7472 2032 7524 2038
rect 7472 1974 7524 1980
rect 7392 898 7420 1974
rect 7576 1834 7604 4082
rect 7668 3058 7696 4490
rect 7760 3398 7788 5034
rect 7944 4486 7972 5510
rect 8036 5370 8064 6015
rect 8116 5840 8168 5846
rect 8116 5782 8168 5788
rect 8024 5364 8076 5370
rect 8024 5306 8076 5312
rect 8024 5228 8076 5234
rect 8024 5170 8076 5176
rect 7840 4480 7892 4486
rect 7840 4422 7892 4428
rect 7932 4480 7984 4486
rect 7932 4422 7984 4428
rect 7852 3738 7880 4422
rect 7932 4208 7984 4214
rect 7932 4150 7984 4156
rect 7944 3738 7972 4150
rect 7840 3732 7892 3738
rect 7840 3674 7892 3680
rect 7932 3732 7984 3738
rect 7932 3674 7984 3680
rect 8036 3534 8064 5170
rect 8128 4214 8156 5782
rect 8220 5642 8248 6038
rect 8208 5636 8260 5642
rect 8208 5578 8260 5584
rect 8208 4684 8260 4690
rect 8208 4626 8260 4632
rect 8116 4208 8168 4214
rect 8116 4150 8168 4156
rect 7840 3528 7892 3534
rect 7840 3470 7892 3476
rect 8024 3528 8076 3534
rect 8024 3470 8076 3476
rect 7748 3392 7800 3398
rect 7748 3334 7800 3340
rect 7852 3194 7880 3470
rect 8024 3392 8076 3398
rect 8128 3369 8156 4150
rect 8220 4010 8248 4626
rect 8208 4004 8260 4010
rect 8208 3946 8260 3952
rect 8220 3670 8248 3946
rect 8208 3664 8260 3670
rect 8208 3606 8260 3612
rect 8312 3602 8340 6054
rect 8404 4146 8432 6666
rect 8496 4758 8524 12566
rect 8680 12238 8708 12786
rect 8956 12782 8984 13262
rect 9036 13184 9088 13190
rect 9508 13138 9536 13806
rect 9588 13796 9640 13802
rect 9588 13738 9640 13744
rect 9600 13190 9628 13738
rect 9036 13126 9088 13132
rect 8944 12776 8996 12782
rect 8944 12718 8996 12724
rect 9048 12628 9076 13126
rect 9416 13110 9536 13138
rect 9588 13184 9640 13190
rect 9588 13126 9640 13132
rect 9416 12986 9444 13110
rect 9404 12980 9456 12986
rect 9404 12922 9456 12928
rect 9404 12640 9456 12646
rect 9048 12600 9260 12628
rect 8747 12540 9055 12549
rect 8747 12538 8753 12540
rect 8809 12538 8833 12540
rect 8889 12538 8913 12540
rect 8969 12538 8993 12540
rect 9049 12538 9055 12540
rect 8809 12486 8811 12538
rect 8991 12486 8993 12538
rect 8747 12484 8753 12486
rect 8809 12484 8833 12486
rect 8889 12484 8913 12486
rect 8969 12484 8993 12486
rect 9049 12484 9055 12486
rect 8747 12475 9055 12484
rect 9232 12442 9260 12600
rect 9404 12582 9456 12588
rect 9586 12608 9642 12617
rect 9220 12436 9272 12442
rect 9220 12378 9272 12384
rect 9416 12306 9444 12582
rect 9586 12543 9642 12552
rect 9496 12436 9548 12442
rect 9496 12378 9548 12384
rect 9508 12306 9536 12378
rect 9404 12300 9456 12306
rect 9404 12242 9456 12248
rect 9496 12300 9548 12306
rect 9496 12242 9548 12248
rect 8668 12232 8720 12238
rect 8588 12192 8668 12220
rect 8588 9110 8616 12192
rect 8668 12174 8720 12180
rect 9312 12096 9364 12102
rect 9312 12038 9364 12044
rect 9404 12096 9456 12102
rect 9404 12038 9456 12044
rect 8668 11892 8720 11898
rect 8668 11834 8720 11840
rect 8680 11286 8708 11834
rect 8852 11756 8904 11762
rect 8852 11698 8904 11704
rect 9128 11756 9180 11762
rect 9128 11698 9180 11704
rect 8864 11558 8892 11698
rect 8852 11552 8904 11558
rect 8852 11494 8904 11500
rect 8747 11452 9055 11461
rect 8747 11450 8753 11452
rect 8809 11450 8833 11452
rect 8889 11450 8913 11452
rect 8969 11450 8993 11452
rect 9049 11450 9055 11452
rect 8809 11398 8811 11450
rect 8991 11398 8993 11450
rect 8747 11396 8753 11398
rect 8809 11396 8833 11398
rect 8889 11396 8913 11398
rect 8969 11396 8993 11398
rect 9049 11396 9055 11398
rect 8747 11387 9055 11396
rect 9140 11286 9168 11698
rect 9220 11552 9272 11558
rect 9218 11520 9220 11529
rect 9272 11520 9274 11529
rect 9218 11455 9274 11464
rect 8668 11280 8720 11286
rect 8668 11222 8720 11228
rect 8944 11280 8996 11286
rect 9128 11280 9180 11286
rect 8944 11222 8996 11228
rect 9034 11248 9090 11257
rect 8668 11008 8720 11014
rect 8668 10950 8720 10956
rect 8680 9926 8708 10950
rect 8956 10452 8984 11222
rect 9128 11222 9180 11228
rect 9034 11183 9090 11192
rect 9048 10826 9076 11183
rect 9140 10985 9168 11222
rect 9126 10976 9182 10985
rect 9126 10911 9182 10920
rect 9048 10798 9260 10826
rect 9232 10452 9260 10798
rect 9324 10588 9352 12038
rect 9416 11218 9444 12038
rect 9600 11937 9628 12543
rect 9586 11928 9642 11937
rect 9586 11863 9642 11872
rect 9404 11212 9456 11218
rect 9404 11154 9456 11160
rect 9692 11098 9720 14742
rect 9784 13734 9812 15370
rect 9968 15162 9996 16594
rect 10060 15314 10088 18176
rect 10232 17876 10284 17882
rect 10232 17818 10284 17824
rect 10140 17196 10192 17202
rect 10140 17138 10192 17144
rect 10152 16658 10180 17138
rect 10140 16652 10192 16658
rect 10140 16594 10192 16600
rect 10152 16250 10180 16594
rect 10140 16244 10192 16250
rect 10140 16186 10192 16192
rect 10152 16114 10180 16186
rect 10140 16108 10192 16114
rect 10140 16050 10192 16056
rect 10060 15286 10180 15314
rect 10046 15192 10102 15201
rect 9956 15156 10008 15162
rect 10046 15127 10102 15136
rect 9956 15098 10008 15104
rect 9956 14544 10008 14550
rect 9956 14486 10008 14492
rect 9968 14278 9996 14486
rect 10060 14482 10088 15127
rect 10048 14476 10100 14482
rect 10048 14418 10100 14424
rect 10152 14362 10180 15286
rect 10060 14334 10180 14362
rect 9956 14272 10008 14278
rect 9956 14214 10008 14220
rect 9772 13728 9824 13734
rect 9968 13705 9996 14214
rect 9772 13670 9824 13676
rect 9954 13696 10010 13705
rect 9954 13631 10010 13640
rect 9770 13560 9826 13569
rect 9770 13495 9826 13504
rect 9784 12918 9812 13495
rect 9772 12912 9824 12918
rect 9772 12854 9824 12860
rect 10060 12850 10088 14334
rect 10140 14272 10192 14278
rect 10244 14260 10272 17818
rect 10324 17604 10376 17610
rect 10324 17546 10376 17552
rect 10416 17604 10468 17610
rect 10416 17546 10468 17552
rect 10336 17513 10364 17546
rect 10322 17504 10378 17513
rect 10322 17439 10378 17448
rect 10428 17134 10456 17546
rect 10416 17128 10468 17134
rect 10416 17070 10468 17076
rect 10428 16590 10456 17070
rect 10416 16584 10468 16590
rect 10416 16526 10468 16532
rect 10520 16402 10548 19502
rect 10612 18970 10640 20470
rect 10692 20460 10744 20466
rect 10692 20402 10744 20408
rect 10600 18964 10652 18970
rect 10600 18906 10652 18912
rect 10600 18760 10652 18766
rect 10600 18702 10652 18708
rect 10612 18601 10640 18702
rect 10598 18592 10654 18601
rect 10598 18527 10654 18536
rect 10704 18426 10732 20402
rect 10784 20392 10836 20398
rect 10782 20360 10784 20369
rect 10836 20360 10838 20369
rect 10782 20295 10838 20304
rect 10968 20324 11020 20330
rect 10968 20266 11020 20272
rect 10876 19848 10928 19854
rect 10876 19790 10928 19796
rect 10888 19446 10916 19790
rect 10980 19786 11008 20266
rect 11152 20256 11204 20262
rect 11152 20198 11204 20204
rect 11060 19916 11112 19922
rect 11060 19858 11112 19864
rect 10968 19780 11020 19786
rect 10968 19722 11020 19728
rect 10876 19440 10928 19446
rect 10782 19408 10838 19417
rect 10876 19382 10928 19388
rect 11072 19378 11100 19858
rect 10782 19343 10838 19352
rect 11060 19372 11112 19378
rect 10796 18766 10824 19343
rect 11060 19314 11112 19320
rect 10874 19272 10930 19281
rect 10874 19207 10930 19216
rect 11060 19236 11112 19242
rect 10784 18760 10836 18766
rect 10784 18702 10836 18708
rect 10692 18420 10744 18426
rect 10692 18362 10744 18368
rect 10784 18148 10836 18154
rect 10784 18090 10836 18096
rect 10692 17876 10744 17882
rect 10692 17818 10744 17824
rect 10598 17504 10654 17513
rect 10598 17439 10654 17448
rect 10612 17202 10640 17439
rect 10600 17196 10652 17202
rect 10600 17138 10652 17144
rect 10704 16998 10732 17818
rect 10692 16992 10744 16998
rect 10692 16934 10744 16940
rect 10600 16788 10652 16794
rect 10600 16730 10652 16736
rect 10612 16590 10640 16730
rect 10600 16584 10652 16590
rect 10600 16526 10652 16532
rect 10520 16374 10732 16402
rect 10506 16280 10562 16289
rect 10506 16215 10562 16224
rect 10324 15972 10376 15978
rect 10324 15914 10376 15920
rect 10336 14550 10364 15914
rect 10416 14952 10468 14958
rect 10416 14894 10468 14900
rect 10324 14544 10376 14550
rect 10324 14486 10376 14492
rect 10324 14408 10376 14414
rect 10322 14376 10324 14385
rect 10376 14376 10378 14385
rect 10322 14311 10378 14320
rect 10244 14232 10364 14260
rect 10140 14214 10192 14220
rect 10152 13977 10180 14214
rect 10230 14104 10286 14113
rect 10230 14039 10286 14048
rect 10138 13968 10194 13977
rect 10138 13903 10194 13912
rect 10244 13870 10272 14039
rect 10232 13864 10284 13870
rect 10232 13806 10284 13812
rect 10138 13696 10194 13705
rect 10138 13631 10194 13640
rect 10048 12844 10100 12850
rect 10048 12786 10100 12792
rect 9772 12708 9824 12714
rect 9772 12650 9824 12656
rect 9784 12617 9812 12650
rect 9770 12608 9826 12617
rect 9770 12543 9826 12552
rect 10060 12442 10088 12786
rect 10152 12628 10180 13631
rect 10230 13560 10286 13569
rect 10230 13495 10286 13504
rect 10244 12918 10272 13495
rect 10232 12912 10284 12918
rect 10232 12854 10284 12860
rect 10152 12600 10272 12628
rect 10048 12436 10100 12442
rect 10048 12378 10100 12384
rect 9956 12232 10008 12238
rect 9956 12174 10008 12180
rect 9862 12064 9918 12073
rect 9862 11999 9918 12008
rect 9770 11928 9826 11937
rect 9770 11863 9826 11872
rect 9600 11082 9720 11098
rect 9588 11076 9720 11082
rect 9640 11070 9720 11076
rect 9588 11018 9640 11024
rect 9680 11008 9732 11014
rect 9586 10976 9642 10985
rect 9680 10950 9732 10956
rect 9586 10911 9642 10920
rect 9324 10560 9444 10588
rect 8956 10424 9168 10452
rect 9232 10441 9352 10452
rect 9232 10432 9366 10441
rect 9232 10424 9310 10432
rect 8747 10364 9055 10373
rect 8747 10362 8753 10364
rect 8809 10362 8833 10364
rect 8889 10362 8913 10364
rect 8969 10362 8993 10364
rect 9049 10362 9055 10364
rect 8809 10310 8811 10362
rect 8991 10310 8993 10362
rect 8747 10308 8753 10310
rect 8809 10308 8833 10310
rect 8889 10308 8913 10310
rect 8969 10308 8993 10310
rect 9049 10308 9055 10310
rect 8747 10299 9055 10308
rect 9140 10282 9168 10424
rect 9310 10367 9366 10376
rect 9140 10254 9260 10282
rect 8852 10124 8904 10130
rect 8852 10066 8904 10072
rect 8864 9994 8892 10066
rect 8852 9988 8904 9994
rect 8852 9930 8904 9936
rect 8668 9920 8720 9926
rect 8944 9920 8996 9926
rect 8720 9880 8800 9908
rect 8668 9862 8720 9868
rect 8772 9625 8800 9880
rect 8942 9888 8944 9897
rect 9128 9920 9180 9926
rect 8996 9888 8998 9897
rect 9128 9862 9180 9868
rect 8942 9823 8998 9832
rect 9140 9761 9168 9862
rect 9126 9752 9182 9761
rect 9126 9687 9182 9696
rect 9128 9648 9180 9654
rect 8758 9616 8814 9625
rect 8659 9580 8711 9586
rect 9128 9590 9180 9596
rect 8758 9551 8814 9560
rect 8659 9522 8711 9528
rect 8680 9178 8708 9522
rect 8747 9276 9055 9285
rect 8747 9274 8753 9276
rect 8809 9274 8833 9276
rect 8889 9274 8913 9276
rect 8969 9274 8993 9276
rect 9049 9274 9055 9276
rect 8809 9222 8811 9274
rect 8991 9222 8993 9274
rect 8747 9220 8753 9222
rect 8809 9220 8833 9222
rect 8889 9220 8913 9222
rect 8969 9220 8993 9222
rect 9049 9220 9055 9222
rect 8747 9211 9055 9220
rect 8668 9172 8720 9178
rect 8668 9114 8720 9120
rect 8576 9104 8628 9110
rect 8576 9046 8628 9052
rect 8680 9042 8708 9114
rect 8668 9036 8720 9042
rect 8668 8978 8720 8984
rect 9036 8900 9088 8906
rect 9036 8842 9088 8848
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8588 8129 8616 8774
rect 9048 8498 9076 8842
rect 9036 8492 9088 8498
rect 9036 8434 9088 8440
rect 9140 8362 9168 9590
rect 9232 8498 9260 10254
rect 9310 10160 9366 10169
rect 9310 10095 9366 10104
rect 9324 8673 9352 10095
rect 9310 8664 9366 8673
rect 9310 8599 9366 8608
rect 9220 8492 9272 8498
rect 9220 8434 9272 8440
rect 9128 8356 9180 8362
rect 9128 8298 9180 8304
rect 8747 8188 9055 8197
rect 8747 8186 8753 8188
rect 8809 8186 8833 8188
rect 8889 8186 8913 8188
rect 8969 8186 8993 8188
rect 9049 8186 9055 8188
rect 8809 8134 8811 8186
rect 8991 8134 8993 8186
rect 8747 8132 8753 8134
rect 8809 8132 8833 8134
rect 8889 8132 8913 8134
rect 8969 8132 8993 8134
rect 9049 8132 9055 8134
rect 8574 8120 8630 8129
rect 8747 8123 9055 8132
rect 8574 8055 8630 8064
rect 9312 8084 9364 8090
rect 9312 8026 9364 8032
rect 8760 7948 8812 7954
rect 8760 7890 8812 7896
rect 8852 7948 8904 7954
rect 8852 7890 8904 7896
rect 8576 7744 8628 7750
rect 8576 7686 8628 7692
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8588 6798 8616 7686
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 8680 6458 8708 7686
rect 8772 7546 8800 7890
rect 8760 7540 8812 7546
rect 8760 7482 8812 7488
rect 8864 7410 8892 7890
rect 9324 7886 9352 8026
rect 9312 7880 9364 7886
rect 9312 7822 9364 7828
rect 8852 7404 8904 7410
rect 8852 7346 8904 7352
rect 9312 7336 9364 7342
rect 9312 7278 9364 7284
rect 9220 7268 9272 7274
rect 9220 7210 9272 7216
rect 8747 7100 9055 7109
rect 8747 7098 8753 7100
rect 8809 7098 8833 7100
rect 8889 7098 8913 7100
rect 8969 7098 8993 7100
rect 9049 7098 9055 7100
rect 8809 7046 8811 7098
rect 8991 7046 8993 7098
rect 8747 7044 8753 7046
rect 8809 7044 8833 7046
rect 8889 7044 8913 7046
rect 8969 7044 8993 7046
rect 9049 7044 9055 7046
rect 8747 7035 9055 7044
rect 8852 6860 8904 6866
rect 8852 6802 8904 6808
rect 8668 6452 8720 6458
rect 8668 6394 8720 6400
rect 8864 6361 8892 6802
rect 8944 6656 8996 6662
rect 8944 6598 8996 6604
rect 8850 6352 8906 6361
rect 8850 6287 8906 6296
rect 8956 6186 8984 6598
rect 9128 6316 9180 6322
rect 9128 6258 9180 6264
rect 8944 6180 8996 6186
rect 8944 6122 8996 6128
rect 8747 6012 9055 6021
rect 8747 6010 8753 6012
rect 8809 6010 8833 6012
rect 8889 6010 8913 6012
rect 8969 6010 8993 6012
rect 9049 6010 9055 6012
rect 8809 5958 8811 6010
rect 8991 5958 8993 6010
rect 8747 5956 8753 5958
rect 8809 5956 8833 5958
rect 8889 5956 8913 5958
rect 8969 5956 8993 5958
rect 9049 5956 9055 5958
rect 8747 5947 9055 5956
rect 8760 5772 8812 5778
rect 8760 5714 8812 5720
rect 8668 5636 8720 5642
rect 8668 5578 8720 5584
rect 8576 5568 8628 5574
rect 8576 5510 8628 5516
rect 8484 4752 8536 4758
rect 8484 4694 8536 4700
rect 8482 4312 8538 4321
rect 8482 4247 8538 4256
rect 8392 4140 8444 4146
rect 8392 4082 8444 4088
rect 8300 3596 8352 3602
rect 8300 3538 8352 3544
rect 8496 3482 8524 4247
rect 8588 4010 8616 5510
rect 8680 4826 8708 5578
rect 8772 5370 8800 5714
rect 8942 5672 8998 5681
rect 8942 5607 8998 5616
rect 8760 5364 8812 5370
rect 8760 5306 8812 5312
rect 8956 5030 8984 5607
rect 8944 5024 8996 5030
rect 8944 4966 8996 4972
rect 8747 4924 9055 4933
rect 8747 4922 8753 4924
rect 8809 4922 8833 4924
rect 8889 4922 8913 4924
rect 8969 4922 8993 4924
rect 9049 4922 9055 4924
rect 8809 4870 8811 4922
rect 8991 4870 8993 4922
rect 8747 4868 8753 4870
rect 8809 4868 8833 4870
rect 8889 4868 8913 4870
rect 8969 4868 8993 4870
rect 9049 4868 9055 4870
rect 8747 4859 9055 4868
rect 8668 4820 8720 4826
rect 8668 4762 8720 4768
rect 9036 4820 9088 4826
rect 9036 4762 9088 4768
rect 8668 4616 8720 4622
rect 8668 4558 8720 4564
rect 8576 4004 8628 4010
rect 8576 3946 8628 3952
rect 8312 3454 8524 3482
rect 8024 3334 8076 3340
rect 8114 3360 8170 3369
rect 7840 3188 7892 3194
rect 7840 3130 7892 3136
rect 7932 3188 7984 3194
rect 7932 3130 7984 3136
rect 7656 3052 7708 3058
rect 7656 2994 7708 3000
rect 7746 2952 7802 2961
rect 7944 2922 7972 3130
rect 7746 2887 7802 2896
rect 7932 2916 7984 2922
rect 7654 2680 7710 2689
rect 7654 2615 7656 2624
rect 7708 2615 7710 2624
rect 7656 2586 7708 2592
rect 7654 2408 7710 2417
rect 7654 2343 7656 2352
rect 7708 2343 7710 2352
rect 7656 2314 7708 2320
rect 7564 1828 7616 1834
rect 7564 1770 7616 1776
rect 7392 870 7512 898
rect 7392 800 7420 870
rect 6380 734 6592 762
rect 6642 0 6698 800
rect 7010 0 7066 800
rect 7378 0 7434 800
rect 7484 134 7512 870
rect 7760 800 7788 2887
rect 7932 2858 7984 2864
rect 7840 2848 7892 2854
rect 7840 2790 7892 2796
rect 7472 128 7524 134
rect 7472 70 7524 76
rect 7746 0 7802 800
rect 7852 762 7880 2790
rect 8036 2650 8064 3334
rect 8114 3295 8170 3304
rect 8312 2990 8340 3454
rect 8392 3392 8444 3398
rect 8680 3380 8708 4558
rect 8944 4480 8996 4486
rect 9048 4457 9076 4762
rect 8944 4422 8996 4428
rect 9034 4448 9090 4457
rect 8956 3942 8984 4422
rect 9034 4383 9090 4392
rect 9034 4312 9090 4321
rect 9034 4247 9090 4256
rect 9048 4214 9076 4247
rect 9036 4208 9088 4214
rect 9036 4150 9088 4156
rect 9048 4049 9076 4150
rect 9034 4040 9090 4049
rect 9034 3975 9090 3984
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 8747 3836 9055 3845
rect 8747 3834 8753 3836
rect 8809 3834 8833 3836
rect 8889 3834 8913 3836
rect 8969 3834 8993 3836
rect 9049 3834 9055 3836
rect 8809 3782 8811 3834
rect 8991 3782 8993 3834
rect 8747 3780 8753 3782
rect 8809 3780 8833 3782
rect 8889 3780 8913 3782
rect 8969 3780 8993 3782
rect 9049 3780 9055 3782
rect 8747 3771 9055 3780
rect 8944 3528 8996 3534
rect 8944 3470 8996 3476
rect 8392 3334 8444 3340
rect 8496 3352 8708 3380
rect 8300 2984 8352 2990
rect 8300 2926 8352 2932
rect 8208 2916 8260 2922
rect 8208 2858 8260 2864
rect 8116 2848 8168 2854
rect 8116 2790 8168 2796
rect 8024 2644 8076 2650
rect 8024 2586 8076 2592
rect 8128 2446 8156 2790
rect 8220 2514 8248 2858
rect 8300 2848 8352 2854
rect 8300 2790 8352 2796
rect 8312 2582 8340 2790
rect 8300 2576 8352 2582
rect 8300 2518 8352 2524
rect 8208 2508 8260 2514
rect 8208 2450 8260 2456
rect 8404 2446 8432 3334
rect 8116 2440 8168 2446
rect 8116 2382 8168 2388
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 8114 2136 8170 2145
rect 8114 2071 8170 2080
rect 8128 1358 8156 2071
rect 8116 1352 8168 1358
rect 8116 1294 8168 1300
rect 8036 870 8156 898
rect 8036 762 8064 870
rect 8128 800 8156 870
rect 8496 800 8524 3352
rect 8956 2990 8984 3470
rect 8576 2984 8628 2990
rect 8576 2926 8628 2932
rect 8944 2984 8996 2990
rect 9140 2972 9168 6258
rect 9232 5409 9260 7210
rect 9218 5400 9274 5409
rect 9218 5335 9274 5344
rect 9232 4486 9260 5335
rect 9324 5234 9352 7278
rect 9416 6186 9444 10560
rect 9496 10464 9548 10470
rect 9496 10406 9548 10412
rect 9508 10062 9536 10406
rect 9600 10130 9628 10911
rect 9692 10810 9720 10950
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9680 10600 9732 10606
rect 9678 10568 9680 10577
rect 9732 10568 9734 10577
rect 9678 10503 9734 10512
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 9496 10056 9548 10062
rect 9496 9998 9548 10004
rect 9784 9926 9812 11863
rect 9772 9920 9824 9926
rect 9772 9862 9824 9868
rect 9586 9752 9642 9761
rect 9586 9687 9642 9696
rect 9600 8634 9628 9687
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 9692 8265 9720 8366
rect 9772 8288 9824 8294
rect 9678 8256 9734 8265
rect 9772 8230 9824 8236
rect 9678 8191 9734 8200
rect 9784 8090 9812 8230
rect 9772 8084 9824 8090
rect 9772 8026 9824 8032
rect 9772 7744 9824 7750
rect 9772 7686 9824 7692
rect 9680 7472 9732 7478
rect 9600 7420 9680 7426
rect 9600 7414 9732 7420
rect 9496 7404 9548 7410
rect 9496 7346 9548 7352
rect 9600 7398 9720 7414
rect 9508 6866 9536 7346
rect 9496 6860 9548 6866
rect 9496 6802 9548 6808
rect 9508 6254 9536 6802
rect 9600 6662 9628 7398
rect 9680 7268 9732 7274
rect 9680 7210 9732 7216
rect 9588 6656 9640 6662
rect 9588 6598 9640 6604
rect 9588 6384 9640 6390
rect 9588 6326 9640 6332
rect 9496 6248 9548 6254
rect 9496 6190 9548 6196
rect 9404 6180 9456 6186
rect 9404 6122 9456 6128
rect 9416 5642 9444 6122
rect 9600 5846 9628 6326
rect 9692 6202 9720 7210
rect 9784 6322 9812 7686
rect 9876 7410 9904 11999
rect 9968 11694 9996 12174
rect 10140 12096 10192 12102
rect 10140 12038 10192 12044
rect 9956 11688 10008 11694
rect 9956 11630 10008 11636
rect 10152 11234 10180 12038
rect 10060 11206 10180 11234
rect 9956 10600 10008 10606
rect 9956 10542 10008 10548
rect 9968 10198 9996 10542
rect 9956 10192 10008 10198
rect 9956 10134 10008 10140
rect 9956 9920 10008 9926
rect 9956 9862 10008 9868
rect 9968 7721 9996 9862
rect 9954 7712 10010 7721
rect 9954 7647 10010 7656
rect 10060 7449 10088 11206
rect 10140 11144 10192 11150
rect 10140 11086 10192 11092
rect 10152 10606 10180 11086
rect 10140 10600 10192 10606
rect 10140 10542 10192 10548
rect 10244 9654 10272 12600
rect 10232 9648 10284 9654
rect 10138 9616 10194 9625
rect 10232 9590 10284 9596
rect 10138 9551 10140 9560
rect 10192 9551 10194 9560
rect 10140 9522 10192 9528
rect 10138 9072 10194 9081
rect 10138 9007 10194 9016
rect 10152 8634 10180 9007
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10152 7546 10180 8570
rect 10230 8392 10286 8401
rect 10230 8327 10232 8336
rect 10284 8327 10286 8336
rect 10232 8298 10284 8304
rect 10232 7744 10284 7750
rect 10232 7686 10284 7692
rect 10140 7540 10192 7546
rect 10140 7482 10192 7488
rect 10046 7440 10102 7449
rect 9864 7404 9916 7410
rect 10046 7375 10102 7384
rect 9864 7346 9916 7352
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9876 6746 9904 7142
rect 10152 6934 10180 7482
rect 10244 7002 10272 7686
rect 10336 7478 10364 14232
rect 10428 9674 10456 14894
rect 10520 14618 10548 16215
rect 10600 15496 10652 15502
rect 10598 15464 10600 15473
rect 10652 15464 10654 15473
rect 10598 15399 10654 15408
rect 10600 15020 10652 15026
rect 10600 14962 10652 14968
rect 10612 14793 10640 14962
rect 10598 14784 10654 14793
rect 10598 14719 10654 14728
rect 10508 14612 10560 14618
rect 10508 14554 10560 14560
rect 10520 14113 10548 14554
rect 10600 14340 10652 14346
rect 10600 14282 10652 14288
rect 10506 14104 10562 14113
rect 10506 14039 10562 14048
rect 10612 13977 10640 14282
rect 10598 13968 10654 13977
rect 10508 13932 10560 13938
rect 10598 13903 10654 13912
rect 10508 13874 10560 13880
rect 10520 13530 10548 13874
rect 10600 13864 10652 13870
rect 10598 13832 10600 13841
rect 10652 13832 10654 13841
rect 10598 13767 10654 13776
rect 10600 13728 10652 13734
rect 10600 13670 10652 13676
rect 10508 13524 10560 13530
rect 10508 13466 10560 13472
rect 10508 13388 10560 13394
rect 10508 13330 10560 13336
rect 10520 12782 10548 13330
rect 10612 12986 10640 13670
rect 10600 12980 10652 12986
rect 10600 12922 10652 12928
rect 10508 12776 10560 12782
rect 10508 12718 10560 12724
rect 10600 12708 10652 12714
rect 10600 12650 10652 12656
rect 10508 12640 10560 12646
rect 10612 12617 10640 12650
rect 10508 12582 10560 12588
rect 10598 12608 10654 12617
rect 10520 11150 10548 12582
rect 10598 12543 10654 12552
rect 10704 12434 10732 16374
rect 10796 16289 10824 18090
rect 10782 16280 10838 16289
rect 10782 16215 10838 16224
rect 10784 16040 10836 16046
rect 10784 15982 10836 15988
rect 10796 15706 10824 15982
rect 10888 15910 10916 19207
rect 11060 19178 11112 19184
rect 10966 17368 11022 17377
rect 11072 17338 11100 19178
rect 10966 17303 11022 17312
rect 11060 17332 11112 17338
rect 10980 16402 11008 17303
rect 11060 17274 11112 17280
rect 11164 16794 11192 20198
rect 11256 20058 11284 22200
rect 11624 20890 11652 22200
rect 11624 20862 11744 20890
rect 11346 20700 11654 20709
rect 11346 20698 11352 20700
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11648 20698 11654 20700
rect 11408 20646 11410 20698
rect 11590 20646 11592 20698
rect 11346 20644 11352 20646
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11648 20644 11654 20646
rect 11346 20635 11654 20644
rect 11716 20602 11744 20862
rect 11992 20602 12020 22200
rect 11704 20596 11756 20602
rect 11704 20538 11756 20544
rect 11980 20596 12032 20602
rect 12360 20584 12388 22200
rect 12728 20602 12756 22200
rect 13096 20602 13124 22200
rect 13464 20602 13492 22200
rect 13832 20602 13860 22200
rect 12440 20596 12492 20602
rect 12360 20556 12440 20584
rect 11980 20538 12032 20544
rect 12440 20538 12492 20544
rect 12716 20596 12768 20602
rect 12716 20538 12768 20544
rect 13084 20596 13136 20602
rect 13084 20538 13136 20544
rect 13452 20596 13504 20602
rect 13452 20538 13504 20544
rect 13820 20596 13872 20602
rect 13820 20538 13872 20544
rect 13634 20496 13690 20505
rect 11796 20460 11848 20466
rect 11796 20402 11848 20408
rect 13084 20460 13136 20466
rect 13634 20431 13690 20440
rect 13084 20402 13136 20408
rect 11244 20052 11296 20058
rect 11244 19994 11296 20000
rect 11244 19848 11296 19854
rect 11244 19790 11296 19796
rect 11256 18426 11284 19790
rect 11704 19712 11756 19718
rect 11704 19654 11756 19660
rect 11346 19612 11654 19621
rect 11346 19610 11352 19612
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11648 19610 11654 19612
rect 11408 19558 11410 19610
rect 11590 19558 11592 19610
rect 11346 19556 11352 19558
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11648 19556 11654 19558
rect 11346 19547 11654 19556
rect 11346 18524 11654 18533
rect 11346 18522 11352 18524
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11648 18522 11654 18524
rect 11408 18470 11410 18522
rect 11590 18470 11592 18522
rect 11346 18468 11352 18470
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11648 18468 11654 18470
rect 11346 18459 11654 18468
rect 11244 18420 11296 18426
rect 11716 18408 11744 19654
rect 11808 18970 11836 20402
rect 11888 20392 11940 20398
rect 11888 20334 11940 20340
rect 11900 19514 11928 20334
rect 12440 19984 12492 19990
rect 12440 19926 12492 19932
rect 11888 19508 11940 19514
rect 11888 19450 11940 19456
rect 12164 19440 12216 19446
rect 12164 19382 12216 19388
rect 11796 18964 11848 18970
rect 11796 18906 11848 18912
rect 12176 18834 12204 19382
rect 12268 18834 12388 18850
rect 11888 18828 11940 18834
rect 11888 18770 11940 18776
rect 12164 18828 12216 18834
rect 12164 18770 12216 18776
rect 12268 18828 12400 18834
rect 12268 18822 12348 18828
rect 11900 18426 11928 18770
rect 11980 18760 12032 18766
rect 11980 18702 12032 18708
rect 11992 18426 12020 18702
rect 12072 18624 12124 18630
rect 12072 18566 12124 18572
rect 11888 18420 11940 18426
rect 11716 18380 11836 18408
rect 11244 18362 11296 18368
rect 11704 18284 11756 18290
rect 11704 18226 11756 18232
rect 11244 18216 11296 18222
rect 11244 18158 11296 18164
rect 11256 18086 11284 18158
rect 11244 18080 11296 18086
rect 11244 18022 11296 18028
rect 11256 17610 11560 17626
rect 11256 17604 11572 17610
rect 11256 17598 11520 17604
rect 11256 17338 11284 17598
rect 11520 17546 11572 17552
rect 11346 17436 11654 17445
rect 11346 17434 11352 17436
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11648 17434 11654 17436
rect 11408 17382 11410 17434
rect 11590 17382 11592 17434
rect 11346 17380 11352 17382
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11648 17380 11654 17382
rect 11346 17371 11654 17380
rect 11244 17332 11296 17338
rect 11244 17274 11296 17280
rect 11716 16998 11744 18226
rect 11704 16992 11756 16998
rect 11704 16934 11756 16940
rect 11808 16946 11836 18380
rect 11888 18362 11940 18368
rect 11980 18420 12032 18426
rect 11980 18362 12032 18368
rect 11978 18320 12034 18329
rect 11978 18255 12034 18264
rect 11888 18080 11940 18086
rect 11886 18048 11888 18057
rect 11940 18048 11942 18057
rect 11992 18034 12020 18255
rect 12084 18154 12112 18566
rect 12176 18290 12204 18770
rect 12164 18284 12216 18290
rect 12164 18226 12216 18232
rect 12072 18148 12124 18154
rect 12072 18090 12124 18096
rect 12268 18086 12296 18822
rect 12348 18770 12400 18776
rect 12348 18352 12400 18358
rect 12348 18294 12400 18300
rect 12256 18080 12308 18086
rect 11992 18006 12204 18034
rect 12256 18022 12308 18028
rect 11886 17983 11942 17992
rect 11980 17740 12032 17746
rect 11980 17682 12032 17688
rect 11888 17672 11940 17678
rect 11888 17614 11940 17620
rect 11900 17338 11928 17614
rect 11888 17332 11940 17338
rect 11888 17274 11940 17280
rect 11992 17270 12020 17682
rect 11980 17264 12032 17270
rect 11980 17206 12032 17212
rect 11152 16788 11204 16794
rect 11152 16730 11204 16736
rect 11060 16720 11112 16726
rect 11060 16662 11112 16668
rect 11072 16522 11100 16662
rect 11716 16658 11744 16934
rect 11808 16918 11928 16946
rect 11796 16788 11848 16794
rect 11796 16730 11848 16736
rect 11152 16652 11204 16658
rect 11152 16594 11204 16600
rect 11704 16652 11756 16658
rect 11704 16594 11756 16600
rect 11060 16516 11112 16522
rect 11060 16458 11112 16464
rect 10980 16374 11100 16402
rect 10968 16040 11020 16046
rect 10968 15982 11020 15988
rect 10876 15904 10928 15910
rect 10876 15846 10928 15852
rect 10784 15700 10836 15706
rect 10784 15642 10836 15648
rect 10784 15564 10836 15570
rect 10784 15506 10836 15512
rect 10796 15162 10824 15506
rect 10980 15366 11008 15982
rect 11072 15638 11100 16374
rect 11060 15632 11112 15638
rect 11060 15574 11112 15580
rect 10968 15360 11020 15366
rect 10968 15302 11020 15308
rect 10784 15156 10836 15162
rect 10784 15098 10836 15104
rect 10876 15088 10928 15094
rect 10876 15030 10928 15036
rect 11060 15088 11112 15094
rect 11060 15030 11112 15036
rect 10782 14920 10838 14929
rect 10782 14855 10838 14864
rect 10796 14074 10824 14855
rect 10784 14068 10836 14074
rect 10784 14010 10836 14016
rect 10782 13560 10838 13569
rect 10782 13495 10838 13504
rect 10796 12986 10824 13495
rect 10784 12980 10836 12986
rect 10784 12922 10836 12928
rect 10704 12406 10824 12434
rect 10600 12164 10652 12170
rect 10600 12106 10652 12112
rect 10612 11354 10640 12106
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10600 11348 10652 11354
rect 10600 11290 10652 11296
rect 10508 11144 10560 11150
rect 10508 11086 10560 11092
rect 10704 11082 10732 12038
rect 10692 11076 10744 11082
rect 10692 11018 10744 11024
rect 10690 10840 10746 10849
rect 10690 10775 10692 10784
rect 10744 10775 10746 10784
rect 10692 10746 10744 10752
rect 10600 10600 10652 10606
rect 10600 10542 10652 10548
rect 10612 10266 10640 10542
rect 10600 10260 10652 10266
rect 10600 10202 10652 10208
rect 10598 10024 10654 10033
rect 10598 9959 10654 9968
rect 10428 9646 10548 9674
rect 10520 9518 10548 9646
rect 10416 9512 10468 9518
rect 10416 9454 10468 9460
rect 10508 9512 10560 9518
rect 10508 9454 10560 9460
rect 10428 9178 10456 9454
rect 10416 9172 10468 9178
rect 10416 9114 10468 9120
rect 10428 8430 10456 9114
rect 10520 8634 10548 9454
rect 10612 8634 10640 9959
rect 10704 9722 10732 10746
rect 10796 9994 10824 12406
rect 10888 12186 10916 15030
rect 11072 14958 11100 15030
rect 11060 14952 11112 14958
rect 11060 14894 11112 14900
rect 11058 14512 11114 14521
rect 11058 14447 11114 14456
rect 10966 14104 11022 14113
rect 11072 14074 11100 14447
rect 10966 14039 11022 14048
rect 11060 14068 11112 14074
rect 10980 13802 11008 14039
rect 11060 14010 11112 14016
rect 10968 13796 11020 13802
rect 10968 13738 11020 13744
rect 11058 13016 11114 13025
rect 11058 12951 11060 12960
rect 11112 12951 11114 12960
rect 11060 12922 11112 12928
rect 11060 12640 11112 12646
rect 11060 12582 11112 12588
rect 11072 12238 11100 12582
rect 11164 12434 11192 16594
rect 11244 16448 11296 16454
rect 11808 16425 11836 16730
rect 11244 16390 11296 16396
rect 11794 16416 11850 16425
rect 11256 15706 11284 16390
rect 11346 16348 11654 16357
rect 11794 16351 11850 16360
rect 11346 16346 11352 16348
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11648 16346 11654 16348
rect 11408 16294 11410 16346
rect 11590 16294 11592 16346
rect 11346 16292 11352 16294
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11648 16292 11654 16294
rect 11346 16283 11654 16292
rect 11336 16244 11388 16250
rect 11900 16232 11928 16918
rect 11980 16448 12032 16454
rect 11980 16390 12032 16396
rect 11336 16186 11388 16192
rect 11716 16204 11928 16232
rect 11348 16017 11376 16186
rect 11610 16144 11666 16153
rect 11610 16079 11612 16088
rect 11664 16079 11666 16088
rect 11612 16050 11664 16056
rect 11520 16040 11572 16046
rect 11334 16008 11390 16017
rect 11334 15943 11390 15952
rect 11518 16008 11520 16017
rect 11572 16008 11574 16017
rect 11518 15943 11574 15952
rect 11244 15700 11296 15706
rect 11244 15642 11296 15648
rect 11348 15348 11376 15943
rect 11256 15320 11376 15348
rect 11256 14056 11284 15320
rect 11346 15260 11654 15269
rect 11346 15258 11352 15260
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11648 15258 11654 15260
rect 11408 15206 11410 15258
rect 11590 15206 11592 15258
rect 11346 15204 11352 15206
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11648 15204 11654 15206
rect 11346 15195 11654 15204
rect 11346 14172 11654 14181
rect 11346 14170 11352 14172
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11648 14170 11654 14172
rect 11408 14118 11410 14170
rect 11590 14118 11592 14170
rect 11346 14116 11352 14118
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11648 14116 11654 14118
rect 11346 14107 11654 14116
rect 11428 14068 11480 14074
rect 11256 14028 11376 14056
rect 11244 13728 11296 13734
rect 11244 13670 11296 13676
rect 11256 12850 11284 13670
rect 11348 13530 11376 14028
rect 11428 14010 11480 14016
rect 11440 13705 11468 14010
rect 11716 13954 11744 16204
rect 11886 16144 11942 16153
rect 11796 16108 11848 16114
rect 11886 16079 11942 16088
rect 11796 16050 11848 16056
rect 11808 14482 11836 16050
rect 11900 15008 11928 16079
rect 11992 15638 12020 16390
rect 12070 16280 12126 16289
rect 12176 16250 12204 18006
rect 12268 16833 12296 18022
rect 12254 16824 12310 16833
rect 12360 16794 12388 18294
rect 12452 18086 12480 19926
rect 12992 19848 13044 19854
rect 12992 19790 13044 19796
rect 13004 19514 13032 19790
rect 13096 19514 13124 20402
rect 13176 19780 13228 19786
rect 13176 19722 13228 19728
rect 12992 19508 13044 19514
rect 12992 19450 13044 19456
rect 13084 19508 13136 19514
rect 13084 19450 13136 19456
rect 12900 19304 12952 19310
rect 12900 19246 12952 19252
rect 12808 19168 12860 19174
rect 12808 19110 12860 19116
rect 12532 18624 12584 18630
rect 12532 18566 12584 18572
rect 12544 18426 12572 18566
rect 12532 18420 12584 18426
rect 12532 18362 12584 18368
rect 12440 18080 12492 18086
rect 12440 18022 12492 18028
rect 12820 17746 12848 19110
rect 12912 18970 12940 19246
rect 13188 19174 13216 19722
rect 13544 19712 13596 19718
rect 13544 19654 13596 19660
rect 13360 19372 13412 19378
rect 13360 19314 13412 19320
rect 13176 19168 13228 19174
rect 13176 19110 13228 19116
rect 12900 18964 12952 18970
rect 12900 18906 12952 18912
rect 13188 18834 13216 19110
rect 13372 18970 13400 19314
rect 13556 19310 13584 19654
rect 13544 19304 13596 19310
rect 13544 19246 13596 19252
rect 13360 18964 13412 18970
rect 13360 18906 13412 18912
rect 12900 18828 12952 18834
rect 12900 18770 12952 18776
rect 13176 18828 13228 18834
rect 13176 18770 13228 18776
rect 12912 18329 12940 18770
rect 13452 18692 13504 18698
rect 13452 18634 13504 18640
rect 13268 18624 13320 18630
rect 13268 18566 13320 18572
rect 12898 18320 12954 18329
rect 12898 18255 12954 18264
rect 13084 18284 13136 18290
rect 13084 18226 13136 18232
rect 13096 18057 13124 18226
rect 13176 18216 13228 18222
rect 13176 18158 13228 18164
rect 13082 18048 13138 18057
rect 13082 17983 13138 17992
rect 13188 17882 13216 18158
rect 13176 17876 13228 17882
rect 13176 17818 13228 17824
rect 13082 17776 13138 17785
rect 12808 17740 12860 17746
rect 13082 17711 13138 17720
rect 12808 17682 12860 17688
rect 12624 17672 12676 17678
rect 12624 17614 12676 17620
rect 12440 17536 12492 17542
rect 12440 17478 12492 17484
rect 12452 17338 12480 17478
rect 12440 17332 12492 17338
rect 12440 17274 12492 17280
rect 12532 17060 12584 17066
rect 12532 17002 12584 17008
rect 12254 16759 12310 16768
rect 12348 16788 12400 16794
rect 12348 16730 12400 16736
rect 12440 16720 12492 16726
rect 12438 16688 12440 16697
rect 12492 16688 12494 16697
rect 12438 16623 12494 16632
rect 12438 16552 12494 16561
rect 12544 16538 12572 17002
rect 12494 16510 12572 16538
rect 12438 16487 12494 16496
rect 12532 16448 12584 16454
rect 12346 16416 12402 16425
rect 12532 16390 12584 16396
rect 12346 16351 12402 16360
rect 12070 16215 12126 16224
rect 12164 16244 12216 16250
rect 12084 16182 12112 16215
rect 12164 16186 12216 16192
rect 12072 16176 12124 16182
rect 12072 16118 12124 16124
rect 12254 16144 12310 16153
rect 12254 16079 12310 16088
rect 12268 15881 12296 16079
rect 12254 15872 12310 15881
rect 12254 15807 12310 15816
rect 11980 15632 12032 15638
rect 11980 15574 12032 15580
rect 11980 15360 12032 15366
rect 11978 15328 11980 15337
rect 12032 15328 12034 15337
rect 11978 15263 12034 15272
rect 12256 15156 12308 15162
rect 12256 15098 12308 15104
rect 11900 14980 12204 15008
rect 12070 14920 12126 14929
rect 12070 14855 12126 14864
rect 11888 14612 11940 14618
rect 11888 14554 11940 14560
rect 11796 14476 11848 14482
rect 11796 14418 11848 14424
rect 11624 13926 11744 13954
rect 11520 13864 11572 13870
rect 11518 13832 11520 13841
rect 11572 13832 11574 13841
rect 11518 13767 11574 13776
rect 11426 13696 11482 13705
rect 11426 13631 11482 13640
rect 11624 13530 11652 13926
rect 11900 13870 11928 14554
rect 11980 14476 12032 14482
rect 11980 14418 12032 14424
rect 11704 13864 11756 13870
rect 11704 13806 11756 13812
rect 11888 13864 11940 13870
rect 11888 13806 11940 13812
rect 11336 13524 11388 13530
rect 11336 13466 11388 13472
rect 11612 13524 11664 13530
rect 11612 13466 11664 13472
rect 11348 13190 11376 13466
rect 11624 13326 11652 13466
rect 11716 13433 11744 13806
rect 11992 13734 12020 14418
rect 11980 13728 12032 13734
rect 11980 13670 12032 13676
rect 11978 13560 12034 13569
rect 11978 13495 11980 13504
rect 12032 13495 12034 13504
rect 11980 13466 12032 13472
rect 11702 13424 11758 13433
rect 12084 13410 12112 14855
rect 11702 13359 11758 13368
rect 11992 13382 12112 13410
rect 11612 13320 11664 13326
rect 11888 13320 11940 13326
rect 11664 13280 11744 13308
rect 11612 13262 11664 13268
rect 11336 13184 11388 13190
rect 11336 13126 11388 13132
rect 11346 13084 11654 13093
rect 11346 13082 11352 13084
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11648 13082 11654 13084
rect 11408 13030 11410 13082
rect 11590 13030 11592 13082
rect 11346 13028 11352 13030
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11648 13028 11654 13030
rect 11346 13019 11654 13028
rect 11244 12844 11296 12850
rect 11244 12786 11296 12792
rect 11716 12764 11744 13280
rect 11888 13262 11940 13268
rect 11796 12844 11848 12850
rect 11796 12786 11848 12792
rect 11624 12736 11744 12764
rect 11164 12406 11284 12434
rect 11060 12232 11112 12238
rect 10888 12158 11008 12186
rect 11060 12174 11112 12180
rect 10876 11280 10928 11286
rect 10876 11222 10928 11228
rect 10888 10674 10916 11222
rect 10876 10668 10928 10674
rect 10876 10610 10928 10616
rect 10980 10033 11008 12158
rect 11072 11218 11100 12174
rect 11060 11212 11112 11218
rect 11060 11154 11112 11160
rect 11256 11098 11284 12406
rect 11624 12170 11652 12736
rect 11808 12434 11836 12786
rect 11716 12406 11836 12434
rect 11612 12164 11664 12170
rect 11612 12106 11664 12112
rect 11346 11996 11654 12005
rect 11346 11994 11352 11996
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11648 11994 11654 11996
rect 11408 11942 11410 11994
rect 11590 11942 11592 11994
rect 11346 11940 11352 11942
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11648 11940 11654 11942
rect 11346 11931 11654 11940
rect 11612 11892 11664 11898
rect 11612 11834 11664 11840
rect 11518 11248 11574 11257
rect 11624 11218 11652 11834
rect 11716 11830 11744 12406
rect 11796 12232 11848 12238
rect 11796 12174 11848 12180
rect 11808 11898 11836 12174
rect 11796 11892 11848 11898
rect 11796 11834 11848 11840
rect 11704 11824 11756 11830
rect 11704 11766 11756 11772
rect 11716 11694 11744 11766
rect 11704 11688 11756 11694
rect 11796 11688 11848 11694
rect 11704 11630 11756 11636
rect 11794 11656 11796 11665
rect 11848 11656 11850 11665
rect 11518 11183 11574 11192
rect 11612 11212 11664 11218
rect 11532 11150 11560 11183
rect 11612 11154 11664 11160
rect 11072 11070 11284 11098
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 10966 10024 11022 10033
rect 10784 9988 10836 9994
rect 10966 9959 11022 9968
rect 10784 9930 10836 9936
rect 10692 9716 10744 9722
rect 10692 9658 10744 9664
rect 10692 9580 10744 9586
rect 10692 9522 10744 9528
rect 10508 8628 10560 8634
rect 10508 8570 10560 8576
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 10520 8498 10548 8570
rect 10508 8492 10560 8498
rect 10508 8434 10560 8440
rect 10416 8424 10468 8430
rect 10416 8366 10468 8372
rect 10414 7984 10470 7993
rect 10414 7919 10470 7928
rect 10324 7472 10376 7478
rect 10324 7414 10376 7420
rect 10232 6996 10284 7002
rect 10232 6938 10284 6944
rect 10140 6928 10192 6934
rect 10336 6905 10364 7414
rect 10428 7041 10456 7919
rect 10414 7032 10470 7041
rect 10414 6967 10470 6976
rect 10140 6870 10192 6876
rect 10322 6896 10378 6905
rect 10322 6831 10378 6840
rect 10048 6792 10100 6798
rect 9876 6718 9996 6746
rect 10048 6734 10100 6740
rect 9864 6656 9916 6662
rect 9864 6598 9916 6604
rect 9772 6316 9824 6322
rect 9772 6258 9824 6264
rect 9692 6174 9812 6202
rect 9680 6112 9732 6118
rect 9680 6054 9732 6060
rect 9588 5840 9640 5846
rect 9588 5782 9640 5788
rect 9692 5778 9720 6054
rect 9680 5772 9732 5778
rect 9680 5714 9732 5720
rect 9404 5636 9456 5642
rect 9784 5624 9812 6174
rect 9876 5778 9904 6598
rect 9864 5772 9916 5778
rect 9864 5714 9916 5720
rect 9404 5578 9456 5584
rect 9692 5596 9812 5624
rect 9864 5636 9916 5642
rect 9692 5522 9720 5596
rect 9864 5578 9916 5584
rect 9600 5494 9720 5522
rect 9312 5228 9364 5234
rect 9312 5170 9364 5176
rect 9600 5001 9628 5494
rect 9680 5296 9732 5302
rect 9680 5238 9732 5244
rect 9586 4992 9642 5001
rect 9586 4927 9642 4936
rect 9692 4690 9720 5238
rect 9876 5001 9904 5578
rect 9862 4992 9918 5001
rect 9862 4927 9918 4936
rect 9968 4826 9996 6718
rect 10060 6390 10088 6734
rect 10416 6656 10468 6662
rect 10416 6598 10468 6604
rect 10048 6384 10100 6390
rect 10048 6326 10100 6332
rect 10060 5234 10088 6326
rect 10324 6316 10376 6322
rect 10324 6258 10376 6264
rect 10336 6225 10364 6258
rect 10322 6216 10378 6225
rect 10322 6151 10378 6160
rect 10140 5568 10192 5574
rect 10140 5510 10192 5516
rect 10230 5536 10286 5545
rect 10152 5370 10180 5510
rect 10230 5471 10286 5480
rect 10140 5364 10192 5370
rect 10140 5306 10192 5312
rect 10138 5264 10194 5273
rect 10048 5228 10100 5234
rect 10138 5199 10194 5208
rect 10048 5170 10100 5176
rect 10152 5030 10180 5199
rect 10140 5024 10192 5030
rect 10140 4966 10192 4972
rect 9956 4820 10008 4826
rect 9956 4762 10008 4768
rect 9680 4684 9732 4690
rect 9680 4626 9732 4632
rect 9772 4684 9824 4690
rect 9772 4626 9824 4632
rect 9220 4480 9272 4486
rect 9220 4422 9272 4428
rect 9586 4312 9642 4321
rect 9586 4247 9642 4256
rect 9600 4146 9628 4247
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 9496 3936 9548 3942
rect 9496 3878 9548 3884
rect 9232 3126 9260 3878
rect 9508 3641 9536 3878
rect 9494 3632 9550 3641
rect 9494 3567 9550 3576
rect 9404 3392 9456 3398
rect 9404 3334 9456 3340
rect 9416 3194 9444 3334
rect 9508 3233 9536 3567
rect 9494 3224 9550 3233
rect 9404 3188 9456 3194
rect 9494 3159 9550 3168
rect 9404 3130 9456 3136
rect 9220 3120 9272 3126
rect 9220 3062 9272 3068
rect 9140 2944 9260 2972
rect 8944 2926 8996 2932
rect 8588 1970 8616 2926
rect 8747 2748 9055 2757
rect 8747 2746 8753 2748
rect 8809 2746 8833 2748
rect 8889 2746 8913 2748
rect 8969 2746 8993 2748
rect 9049 2746 9055 2748
rect 8809 2694 8811 2746
rect 8991 2694 8993 2746
rect 8747 2692 8753 2694
rect 8809 2692 8833 2694
rect 8889 2692 8913 2694
rect 8969 2692 8993 2694
rect 9049 2692 9055 2694
rect 8747 2683 9055 2692
rect 8668 2576 8720 2582
rect 8668 2518 8720 2524
rect 8680 2446 8708 2518
rect 8668 2440 8720 2446
rect 8668 2382 8720 2388
rect 8576 1964 8628 1970
rect 8576 1906 8628 1912
rect 8852 1896 8904 1902
rect 8852 1838 8904 1844
rect 8864 800 8892 1838
rect 9232 800 9260 2944
rect 9310 2680 9366 2689
rect 9310 2615 9366 2624
rect 9324 2310 9352 2615
rect 9402 2544 9458 2553
rect 9402 2479 9458 2488
rect 9416 2446 9444 2479
rect 9404 2440 9456 2446
rect 9404 2382 9456 2388
rect 9312 2304 9364 2310
rect 9312 2246 9364 2252
rect 9496 2304 9548 2310
rect 9496 2246 9548 2252
rect 9324 1465 9352 2246
rect 9508 1601 9536 2246
rect 9494 1592 9550 1601
rect 9494 1527 9550 1536
rect 9310 1456 9366 1465
rect 9310 1391 9366 1400
rect 9600 800 9628 4082
rect 9692 4078 9720 4626
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 9692 1698 9720 3878
rect 9784 3126 9812 4626
rect 10244 4622 10272 5471
rect 10324 5024 10376 5030
rect 10324 4966 10376 4972
rect 10232 4616 10284 4622
rect 10232 4558 10284 4564
rect 9954 4448 10010 4457
rect 9954 4383 10010 4392
rect 9862 3632 9918 3641
rect 9862 3567 9918 3576
rect 9876 3369 9904 3567
rect 9862 3360 9918 3369
rect 9862 3295 9918 3304
rect 9772 3120 9824 3126
rect 9772 3062 9824 3068
rect 9784 2582 9812 3062
rect 9864 2984 9916 2990
rect 9864 2926 9916 2932
rect 9876 2650 9904 2926
rect 9864 2644 9916 2650
rect 9864 2586 9916 2592
rect 9772 2576 9824 2582
rect 9772 2518 9824 2524
rect 9968 2446 9996 4383
rect 10336 4146 10364 4966
rect 10324 4140 10376 4146
rect 10324 4082 10376 4088
rect 10232 4072 10284 4078
rect 10232 4014 10284 4020
rect 10140 3460 10192 3466
rect 10140 3402 10192 3408
rect 9956 2440 10008 2446
rect 10152 2417 10180 3402
rect 10244 3398 10272 4014
rect 10322 3768 10378 3777
rect 10322 3703 10324 3712
rect 10376 3703 10378 3712
rect 10324 3674 10376 3680
rect 10232 3392 10284 3398
rect 10232 3334 10284 3340
rect 10244 3058 10272 3334
rect 10324 3188 10376 3194
rect 10324 3130 10376 3136
rect 10232 3052 10284 3058
rect 10232 2994 10284 3000
rect 10336 2825 10364 3130
rect 10322 2816 10378 2825
rect 10322 2751 10378 2760
rect 10428 2774 10456 6598
rect 10520 6361 10548 8434
rect 10600 7880 10652 7886
rect 10600 7822 10652 7828
rect 10612 6798 10640 7822
rect 10704 7449 10732 9522
rect 10796 8922 10824 9930
rect 10876 9648 10928 9654
rect 10876 9590 10928 9596
rect 10888 9489 10916 9590
rect 11072 9518 11100 11070
rect 11150 10976 11206 10985
rect 11150 10911 11206 10920
rect 11060 9512 11112 9518
rect 10874 9480 10930 9489
rect 11060 9454 11112 9460
rect 10874 9415 10930 9424
rect 10966 9344 11022 9353
rect 10966 9279 11022 9288
rect 10980 9178 11008 9279
rect 10968 9172 11020 9178
rect 10968 9114 11020 9120
rect 10796 8894 10916 8922
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10796 7886 10824 8774
rect 10784 7880 10836 7886
rect 10784 7822 10836 7828
rect 10888 7818 10916 8894
rect 11060 8832 11112 8838
rect 11060 8774 11112 8780
rect 11072 8294 11100 8774
rect 11060 8288 11112 8294
rect 11060 8230 11112 8236
rect 11164 7936 11192 10911
rect 11346 10908 11654 10917
rect 11346 10906 11352 10908
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11648 10906 11654 10908
rect 11408 10854 11410 10906
rect 11590 10854 11592 10906
rect 11346 10852 11352 10854
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11648 10852 11654 10854
rect 11346 10843 11654 10852
rect 11242 10704 11298 10713
rect 11242 10639 11244 10648
rect 11296 10639 11298 10648
rect 11244 10610 11296 10616
rect 11716 10606 11744 11630
rect 11794 11591 11850 11600
rect 11796 11552 11848 11558
rect 11796 11494 11848 11500
rect 11808 11150 11836 11494
rect 11796 11144 11848 11150
rect 11796 11086 11848 11092
rect 11704 10600 11756 10606
rect 11704 10542 11756 10548
rect 11518 10160 11574 10169
rect 11518 10095 11574 10104
rect 11704 10124 11756 10130
rect 11532 9994 11560 10095
rect 11704 10066 11756 10072
rect 11716 9994 11744 10066
rect 11244 9988 11296 9994
rect 11244 9930 11296 9936
rect 11520 9988 11572 9994
rect 11520 9930 11572 9936
rect 11704 9988 11756 9994
rect 11704 9930 11756 9936
rect 11256 8022 11284 9930
rect 11346 9820 11654 9829
rect 11346 9818 11352 9820
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11648 9818 11654 9820
rect 11408 9766 11410 9818
rect 11590 9766 11592 9818
rect 11346 9764 11352 9766
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11648 9764 11654 9766
rect 11346 9755 11654 9764
rect 11336 9580 11388 9586
rect 11336 9522 11388 9528
rect 11612 9580 11664 9586
rect 11612 9522 11664 9528
rect 11348 9178 11376 9522
rect 11520 9512 11572 9518
rect 11520 9454 11572 9460
rect 11336 9172 11388 9178
rect 11336 9114 11388 9120
rect 11532 9092 11560 9454
rect 11624 9217 11652 9522
rect 11716 9518 11744 9930
rect 11794 9616 11850 9625
rect 11794 9551 11850 9560
rect 11704 9512 11756 9518
rect 11704 9454 11756 9460
rect 11808 9217 11836 9551
rect 11610 9208 11666 9217
rect 11610 9143 11666 9152
rect 11794 9208 11850 9217
rect 11794 9143 11850 9152
rect 11532 9064 11836 9092
rect 11704 8900 11756 8906
rect 11704 8842 11756 8848
rect 11346 8732 11654 8741
rect 11346 8730 11352 8732
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11648 8730 11654 8732
rect 11408 8678 11410 8730
rect 11590 8678 11592 8730
rect 11346 8676 11352 8678
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11648 8676 11654 8678
rect 11346 8667 11654 8676
rect 11612 8424 11664 8430
rect 11612 8366 11664 8372
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 11244 8016 11296 8022
rect 11244 7958 11296 7964
rect 11072 7908 11192 7936
rect 10876 7812 10928 7818
rect 10876 7754 10928 7760
rect 10782 7576 10838 7585
rect 10782 7511 10838 7520
rect 10690 7440 10746 7449
rect 10690 7375 10746 7384
rect 10796 7177 10824 7511
rect 10888 7478 10916 7754
rect 10876 7472 10928 7478
rect 10876 7414 10928 7420
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 10980 7290 11008 7346
rect 10888 7274 11008 7290
rect 10876 7268 11008 7274
rect 10928 7262 11008 7268
rect 10876 7210 10928 7216
rect 10968 7200 11020 7206
rect 10782 7168 10838 7177
rect 10968 7142 11020 7148
rect 10782 7103 10838 7112
rect 10876 6996 10928 7002
rect 10876 6938 10928 6944
rect 10600 6792 10652 6798
rect 10600 6734 10652 6740
rect 10692 6724 10744 6730
rect 10692 6666 10744 6672
rect 10600 6384 10652 6390
rect 10506 6352 10562 6361
rect 10600 6326 10652 6332
rect 10506 6287 10562 6296
rect 10612 5914 10640 6326
rect 10704 6118 10732 6666
rect 10888 6497 10916 6938
rect 10980 6633 11008 7142
rect 10966 6624 11022 6633
rect 10966 6559 11022 6568
rect 10874 6488 10930 6497
rect 10874 6423 10930 6432
rect 10784 6180 10836 6186
rect 10784 6122 10836 6128
rect 10692 6112 10744 6118
rect 10692 6054 10744 6060
rect 10600 5908 10652 5914
rect 10600 5850 10652 5856
rect 10600 5704 10652 5710
rect 10600 5646 10652 5652
rect 10508 5568 10560 5574
rect 10508 5510 10560 5516
rect 10520 5234 10548 5510
rect 10508 5228 10560 5234
rect 10508 5170 10560 5176
rect 10612 4826 10640 5646
rect 10704 5166 10732 6054
rect 10796 5370 10824 6122
rect 10876 6112 10928 6118
rect 10876 6054 10928 6060
rect 10888 5914 10916 6054
rect 10980 5953 11008 6559
rect 10966 5944 11022 5953
rect 10876 5908 10928 5914
rect 10966 5879 11022 5888
rect 10876 5850 10928 5856
rect 10968 5840 11020 5846
rect 10968 5782 11020 5788
rect 10876 5772 10928 5778
rect 10876 5714 10928 5720
rect 10784 5364 10836 5370
rect 10784 5306 10836 5312
rect 10692 5160 10744 5166
rect 10692 5102 10744 5108
rect 10600 4820 10652 4826
rect 10600 4762 10652 4768
rect 10784 4820 10836 4826
rect 10784 4762 10836 4768
rect 10508 4004 10560 4010
rect 10508 3946 10560 3952
rect 10520 3534 10548 3946
rect 10692 3936 10744 3942
rect 10692 3878 10744 3884
rect 10508 3528 10560 3534
rect 10508 3470 10560 3476
rect 10704 3466 10732 3878
rect 10692 3460 10744 3466
rect 10692 3402 10744 3408
rect 10138 2408 10194 2417
rect 9956 2382 10008 2388
rect 10060 2366 10138 2394
rect 10060 1714 10088 2366
rect 10138 2343 10194 2352
rect 10232 2304 10284 2310
rect 10232 2246 10284 2252
rect 10244 2106 10272 2246
rect 10232 2100 10284 2106
rect 10232 2042 10284 2048
rect 9680 1692 9732 1698
rect 9680 1634 9732 1640
rect 9968 1686 10088 1714
rect 9968 800 9996 1686
rect 10336 800 10364 2751
rect 10428 2746 10732 2774
rect 10600 2304 10652 2310
rect 10600 2246 10652 2252
rect 10612 1358 10640 2246
rect 10600 1352 10652 1358
rect 10600 1294 10652 1300
rect 10704 800 10732 2746
rect 10796 1902 10824 4762
rect 10888 3670 10916 5714
rect 10980 4622 11008 5782
rect 10968 4616 11020 4622
rect 10968 4558 11020 4564
rect 11072 4570 11100 7908
rect 11256 7868 11284 7958
rect 11348 7954 11376 8230
rect 11624 7993 11652 8366
rect 11716 8294 11744 8842
rect 11808 8430 11836 9064
rect 11796 8424 11848 8430
rect 11796 8366 11848 8372
rect 11704 8288 11756 8294
rect 11704 8230 11756 8236
rect 11610 7984 11666 7993
rect 11336 7948 11388 7954
rect 11610 7919 11666 7928
rect 11336 7890 11388 7896
rect 11164 7840 11284 7868
rect 11164 7410 11192 7840
rect 11244 7744 11296 7750
rect 11244 7686 11296 7692
rect 11256 7546 11284 7686
rect 11346 7644 11654 7653
rect 11346 7642 11352 7644
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11648 7642 11654 7644
rect 11408 7590 11410 7642
rect 11590 7590 11592 7642
rect 11346 7588 11352 7590
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11648 7588 11654 7590
rect 11346 7579 11654 7588
rect 11244 7540 11296 7546
rect 11244 7482 11296 7488
rect 11152 7404 11204 7410
rect 11152 7346 11204 7352
rect 11716 7342 11744 8230
rect 11796 8084 11848 8090
rect 11796 8026 11848 8032
rect 11704 7336 11756 7342
rect 11704 7278 11756 7284
rect 11244 7268 11296 7274
rect 11244 7210 11296 7216
rect 11256 6440 11284 7210
rect 11612 7200 11664 7206
rect 11612 7142 11664 7148
rect 11624 6934 11652 7142
rect 11612 6928 11664 6934
rect 11612 6870 11664 6876
rect 11808 6848 11836 8026
rect 11716 6820 11836 6848
rect 11334 6760 11390 6769
rect 11334 6695 11390 6704
rect 11348 6662 11376 6695
rect 11336 6656 11388 6662
rect 11336 6598 11388 6604
rect 11346 6556 11654 6565
rect 11346 6554 11352 6556
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11648 6554 11654 6556
rect 11408 6502 11410 6554
rect 11590 6502 11592 6554
rect 11346 6500 11352 6502
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11648 6500 11654 6502
rect 11346 6491 11654 6500
rect 11256 6412 11376 6440
rect 11150 6216 11206 6225
rect 11150 6151 11206 6160
rect 11164 5166 11192 6151
rect 11244 6112 11296 6118
rect 11242 6080 11244 6089
rect 11296 6080 11298 6089
rect 11242 6015 11298 6024
rect 11256 5574 11284 6015
rect 11348 5953 11376 6412
rect 11610 6216 11666 6225
rect 11610 6151 11612 6160
rect 11664 6151 11666 6160
rect 11612 6122 11664 6128
rect 11610 6080 11666 6089
rect 11610 6015 11666 6024
rect 11334 5944 11390 5953
rect 11334 5879 11390 5888
rect 11348 5642 11376 5879
rect 11336 5636 11388 5642
rect 11336 5578 11388 5584
rect 11624 5574 11652 6015
rect 11244 5568 11296 5574
rect 11244 5510 11296 5516
rect 11612 5568 11664 5574
rect 11612 5510 11664 5516
rect 11346 5468 11654 5477
rect 11346 5466 11352 5468
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11648 5466 11654 5468
rect 11408 5414 11410 5466
rect 11590 5414 11592 5466
rect 11346 5412 11352 5414
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11648 5412 11654 5414
rect 11346 5403 11654 5412
rect 11612 5364 11664 5370
rect 11612 5306 11664 5312
rect 11624 5234 11652 5306
rect 11612 5228 11664 5234
rect 11612 5170 11664 5176
rect 11152 5160 11204 5166
rect 11152 5102 11204 5108
rect 11164 4690 11192 5102
rect 11152 4684 11204 4690
rect 11152 4626 11204 4632
rect 11072 4542 11192 4570
rect 10876 3664 10928 3670
rect 10876 3606 10928 3612
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 10888 2650 10916 3470
rect 11058 3224 11114 3233
rect 11058 3159 11114 3168
rect 11072 2990 11100 3159
rect 11060 2984 11112 2990
rect 11060 2926 11112 2932
rect 10968 2916 11020 2922
rect 10968 2858 11020 2864
rect 10876 2644 10928 2650
rect 10876 2586 10928 2592
rect 10980 2009 11008 2858
rect 11164 2650 11192 4542
rect 11346 4380 11654 4389
rect 11346 4378 11352 4380
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11648 4378 11654 4380
rect 11408 4326 11410 4378
rect 11590 4326 11592 4378
rect 11346 4324 11352 4326
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11648 4324 11654 4326
rect 11346 4315 11654 4324
rect 11244 4208 11296 4214
rect 11244 4150 11296 4156
rect 11256 2854 11284 4150
rect 11612 4140 11664 4146
rect 11612 4082 11664 4088
rect 11624 3738 11652 4082
rect 11612 3732 11664 3738
rect 11612 3674 11664 3680
rect 11346 3292 11654 3301
rect 11346 3290 11352 3292
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11648 3290 11654 3292
rect 11408 3238 11410 3290
rect 11590 3238 11592 3290
rect 11346 3236 11352 3238
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11648 3236 11654 3238
rect 11346 3227 11654 3236
rect 11244 2848 11296 2854
rect 11244 2790 11296 2796
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 11716 2446 11744 6820
rect 11796 6724 11848 6730
rect 11796 6666 11848 6672
rect 11808 2774 11836 6666
rect 11900 6458 11928 13262
rect 11992 11286 12020 13382
rect 12072 13184 12124 13190
rect 12072 13126 12124 13132
rect 12084 12986 12112 13126
rect 12072 12980 12124 12986
rect 12072 12922 12124 12928
rect 12176 11937 12204 14980
rect 12268 14958 12296 15098
rect 12256 14952 12308 14958
rect 12360 14929 12388 16351
rect 12438 15736 12494 15745
rect 12438 15671 12494 15680
rect 12256 14894 12308 14900
rect 12346 14920 12402 14929
rect 12346 14855 12402 14864
rect 12256 14816 12308 14822
rect 12256 14758 12308 14764
rect 12268 13870 12296 14758
rect 12256 13864 12308 13870
rect 12256 13806 12308 13812
rect 12452 13258 12480 15671
rect 12544 14929 12572 16390
rect 12636 16153 12664 17614
rect 12900 17264 12952 17270
rect 12900 17206 12952 17212
rect 12716 16720 12768 16726
rect 12714 16688 12716 16697
rect 12768 16688 12770 16697
rect 12912 16658 12940 17206
rect 12992 16788 13044 16794
rect 12992 16730 13044 16736
rect 12714 16623 12770 16632
rect 12900 16652 12952 16658
rect 12900 16594 12952 16600
rect 12716 16584 12768 16590
rect 12716 16526 12768 16532
rect 12808 16584 12860 16590
rect 12860 16532 12940 16538
rect 12808 16526 12940 16532
rect 12728 16250 12756 16526
rect 12820 16510 12940 16526
rect 12716 16244 12768 16250
rect 12768 16204 12848 16232
rect 12716 16186 12768 16192
rect 12622 16144 12678 16153
rect 12622 16079 12678 16088
rect 12716 15360 12768 15366
rect 12716 15302 12768 15308
rect 12530 14920 12586 14929
rect 12530 14855 12586 14864
rect 12624 14884 12676 14890
rect 12624 14826 12676 14832
rect 12532 14816 12584 14822
rect 12532 14758 12584 14764
rect 12544 14074 12572 14758
rect 12636 14618 12664 14826
rect 12624 14612 12676 14618
rect 12624 14554 12676 14560
rect 12636 14414 12664 14554
rect 12624 14408 12676 14414
rect 12624 14350 12676 14356
rect 12728 14074 12756 15302
rect 12820 14958 12848 16204
rect 12912 15910 12940 16510
rect 13004 16454 13032 16730
rect 12992 16448 13044 16454
rect 12992 16390 13044 16396
rect 12900 15904 12952 15910
rect 12900 15846 12952 15852
rect 12900 15700 12952 15706
rect 12900 15642 12952 15648
rect 12912 15201 12940 15642
rect 12898 15192 12954 15201
rect 13096 15162 13124 17711
rect 13176 16992 13228 16998
rect 13176 16934 13228 16940
rect 13188 16697 13216 16934
rect 13174 16688 13230 16697
rect 13174 16623 13230 16632
rect 13280 16522 13308 18566
rect 13464 17814 13492 18634
rect 13648 18426 13676 20431
rect 14200 20330 14228 22200
rect 14462 21448 14518 21457
rect 14462 21383 14518 21392
rect 14280 21208 14332 21214
rect 14280 21150 14332 21156
rect 14188 20324 14240 20330
rect 14188 20266 14240 20272
rect 13820 20256 13872 20262
rect 13820 20198 13872 20204
rect 13832 19718 13860 20198
rect 13945 20156 14253 20165
rect 13945 20154 13951 20156
rect 14007 20154 14031 20156
rect 14087 20154 14111 20156
rect 14167 20154 14191 20156
rect 14247 20154 14253 20156
rect 14007 20102 14009 20154
rect 14189 20102 14191 20154
rect 13945 20100 13951 20102
rect 14007 20100 14031 20102
rect 14087 20100 14111 20102
rect 14167 20100 14191 20102
rect 14247 20100 14253 20102
rect 13945 20091 14253 20100
rect 14188 19848 14240 19854
rect 14188 19790 14240 19796
rect 14292 19802 14320 21150
rect 14372 20460 14424 20466
rect 14372 20402 14424 20408
rect 14384 19990 14412 20402
rect 14372 19984 14424 19990
rect 14372 19926 14424 19932
rect 13820 19712 13872 19718
rect 13820 19654 13872 19660
rect 13912 19712 13964 19718
rect 13912 19654 13964 19660
rect 13728 18624 13780 18630
rect 13728 18566 13780 18572
rect 13636 18420 13688 18426
rect 13636 18362 13688 18368
rect 13636 18148 13688 18154
rect 13636 18090 13688 18096
rect 13452 17808 13504 17814
rect 13452 17750 13504 17756
rect 13452 17672 13504 17678
rect 13452 17614 13504 17620
rect 13360 17536 13412 17542
rect 13360 17478 13412 17484
rect 13372 16590 13400 17478
rect 13464 17202 13492 17614
rect 13648 17338 13676 18090
rect 13740 17921 13768 18566
rect 13726 17912 13782 17921
rect 13726 17847 13782 17856
rect 13832 17728 13860 19654
rect 13924 19446 13952 19654
rect 14200 19514 14228 19790
rect 14292 19774 14412 19802
rect 14188 19508 14240 19514
rect 14188 19450 14240 19456
rect 13912 19440 13964 19446
rect 13912 19382 13964 19388
rect 14096 19372 14148 19378
rect 14148 19332 14320 19360
rect 14096 19314 14148 19320
rect 13945 19068 14253 19077
rect 13945 19066 13951 19068
rect 14007 19066 14031 19068
rect 14087 19066 14111 19068
rect 14167 19066 14191 19068
rect 14247 19066 14253 19068
rect 14007 19014 14009 19066
rect 14189 19014 14191 19066
rect 13945 19012 13951 19014
rect 14007 19012 14031 19014
rect 14087 19012 14111 19014
rect 14167 19012 14191 19014
rect 14247 19012 14253 19014
rect 13945 19003 14253 19012
rect 14292 18630 14320 19332
rect 14280 18624 14332 18630
rect 14280 18566 14332 18572
rect 14292 18358 14320 18566
rect 14280 18352 14332 18358
rect 14280 18294 14332 18300
rect 13945 17980 14253 17989
rect 13945 17978 13951 17980
rect 14007 17978 14031 17980
rect 14087 17978 14111 17980
rect 14167 17978 14191 17980
rect 14247 17978 14253 17980
rect 14007 17926 14009 17978
rect 14189 17926 14191 17978
rect 13945 17924 13951 17926
rect 14007 17924 14031 17926
rect 14087 17924 14111 17926
rect 14167 17924 14191 17926
rect 14247 17924 14253 17926
rect 13945 17915 14253 17924
rect 14280 17740 14332 17746
rect 13832 17700 13952 17728
rect 13818 17640 13874 17649
rect 13818 17575 13820 17584
rect 13872 17575 13874 17584
rect 13820 17546 13872 17552
rect 13636 17332 13688 17338
rect 13636 17274 13688 17280
rect 13452 17196 13504 17202
rect 13452 17138 13504 17144
rect 13360 16584 13412 16590
rect 13360 16526 13412 16532
rect 13268 16516 13320 16522
rect 13268 16458 13320 16464
rect 13176 16448 13228 16454
rect 13176 16390 13228 16396
rect 13188 16114 13216 16390
rect 13372 16182 13400 16526
rect 13360 16176 13412 16182
rect 13360 16118 13412 16124
rect 13176 16108 13228 16114
rect 13176 16050 13228 16056
rect 13452 15904 13504 15910
rect 13452 15846 13504 15852
rect 13268 15564 13320 15570
rect 13268 15506 13320 15512
rect 13176 15496 13228 15502
rect 13176 15438 13228 15444
rect 12898 15127 12954 15136
rect 13084 15156 13136 15162
rect 13084 15098 13136 15104
rect 12808 14952 12860 14958
rect 12808 14894 12860 14900
rect 12898 14920 12954 14929
rect 12820 14346 12848 14894
rect 12898 14855 12954 14864
rect 12808 14340 12860 14346
rect 12808 14282 12860 14288
rect 12532 14068 12584 14074
rect 12532 14010 12584 14016
rect 12716 14068 12768 14074
rect 12716 14010 12768 14016
rect 12532 13932 12584 13938
rect 12532 13874 12584 13880
rect 12440 13252 12492 13258
rect 12440 13194 12492 13200
rect 12256 13184 12308 13190
rect 12256 13126 12308 13132
rect 12162 11928 12218 11937
rect 12268 11898 12296 13126
rect 12348 12096 12400 12102
rect 12348 12038 12400 12044
rect 12162 11863 12218 11872
rect 12256 11892 12308 11898
rect 12256 11834 12308 11840
rect 12360 11830 12388 12038
rect 12438 11928 12494 11937
rect 12438 11863 12494 11872
rect 12348 11824 12400 11830
rect 12348 11766 12400 11772
rect 12072 11688 12124 11694
rect 12072 11630 12124 11636
rect 12084 11354 12112 11630
rect 12348 11552 12400 11558
rect 12348 11494 12400 11500
rect 12072 11348 12124 11354
rect 12124 11308 12204 11336
rect 12072 11290 12124 11296
rect 11980 11280 12032 11286
rect 11980 11222 12032 11228
rect 12070 11248 12126 11257
rect 12176 11234 12204 11308
rect 12176 11206 12296 11234
rect 12070 11183 12126 11192
rect 11980 11008 12032 11014
rect 11980 10950 12032 10956
rect 11992 10810 12020 10950
rect 11980 10804 12032 10810
rect 11980 10746 12032 10752
rect 11980 10668 12032 10674
rect 11980 10610 12032 10616
rect 11992 9761 12020 10610
rect 12084 10130 12112 11183
rect 12164 11076 12216 11082
rect 12164 11018 12216 11024
rect 12072 10124 12124 10130
rect 12072 10066 12124 10072
rect 12072 9920 12124 9926
rect 12072 9862 12124 9868
rect 11978 9752 12034 9761
rect 11978 9687 12034 9696
rect 11978 9616 12034 9625
rect 11978 9551 12034 9560
rect 11992 7410 12020 9551
rect 12084 7528 12112 9862
rect 12176 7834 12204 11018
rect 12268 7993 12296 11206
rect 12360 11014 12388 11494
rect 12348 11008 12400 11014
rect 12348 10950 12400 10956
rect 12452 10690 12480 11863
rect 12544 11234 12572 13874
rect 12820 13870 12848 14282
rect 12808 13864 12860 13870
rect 12808 13806 12860 13812
rect 12716 13728 12768 13734
rect 12716 13670 12768 13676
rect 12622 13424 12678 13433
rect 12622 13359 12624 13368
rect 12676 13359 12678 13368
rect 12624 13330 12676 13336
rect 12624 13252 12676 13258
rect 12624 13194 12676 13200
rect 12636 12617 12664 13194
rect 12622 12608 12678 12617
rect 12622 12543 12678 12552
rect 12728 12209 12756 13670
rect 12808 13184 12860 13190
rect 12808 13126 12860 13132
rect 12820 12889 12848 13126
rect 12806 12880 12862 12889
rect 12806 12815 12862 12824
rect 12808 12436 12860 12442
rect 12808 12378 12860 12384
rect 12820 12238 12848 12378
rect 12808 12232 12860 12238
rect 12714 12200 12770 12209
rect 12808 12174 12860 12180
rect 12714 12135 12770 12144
rect 12728 11898 12756 12135
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 12714 11792 12770 11801
rect 12714 11727 12716 11736
rect 12768 11727 12770 11736
rect 12716 11698 12768 11704
rect 12808 11552 12860 11558
rect 12912 11540 12940 14855
rect 13096 13326 13124 15098
rect 13188 14929 13216 15438
rect 13174 14920 13230 14929
rect 13174 14855 13230 14864
rect 13280 14618 13308 15506
rect 13360 15360 13412 15366
rect 13360 15302 13412 15308
rect 13372 15162 13400 15302
rect 13360 15156 13412 15162
rect 13360 15098 13412 15104
rect 13360 15020 13412 15026
rect 13360 14962 13412 14968
rect 13268 14612 13320 14618
rect 13268 14554 13320 14560
rect 13372 14498 13400 14962
rect 13188 14470 13400 14498
rect 13084 13320 13136 13326
rect 13084 13262 13136 13268
rect 13188 13172 13216 14470
rect 13464 14396 13492 15846
rect 13372 14368 13492 14396
rect 13268 13864 13320 13870
rect 13268 13806 13320 13812
rect 13004 13144 13216 13172
rect 13004 11642 13032 13144
rect 13280 12918 13308 13806
rect 13372 13734 13400 14368
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 13464 13841 13492 14214
rect 13544 13932 13596 13938
rect 13544 13874 13596 13880
rect 13450 13832 13506 13841
rect 13450 13767 13506 13776
rect 13556 13734 13584 13874
rect 13360 13728 13412 13734
rect 13544 13728 13596 13734
rect 13360 13670 13412 13676
rect 13542 13696 13544 13705
rect 13596 13696 13598 13705
rect 13542 13631 13598 13640
rect 13648 13410 13676 17274
rect 13728 16992 13780 16998
rect 13726 16960 13728 16969
rect 13924 16980 13952 17700
rect 14280 17682 14332 17688
rect 13780 16960 13782 16969
rect 13726 16895 13782 16904
rect 13832 16952 13952 16980
rect 13832 15502 13860 16952
rect 13945 16892 14253 16901
rect 13945 16890 13951 16892
rect 14007 16890 14031 16892
rect 14087 16890 14111 16892
rect 14167 16890 14191 16892
rect 14247 16890 14253 16892
rect 14007 16838 14009 16890
rect 14189 16838 14191 16890
rect 13945 16836 13951 16838
rect 14007 16836 14031 16838
rect 14087 16836 14111 16838
rect 14167 16836 14191 16838
rect 14247 16836 14253 16838
rect 13945 16827 14253 16836
rect 14292 16794 14320 17682
rect 14280 16788 14332 16794
rect 14280 16730 14332 16736
rect 14292 16182 14320 16730
rect 14280 16176 14332 16182
rect 14280 16118 14332 16124
rect 13945 15804 14253 15813
rect 13945 15802 13951 15804
rect 14007 15802 14031 15804
rect 14087 15802 14111 15804
rect 14167 15802 14191 15804
rect 14247 15802 14253 15804
rect 14007 15750 14009 15802
rect 14189 15750 14191 15802
rect 13945 15748 13951 15750
rect 14007 15748 14031 15750
rect 14087 15748 14111 15750
rect 14167 15748 14191 15750
rect 14247 15748 14253 15750
rect 13945 15739 14253 15748
rect 13820 15496 13872 15502
rect 13820 15438 13872 15444
rect 13912 15428 13964 15434
rect 13912 15370 13964 15376
rect 13728 15360 13780 15366
rect 13728 15302 13780 15308
rect 13740 14657 13768 15302
rect 13924 15162 13952 15370
rect 14186 15192 14242 15201
rect 13912 15156 13964 15162
rect 14186 15127 14242 15136
rect 13912 15098 13964 15104
rect 14200 15094 14228 15127
rect 14188 15088 14240 15094
rect 14188 15030 14240 15036
rect 14280 15020 14332 15026
rect 14280 14962 14332 14968
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13726 14648 13782 14657
rect 13726 14583 13782 14592
rect 13832 14414 13860 14758
rect 13945 14716 14253 14725
rect 13945 14714 13951 14716
rect 14007 14714 14031 14716
rect 14087 14714 14111 14716
rect 14167 14714 14191 14716
rect 14247 14714 14253 14716
rect 14007 14662 14009 14714
rect 14189 14662 14191 14714
rect 13945 14660 13951 14662
rect 14007 14660 14031 14662
rect 14087 14660 14111 14662
rect 14167 14660 14191 14662
rect 14247 14660 14253 14662
rect 13945 14651 14253 14660
rect 14002 14512 14058 14521
rect 14002 14447 14058 14456
rect 13820 14408 13872 14414
rect 13820 14350 13872 14356
rect 14016 13870 14044 14447
rect 14096 14272 14148 14278
rect 14096 14214 14148 14220
rect 14108 13938 14136 14214
rect 14292 14074 14320 14962
rect 14280 14068 14332 14074
rect 14280 14010 14332 14016
rect 14278 13968 14334 13977
rect 14096 13932 14148 13938
rect 14278 13903 14334 13912
rect 14096 13874 14148 13880
rect 14004 13864 14056 13870
rect 13726 13832 13782 13841
rect 14004 13806 14056 13812
rect 13726 13767 13782 13776
rect 13740 13530 13768 13767
rect 13945 13628 14253 13637
rect 13945 13626 13951 13628
rect 14007 13626 14031 13628
rect 14087 13626 14111 13628
rect 14167 13626 14191 13628
rect 14247 13626 14253 13628
rect 14007 13574 14009 13626
rect 14189 13574 14191 13626
rect 13945 13572 13951 13574
rect 14007 13572 14031 13574
rect 14087 13572 14111 13574
rect 14167 13572 14191 13574
rect 14247 13572 14253 13574
rect 13945 13563 14253 13572
rect 13728 13524 13780 13530
rect 14292 13512 14320 13903
rect 14384 13530 14412 19774
rect 14476 15178 14504 21383
rect 14568 20602 14596 22200
rect 14648 21276 14700 21282
rect 14648 21218 14700 21224
rect 14556 20596 14608 20602
rect 14556 20538 14608 20544
rect 14660 20482 14688 21218
rect 14936 20584 14964 22200
rect 15200 20596 15252 20602
rect 14936 20556 15200 20584
rect 15304 20584 15332 22200
rect 15384 20596 15436 20602
rect 15304 20556 15384 20584
rect 15200 20538 15252 20544
rect 15672 20584 15700 22200
rect 15936 21140 15988 21146
rect 15936 21082 15988 21088
rect 15752 20596 15804 20602
rect 15672 20556 15752 20584
rect 15384 20538 15436 20544
rect 15752 20538 15804 20544
rect 14568 20454 14688 20482
rect 14740 20460 14792 20466
rect 14568 16096 14596 20454
rect 14740 20402 14792 20408
rect 15476 20460 15528 20466
rect 15476 20402 15528 20408
rect 15844 20460 15896 20466
rect 15844 20402 15896 20408
rect 14752 19514 14780 20402
rect 15200 19712 15252 19718
rect 15200 19654 15252 19660
rect 14740 19508 14792 19514
rect 14740 19450 14792 19456
rect 15016 18760 15068 18766
rect 15016 18702 15068 18708
rect 15108 18760 15160 18766
rect 15108 18702 15160 18708
rect 14648 18624 14700 18630
rect 14648 18566 14700 18572
rect 14660 18426 14688 18566
rect 14648 18420 14700 18426
rect 14648 18362 14700 18368
rect 14924 18216 14976 18222
rect 14924 18158 14976 18164
rect 14936 17762 14964 18158
rect 15028 17882 15056 18702
rect 15120 17921 15148 18702
rect 15106 17912 15162 17921
rect 15016 17876 15068 17882
rect 15106 17847 15162 17856
rect 15016 17818 15068 17824
rect 14936 17734 15148 17762
rect 15120 17542 15148 17734
rect 15212 17678 15240 19654
rect 15488 18970 15516 20402
rect 15568 20392 15620 20398
rect 15568 20334 15620 20340
rect 15580 20058 15608 20334
rect 15660 20256 15712 20262
rect 15660 20198 15712 20204
rect 15568 20052 15620 20058
rect 15568 19994 15620 20000
rect 15672 19854 15700 20198
rect 15856 19990 15884 20402
rect 15844 19984 15896 19990
rect 15844 19926 15896 19932
rect 15752 19916 15804 19922
rect 15752 19858 15804 19864
rect 15660 19848 15712 19854
rect 15660 19790 15712 19796
rect 15764 19378 15792 19858
rect 15844 19508 15896 19514
rect 15844 19450 15896 19456
rect 15752 19372 15804 19378
rect 15752 19314 15804 19320
rect 15660 19168 15712 19174
rect 15660 19110 15712 19116
rect 15476 18964 15528 18970
rect 15476 18906 15528 18912
rect 15568 18760 15620 18766
rect 15566 18728 15568 18737
rect 15620 18728 15622 18737
rect 15566 18663 15622 18672
rect 15672 18630 15700 19110
rect 15660 18624 15712 18630
rect 15660 18566 15712 18572
rect 15382 18456 15438 18465
rect 15382 18391 15384 18400
rect 15436 18391 15438 18400
rect 15384 18362 15436 18368
rect 15476 18284 15528 18290
rect 15476 18226 15528 18232
rect 15292 18080 15344 18086
rect 15292 18022 15344 18028
rect 15304 17785 15332 18022
rect 15290 17776 15346 17785
rect 15290 17711 15346 17720
rect 15200 17672 15252 17678
rect 15200 17614 15252 17620
rect 14924 17536 14976 17542
rect 14924 17478 14976 17484
rect 15108 17536 15160 17542
rect 15108 17478 15160 17484
rect 14936 17338 14964 17478
rect 14924 17332 14976 17338
rect 14924 17274 14976 17280
rect 15016 17332 15068 17338
rect 15016 17274 15068 17280
rect 15028 17134 15056 17274
rect 15120 17202 15148 17478
rect 15304 17354 15332 17711
rect 15212 17326 15332 17354
rect 15212 17241 15240 17326
rect 15198 17232 15254 17241
rect 15108 17196 15160 17202
rect 15198 17167 15254 17176
rect 15292 17196 15344 17202
rect 15108 17138 15160 17144
rect 15292 17138 15344 17144
rect 15016 17128 15068 17134
rect 15016 17070 15068 17076
rect 15120 16998 15148 17138
rect 15200 17060 15252 17066
rect 15200 17002 15252 17008
rect 15108 16992 15160 16998
rect 14936 16952 15108 16980
rect 14568 16068 14688 16096
rect 14476 15150 14596 15178
rect 14464 14816 14516 14822
rect 14464 14758 14516 14764
rect 13728 13466 13780 13472
rect 14016 13484 14320 13512
rect 14372 13524 14424 13530
rect 13648 13382 13768 13410
rect 13636 13252 13688 13258
rect 13636 13194 13688 13200
rect 13360 13184 13412 13190
rect 13360 13126 13412 13132
rect 13544 13184 13596 13190
rect 13544 13126 13596 13132
rect 13268 12912 13320 12918
rect 13372 12889 13400 13126
rect 13452 12912 13504 12918
rect 13268 12854 13320 12860
rect 13358 12880 13414 12889
rect 13176 12844 13228 12850
rect 13452 12854 13504 12860
rect 13358 12815 13414 12824
rect 13176 12786 13228 12792
rect 13084 12776 13136 12782
rect 13084 12718 13136 12724
rect 13096 12306 13124 12718
rect 13084 12300 13136 12306
rect 13084 12242 13136 12248
rect 13188 11762 13216 12786
rect 13266 12448 13322 12457
rect 13322 12406 13400 12434
rect 13266 12383 13322 12392
rect 13372 12238 13400 12406
rect 13464 12345 13492 12854
rect 13556 12753 13584 13126
rect 13648 13025 13676 13194
rect 13634 13016 13690 13025
rect 13634 12951 13690 12960
rect 13740 12782 13768 13382
rect 13728 12776 13780 12782
rect 13542 12744 13598 12753
rect 13728 12718 13780 12724
rect 13542 12679 13598 12688
rect 14016 12646 14044 13484
rect 14372 13466 14424 13472
rect 14476 13394 14504 14758
rect 14568 14278 14596 15150
rect 14556 14272 14608 14278
rect 14556 14214 14608 14220
rect 14556 14068 14608 14074
rect 14556 14010 14608 14016
rect 14464 13388 14516 13394
rect 14464 13330 14516 13336
rect 14568 13274 14596 14010
rect 14476 13246 14596 13274
rect 14660 13258 14688 16068
rect 14936 16046 14964 16952
rect 15108 16934 15160 16940
rect 15212 16590 15240 17002
rect 15304 16794 15332 17138
rect 15384 17128 15436 17134
rect 15384 17070 15436 17076
rect 15292 16788 15344 16794
rect 15292 16730 15344 16736
rect 15200 16584 15252 16590
rect 15200 16526 15252 16532
rect 15396 16250 15424 17070
rect 15488 16454 15516 18226
rect 15568 18080 15620 18086
rect 15566 18048 15568 18057
rect 15620 18048 15622 18057
rect 15566 17983 15622 17992
rect 15672 17678 15700 18566
rect 15764 17882 15792 19314
rect 15752 17876 15804 17882
rect 15752 17818 15804 17824
rect 15660 17672 15712 17678
rect 15660 17614 15712 17620
rect 15672 16726 15700 17614
rect 15752 17604 15804 17610
rect 15752 17546 15804 17552
rect 15764 17066 15792 17546
rect 15752 17060 15804 17066
rect 15752 17002 15804 17008
rect 15660 16720 15712 16726
rect 15660 16662 15712 16668
rect 15476 16448 15528 16454
rect 15476 16390 15528 16396
rect 15384 16244 15436 16250
rect 15384 16186 15436 16192
rect 15752 16244 15804 16250
rect 15752 16186 15804 16192
rect 15108 16108 15160 16114
rect 15108 16050 15160 16056
rect 14924 16040 14976 16046
rect 14924 15982 14976 15988
rect 15016 16040 15068 16046
rect 15016 15982 15068 15988
rect 14924 15632 14976 15638
rect 14924 15574 14976 15580
rect 14832 15020 14884 15026
rect 14832 14962 14884 14968
rect 14740 13864 14792 13870
rect 14740 13806 14792 13812
rect 14752 13326 14780 13806
rect 14740 13320 14792 13326
rect 14740 13262 14792 13268
rect 14648 13252 14700 13258
rect 14188 13184 14240 13190
rect 14094 13152 14150 13161
rect 14188 13126 14240 13132
rect 14094 13087 14150 13096
rect 14108 12986 14136 13087
rect 14096 12980 14148 12986
rect 14096 12922 14148 12928
rect 14200 12889 14228 13126
rect 14186 12880 14242 12889
rect 14186 12815 14242 12824
rect 14372 12844 14424 12850
rect 14372 12786 14424 12792
rect 14280 12776 14332 12782
rect 14384 12753 14412 12786
rect 14280 12718 14332 12724
rect 14370 12744 14426 12753
rect 13544 12640 13596 12646
rect 13544 12582 13596 12588
rect 13728 12640 13780 12646
rect 13728 12582 13780 12588
rect 13820 12640 13872 12646
rect 13820 12582 13872 12588
rect 14004 12640 14056 12646
rect 14004 12582 14056 12588
rect 13450 12336 13506 12345
rect 13450 12271 13506 12280
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 13452 12096 13504 12102
rect 13452 12038 13504 12044
rect 13464 11898 13492 12038
rect 13268 11892 13320 11898
rect 13268 11834 13320 11840
rect 13452 11892 13504 11898
rect 13452 11834 13504 11840
rect 13176 11756 13228 11762
rect 13176 11698 13228 11704
rect 13004 11614 13216 11642
rect 12912 11512 13124 11540
rect 12808 11494 12860 11500
rect 12544 11206 12756 11234
rect 12360 10662 12480 10690
rect 12360 8344 12388 10662
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12452 10130 12480 10406
rect 12440 10124 12492 10130
rect 12440 10066 12492 10072
rect 12452 9586 12480 10066
rect 12532 9716 12584 9722
rect 12532 9658 12584 9664
rect 12544 9625 12572 9658
rect 12530 9616 12586 9625
rect 12440 9580 12492 9586
rect 12530 9551 12586 9560
rect 12440 9522 12492 9528
rect 12624 9512 12676 9518
rect 12438 9480 12494 9489
rect 12624 9454 12676 9460
rect 12438 9415 12494 9424
rect 12452 9058 12480 9415
rect 12530 9072 12586 9081
rect 12452 9030 12530 9058
rect 12530 9007 12586 9016
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 12360 8316 12480 8344
rect 12452 8090 12480 8316
rect 12440 8084 12492 8090
rect 12440 8026 12492 8032
rect 12254 7984 12310 7993
rect 12254 7919 12310 7928
rect 12544 7886 12572 8774
rect 12636 8498 12664 9454
rect 12728 8537 12756 11206
rect 12820 11150 12848 11494
rect 12808 11144 12860 11150
rect 12808 11086 12860 11092
rect 12808 11008 12860 11014
rect 12808 10950 12860 10956
rect 12900 11008 12952 11014
rect 12900 10950 12952 10956
rect 12820 10062 12848 10950
rect 12912 10130 12940 10950
rect 12990 10568 13046 10577
rect 12990 10503 13046 10512
rect 12900 10124 12952 10130
rect 12900 10066 12952 10072
rect 12808 10056 12860 10062
rect 12808 9998 12860 10004
rect 13004 9654 13032 10503
rect 12992 9648 13044 9654
rect 12992 9590 13044 9596
rect 12820 9438 13032 9466
rect 12820 9382 12848 9438
rect 12808 9376 12860 9382
rect 12808 9318 12860 9324
rect 12900 9376 12952 9382
rect 12900 9318 12952 9324
rect 12912 8974 12940 9318
rect 12900 8968 12952 8974
rect 12900 8910 12952 8916
rect 12808 8900 12860 8906
rect 12808 8842 12860 8848
rect 12714 8528 12770 8537
rect 12624 8492 12676 8498
rect 12820 8498 12848 8842
rect 12900 8832 12952 8838
rect 12900 8774 12952 8780
rect 12912 8634 12940 8774
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 13004 8514 13032 9438
rect 12714 8463 12770 8472
rect 12808 8492 12860 8498
rect 12624 8434 12676 8440
rect 12808 8434 12860 8440
rect 12912 8486 13032 8514
rect 12636 8022 12664 8434
rect 12912 8362 12940 8486
rect 12992 8424 13044 8430
rect 12992 8366 13044 8372
rect 12900 8356 12952 8362
rect 12900 8298 12952 8304
rect 12714 8120 12770 8129
rect 12714 8055 12770 8064
rect 12624 8016 12676 8022
rect 12624 7958 12676 7964
rect 12532 7880 12584 7886
rect 12176 7806 12480 7834
rect 12532 7822 12584 7828
rect 12256 7744 12308 7750
rect 12256 7686 12308 7692
rect 12084 7500 12204 7528
rect 11980 7404 12032 7410
rect 11980 7346 12032 7352
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 11978 7032 12034 7041
rect 11978 6967 12034 6976
rect 11992 6934 12020 6967
rect 11980 6928 12032 6934
rect 11980 6870 12032 6876
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 11980 6248 12032 6254
rect 11886 6216 11942 6225
rect 11980 6190 12032 6196
rect 11886 6151 11942 6160
rect 11900 5953 11928 6151
rect 11886 5944 11942 5953
rect 11886 5879 11942 5888
rect 11900 5370 11928 5879
rect 11992 5817 12020 6190
rect 11978 5808 12034 5817
rect 11978 5743 12034 5752
rect 11980 5636 12032 5642
rect 11980 5578 12032 5584
rect 11888 5364 11940 5370
rect 11888 5306 11940 5312
rect 11992 5234 12020 5578
rect 11888 5228 11940 5234
rect 11888 5170 11940 5176
rect 11980 5228 12032 5234
rect 11980 5170 12032 5176
rect 11900 5030 11928 5170
rect 11888 5024 11940 5030
rect 11888 4966 11940 4972
rect 11900 4185 11928 4966
rect 11992 4690 12020 5170
rect 11980 4684 12032 4690
rect 11980 4626 12032 4632
rect 11980 4480 12032 4486
rect 11978 4448 11980 4457
rect 12032 4448 12034 4457
rect 11978 4383 12034 4392
rect 11978 4312 12034 4321
rect 11978 4247 11980 4256
rect 12032 4247 12034 4256
rect 11980 4218 12032 4224
rect 11886 4176 11942 4185
rect 11886 4111 11942 4120
rect 11888 3040 11940 3042
rect 11992 3040 12020 4218
rect 12084 4146 12112 7346
rect 12176 7313 12204 7500
rect 12268 7410 12296 7686
rect 12256 7404 12308 7410
rect 12256 7346 12308 7352
rect 12162 7304 12218 7313
rect 12162 7239 12218 7248
rect 12256 7200 12308 7206
rect 12256 7142 12308 7148
rect 12164 6860 12216 6866
rect 12164 6802 12216 6808
rect 12176 5710 12204 6802
rect 12164 5704 12216 5710
rect 12164 5646 12216 5652
rect 12164 5568 12216 5574
rect 12164 5510 12216 5516
rect 12176 5370 12204 5510
rect 12268 5370 12296 7142
rect 12348 6724 12400 6730
rect 12348 6666 12400 6672
rect 12164 5364 12216 5370
rect 12164 5306 12216 5312
rect 12256 5364 12308 5370
rect 12256 5306 12308 5312
rect 12256 5228 12308 5234
rect 12256 5170 12308 5176
rect 12072 4140 12124 4146
rect 12072 4082 12124 4088
rect 12072 3936 12124 3942
rect 12072 3878 12124 3884
rect 11888 3036 12020 3040
rect 11940 3012 12020 3036
rect 11888 2978 11940 2984
rect 11808 2746 11928 2774
rect 11900 2446 11928 2746
rect 12084 2514 12112 3878
rect 12164 3732 12216 3738
rect 12164 3674 12216 3680
rect 12072 2508 12124 2514
rect 12072 2450 12124 2456
rect 11704 2440 11756 2446
rect 11704 2382 11756 2388
rect 11888 2440 11940 2446
rect 11888 2382 11940 2388
rect 11346 2204 11654 2213
rect 11346 2202 11352 2204
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11648 2202 11654 2204
rect 11408 2150 11410 2202
rect 11590 2150 11592 2202
rect 11346 2148 11352 2150
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11648 2148 11654 2150
rect 11346 2139 11654 2148
rect 11060 2100 11112 2106
rect 11060 2042 11112 2048
rect 10966 2000 11022 2009
rect 10966 1935 11022 1944
rect 10784 1896 10836 1902
rect 10784 1838 10836 1844
rect 11072 800 11100 2042
rect 11242 1184 11298 1193
rect 11242 1119 11298 1128
rect 11256 921 11284 1119
rect 11242 912 11298 921
rect 11242 847 11298 856
rect 11440 870 11560 898
rect 11440 800 11468 870
rect 7852 734 8064 762
rect 8114 0 8170 800
rect 8482 0 8538 800
rect 8850 0 8906 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 9954 0 10010 800
rect 10322 0 10378 800
rect 10690 0 10746 800
rect 11058 0 11114 800
rect 11426 0 11482 800
rect 11532 762 11560 870
rect 11716 762 11744 2382
rect 11900 1714 11928 2382
rect 12072 2304 12124 2310
rect 12072 2246 12124 2252
rect 12084 1737 12112 2246
rect 11808 1686 11928 1714
rect 12070 1728 12126 1737
rect 11808 800 11836 1686
rect 12070 1663 12126 1672
rect 12176 800 12204 3674
rect 12268 2038 12296 5170
rect 12360 5030 12388 6666
rect 12452 6610 12480 7806
rect 12624 7812 12676 7818
rect 12624 7754 12676 7760
rect 12636 7342 12664 7754
rect 12728 7410 12756 8055
rect 13004 7886 13032 8366
rect 12992 7880 13044 7886
rect 12992 7822 13044 7828
rect 12808 7812 12860 7818
rect 12808 7754 12860 7760
rect 12716 7404 12768 7410
rect 12716 7346 12768 7352
rect 12624 7336 12676 7342
rect 12624 7278 12676 7284
rect 12636 6866 12664 7278
rect 12820 7177 12848 7754
rect 12992 7744 13044 7750
rect 12992 7686 13044 7692
rect 13004 7546 13032 7686
rect 12992 7540 13044 7546
rect 12992 7482 13044 7488
rect 12992 7200 13044 7206
rect 12806 7168 12862 7177
rect 12992 7142 13044 7148
rect 12806 7103 12862 7112
rect 12806 7032 12862 7041
rect 12806 6967 12808 6976
rect 12860 6967 12862 6976
rect 12808 6938 12860 6944
rect 12624 6860 12676 6866
rect 12624 6802 12676 6808
rect 12452 6582 12572 6610
rect 12440 6452 12492 6458
rect 12440 6394 12492 6400
rect 12348 5024 12400 5030
rect 12348 4966 12400 4972
rect 12452 4826 12480 6394
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 12438 4720 12494 4729
rect 12438 4655 12494 4664
rect 12452 4214 12480 4655
rect 12544 4554 12572 6582
rect 12636 5692 12664 6802
rect 12820 5760 12848 6938
rect 13004 6633 13032 7142
rect 13096 6866 13124 11512
rect 13188 7018 13216 11614
rect 13280 11354 13308 11834
rect 13360 11552 13412 11558
rect 13360 11494 13412 11500
rect 13268 11348 13320 11354
rect 13268 11290 13320 11296
rect 13372 11218 13400 11494
rect 13556 11218 13584 12582
rect 13636 12232 13688 12238
rect 13636 12174 13688 12180
rect 13360 11212 13412 11218
rect 13360 11154 13412 11160
rect 13544 11212 13596 11218
rect 13544 11154 13596 11160
rect 13452 11144 13504 11150
rect 13452 11086 13504 11092
rect 13268 11008 13320 11014
rect 13268 10950 13320 10956
rect 13360 11008 13412 11014
rect 13360 10950 13412 10956
rect 13280 10810 13308 10950
rect 13268 10804 13320 10810
rect 13268 10746 13320 10752
rect 13268 10124 13320 10130
rect 13268 10066 13320 10072
rect 13280 9722 13308 10066
rect 13268 9716 13320 9722
rect 13268 9658 13320 9664
rect 13372 9353 13400 10950
rect 13358 9344 13414 9353
rect 13358 9279 13414 9288
rect 13358 9208 13414 9217
rect 13358 9143 13414 9152
rect 13372 9042 13400 9143
rect 13360 9036 13412 9042
rect 13360 8978 13412 8984
rect 13360 8900 13412 8906
rect 13360 8842 13412 8848
rect 13268 8628 13320 8634
rect 13268 8570 13320 8576
rect 13280 8242 13308 8570
rect 13372 8537 13400 8842
rect 13358 8528 13414 8537
rect 13358 8463 13414 8472
rect 13280 8214 13400 8242
rect 13268 8084 13320 8090
rect 13268 8026 13320 8032
rect 13280 7274 13308 8026
rect 13372 7886 13400 8214
rect 13360 7880 13412 7886
rect 13360 7822 13412 7828
rect 13360 7336 13412 7342
rect 13360 7278 13412 7284
rect 13268 7268 13320 7274
rect 13268 7210 13320 7216
rect 13188 6990 13308 7018
rect 13372 7002 13400 7278
rect 13084 6860 13136 6866
rect 13136 6820 13216 6848
rect 13084 6802 13136 6808
rect 13084 6656 13136 6662
rect 12990 6624 13046 6633
rect 13084 6598 13136 6604
rect 12990 6559 13046 6568
rect 12900 6248 12952 6254
rect 12900 6190 12952 6196
rect 12912 6089 12940 6190
rect 12992 6112 13044 6118
rect 12898 6080 12954 6089
rect 12992 6054 13044 6060
rect 12898 6015 12954 6024
rect 12820 5732 12940 5760
rect 12636 5664 12848 5692
rect 12716 5568 12768 5574
rect 12716 5510 12768 5516
rect 12624 5364 12676 5370
rect 12624 5306 12676 5312
rect 12532 4548 12584 4554
rect 12532 4490 12584 4496
rect 12544 4282 12572 4490
rect 12532 4276 12584 4282
rect 12532 4218 12584 4224
rect 12440 4208 12492 4214
rect 12440 4150 12492 4156
rect 12348 3936 12400 3942
rect 12348 3878 12400 3884
rect 12360 3448 12388 3878
rect 12452 3670 12480 4150
rect 12530 3768 12586 3777
rect 12530 3703 12586 3712
rect 12440 3664 12492 3670
rect 12440 3606 12492 3612
rect 12360 3420 12480 3448
rect 12346 3360 12402 3369
rect 12346 3295 12402 3304
rect 12360 3194 12388 3295
rect 12452 3233 12480 3420
rect 12438 3224 12494 3233
rect 12348 3188 12400 3194
rect 12438 3159 12494 3168
rect 12348 3130 12400 3136
rect 12544 3126 12572 3703
rect 12532 3120 12584 3126
rect 12532 3062 12584 3068
rect 12348 3052 12400 3058
rect 12348 2994 12400 3000
rect 12360 2825 12388 2994
rect 12530 2952 12586 2961
rect 12530 2887 12586 2896
rect 12544 2854 12572 2887
rect 12532 2848 12584 2854
rect 12346 2816 12402 2825
rect 12532 2790 12584 2796
rect 12346 2751 12402 2760
rect 12348 2576 12400 2582
rect 12346 2544 12348 2553
rect 12400 2544 12402 2553
rect 12346 2479 12402 2488
rect 12348 2440 12400 2446
rect 12348 2382 12400 2388
rect 12360 2106 12388 2382
rect 12532 2304 12584 2310
rect 12532 2246 12584 2252
rect 12348 2100 12400 2106
rect 12348 2042 12400 2048
rect 12256 2032 12308 2038
rect 12256 1974 12308 1980
rect 12544 800 12572 2246
rect 12636 2038 12664 5306
rect 12728 5234 12756 5510
rect 12716 5228 12768 5234
rect 12716 5170 12768 5176
rect 12714 4720 12770 4729
rect 12714 4655 12716 4664
rect 12768 4655 12770 4664
rect 12716 4626 12768 4632
rect 12716 4548 12768 4554
rect 12716 4490 12768 4496
rect 12728 3097 12756 4490
rect 12714 3088 12770 3097
rect 12714 3023 12770 3032
rect 12820 2990 12848 5664
rect 12912 4622 12940 5732
rect 13004 5273 13032 6054
rect 13096 5817 13124 6598
rect 13082 5808 13138 5817
rect 13188 5778 13216 6820
rect 13082 5743 13138 5752
rect 13176 5772 13228 5778
rect 13096 5710 13124 5743
rect 13176 5714 13228 5720
rect 13084 5704 13136 5710
rect 13280 5658 13308 6990
rect 13360 6996 13412 7002
rect 13360 6938 13412 6944
rect 13360 6656 13412 6662
rect 13360 6598 13412 6604
rect 13084 5646 13136 5652
rect 13188 5630 13308 5658
rect 12990 5264 13046 5273
rect 12990 5199 13046 5208
rect 13084 5228 13136 5234
rect 13084 5170 13136 5176
rect 12990 4856 13046 4865
rect 12990 4791 12992 4800
rect 13044 4791 13046 4800
rect 12992 4762 13044 4768
rect 13096 4758 13124 5170
rect 13084 4752 13136 4758
rect 13084 4694 13136 4700
rect 12992 4684 13044 4690
rect 12992 4626 13044 4632
rect 12900 4616 12952 4622
rect 12900 4558 12952 4564
rect 13004 4078 13032 4626
rect 13084 4616 13136 4622
rect 13188 4604 13216 5630
rect 13372 5545 13400 6598
rect 13358 5536 13414 5545
rect 13358 5471 13414 5480
rect 13464 5114 13492 11086
rect 13556 10742 13584 11154
rect 13544 10736 13596 10742
rect 13544 10678 13596 10684
rect 13648 10554 13676 12174
rect 13740 11830 13768 12582
rect 13832 12442 13860 12582
rect 13945 12540 14253 12549
rect 13945 12538 13951 12540
rect 14007 12538 14031 12540
rect 14087 12538 14111 12540
rect 14167 12538 14191 12540
rect 14247 12538 14253 12540
rect 14007 12486 14009 12538
rect 14189 12486 14191 12538
rect 13945 12484 13951 12486
rect 14007 12484 14031 12486
rect 14087 12484 14111 12486
rect 14167 12484 14191 12486
rect 14247 12484 14253 12486
rect 13945 12475 14253 12484
rect 13820 12436 13872 12442
rect 13820 12378 13872 12384
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 13728 11824 13780 11830
rect 13728 11766 13780 11772
rect 13728 11552 13780 11558
rect 13728 11494 13780 11500
rect 13740 10810 13768 11494
rect 13832 11082 13860 12174
rect 13912 12096 13964 12102
rect 13910 12064 13912 12073
rect 13964 12064 13966 12073
rect 13910 11999 13966 12008
rect 13924 11830 13952 11999
rect 14096 11892 14148 11898
rect 14096 11834 14148 11840
rect 13912 11824 13964 11830
rect 14108 11801 14136 11834
rect 13912 11766 13964 11772
rect 14094 11792 14150 11801
rect 14094 11727 14150 11736
rect 13945 11452 14253 11461
rect 13945 11450 13951 11452
rect 14007 11450 14031 11452
rect 14087 11450 14111 11452
rect 14167 11450 14191 11452
rect 14247 11450 14253 11452
rect 14007 11398 14009 11450
rect 14189 11398 14191 11450
rect 13945 11396 13951 11398
rect 14007 11396 14031 11398
rect 14087 11396 14111 11398
rect 14167 11396 14191 11398
rect 14247 11396 14253 11398
rect 13945 11387 14253 11396
rect 14292 11218 14320 12718
rect 14370 12679 14426 12688
rect 14476 12594 14504 13246
rect 14648 13194 14700 13200
rect 14556 13184 14608 13190
rect 14556 13126 14608 13132
rect 14384 12566 14504 12594
rect 14384 11626 14412 12566
rect 14568 12458 14596 13126
rect 14476 12430 14596 12458
rect 14372 11620 14424 11626
rect 14372 11562 14424 11568
rect 14476 11506 14504 12430
rect 14752 12306 14780 13262
rect 14844 13190 14872 14962
rect 14936 14074 14964 15574
rect 15028 15366 15056 15982
rect 15120 15638 15148 16050
rect 15384 16040 15436 16046
rect 15384 15982 15436 15988
rect 15108 15632 15160 15638
rect 15108 15574 15160 15580
rect 15016 15360 15068 15366
rect 15016 15302 15068 15308
rect 15106 14240 15162 14249
rect 15106 14175 15162 14184
rect 14924 14068 14976 14074
rect 14924 14010 14976 14016
rect 14832 13184 14884 13190
rect 14832 13126 14884 13132
rect 14924 12776 14976 12782
rect 14924 12718 14976 12724
rect 14832 12640 14884 12646
rect 14832 12582 14884 12588
rect 14844 12442 14872 12582
rect 14936 12442 14964 12718
rect 14832 12436 14884 12442
rect 14832 12378 14884 12384
rect 14924 12436 14976 12442
rect 14924 12378 14976 12384
rect 14740 12300 14792 12306
rect 14740 12242 14792 12248
rect 14646 12200 14702 12209
rect 15120 12186 15148 14175
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 15200 13184 15252 13190
rect 15200 13126 15252 13132
rect 15212 12850 15240 13126
rect 15304 12918 15332 13262
rect 15292 12912 15344 12918
rect 15292 12854 15344 12860
rect 15200 12844 15252 12850
rect 15200 12786 15252 12792
rect 15200 12300 15252 12306
rect 15200 12242 15252 12248
rect 14646 12135 14702 12144
rect 14936 12158 15148 12186
rect 14556 12096 14608 12102
rect 14556 12038 14608 12044
rect 14568 11937 14596 12038
rect 14554 11928 14610 11937
rect 14554 11863 14610 11872
rect 14556 11688 14608 11694
rect 14556 11630 14608 11636
rect 14384 11478 14504 11506
rect 14280 11212 14332 11218
rect 14280 11154 14332 11160
rect 13820 11076 13872 11082
rect 13820 11018 13872 11024
rect 14186 10840 14242 10849
rect 13728 10804 13780 10810
rect 14186 10775 14242 10784
rect 13728 10746 13780 10752
rect 14200 10674 14228 10775
rect 14292 10742 14320 11154
rect 14280 10736 14332 10742
rect 14280 10678 14332 10684
rect 14188 10668 14240 10674
rect 14188 10610 14240 10616
rect 13556 10526 13676 10554
rect 13820 10532 13872 10538
rect 13556 9058 13584 10526
rect 13820 10474 13872 10480
rect 13832 10266 13860 10474
rect 13945 10364 14253 10373
rect 13945 10362 13951 10364
rect 14007 10362 14031 10364
rect 14087 10362 14111 10364
rect 14167 10362 14191 10364
rect 14247 10362 14253 10364
rect 14007 10310 14009 10362
rect 14189 10310 14191 10362
rect 13945 10308 13951 10310
rect 14007 10308 14031 10310
rect 14087 10308 14111 10310
rect 14167 10308 14191 10310
rect 14247 10308 14253 10310
rect 13945 10299 14253 10308
rect 14292 10266 14320 10678
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 14280 10260 14332 10266
rect 14280 10202 14332 10208
rect 14004 10192 14056 10198
rect 13818 10160 13874 10169
rect 13818 10095 13874 10104
rect 14002 10160 14004 10169
rect 14056 10160 14058 10169
rect 14002 10095 14058 10104
rect 13636 9988 13688 9994
rect 13636 9930 13688 9936
rect 13648 9897 13676 9930
rect 13728 9920 13780 9926
rect 13634 9888 13690 9897
rect 13728 9862 13780 9868
rect 13634 9823 13690 9832
rect 13740 9761 13768 9862
rect 13726 9752 13782 9761
rect 13726 9687 13782 9696
rect 13636 9648 13688 9654
rect 13636 9590 13688 9596
rect 13648 9178 13676 9590
rect 13728 9580 13780 9586
rect 13728 9522 13780 9528
rect 13636 9172 13688 9178
rect 13636 9114 13688 9120
rect 13556 9030 13676 9058
rect 13544 8832 13596 8838
rect 13544 8774 13596 8780
rect 13556 7410 13584 8774
rect 13648 8566 13676 9030
rect 13740 8906 13768 9522
rect 13832 9160 13860 10095
rect 14280 9376 14332 9382
rect 14280 9318 14332 9324
rect 13945 9276 14253 9285
rect 13945 9274 13951 9276
rect 14007 9274 14031 9276
rect 14087 9274 14111 9276
rect 14167 9274 14191 9276
rect 14247 9274 14253 9276
rect 14007 9222 14009 9274
rect 14189 9222 14191 9274
rect 13945 9220 13951 9222
rect 14007 9220 14031 9222
rect 14087 9220 14111 9222
rect 14167 9220 14191 9222
rect 14247 9220 14253 9222
rect 13945 9211 14253 9220
rect 14096 9172 14148 9178
rect 13832 9132 13952 9160
rect 13820 9036 13872 9042
rect 13820 8978 13872 8984
rect 13728 8900 13780 8906
rect 13728 8842 13780 8848
rect 13832 8634 13860 8978
rect 13820 8628 13872 8634
rect 13820 8570 13872 8576
rect 13636 8560 13688 8566
rect 13636 8502 13688 8508
rect 13648 8430 13676 8502
rect 13636 8424 13688 8430
rect 13636 8366 13688 8372
rect 13820 8288 13872 8294
rect 13924 8276 13952 9132
rect 14096 9114 14148 9120
rect 14108 8974 14136 9114
rect 14096 8968 14148 8974
rect 14096 8910 14148 8916
rect 14004 8560 14056 8566
rect 14004 8502 14056 8508
rect 14094 8528 14150 8537
rect 14016 8362 14044 8502
rect 14094 8463 14096 8472
rect 14148 8463 14150 8472
rect 14096 8434 14148 8440
rect 14186 8392 14242 8401
rect 14004 8356 14056 8362
rect 14186 8327 14188 8336
rect 14004 8298 14056 8304
rect 14240 8327 14242 8336
rect 14188 8298 14240 8304
rect 13872 8248 13952 8276
rect 13820 8230 13872 8236
rect 13728 7948 13780 7954
rect 13728 7890 13780 7896
rect 13636 7744 13688 7750
rect 13636 7686 13688 7692
rect 13648 7546 13676 7686
rect 13636 7540 13688 7546
rect 13636 7482 13688 7488
rect 13544 7404 13596 7410
rect 13544 7346 13596 7352
rect 13634 7304 13690 7313
rect 13544 7268 13596 7274
rect 13740 7274 13768 7890
rect 13832 7585 13860 8230
rect 13945 8188 14253 8197
rect 13945 8186 13951 8188
rect 14007 8186 14031 8188
rect 14087 8186 14111 8188
rect 14167 8186 14191 8188
rect 14247 8186 14253 8188
rect 14007 8134 14009 8186
rect 14189 8134 14191 8186
rect 13945 8132 13951 8134
rect 14007 8132 14031 8134
rect 14087 8132 14111 8134
rect 14167 8132 14191 8134
rect 14247 8132 14253 8134
rect 13945 8123 14253 8132
rect 13912 8084 13964 8090
rect 13912 8026 13964 8032
rect 13818 7576 13874 7585
rect 13818 7511 13874 7520
rect 13924 7460 13952 8026
rect 13832 7432 13952 7460
rect 13634 7239 13690 7248
rect 13728 7268 13780 7274
rect 13544 7210 13596 7216
rect 13556 6730 13584 7210
rect 13544 6724 13596 6730
rect 13544 6666 13596 6672
rect 13648 6662 13676 7239
rect 13728 7210 13780 7216
rect 13832 7041 13860 7432
rect 13945 7100 14253 7109
rect 13945 7098 13951 7100
rect 14007 7098 14031 7100
rect 14087 7098 14111 7100
rect 14167 7098 14191 7100
rect 14247 7098 14253 7100
rect 14007 7046 14009 7098
rect 14189 7046 14191 7098
rect 13945 7044 13951 7046
rect 14007 7044 14031 7046
rect 14087 7044 14111 7046
rect 14167 7044 14191 7046
rect 14247 7044 14253 7046
rect 13818 7032 13874 7041
rect 13945 7035 14253 7044
rect 13818 6967 13874 6976
rect 14292 6882 14320 9318
rect 14384 7818 14412 11478
rect 14464 10804 14516 10810
rect 14464 10746 14516 10752
rect 14476 9178 14504 10746
rect 14568 9994 14596 11630
rect 14660 11257 14688 12135
rect 14832 11552 14884 11558
rect 14752 11512 14832 11540
rect 14646 11248 14702 11257
rect 14646 11183 14702 11192
rect 14648 11076 14700 11082
rect 14648 11018 14700 11024
rect 14660 10742 14688 11018
rect 14648 10736 14700 10742
rect 14648 10678 14700 10684
rect 14660 10606 14688 10678
rect 14648 10600 14700 10606
rect 14648 10542 14700 10548
rect 14556 9988 14608 9994
rect 14556 9930 14608 9936
rect 14554 9888 14610 9897
rect 14554 9823 14610 9832
rect 14464 9172 14516 9178
rect 14464 9114 14516 9120
rect 14462 7984 14518 7993
rect 14462 7919 14518 7928
rect 14476 7886 14504 7919
rect 14464 7880 14516 7886
rect 14464 7822 14516 7828
rect 14372 7812 14424 7818
rect 14372 7754 14424 7760
rect 14476 7002 14504 7822
rect 14568 7546 14596 9823
rect 14648 9376 14700 9382
rect 14646 9344 14648 9353
rect 14700 9344 14702 9353
rect 14646 9279 14702 9288
rect 14660 8129 14688 9279
rect 14752 8786 14780 11512
rect 14832 11494 14884 11500
rect 14832 10600 14884 10606
rect 14832 10542 14884 10548
rect 14844 9625 14872 10542
rect 14830 9616 14886 9625
rect 14830 9551 14886 9560
rect 14936 9518 14964 12158
rect 15016 12096 15068 12102
rect 15016 12038 15068 12044
rect 15106 12064 15162 12073
rect 14924 9512 14976 9518
rect 14924 9454 14976 9460
rect 14752 8758 14872 8786
rect 14738 8664 14794 8673
rect 14738 8599 14794 8608
rect 14752 8430 14780 8599
rect 14740 8424 14792 8430
rect 14740 8366 14792 8372
rect 14844 8294 14872 8758
rect 14936 8498 14964 9454
rect 15028 8945 15056 12038
rect 15106 11999 15162 12008
rect 15120 11898 15148 11999
rect 15212 11898 15240 12242
rect 15108 11892 15160 11898
rect 15108 11834 15160 11840
rect 15200 11892 15252 11898
rect 15200 11834 15252 11840
rect 15198 11792 15254 11801
rect 15198 11727 15254 11736
rect 15212 11642 15240 11727
rect 15120 11614 15240 11642
rect 15120 11370 15148 11614
rect 15200 11552 15252 11558
rect 15198 11520 15200 11529
rect 15252 11520 15254 11529
rect 15198 11455 15254 11464
rect 15120 11342 15240 11370
rect 15108 10736 15160 10742
rect 15108 10678 15160 10684
rect 15120 10198 15148 10678
rect 15108 10192 15160 10198
rect 15108 10134 15160 10140
rect 15108 9376 15160 9382
rect 15108 9318 15160 9324
rect 15014 8936 15070 8945
rect 15014 8871 15070 8880
rect 14924 8492 14976 8498
rect 14924 8434 14976 8440
rect 14832 8288 14884 8294
rect 14738 8256 14794 8265
rect 14832 8230 14884 8236
rect 14738 8191 14794 8200
rect 14646 8120 14702 8129
rect 14646 8055 14702 8064
rect 14752 7954 14780 8191
rect 14740 7948 14792 7954
rect 14740 7890 14792 7896
rect 14648 7880 14700 7886
rect 14648 7822 14700 7828
rect 14556 7540 14608 7546
rect 14556 7482 14608 7488
rect 14556 7404 14608 7410
rect 14556 7346 14608 7352
rect 14464 6996 14516 7002
rect 14464 6938 14516 6944
rect 14016 6854 14320 6882
rect 13820 6724 13872 6730
rect 13820 6666 13872 6672
rect 13636 6656 13688 6662
rect 13636 6598 13688 6604
rect 13832 6390 13860 6666
rect 13820 6384 13872 6390
rect 13820 6326 13872 6332
rect 14016 6322 14044 6854
rect 14096 6792 14148 6798
rect 14096 6734 14148 6740
rect 14108 6322 14136 6734
rect 14188 6656 14240 6662
rect 14240 6616 14320 6644
rect 14188 6598 14240 6604
rect 14004 6316 14056 6322
rect 14004 6258 14056 6264
rect 14096 6316 14148 6322
rect 14096 6258 14148 6264
rect 13820 6248 13872 6254
rect 13820 6190 13872 6196
rect 13544 6112 13596 6118
rect 13544 6054 13596 6060
rect 13556 5658 13584 6054
rect 13636 5772 13688 5778
rect 13688 5732 13768 5760
rect 13636 5714 13688 5720
rect 13556 5630 13676 5658
rect 13544 5568 13596 5574
rect 13544 5510 13596 5516
rect 13556 5137 13584 5510
rect 13372 5086 13492 5114
rect 13542 5128 13598 5137
rect 13268 5024 13320 5030
rect 13268 4966 13320 4972
rect 13136 4576 13216 4604
rect 13084 4558 13136 4564
rect 12992 4072 13044 4078
rect 12992 4014 13044 4020
rect 12992 3936 13044 3942
rect 13096 3924 13124 4558
rect 13176 4480 13228 4486
rect 13176 4422 13228 4428
rect 13188 4282 13216 4422
rect 13176 4276 13228 4282
rect 13280 4264 13308 4966
rect 13372 4690 13400 5086
rect 13542 5063 13598 5072
rect 13452 5024 13504 5030
rect 13452 4966 13504 4972
rect 13544 5024 13596 5030
rect 13544 4966 13596 4972
rect 13360 4684 13412 4690
rect 13360 4626 13412 4632
rect 13464 4282 13492 4966
rect 13452 4276 13504 4282
rect 13280 4236 13400 4264
rect 13176 4218 13228 4224
rect 13268 4140 13320 4146
rect 13268 4082 13320 4088
rect 13176 4072 13228 4078
rect 13176 4014 13228 4020
rect 13044 3896 13124 3924
rect 12992 3878 13044 3884
rect 12808 2984 12860 2990
rect 12808 2926 12860 2932
rect 12900 2304 12952 2310
rect 12900 2246 12952 2252
rect 12624 2032 12676 2038
rect 12624 1974 12676 1980
rect 12912 800 12940 2246
rect 13004 1329 13032 3878
rect 13188 3466 13216 4014
rect 13280 3738 13308 4082
rect 13268 3732 13320 3738
rect 13268 3674 13320 3680
rect 13268 3528 13320 3534
rect 13268 3470 13320 3476
rect 13176 3460 13228 3466
rect 13176 3402 13228 3408
rect 13188 2514 13216 3402
rect 13280 3097 13308 3470
rect 13266 3088 13322 3097
rect 13266 3023 13322 3032
rect 13176 2508 13228 2514
rect 13176 2450 13228 2456
rect 13372 2446 13400 4236
rect 13452 4218 13504 4224
rect 13556 4185 13584 4966
rect 13648 4457 13676 5630
rect 13740 5302 13768 5732
rect 13832 5574 13860 6190
rect 14016 6118 14044 6258
rect 14004 6112 14056 6118
rect 14004 6054 14056 6060
rect 13945 6012 14253 6021
rect 13945 6010 13951 6012
rect 14007 6010 14031 6012
rect 14087 6010 14111 6012
rect 14167 6010 14191 6012
rect 14247 6010 14253 6012
rect 14007 5958 14009 6010
rect 14189 5958 14191 6010
rect 13945 5956 13951 5958
rect 14007 5956 14031 5958
rect 14087 5956 14111 5958
rect 14167 5956 14191 5958
rect 14247 5956 14253 5958
rect 13945 5947 14253 5956
rect 14186 5808 14242 5817
rect 14292 5778 14320 6616
rect 14464 6180 14516 6186
rect 14464 6122 14516 6128
rect 14372 6112 14424 6118
rect 14372 6054 14424 6060
rect 14186 5743 14242 5752
rect 14280 5772 14332 5778
rect 13912 5636 13964 5642
rect 13912 5578 13964 5584
rect 13820 5568 13872 5574
rect 13820 5510 13872 5516
rect 13728 5296 13780 5302
rect 13728 5238 13780 5244
rect 13740 4729 13768 5238
rect 13924 5012 13952 5578
rect 14200 5574 14228 5743
rect 14280 5714 14332 5720
rect 14188 5568 14240 5574
rect 14188 5510 14240 5516
rect 14292 5250 14320 5714
rect 14384 5370 14412 6054
rect 14476 5778 14504 6122
rect 14464 5772 14516 5778
rect 14464 5714 14516 5720
rect 14464 5568 14516 5574
rect 14464 5510 14516 5516
rect 14476 5409 14504 5510
rect 14462 5400 14518 5409
rect 14372 5364 14424 5370
rect 14462 5335 14518 5344
rect 14372 5306 14424 5312
rect 14292 5222 14412 5250
rect 13832 5001 13952 5012
rect 13818 4992 13952 5001
rect 13874 4984 13952 4992
rect 13818 4927 13874 4936
rect 13945 4924 14253 4933
rect 13945 4922 13951 4924
rect 14007 4922 14031 4924
rect 14087 4922 14111 4924
rect 14167 4922 14191 4924
rect 14247 4922 14253 4924
rect 14007 4870 14009 4922
rect 14189 4870 14191 4922
rect 13945 4868 13951 4870
rect 14007 4868 14031 4870
rect 14087 4868 14111 4870
rect 14167 4868 14191 4870
rect 14247 4868 14253 4870
rect 13945 4859 14253 4868
rect 13726 4720 13782 4729
rect 13726 4655 13728 4664
rect 13780 4655 13782 4664
rect 13728 4626 13780 4632
rect 13740 4595 13768 4626
rect 13634 4448 13690 4457
rect 13634 4383 13690 4392
rect 13542 4176 13598 4185
rect 13542 4111 13598 4120
rect 13556 4078 13584 4111
rect 13544 4072 13596 4078
rect 13544 4014 13596 4020
rect 13544 3664 13596 3670
rect 13544 3606 13596 3612
rect 13556 3398 13584 3606
rect 13648 3534 13676 4383
rect 14280 4072 14332 4078
rect 14280 4014 14332 4020
rect 13728 4004 13780 4010
rect 13728 3946 13780 3952
rect 13636 3528 13688 3534
rect 13636 3470 13688 3476
rect 13544 3392 13596 3398
rect 13544 3334 13596 3340
rect 13556 3194 13584 3334
rect 13544 3188 13596 3194
rect 13544 3130 13596 3136
rect 13636 2576 13688 2582
rect 13636 2518 13688 2524
rect 13360 2440 13412 2446
rect 13360 2382 13412 2388
rect 13268 2304 13320 2310
rect 13268 2246 13320 2252
rect 12990 1320 13046 1329
rect 12990 1255 13046 1264
rect 13280 800 13308 2246
rect 13648 800 13676 2518
rect 13740 2446 13768 3946
rect 13945 3836 14253 3845
rect 13945 3834 13951 3836
rect 14007 3834 14031 3836
rect 14087 3834 14111 3836
rect 14167 3834 14191 3836
rect 14247 3834 14253 3836
rect 14007 3782 14009 3834
rect 14189 3782 14191 3834
rect 13945 3780 13951 3782
rect 14007 3780 14031 3782
rect 14087 3780 14111 3782
rect 14167 3780 14191 3782
rect 14247 3780 14253 3782
rect 13945 3771 14253 3780
rect 14292 3720 14320 4014
rect 14200 3692 14320 3720
rect 13818 3632 13874 3641
rect 13818 3567 13874 3576
rect 13728 2440 13780 2446
rect 13728 2382 13780 2388
rect 13832 2310 13860 3567
rect 14200 3398 14228 3692
rect 13912 3392 13964 3398
rect 13912 3334 13964 3340
rect 14188 3392 14240 3398
rect 14188 3334 14240 3340
rect 14280 3392 14332 3398
rect 14280 3334 14332 3340
rect 13924 3058 13952 3334
rect 14200 3074 14228 3334
rect 14292 3194 14320 3334
rect 14280 3188 14332 3194
rect 14280 3130 14332 3136
rect 14384 3074 14412 5222
rect 14462 4720 14518 4729
rect 14462 4655 14464 4664
rect 14516 4655 14518 4664
rect 14464 4626 14516 4632
rect 14568 4622 14596 7346
rect 14660 5914 14688 7822
rect 14648 5908 14700 5914
rect 14648 5850 14700 5856
rect 14556 4616 14608 4622
rect 14556 4558 14608 4564
rect 14556 4480 14608 4486
rect 14554 4448 14556 4457
rect 14608 4448 14610 4457
rect 14554 4383 14610 4392
rect 14464 3936 14516 3942
rect 14464 3878 14516 3884
rect 14556 3936 14608 3942
rect 14556 3878 14608 3884
rect 14476 3194 14504 3878
rect 14568 3602 14596 3878
rect 14752 3641 14780 7890
rect 14936 7857 14964 8434
rect 15016 8356 15068 8362
rect 15016 8298 15068 8304
rect 15028 7970 15056 8298
rect 15120 8090 15148 9318
rect 15212 9058 15240 11342
rect 15292 11076 15344 11082
rect 15292 11018 15344 11024
rect 15304 10810 15332 11018
rect 15292 10804 15344 10810
rect 15292 10746 15344 10752
rect 15396 9722 15424 15982
rect 15568 15360 15620 15366
rect 15568 15302 15620 15308
rect 15660 15360 15712 15366
rect 15660 15302 15712 15308
rect 15474 14376 15530 14385
rect 15474 14311 15530 14320
rect 15488 13258 15516 14311
rect 15580 13870 15608 15302
rect 15568 13864 15620 13870
rect 15568 13806 15620 13812
rect 15476 13252 15528 13258
rect 15476 13194 15528 13200
rect 15672 12986 15700 15302
rect 15764 15162 15792 16186
rect 15856 15706 15884 19450
rect 15948 19242 15976 21082
rect 16040 20330 16068 22200
rect 16120 21004 16172 21010
rect 16120 20946 16172 20952
rect 16028 20324 16080 20330
rect 16028 20266 16080 20272
rect 16132 20262 16160 20946
rect 16408 20584 16436 22200
rect 16776 20890 16804 22200
rect 16776 20862 16988 20890
rect 16544 20700 16852 20709
rect 16544 20698 16550 20700
rect 16606 20698 16630 20700
rect 16686 20698 16710 20700
rect 16766 20698 16790 20700
rect 16846 20698 16852 20700
rect 16606 20646 16608 20698
rect 16788 20646 16790 20698
rect 16544 20644 16550 20646
rect 16606 20644 16630 20646
rect 16686 20644 16710 20646
rect 16766 20644 16790 20646
rect 16846 20644 16852 20646
rect 16544 20635 16852 20644
rect 16580 20596 16632 20602
rect 16408 20556 16580 20584
rect 16580 20538 16632 20544
rect 16304 20528 16356 20534
rect 16304 20470 16356 20476
rect 16212 20460 16264 20466
rect 16212 20402 16264 20408
rect 16120 20256 16172 20262
rect 16120 20198 16172 20204
rect 16224 20058 16252 20402
rect 16212 20052 16264 20058
rect 16212 19994 16264 20000
rect 16316 19718 16344 20470
rect 16960 20330 16988 20862
rect 17144 20584 17172 22200
rect 17512 20602 17540 22200
rect 17774 21040 17830 21049
rect 17774 20975 17830 20984
rect 17684 20800 17736 20806
rect 17684 20742 17736 20748
rect 17500 20596 17552 20602
rect 17144 20556 17264 20584
rect 17040 20460 17092 20466
rect 17040 20402 17092 20408
rect 17132 20460 17184 20466
rect 17132 20402 17184 20408
rect 16948 20324 17000 20330
rect 16948 20266 17000 20272
rect 16394 20088 16450 20097
rect 16394 20023 16450 20032
rect 16408 19922 16436 20023
rect 16396 19916 16448 19922
rect 16396 19858 16448 19864
rect 16948 19848 17000 19854
rect 16948 19790 17000 19796
rect 16396 19780 16448 19786
rect 16396 19722 16448 19728
rect 16304 19712 16356 19718
rect 16304 19654 16356 19660
rect 16120 19304 16172 19310
rect 16120 19246 16172 19252
rect 15936 19236 15988 19242
rect 15936 19178 15988 19184
rect 16028 18828 16080 18834
rect 16028 18770 16080 18776
rect 15936 16448 15988 16454
rect 15936 16390 15988 16396
rect 15948 16182 15976 16390
rect 15936 16176 15988 16182
rect 15936 16118 15988 16124
rect 15844 15700 15896 15706
rect 15844 15642 15896 15648
rect 15752 15156 15804 15162
rect 15804 15116 15884 15144
rect 15752 15098 15804 15104
rect 15752 14816 15804 14822
rect 15752 14758 15804 14764
rect 15764 14414 15792 14758
rect 15752 14408 15804 14414
rect 15752 14350 15804 14356
rect 15856 14056 15884 15116
rect 15764 14028 15884 14056
rect 15660 12980 15712 12986
rect 15660 12922 15712 12928
rect 15476 12844 15528 12850
rect 15476 12786 15528 12792
rect 15660 12844 15712 12850
rect 15660 12786 15712 12792
rect 15488 12306 15516 12786
rect 15568 12776 15620 12782
rect 15568 12718 15620 12724
rect 15580 12434 15608 12718
rect 15672 12714 15700 12786
rect 15660 12708 15712 12714
rect 15660 12650 15712 12656
rect 15580 12406 15700 12434
rect 15476 12300 15528 12306
rect 15476 12242 15528 12248
rect 15568 11756 15620 11762
rect 15568 11698 15620 11704
rect 15476 11552 15528 11558
rect 15476 11494 15528 11500
rect 15488 10713 15516 11494
rect 15580 11354 15608 11698
rect 15672 11694 15700 12406
rect 15660 11688 15712 11694
rect 15660 11630 15712 11636
rect 15568 11348 15620 11354
rect 15568 11290 15620 11296
rect 15566 11112 15622 11121
rect 15566 11047 15622 11056
rect 15474 10704 15530 10713
rect 15474 10639 15530 10648
rect 15384 9716 15436 9722
rect 15384 9658 15436 9664
rect 15580 9654 15608 11047
rect 15660 10600 15712 10606
rect 15660 10542 15712 10548
rect 15672 10266 15700 10542
rect 15660 10260 15712 10266
rect 15660 10202 15712 10208
rect 15660 10124 15712 10130
rect 15660 10066 15712 10072
rect 15568 9648 15620 9654
rect 15290 9616 15346 9625
rect 15568 9590 15620 9596
rect 15290 9551 15346 9560
rect 15476 9580 15528 9586
rect 15304 9450 15332 9551
rect 15476 9522 15528 9528
rect 15292 9444 15344 9450
rect 15292 9386 15344 9392
rect 15488 9353 15516 9522
rect 15568 9376 15620 9382
rect 15474 9344 15530 9353
rect 15568 9318 15620 9324
rect 15474 9279 15530 9288
rect 15474 9208 15530 9217
rect 15474 9143 15530 9152
rect 15212 9030 15424 9058
rect 15200 8900 15252 8906
rect 15200 8842 15252 8848
rect 15212 8430 15240 8842
rect 15292 8832 15344 8838
rect 15292 8774 15344 8780
rect 15200 8424 15252 8430
rect 15200 8366 15252 8372
rect 15108 8084 15160 8090
rect 15108 8026 15160 8032
rect 15028 7942 15148 7970
rect 15212 7954 15240 8366
rect 15304 7954 15332 8774
rect 14922 7848 14978 7857
rect 14922 7783 14978 7792
rect 14832 7540 14884 7546
rect 14832 7482 14884 7488
rect 15016 7540 15068 7546
rect 15016 7482 15068 7488
rect 14844 7206 14872 7482
rect 14924 7336 14976 7342
rect 14924 7278 14976 7284
rect 14832 7200 14884 7206
rect 14832 7142 14884 7148
rect 14832 6112 14884 6118
rect 14832 6054 14884 6060
rect 14844 5234 14872 6054
rect 14936 5710 14964 7278
rect 14924 5704 14976 5710
rect 14924 5646 14976 5652
rect 14832 5228 14884 5234
rect 14832 5170 14884 5176
rect 14738 3632 14794 3641
rect 14556 3596 14608 3602
rect 14738 3567 14794 3576
rect 14556 3538 14608 3544
rect 14740 3528 14792 3534
rect 14740 3470 14792 3476
rect 14752 3233 14780 3470
rect 14738 3224 14794 3233
rect 14464 3188 14516 3194
rect 14738 3159 14794 3168
rect 14464 3130 14516 3136
rect 14844 3126 14872 5170
rect 14832 3120 14884 3126
rect 14830 3088 14832 3097
rect 14884 3088 14886 3097
rect 13912 3052 13964 3058
rect 14200 3046 14320 3074
rect 14384 3046 14596 3074
rect 13912 2994 13964 3000
rect 14292 2990 14320 3046
rect 14280 2984 14332 2990
rect 14280 2926 14332 2932
rect 14372 2848 14424 2854
rect 14372 2790 14424 2796
rect 13945 2748 14253 2757
rect 13945 2746 13951 2748
rect 14007 2746 14031 2748
rect 14087 2746 14111 2748
rect 14167 2746 14191 2748
rect 14247 2746 14253 2748
rect 14007 2694 14009 2746
rect 14189 2694 14191 2746
rect 13945 2692 13951 2694
rect 14007 2692 14031 2694
rect 14087 2692 14111 2694
rect 14167 2692 14191 2694
rect 14247 2692 14253 2694
rect 13945 2683 14253 2692
rect 14004 2372 14056 2378
rect 14004 2314 14056 2320
rect 13820 2304 13872 2310
rect 13820 2246 13872 2252
rect 14016 800 14044 2314
rect 14384 800 14412 2790
rect 14464 2304 14516 2310
rect 14464 2246 14516 2252
rect 14476 1834 14504 2246
rect 14568 1970 14596 3046
rect 14648 3052 14700 3058
rect 14830 3023 14886 3032
rect 14648 2994 14700 3000
rect 14660 2650 14688 2994
rect 14648 2644 14700 2650
rect 14648 2586 14700 2592
rect 14740 2372 14792 2378
rect 14740 2314 14792 2320
rect 14556 1964 14608 1970
rect 14556 1906 14608 1912
rect 14464 1828 14516 1834
rect 14464 1770 14516 1776
rect 14752 800 14780 2314
rect 14936 1902 14964 5646
rect 15028 4321 15056 7482
rect 15120 7002 15148 7942
rect 15200 7948 15252 7954
rect 15200 7890 15252 7896
rect 15292 7948 15344 7954
rect 15292 7890 15344 7896
rect 15304 7834 15332 7890
rect 15212 7806 15332 7834
rect 15212 7342 15240 7806
rect 15292 7744 15344 7750
rect 15292 7686 15344 7692
rect 15304 7546 15332 7686
rect 15292 7540 15344 7546
rect 15292 7482 15344 7488
rect 15200 7336 15252 7342
rect 15396 7313 15424 9030
rect 15488 8974 15516 9143
rect 15476 8968 15528 8974
rect 15476 8910 15528 8916
rect 15580 8430 15608 9318
rect 15568 8424 15620 8430
rect 15568 8366 15620 8372
rect 15672 8362 15700 10066
rect 15764 9674 15792 14028
rect 15844 13932 15896 13938
rect 15844 13874 15896 13880
rect 15856 13530 15884 13874
rect 15844 13524 15896 13530
rect 15844 13466 15896 13472
rect 15936 13320 15988 13326
rect 15936 13262 15988 13268
rect 15948 12646 15976 13262
rect 15936 12640 15988 12646
rect 15936 12582 15988 12588
rect 15844 12096 15896 12102
rect 15844 12038 15896 12044
rect 15856 11150 15884 12038
rect 15936 11892 15988 11898
rect 15936 11834 15988 11840
rect 15844 11144 15896 11150
rect 15844 11086 15896 11092
rect 15856 11014 15884 11086
rect 15844 11008 15896 11014
rect 15844 10950 15896 10956
rect 15856 10674 15884 10950
rect 15844 10668 15896 10674
rect 15844 10610 15896 10616
rect 15764 9646 15884 9674
rect 15752 9580 15804 9586
rect 15752 9522 15804 9528
rect 15764 8838 15792 9522
rect 15752 8832 15804 8838
rect 15752 8774 15804 8780
rect 15856 8566 15884 9646
rect 15844 8560 15896 8566
rect 15844 8502 15896 8508
rect 15752 8424 15804 8430
rect 15752 8366 15804 8372
rect 15660 8356 15712 8362
rect 15660 8298 15712 8304
rect 15566 8120 15622 8129
rect 15566 8055 15622 8064
rect 15474 7576 15530 7585
rect 15474 7511 15530 7520
rect 15488 7410 15516 7511
rect 15476 7404 15528 7410
rect 15476 7346 15528 7352
rect 15200 7278 15252 7284
rect 15382 7304 15438 7313
rect 15108 6996 15160 7002
rect 15108 6938 15160 6944
rect 15106 6896 15162 6905
rect 15106 6831 15162 6840
rect 15120 6798 15148 6831
rect 15108 6792 15160 6798
rect 15108 6734 15160 6740
rect 15120 5234 15148 6734
rect 15212 6730 15240 7278
rect 15292 7268 15344 7274
rect 15382 7239 15438 7248
rect 15292 7210 15344 7216
rect 15200 6724 15252 6730
rect 15200 6666 15252 6672
rect 15108 5228 15160 5234
rect 15108 5170 15160 5176
rect 15212 5166 15240 6666
rect 15200 5160 15252 5166
rect 15200 5102 15252 5108
rect 15200 5024 15252 5030
rect 15200 4966 15252 4972
rect 15108 4548 15160 4554
rect 15108 4490 15160 4496
rect 15014 4312 15070 4321
rect 15120 4282 15148 4490
rect 15014 4247 15070 4256
rect 15108 4276 15160 4282
rect 15108 4218 15160 4224
rect 15212 4049 15240 4966
rect 15304 4622 15332 7210
rect 15384 7200 15436 7206
rect 15384 7142 15436 7148
rect 15396 5710 15424 7142
rect 15580 7041 15608 8055
rect 15566 7032 15622 7041
rect 15566 6967 15622 6976
rect 15568 6860 15620 6866
rect 15488 6820 15568 6848
rect 15488 6662 15516 6820
rect 15568 6802 15620 6808
rect 15476 6656 15528 6662
rect 15476 6598 15528 6604
rect 15568 6656 15620 6662
rect 15568 6598 15620 6604
rect 15488 6322 15516 6598
rect 15476 6316 15528 6322
rect 15476 6258 15528 6264
rect 15476 5840 15528 5846
rect 15476 5782 15528 5788
rect 15384 5704 15436 5710
rect 15384 5646 15436 5652
rect 15384 5568 15436 5574
rect 15384 5510 15436 5516
rect 15292 4616 15344 4622
rect 15292 4558 15344 4564
rect 15290 4176 15346 4185
rect 15290 4111 15346 4120
rect 15304 4078 15332 4111
rect 15292 4072 15344 4078
rect 15198 4040 15254 4049
rect 15016 4004 15068 4010
rect 15292 4014 15344 4020
rect 15198 3975 15254 3984
rect 15016 3946 15068 3952
rect 15028 3777 15056 3946
rect 15014 3768 15070 3777
rect 15014 3703 15070 3712
rect 15292 3664 15344 3670
rect 15292 3606 15344 3612
rect 15016 3460 15068 3466
rect 15016 3402 15068 3408
rect 15028 2990 15056 3402
rect 15200 3392 15252 3398
rect 15200 3334 15252 3340
rect 15016 2984 15068 2990
rect 15016 2926 15068 2932
rect 15212 2666 15240 3334
rect 15028 2638 15240 2666
rect 15028 2446 15056 2638
rect 15108 2576 15160 2582
rect 15108 2518 15160 2524
rect 15016 2440 15068 2446
rect 15016 2382 15068 2388
rect 14924 1896 14976 1902
rect 14924 1838 14976 1844
rect 15120 800 15148 2518
rect 15304 2446 15332 3606
rect 15396 2922 15424 5510
rect 15488 3058 15516 5782
rect 15580 4622 15608 6598
rect 15672 6100 15700 8298
rect 15764 6254 15792 8366
rect 15844 8288 15896 8294
rect 15844 8230 15896 8236
rect 15856 7342 15884 8230
rect 15948 7834 15976 11834
rect 16040 10130 16068 18770
rect 16132 18630 16160 19246
rect 16408 18630 16436 19722
rect 16544 19612 16852 19621
rect 16544 19610 16550 19612
rect 16606 19610 16630 19612
rect 16686 19610 16710 19612
rect 16766 19610 16790 19612
rect 16846 19610 16852 19612
rect 16606 19558 16608 19610
rect 16788 19558 16790 19610
rect 16544 19556 16550 19558
rect 16606 19556 16630 19558
rect 16686 19556 16710 19558
rect 16766 19556 16790 19558
rect 16846 19556 16852 19558
rect 16544 19547 16852 19556
rect 16854 19408 16910 19417
rect 16854 19343 16856 19352
rect 16908 19343 16910 19352
rect 16856 19314 16908 19320
rect 16960 18902 16988 19790
rect 17052 18970 17080 20402
rect 17144 20058 17172 20402
rect 17236 20262 17264 20556
rect 17500 20538 17552 20544
rect 17408 20460 17460 20466
rect 17408 20402 17460 20408
rect 17592 20460 17644 20466
rect 17592 20402 17644 20408
rect 17224 20256 17276 20262
rect 17224 20198 17276 20204
rect 17132 20052 17184 20058
rect 17132 19994 17184 20000
rect 17224 19848 17276 19854
rect 17224 19790 17276 19796
rect 17132 19780 17184 19786
rect 17132 19722 17184 19728
rect 17040 18964 17092 18970
rect 17040 18906 17092 18912
rect 16948 18896 17000 18902
rect 16948 18838 17000 18844
rect 16120 18624 16172 18630
rect 16120 18566 16172 18572
rect 16396 18624 16448 18630
rect 17144 18612 17172 19722
rect 17236 19394 17264 19790
rect 17420 19514 17448 20402
rect 17604 20058 17632 20402
rect 17696 20058 17724 20742
rect 17592 20052 17644 20058
rect 17592 19994 17644 20000
rect 17684 20052 17736 20058
rect 17684 19994 17736 20000
rect 17684 19916 17736 19922
rect 17684 19858 17736 19864
rect 17408 19508 17460 19514
rect 17408 19450 17460 19456
rect 17236 19366 17448 19394
rect 17316 19236 17368 19242
rect 17316 19178 17368 19184
rect 17224 18624 17276 18630
rect 17144 18584 17224 18612
rect 16396 18566 16448 18572
rect 17224 18566 17276 18572
rect 16132 18222 16160 18566
rect 16120 18216 16172 18222
rect 16120 18158 16172 18164
rect 16212 18148 16264 18154
rect 16212 18090 16264 18096
rect 16224 17134 16252 18090
rect 16212 17128 16264 17134
rect 16212 17070 16264 17076
rect 16408 17066 16436 18566
rect 16544 18524 16852 18533
rect 16544 18522 16550 18524
rect 16606 18522 16630 18524
rect 16686 18522 16710 18524
rect 16766 18522 16790 18524
rect 16846 18522 16852 18524
rect 16606 18470 16608 18522
rect 16788 18470 16790 18522
rect 16544 18468 16550 18470
rect 16606 18468 16630 18470
rect 16686 18468 16710 18470
rect 16766 18468 16790 18470
rect 16846 18468 16852 18470
rect 16544 18459 16852 18468
rect 17236 18057 17264 18566
rect 17222 18048 17278 18057
rect 17222 17983 17278 17992
rect 17040 17876 17092 17882
rect 17040 17818 17092 17824
rect 16948 17604 17000 17610
rect 16948 17546 17000 17552
rect 16544 17436 16852 17445
rect 16544 17434 16550 17436
rect 16606 17434 16630 17436
rect 16686 17434 16710 17436
rect 16766 17434 16790 17436
rect 16846 17434 16852 17436
rect 16606 17382 16608 17434
rect 16788 17382 16790 17434
rect 16544 17380 16550 17382
rect 16606 17380 16630 17382
rect 16686 17380 16710 17382
rect 16766 17380 16790 17382
rect 16846 17380 16852 17382
rect 16544 17371 16852 17380
rect 16396 17060 16448 17066
rect 16396 17002 16448 17008
rect 16210 16688 16266 16697
rect 16210 16623 16212 16632
rect 16264 16623 16266 16632
rect 16212 16594 16264 16600
rect 16396 16584 16448 16590
rect 16396 16526 16448 16532
rect 16120 16448 16172 16454
rect 16120 16390 16172 16396
rect 16132 16289 16160 16390
rect 16118 16280 16174 16289
rect 16118 16215 16174 16224
rect 16120 16108 16172 16114
rect 16120 16050 16172 16056
rect 16132 15706 16160 16050
rect 16408 15910 16436 16526
rect 16960 16522 16988 17546
rect 17052 17338 17080 17818
rect 17040 17332 17092 17338
rect 17040 17274 17092 17280
rect 17132 17128 17184 17134
rect 17132 17070 17184 17076
rect 17224 17128 17276 17134
rect 17224 17070 17276 17076
rect 17144 16794 17172 17070
rect 17236 16998 17264 17070
rect 17224 16992 17276 16998
rect 17224 16934 17276 16940
rect 17132 16788 17184 16794
rect 17132 16730 17184 16736
rect 17236 16658 17264 16934
rect 17224 16652 17276 16658
rect 17224 16594 17276 16600
rect 16948 16516 17000 16522
rect 16948 16458 17000 16464
rect 16544 16348 16852 16357
rect 16544 16346 16550 16348
rect 16606 16346 16630 16348
rect 16686 16346 16710 16348
rect 16766 16346 16790 16348
rect 16846 16346 16852 16348
rect 16606 16294 16608 16346
rect 16788 16294 16790 16346
rect 16544 16292 16550 16294
rect 16606 16292 16630 16294
rect 16686 16292 16710 16294
rect 16766 16292 16790 16294
rect 16846 16292 16852 16294
rect 16544 16283 16852 16292
rect 17132 16040 17184 16046
rect 17132 15982 17184 15988
rect 16396 15904 16448 15910
rect 16396 15846 16448 15852
rect 16120 15700 16172 15706
rect 16120 15642 16172 15648
rect 17144 15570 17172 15982
rect 16120 15564 16172 15570
rect 16120 15506 16172 15512
rect 17132 15564 17184 15570
rect 17132 15506 17184 15512
rect 16132 15162 16160 15506
rect 16304 15496 16356 15502
rect 16304 15438 16356 15444
rect 16948 15496 17000 15502
rect 16948 15438 17000 15444
rect 17038 15464 17094 15473
rect 16120 15156 16172 15162
rect 16120 15098 16172 15104
rect 16132 14346 16160 15098
rect 16120 14340 16172 14346
rect 16120 14282 16172 14288
rect 16316 14006 16344 15438
rect 16396 15360 16448 15366
rect 16396 15302 16448 15308
rect 16408 14618 16436 15302
rect 16544 15260 16852 15269
rect 16544 15258 16550 15260
rect 16606 15258 16630 15260
rect 16686 15258 16710 15260
rect 16766 15258 16790 15260
rect 16846 15258 16852 15260
rect 16606 15206 16608 15258
rect 16788 15206 16790 15258
rect 16544 15204 16550 15206
rect 16606 15204 16630 15206
rect 16686 15204 16710 15206
rect 16766 15204 16790 15206
rect 16846 15204 16852 15206
rect 16544 15195 16852 15204
rect 16856 14952 16908 14958
rect 16856 14894 16908 14900
rect 16396 14612 16448 14618
rect 16396 14554 16448 14560
rect 16868 14414 16896 14894
rect 16856 14408 16908 14414
rect 16856 14350 16908 14356
rect 16544 14172 16852 14181
rect 16544 14170 16550 14172
rect 16606 14170 16630 14172
rect 16686 14170 16710 14172
rect 16766 14170 16790 14172
rect 16846 14170 16852 14172
rect 16606 14118 16608 14170
rect 16788 14118 16790 14170
rect 16544 14116 16550 14118
rect 16606 14116 16630 14118
rect 16686 14116 16710 14118
rect 16766 14116 16790 14118
rect 16846 14116 16852 14118
rect 16544 14107 16852 14116
rect 16960 14074 16988 15438
rect 17038 15399 17094 15408
rect 16948 14068 17000 14074
rect 16948 14010 17000 14016
rect 16212 14000 16264 14006
rect 16212 13942 16264 13948
rect 16304 14000 16356 14006
rect 16304 13942 16356 13948
rect 16120 13796 16172 13802
rect 16120 13738 16172 13744
rect 16132 13190 16160 13738
rect 16120 13184 16172 13190
rect 16120 13126 16172 13132
rect 16224 12434 16252 13942
rect 16316 13462 16344 13942
rect 16304 13456 16356 13462
rect 16304 13398 16356 13404
rect 16948 13388 17000 13394
rect 16948 13330 17000 13336
rect 16544 13084 16852 13093
rect 16544 13082 16550 13084
rect 16606 13082 16630 13084
rect 16686 13082 16710 13084
rect 16766 13082 16790 13084
rect 16846 13082 16852 13084
rect 16606 13030 16608 13082
rect 16788 13030 16790 13082
rect 16544 13028 16550 13030
rect 16606 13028 16630 13030
rect 16686 13028 16710 13030
rect 16766 13028 16790 13030
rect 16846 13028 16852 13030
rect 16544 13019 16852 13028
rect 16960 12986 16988 13330
rect 17052 13308 17080 15399
rect 17144 15026 17172 15506
rect 17132 15020 17184 15026
rect 17132 14962 17184 14968
rect 17144 14550 17172 14962
rect 17132 14544 17184 14550
rect 17132 14486 17184 14492
rect 17224 14476 17276 14482
rect 17224 14418 17276 14424
rect 17132 13932 17184 13938
rect 17132 13874 17184 13880
rect 17144 13734 17172 13874
rect 17236 13870 17264 14418
rect 17328 13938 17356 19178
rect 17420 19174 17448 19366
rect 17696 19174 17724 19858
rect 17788 19378 17816 20975
rect 17880 20584 17908 22200
rect 18052 20800 18104 20806
rect 18052 20742 18104 20748
rect 17880 20556 18000 20584
rect 17972 20398 18000 20556
rect 17960 20392 18012 20398
rect 17960 20334 18012 20340
rect 17960 19984 18012 19990
rect 17958 19952 17960 19961
rect 18012 19952 18014 19961
rect 17958 19887 18014 19896
rect 17776 19372 17828 19378
rect 17776 19314 17828 19320
rect 17408 19168 17460 19174
rect 17684 19168 17736 19174
rect 17408 19110 17460 19116
rect 17682 19136 17684 19145
rect 17736 19136 17738 19145
rect 17420 18834 17448 19110
rect 17682 19071 17738 19080
rect 17408 18828 17460 18834
rect 17408 18770 17460 18776
rect 17788 17882 17816 19314
rect 18064 18970 18092 20742
rect 18144 20460 18196 20466
rect 18144 20402 18196 20408
rect 18156 19446 18184 20402
rect 18248 20058 18276 22200
rect 18510 21856 18566 21865
rect 18510 21791 18566 21800
rect 18328 20460 18380 20466
rect 18328 20402 18380 20408
rect 18236 20052 18288 20058
rect 18236 19994 18288 20000
rect 18234 19816 18290 19825
rect 18234 19751 18290 19760
rect 18144 19440 18196 19446
rect 18144 19382 18196 19388
rect 18248 19378 18276 19751
rect 18340 19514 18368 20402
rect 18420 19848 18472 19854
rect 18420 19790 18472 19796
rect 18328 19508 18380 19514
rect 18328 19450 18380 19456
rect 18236 19372 18288 19378
rect 18236 19314 18288 19320
rect 18052 18964 18104 18970
rect 18052 18906 18104 18912
rect 18050 18864 18106 18873
rect 18050 18799 18106 18808
rect 18064 18766 18092 18799
rect 18432 18766 18460 19790
rect 18524 18970 18552 21791
rect 18616 19310 18644 22200
rect 18786 22128 18842 22137
rect 18786 22063 18842 22072
rect 18696 20052 18748 20058
rect 18696 19994 18748 20000
rect 18708 19378 18736 19994
rect 18800 19990 18828 22063
rect 18984 20466 19012 22200
rect 18972 20460 19024 20466
rect 18972 20402 19024 20408
rect 18880 20324 18932 20330
rect 18880 20266 18932 20272
rect 18788 19984 18840 19990
rect 18788 19926 18840 19932
rect 18788 19848 18840 19854
rect 18788 19790 18840 19796
rect 18800 19514 18828 19790
rect 18788 19508 18840 19514
rect 18788 19450 18840 19456
rect 18696 19372 18748 19378
rect 18696 19314 18748 19320
rect 18604 19304 18656 19310
rect 18604 19246 18656 19252
rect 18786 19272 18842 19281
rect 18512 18964 18564 18970
rect 18512 18906 18564 18912
rect 18052 18760 18104 18766
rect 18052 18702 18104 18708
rect 18420 18760 18472 18766
rect 18420 18702 18472 18708
rect 18432 18154 18460 18702
rect 18616 18426 18644 19246
rect 18786 19207 18842 19216
rect 18800 18766 18828 19207
rect 18788 18760 18840 18766
rect 18788 18702 18840 18708
rect 18892 18630 18920 20266
rect 18984 19514 19012 20402
rect 19064 20392 19116 20398
rect 19064 20334 19116 20340
rect 19076 19990 19104 20334
rect 19352 20244 19380 22200
rect 19522 21040 19578 21049
rect 19522 20975 19578 20984
rect 19536 20602 19564 20975
rect 19720 20806 19748 22200
rect 19708 20800 19760 20806
rect 19760 20760 19932 20788
rect 19708 20742 19760 20748
rect 19524 20596 19576 20602
rect 19524 20538 19576 20544
rect 19708 20460 19760 20466
rect 19708 20402 19760 20408
rect 19800 20460 19852 20466
rect 19800 20402 19852 20408
rect 19352 20216 19564 20244
rect 19143 20156 19451 20165
rect 19143 20154 19149 20156
rect 19205 20154 19229 20156
rect 19285 20154 19309 20156
rect 19365 20154 19389 20156
rect 19445 20154 19451 20156
rect 19205 20102 19207 20154
rect 19387 20102 19389 20154
rect 19143 20100 19149 20102
rect 19205 20100 19229 20102
rect 19285 20100 19309 20102
rect 19365 20100 19389 20102
rect 19445 20100 19451 20102
rect 19143 20091 19451 20100
rect 19340 20052 19392 20058
rect 19340 19994 19392 20000
rect 19064 19984 19116 19990
rect 19064 19926 19116 19932
rect 19076 19514 19104 19926
rect 19154 19816 19210 19825
rect 19154 19751 19210 19760
rect 18972 19508 19024 19514
rect 18972 19450 19024 19456
rect 19064 19508 19116 19514
rect 19064 19450 19116 19456
rect 19168 19378 19196 19751
rect 19156 19372 19208 19378
rect 19156 19314 19208 19320
rect 19352 19258 19380 19994
rect 19536 19938 19564 20216
rect 19444 19910 19564 19938
rect 19614 19952 19670 19961
rect 19444 19378 19472 19910
rect 19614 19887 19616 19896
rect 19668 19887 19670 19896
rect 19616 19858 19668 19864
rect 19524 19848 19576 19854
rect 19524 19790 19576 19796
rect 19432 19372 19484 19378
rect 19432 19314 19484 19320
rect 19536 19258 19564 19790
rect 19616 19780 19668 19786
rect 19616 19722 19668 19728
rect 19628 19281 19656 19722
rect 19076 19230 19380 19258
rect 19444 19230 19564 19258
rect 19614 19272 19670 19281
rect 18972 19168 19024 19174
rect 18972 19110 19024 19116
rect 18984 18766 19012 19110
rect 19076 18850 19104 19230
rect 19444 19156 19472 19230
rect 19614 19207 19670 19216
rect 19444 19128 19503 19156
rect 19475 19122 19503 19128
rect 19614 19136 19670 19145
rect 19475 19094 19555 19122
rect 19143 19068 19451 19077
rect 19143 19066 19149 19068
rect 19205 19066 19229 19068
rect 19285 19066 19309 19068
rect 19365 19066 19389 19068
rect 19445 19066 19451 19068
rect 19205 19014 19207 19066
rect 19387 19014 19389 19066
rect 19143 19012 19149 19014
rect 19205 19012 19229 19014
rect 19285 19012 19309 19014
rect 19365 19012 19389 19014
rect 19445 19012 19451 19014
rect 19143 19003 19451 19012
rect 19527 18986 19555 19094
rect 19614 19071 19670 19080
rect 19527 18958 19564 18986
rect 19076 18822 19196 18850
rect 18972 18760 19024 18766
rect 18972 18702 19024 18708
rect 19168 18630 19196 18822
rect 19294 18828 19346 18834
rect 19294 18770 19346 18776
rect 19432 18828 19484 18834
rect 19432 18770 19484 18776
rect 19306 18737 19334 18770
rect 19444 18737 19472 18770
rect 19292 18728 19348 18737
rect 19292 18663 19348 18672
rect 19430 18728 19486 18737
rect 19430 18663 19486 18672
rect 19536 18630 19564 18958
rect 19628 18698 19656 19071
rect 19616 18692 19668 18698
rect 19616 18634 19668 18640
rect 18880 18624 18932 18630
rect 18880 18566 18932 18572
rect 19156 18624 19208 18630
rect 19156 18566 19208 18572
rect 19340 18624 19392 18630
rect 19340 18566 19392 18572
rect 19524 18624 19576 18630
rect 19524 18566 19576 18572
rect 19352 18442 19380 18566
rect 19614 18456 19670 18465
rect 18604 18420 18656 18426
rect 19352 18414 19564 18442
rect 18604 18362 18656 18368
rect 18512 18352 18564 18358
rect 18512 18294 18564 18300
rect 18420 18148 18472 18154
rect 18420 18090 18472 18096
rect 17776 17876 17828 17882
rect 17776 17818 17828 17824
rect 17500 16992 17552 16998
rect 17500 16934 17552 16940
rect 17512 16454 17540 16934
rect 17774 16688 17830 16697
rect 17774 16623 17776 16632
rect 17828 16623 17830 16632
rect 17776 16594 17828 16600
rect 18052 16584 18104 16590
rect 18052 16526 18104 16532
rect 17500 16448 17552 16454
rect 17500 16390 17552 16396
rect 17408 14340 17460 14346
rect 17408 14282 17460 14288
rect 17316 13932 17368 13938
rect 17316 13874 17368 13880
rect 17224 13864 17276 13870
rect 17224 13806 17276 13812
rect 17132 13728 17184 13734
rect 17132 13670 17184 13676
rect 17052 13280 17172 13308
rect 17040 13184 17092 13190
rect 17038 13152 17040 13161
rect 17092 13152 17094 13161
rect 17038 13087 17094 13096
rect 16948 12980 17000 12986
rect 16948 12922 17000 12928
rect 16488 12912 16540 12918
rect 16488 12854 16540 12860
rect 16500 12434 16528 12854
rect 16856 12844 16908 12850
rect 16856 12786 16908 12792
rect 16868 12442 16896 12786
rect 16948 12640 17000 12646
rect 16948 12582 17000 12588
rect 16960 12442 16988 12582
rect 16224 12406 16344 12434
rect 16212 12164 16264 12170
rect 16212 12106 16264 12112
rect 16224 12073 16252 12106
rect 16210 12064 16266 12073
rect 16210 11999 16266 12008
rect 16210 11928 16266 11937
rect 16210 11863 16266 11872
rect 16120 11756 16172 11762
rect 16120 11698 16172 11704
rect 16132 10810 16160 11698
rect 16224 11082 16252 11863
rect 16316 11540 16344 12406
rect 16408 12406 16528 12434
rect 16856 12436 16908 12442
rect 16408 11898 16436 12406
rect 16856 12378 16908 12384
rect 16948 12436 17000 12442
rect 16948 12378 17000 12384
rect 16544 11996 16852 12005
rect 16544 11994 16550 11996
rect 16606 11994 16630 11996
rect 16686 11994 16710 11996
rect 16766 11994 16790 11996
rect 16846 11994 16852 11996
rect 16606 11942 16608 11994
rect 16788 11942 16790 11994
rect 16544 11940 16550 11942
rect 16606 11940 16630 11942
rect 16686 11940 16710 11942
rect 16766 11940 16790 11942
rect 16846 11940 16852 11942
rect 16544 11931 16852 11940
rect 16946 11928 17002 11937
rect 16396 11892 16448 11898
rect 16946 11863 16948 11872
rect 16396 11834 16448 11840
rect 17000 11863 17002 11872
rect 16948 11834 17000 11840
rect 16854 11656 16910 11665
rect 16854 11591 16910 11600
rect 16948 11620 17000 11626
rect 16396 11552 16448 11558
rect 16316 11512 16396 11540
rect 16396 11494 16448 11500
rect 16212 11076 16264 11082
rect 16212 11018 16264 11024
rect 16120 10804 16172 10810
rect 16120 10746 16172 10752
rect 16210 10296 16266 10305
rect 16210 10231 16266 10240
rect 16028 10124 16080 10130
rect 16028 10066 16080 10072
rect 16118 10024 16174 10033
rect 16224 10010 16252 10231
rect 16174 9982 16252 10010
rect 16118 9959 16174 9968
rect 16028 9920 16080 9926
rect 16120 9920 16172 9926
rect 16028 9862 16080 9868
rect 16118 9888 16120 9897
rect 16172 9888 16174 9897
rect 16040 9654 16068 9862
rect 16118 9823 16174 9832
rect 16224 9654 16252 9982
rect 16304 9988 16356 9994
rect 16304 9930 16356 9936
rect 16316 9722 16344 9930
rect 16304 9716 16356 9722
rect 16304 9658 16356 9664
rect 16028 9648 16080 9654
rect 16028 9590 16080 9596
rect 16212 9648 16264 9654
rect 16212 9590 16264 9596
rect 16316 9586 16344 9658
rect 16304 9580 16356 9586
rect 16304 9522 16356 9528
rect 16028 8900 16080 8906
rect 16028 8842 16080 8848
rect 16040 8090 16068 8842
rect 16120 8832 16172 8838
rect 16120 8774 16172 8780
rect 16132 8090 16160 8774
rect 16212 8560 16264 8566
rect 16212 8502 16264 8508
rect 16224 8294 16252 8502
rect 16304 8356 16356 8362
rect 16304 8298 16356 8304
rect 16212 8288 16264 8294
rect 16212 8230 16264 8236
rect 16028 8084 16080 8090
rect 16028 8026 16080 8032
rect 16120 8084 16172 8090
rect 16120 8026 16172 8032
rect 16118 7848 16174 7857
rect 15948 7806 16118 7834
rect 16224 7818 16252 8230
rect 16118 7783 16174 7792
rect 16212 7812 16264 7818
rect 15936 7744 15988 7750
rect 15936 7686 15988 7692
rect 15844 7336 15896 7342
rect 15844 7278 15896 7284
rect 15856 6322 15884 7278
rect 15948 6730 15976 7686
rect 16028 7336 16080 7342
rect 16026 7304 16028 7313
rect 16080 7304 16082 7313
rect 16026 7239 16082 7248
rect 15936 6724 15988 6730
rect 15936 6666 15988 6672
rect 16028 6656 16080 6662
rect 16028 6598 16080 6604
rect 15934 6488 15990 6497
rect 16040 6458 16068 6598
rect 15934 6423 15990 6432
rect 16028 6452 16080 6458
rect 15844 6316 15896 6322
rect 15844 6258 15896 6264
rect 15752 6248 15804 6254
rect 15752 6190 15804 6196
rect 15672 6072 15884 6100
rect 15660 5228 15712 5234
rect 15660 5170 15712 5176
rect 15568 4616 15620 4622
rect 15568 4558 15620 4564
rect 15672 3913 15700 5170
rect 15752 4480 15804 4486
rect 15752 4422 15804 4428
rect 15658 3904 15714 3913
rect 15658 3839 15714 3848
rect 15764 3398 15792 4422
rect 15856 4078 15884 6072
rect 15948 4282 15976 6423
rect 16028 6394 16080 6400
rect 16028 6316 16080 6322
rect 16028 6258 16080 6264
rect 15936 4276 15988 4282
rect 15936 4218 15988 4224
rect 16040 4185 16068 6258
rect 16132 6118 16160 7783
rect 16212 7754 16264 7760
rect 16212 7404 16264 7410
rect 16212 7346 16264 7352
rect 16224 7206 16252 7346
rect 16212 7200 16264 7206
rect 16210 7168 16212 7177
rect 16264 7168 16266 7177
rect 16210 7103 16266 7112
rect 16316 6390 16344 8298
rect 16408 8265 16436 11494
rect 16868 11286 16896 11591
rect 16948 11562 17000 11568
rect 16856 11280 16908 11286
rect 16856 11222 16908 11228
rect 16960 11218 16988 11562
rect 17040 11552 17092 11558
rect 17040 11494 17092 11500
rect 16948 11212 17000 11218
rect 16948 11154 17000 11160
rect 16948 11008 17000 11014
rect 16948 10950 17000 10956
rect 16544 10908 16852 10917
rect 16544 10906 16550 10908
rect 16606 10906 16630 10908
rect 16686 10906 16710 10908
rect 16766 10906 16790 10908
rect 16846 10906 16852 10908
rect 16606 10854 16608 10906
rect 16788 10854 16790 10906
rect 16544 10852 16550 10854
rect 16606 10852 16630 10854
rect 16686 10852 16710 10854
rect 16766 10852 16790 10854
rect 16846 10852 16852 10854
rect 16544 10843 16852 10852
rect 16960 10810 16988 10950
rect 16948 10804 17000 10810
rect 16948 10746 17000 10752
rect 16764 10736 16816 10742
rect 16764 10678 16816 10684
rect 16776 10577 16804 10678
rect 16762 10568 16818 10577
rect 16762 10503 16818 10512
rect 16776 10198 16804 10503
rect 16764 10192 16816 10198
rect 16764 10134 16816 10140
rect 16948 10056 17000 10062
rect 16948 9998 17000 10004
rect 16960 9926 16988 9998
rect 16948 9920 17000 9926
rect 16948 9862 17000 9868
rect 16544 9820 16852 9829
rect 16544 9818 16550 9820
rect 16606 9818 16630 9820
rect 16686 9818 16710 9820
rect 16766 9818 16790 9820
rect 16846 9818 16852 9820
rect 16606 9766 16608 9818
rect 16788 9766 16790 9818
rect 16544 9764 16550 9766
rect 16606 9764 16630 9766
rect 16686 9764 16710 9766
rect 16766 9764 16790 9766
rect 16846 9764 16852 9766
rect 16544 9755 16852 9764
rect 16960 9674 16988 9862
rect 16868 9646 16988 9674
rect 16868 9178 16896 9646
rect 16948 9512 17000 9518
rect 16948 9454 17000 9460
rect 16856 9172 16908 9178
rect 16856 9114 16908 9120
rect 16544 8732 16852 8741
rect 16544 8730 16550 8732
rect 16606 8730 16630 8732
rect 16686 8730 16710 8732
rect 16766 8730 16790 8732
rect 16846 8730 16852 8732
rect 16606 8678 16608 8730
rect 16788 8678 16790 8730
rect 16544 8676 16550 8678
rect 16606 8676 16630 8678
rect 16686 8676 16710 8678
rect 16766 8676 16790 8678
rect 16846 8676 16852 8678
rect 16544 8667 16852 8676
rect 16580 8424 16632 8430
rect 16580 8366 16632 8372
rect 16394 8256 16450 8265
rect 16394 8191 16450 8200
rect 16408 7721 16436 8191
rect 16592 8022 16620 8366
rect 16960 8362 16988 9454
rect 16948 8356 17000 8362
rect 16948 8298 17000 8304
rect 16580 8016 16632 8022
rect 16580 7958 16632 7964
rect 16394 7712 16450 7721
rect 16394 7647 16450 7656
rect 16544 7644 16852 7653
rect 16544 7642 16550 7644
rect 16606 7642 16630 7644
rect 16686 7642 16710 7644
rect 16766 7642 16790 7644
rect 16846 7642 16852 7644
rect 16606 7590 16608 7642
rect 16788 7590 16790 7642
rect 16544 7588 16550 7590
rect 16606 7588 16630 7590
rect 16686 7588 16710 7590
rect 16766 7588 16790 7590
rect 16846 7588 16852 7590
rect 16544 7579 16852 7588
rect 16396 7404 16448 7410
rect 16396 7346 16448 7352
rect 16304 6384 16356 6390
rect 16304 6326 16356 6332
rect 16212 6180 16264 6186
rect 16264 6140 16344 6168
rect 16212 6122 16264 6128
rect 16120 6112 16172 6118
rect 16120 6054 16172 6060
rect 16316 5642 16344 6140
rect 16304 5636 16356 5642
rect 16304 5578 16356 5584
rect 16210 5536 16266 5545
rect 16210 5471 16266 5480
rect 16118 4720 16174 4729
rect 16118 4655 16174 4664
rect 16132 4554 16160 4655
rect 16120 4548 16172 4554
rect 16120 4490 16172 4496
rect 16026 4176 16082 4185
rect 16026 4111 16082 4120
rect 15844 4072 15896 4078
rect 15844 4014 15896 4020
rect 15752 3392 15804 3398
rect 15856 3369 15884 4014
rect 16132 3738 16160 4490
rect 16120 3732 16172 3738
rect 16120 3674 16172 3680
rect 16028 3460 16080 3466
rect 16028 3402 16080 3408
rect 15752 3334 15804 3340
rect 15842 3360 15898 3369
rect 15842 3295 15898 3304
rect 15660 3120 15712 3126
rect 15660 3062 15712 3068
rect 15476 3052 15528 3058
rect 15476 2994 15528 3000
rect 15672 2922 15700 3062
rect 15384 2916 15436 2922
rect 15384 2858 15436 2864
rect 15660 2916 15712 2922
rect 15660 2858 15712 2864
rect 15476 2848 15528 2854
rect 15476 2790 15528 2796
rect 15936 2848 15988 2854
rect 15936 2790 15988 2796
rect 16040 2802 16068 3402
rect 16132 3058 16160 3674
rect 16224 3074 16252 5471
rect 16316 4690 16344 5578
rect 16408 5098 16436 7346
rect 16488 7336 16540 7342
rect 16488 7278 16540 7284
rect 16500 6866 16528 7278
rect 16488 6860 16540 6866
rect 16488 6802 16540 6808
rect 16960 6798 16988 8298
rect 16948 6792 17000 6798
rect 16948 6734 17000 6740
rect 16856 6656 16908 6662
rect 16908 6616 16988 6644
rect 17052 6633 17080 11494
rect 17144 10742 17172 13280
rect 17224 13252 17276 13258
rect 17224 13194 17276 13200
rect 17316 13252 17368 13258
rect 17316 13194 17368 13200
rect 17236 11762 17264 13194
rect 17328 12170 17356 13194
rect 17316 12164 17368 12170
rect 17316 12106 17368 12112
rect 17224 11756 17276 11762
rect 17224 11698 17276 11704
rect 17316 11552 17368 11558
rect 17316 11494 17368 11500
rect 17224 11212 17276 11218
rect 17224 11154 17276 11160
rect 17132 10736 17184 10742
rect 17132 10678 17184 10684
rect 17236 10606 17264 11154
rect 17224 10600 17276 10606
rect 17130 10568 17186 10577
rect 17224 10542 17276 10548
rect 17130 10503 17186 10512
rect 17144 10146 17172 10503
rect 17236 10266 17264 10542
rect 17224 10260 17276 10266
rect 17224 10202 17276 10208
rect 17144 10118 17264 10146
rect 17132 9580 17184 9586
rect 17132 9522 17184 9528
rect 17144 9178 17172 9522
rect 17132 9172 17184 9178
rect 17132 9114 17184 9120
rect 17132 9036 17184 9042
rect 17132 8978 17184 8984
rect 17144 8566 17172 8978
rect 17132 8560 17184 8566
rect 17132 8502 17184 8508
rect 17236 8344 17264 10118
rect 17328 9178 17356 11494
rect 17420 9602 17448 14282
rect 17512 13326 17540 16390
rect 17868 16176 17920 16182
rect 17868 16118 17920 16124
rect 17960 16176 18012 16182
rect 17960 16118 18012 16124
rect 17684 16108 17736 16114
rect 17684 16050 17736 16056
rect 17592 15904 17644 15910
rect 17592 15846 17644 15852
rect 17604 15609 17632 15846
rect 17590 15600 17646 15609
rect 17590 15535 17646 15544
rect 17500 13320 17552 13326
rect 17500 13262 17552 13268
rect 17592 13184 17644 13190
rect 17592 13126 17644 13132
rect 17604 12481 17632 13126
rect 17590 12472 17646 12481
rect 17590 12407 17592 12416
rect 17644 12407 17646 12416
rect 17592 12378 17644 12384
rect 17604 12347 17632 12378
rect 17592 12232 17644 12238
rect 17592 12174 17644 12180
rect 17500 11756 17552 11762
rect 17500 11698 17552 11704
rect 17512 9761 17540 11698
rect 17498 9752 17554 9761
rect 17498 9687 17554 9696
rect 17420 9574 17540 9602
rect 17408 9444 17460 9450
rect 17408 9386 17460 9392
rect 17316 9172 17368 9178
rect 17316 9114 17368 9120
rect 17420 9110 17448 9386
rect 17408 9104 17460 9110
rect 17408 9046 17460 9052
rect 17144 8316 17264 8344
rect 17144 7313 17172 8316
rect 17316 8084 17368 8090
rect 17316 8026 17368 8032
rect 17224 7948 17276 7954
rect 17224 7890 17276 7896
rect 17236 7324 17264 7890
rect 17328 7721 17356 8026
rect 17408 7880 17460 7886
rect 17408 7822 17460 7828
rect 17314 7712 17370 7721
rect 17314 7647 17370 7656
rect 17316 7336 17368 7342
rect 17130 7304 17186 7313
rect 17130 7239 17186 7248
rect 17236 7296 17316 7324
rect 16856 6598 16908 6604
rect 16544 6556 16852 6565
rect 16544 6554 16550 6556
rect 16606 6554 16630 6556
rect 16686 6554 16710 6556
rect 16766 6554 16790 6556
rect 16846 6554 16852 6556
rect 16606 6502 16608 6554
rect 16788 6502 16790 6554
rect 16544 6500 16550 6502
rect 16606 6500 16630 6502
rect 16686 6500 16710 6502
rect 16766 6500 16790 6502
rect 16846 6500 16852 6502
rect 16544 6491 16852 6500
rect 16580 6452 16632 6458
rect 16580 6394 16632 6400
rect 16592 5778 16620 6394
rect 16764 6384 16816 6390
rect 16764 6326 16816 6332
rect 16580 5772 16632 5778
rect 16580 5714 16632 5720
rect 16776 5710 16804 6326
rect 16764 5704 16816 5710
rect 16764 5646 16816 5652
rect 16776 5574 16804 5646
rect 16764 5568 16816 5574
rect 16764 5510 16816 5516
rect 16544 5468 16852 5477
rect 16544 5466 16550 5468
rect 16606 5466 16630 5468
rect 16686 5466 16710 5468
rect 16766 5466 16790 5468
rect 16846 5466 16852 5468
rect 16606 5414 16608 5466
rect 16788 5414 16790 5466
rect 16544 5412 16550 5414
rect 16606 5412 16630 5414
rect 16686 5412 16710 5414
rect 16766 5412 16790 5414
rect 16846 5412 16852 5414
rect 16544 5403 16852 5412
rect 16960 5302 16988 6616
rect 17038 6624 17094 6633
rect 17038 6559 17094 6568
rect 17040 6452 17092 6458
rect 17040 6394 17092 6400
rect 17052 6322 17080 6394
rect 17040 6316 17092 6322
rect 17040 6258 17092 6264
rect 17144 6186 17172 7239
rect 17040 6180 17092 6186
rect 17040 6122 17092 6128
rect 17132 6180 17184 6186
rect 17132 6122 17184 6128
rect 17052 5710 17080 6122
rect 17040 5704 17092 5710
rect 17040 5646 17092 5652
rect 16948 5296 17000 5302
rect 16578 5264 16634 5273
rect 16948 5238 17000 5244
rect 16578 5199 16634 5208
rect 16488 5160 16540 5166
rect 16486 5128 16488 5137
rect 16540 5128 16542 5137
rect 16396 5092 16448 5098
rect 16486 5063 16542 5072
rect 16396 5034 16448 5040
rect 16304 4684 16356 4690
rect 16304 4626 16356 4632
rect 16592 4622 16620 5199
rect 16960 4690 16988 5238
rect 16948 4684 17000 4690
rect 16948 4626 17000 4632
rect 16396 4616 16448 4622
rect 16316 4564 16396 4570
rect 16316 4558 16448 4564
rect 16580 4616 16632 4622
rect 16580 4558 16632 4564
rect 16762 4584 16818 4593
rect 16316 4542 16436 4558
rect 16316 4457 16344 4542
rect 16762 4519 16818 4528
rect 16948 4548 17000 4554
rect 16776 4486 16804 4519
rect 16948 4490 17000 4496
rect 16396 4480 16448 4486
rect 16302 4448 16358 4457
rect 16396 4422 16448 4428
rect 16764 4480 16816 4486
rect 16764 4422 16816 4428
rect 16302 4383 16358 4392
rect 16316 4026 16344 4383
rect 16408 4214 16436 4422
rect 16544 4380 16852 4389
rect 16544 4378 16550 4380
rect 16606 4378 16630 4380
rect 16686 4378 16710 4380
rect 16766 4378 16790 4380
rect 16846 4378 16852 4380
rect 16606 4326 16608 4378
rect 16788 4326 16790 4378
rect 16544 4324 16550 4326
rect 16606 4324 16630 4326
rect 16686 4324 16710 4326
rect 16766 4324 16790 4326
rect 16846 4324 16852 4326
rect 16544 4315 16852 4324
rect 16396 4208 16448 4214
rect 16396 4150 16448 4156
rect 16396 4072 16448 4078
rect 16316 4020 16396 4026
rect 16316 4014 16448 4020
rect 16316 3998 16436 4014
rect 16304 3936 16356 3942
rect 16304 3878 16356 3884
rect 16316 3738 16344 3878
rect 16304 3732 16356 3738
rect 16304 3674 16356 3680
rect 16408 3466 16436 3998
rect 16856 3936 16908 3942
rect 16856 3878 16908 3884
rect 16868 3466 16896 3878
rect 16396 3460 16448 3466
rect 16396 3402 16448 3408
rect 16856 3460 16908 3466
rect 16856 3402 16908 3408
rect 16304 3392 16356 3398
rect 16304 3334 16356 3340
rect 16316 3210 16344 3334
rect 16544 3292 16852 3301
rect 16544 3290 16550 3292
rect 16606 3290 16630 3292
rect 16686 3290 16710 3292
rect 16766 3290 16790 3292
rect 16846 3290 16852 3292
rect 16606 3238 16608 3290
rect 16788 3238 16790 3290
rect 16544 3236 16550 3238
rect 16606 3236 16630 3238
rect 16686 3236 16710 3238
rect 16766 3236 16790 3238
rect 16846 3236 16852 3238
rect 16544 3227 16852 3236
rect 16960 3210 16988 4490
rect 17052 4298 17080 5646
rect 17132 5568 17184 5574
rect 17132 5510 17184 5516
rect 17144 4978 17172 5510
rect 17236 5302 17264 7296
rect 17316 7278 17368 7284
rect 17316 5840 17368 5846
rect 17316 5782 17368 5788
rect 17224 5296 17276 5302
rect 17224 5238 17276 5244
rect 17328 5166 17356 5782
rect 17316 5160 17368 5166
rect 17316 5102 17368 5108
rect 17144 4950 17356 4978
rect 17222 4584 17278 4593
rect 17222 4519 17224 4528
rect 17276 4519 17278 4528
rect 17224 4490 17276 4496
rect 17052 4270 17172 4298
rect 17040 4208 17092 4214
rect 17040 4150 17092 4156
rect 17052 3534 17080 4150
rect 17040 3528 17092 3534
rect 17040 3470 17092 3476
rect 17144 3398 17172 4270
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 17236 3602 17264 4082
rect 17328 3641 17356 4950
rect 17314 3632 17370 3641
rect 17224 3596 17276 3602
rect 17314 3567 17370 3576
rect 17224 3538 17276 3544
rect 17132 3392 17184 3398
rect 17132 3334 17184 3340
rect 17314 3360 17370 3369
rect 17314 3295 17370 3304
rect 16316 3194 16436 3210
rect 16316 3188 16448 3194
rect 16316 3182 16396 3188
rect 16960 3182 17172 3210
rect 16396 3130 16448 3136
rect 16762 3088 16818 3097
rect 16224 3058 16528 3074
rect 16120 3052 16172 3058
rect 16224 3052 16540 3058
rect 16224 3046 16488 3052
rect 16120 2994 16172 3000
rect 16762 3023 16818 3032
rect 16946 3088 17002 3097
rect 16946 3023 16948 3032
rect 16488 2994 16540 3000
rect 16776 2990 16804 3023
rect 17000 3023 17002 3032
rect 16948 2994 17000 3000
rect 16764 2984 16816 2990
rect 16764 2926 16816 2932
rect 16672 2848 16724 2854
rect 16118 2816 16174 2825
rect 15292 2440 15344 2446
rect 15292 2382 15344 2388
rect 15488 800 15516 2790
rect 15844 2644 15896 2650
rect 15844 2586 15896 2592
rect 15660 2440 15712 2446
rect 15660 2382 15712 2388
rect 15672 2038 15700 2382
rect 15660 2032 15712 2038
rect 15660 1974 15712 1980
rect 15856 800 15884 2586
rect 15948 2514 15976 2790
rect 16040 2774 16118 2802
rect 16672 2790 16724 2796
rect 16118 2751 16174 2760
rect 15936 2508 15988 2514
rect 15936 2450 15988 2456
rect 16132 1290 16160 2751
rect 16212 2576 16264 2582
rect 16212 2518 16264 2524
rect 16120 1284 16172 1290
rect 16120 1226 16172 1232
rect 16224 800 16252 2518
rect 16684 2446 16712 2790
rect 16672 2440 16724 2446
rect 16672 2382 16724 2388
rect 17040 2372 17092 2378
rect 17040 2314 17092 2320
rect 16396 2304 16448 2310
rect 16396 2246 16448 2252
rect 16948 2304 17000 2310
rect 16948 2246 17000 2252
rect 16408 2106 16436 2246
rect 16544 2204 16852 2213
rect 16544 2202 16550 2204
rect 16606 2202 16630 2204
rect 16686 2202 16710 2204
rect 16766 2202 16790 2204
rect 16846 2202 16852 2204
rect 16606 2150 16608 2202
rect 16788 2150 16790 2202
rect 16544 2148 16550 2150
rect 16606 2148 16630 2150
rect 16686 2148 16710 2150
rect 16766 2148 16790 2150
rect 16846 2148 16852 2150
rect 16544 2139 16852 2148
rect 16396 2100 16448 2106
rect 16396 2042 16448 2048
rect 16960 1170 16988 2246
rect 16868 1142 16988 1170
rect 16592 870 16712 898
rect 16592 800 16620 870
rect 11532 734 11744 762
rect 11794 0 11850 800
rect 12162 0 12218 800
rect 12530 0 12586 800
rect 12898 0 12954 800
rect 13266 0 13322 800
rect 13634 0 13690 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15106 0 15162 800
rect 15474 0 15530 800
rect 15842 0 15898 800
rect 16210 0 16266 800
rect 16578 0 16634 800
rect 16684 762 16712 870
rect 16868 762 16896 1142
rect 17052 898 17080 2314
rect 17144 1358 17172 3182
rect 17328 3058 17356 3295
rect 17316 3052 17368 3058
rect 17316 2994 17368 3000
rect 17224 2848 17276 2854
rect 17224 2790 17276 2796
rect 17236 2446 17264 2790
rect 17316 2576 17368 2582
rect 17316 2518 17368 2524
rect 17224 2440 17276 2446
rect 17224 2382 17276 2388
rect 17132 1352 17184 1358
rect 17132 1294 17184 1300
rect 16960 870 17080 898
rect 16960 800 16988 870
rect 17328 800 17356 2518
rect 17420 2417 17448 7822
rect 17512 7290 17540 9574
rect 17604 8922 17632 12174
rect 17696 9382 17724 16050
rect 17776 15360 17828 15366
rect 17776 15302 17828 15308
rect 17788 14822 17816 15302
rect 17776 14816 17828 14822
rect 17776 14758 17828 14764
rect 17776 12368 17828 12374
rect 17776 12310 17828 12316
rect 17788 11830 17816 12310
rect 17880 12209 17908 16118
rect 17972 14074 18000 16118
rect 18064 15065 18092 16526
rect 18524 15638 18552 18294
rect 19340 18284 19392 18290
rect 19260 18244 19340 18272
rect 19260 18154 19288 18244
rect 19340 18226 19392 18232
rect 19248 18148 19300 18154
rect 19248 18090 19300 18096
rect 19143 17980 19451 17989
rect 19143 17978 19149 17980
rect 19205 17978 19229 17980
rect 19285 17978 19309 17980
rect 19365 17978 19389 17980
rect 19445 17978 19451 17980
rect 19205 17926 19207 17978
rect 19387 17926 19389 17978
rect 19143 17924 19149 17926
rect 19205 17924 19229 17926
rect 19285 17924 19309 17926
rect 19365 17924 19389 17926
rect 19445 17924 19451 17926
rect 19143 17915 19451 17924
rect 18788 17876 18840 17882
rect 19536 17864 19564 18414
rect 19614 18391 19616 18400
rect 19668 18391 19670 18400
rect 19616 18362 19668 18368
rect 19616 17876 19668 17882
rect 19536 17836 19616 17864
rect 18788 17818 18840 17824
rect 19616 17818 19668 17824
rect 18144 15632 18196 15638
rect 18142 15600 18144 15609
rect 18512 15632 18564 15638
rect 18196 15600 18198 15609
rect 18512 15574 18564 15580
rect 18142 15535 18198 15544
rect 18512 15496 18564 15502
rect 18326 15464 18382 15473
rect 18512 15438 18564 15444
rect 18604 15496 18656 15502
rect 18604 15438 18656 15444
rect 18326 15399 18382 15408
rect 18340 15366 18368 15399
rect 18328 15360 18380 15366
rect 18328 15302 18380 15308
rect 18524 15094 18552 15438
rect 18512 15088 18564 15094
rect 18050 15056 18106 15065
rect 18512 15030 18564 15036
rect 18050 14991 18106 15000
rect 18328 15020 18380 15026
rect 18328 14962 18380 14968
rect 18340 14822 18368 14962
rect 18524 14958 18552 15030
rect 18512 14952 18564 14958
rect 18512 14894 18564 14900
rect 18328 14816 18380 14822
rect 18328 14758 18380 14764
rect 17960 14068 18012 14074
rect 17960 14010 18012 14016
rect 18236 13932 18288 13938
rect 18236 13874 18288 13880
rect 18052 13864 18104 13870
rect 18052 13806 18104 13812
rect 18064 12986 18092 13806
rect 18248 13530 18276 13874
rect 18236 13524 18288 13530
rect 18236 13466 18288 13472
rect 18340 13410 18368 14758
rect 18524 14618 18552 14894
rect 18512 14612 18564 14618
rect 18512 14554 18564 14560
rect 18420 14408 18472 14414
rect 18420 14350 18472 14356
rect 18432 14278 18460 14350
rect 18420 14272 18472 14278
rect 18420 14214 18472 14220
rect 18248 13394 18368 13410
rect 18236 13388 18368 13394
rect 18288 13382 18368 13388
rect 18236 13330 18288 13336
rect 18052 12980 18104 12986
rect 18052 12922 18104 12928
rect 18142 12744 18198 12753
rect 18248 12714 18276 13330
rect 18328 13184 18380 13190
rect 18328 13126 18380 13132
rect 18340 12918 18368 13126
rect 18328 12912 18380 12918
rect 18328 12854 18380 12860
rect 18432 12782 18460 14214
rect 18420 12776 18472 12782
rect 18420 12718 18472 12724
rect 18142 12679 18198 12688
rect 18236 12708 18288 12714
rect 18156 12434 18184 12679
rect 18236 12650 18288 12656
rect 17972 12406 18184 12434
rect 17866 12200 17922 12209
rect 17866 12135 17922 12144
rect 17776 11824 17828 11830
rect 17776 11766 17828 11772
rect 17866 11656 17922 11665
rect 17866 11591 17922 11600
rect 17776 11552 17828 11558
rect 17776 11494 17828 11500
rect 17788 10742 17816 11494
rect 17880 10810 17908 11591
rect 17868 10804 17920 10810
rect 17868 10746 17920 10752
rect 17776 10736 17828 10742
rect 17776 10678 17828 10684
rect 17866 10704 17922 10713
rect 17866 10639 17922 10648
rect 17776 10600 17828 10606
rect 17776 10542 17828 10548
rect 17788 10033 17816 10542
rect 17774 10024 17830 10033
rect 17774 9959 17830 9968
rect 17776 9512 17828 9518
rect 17774 9480 17776 9489
rect 17828 9480 17830 9489
rect 17774 9415 17830 9424
rect 17684 9376 17736 9382
rect 17684 9318 17736 9324
rect 17776 9376 17828 9382
rect 17776 9318 17828 9324
rect 17604 8894 17724 8922
rect 17590 7848 17646 7857
rect 17590 7783 17646 7792
rect 17604 7750 17632 7783
rect 17592 7744 17644 7750
rect 17592 7686 17644 7692
rect 17512 7262 17632 7290
rect 17500 7200 17552 7206
rect 17500 7142 17552 7148
rect 17512 5370 17540 7142
rect 17604 6440 17632 7262
rect 17696 7206 17724 8894
rect 17788 7274 17816 9318
rect 17880 7834 17908 10639
rect 17972 9738 18000 12406
rect 18248 12306 18276 12650
rect 18328 12640 18380 12646
rect 18328 12582 18380 12588
rect 18340 12442 18368 12582
rect 18328 12436 18380 12442
rect 18616 12434 18644 15438
rect 18696 15360 18748 15366
rect 18696 15302 18748 15308
rect 18708 13297 18736 15302
rect 18800 14550 18828 17818
rect 19628 17338 19656 17818
rect 19720 17814 19748 20402
rect 19812 19009 19840 20402
rect 19904 19496 19932 20760
rect 19984 20596 20036 20602
rect 19984 20538 20036 20544
rect 19996 20505 20024 20538
rect 19982 20496 20038 20505
rect 19982 20431 20038 20440
rect 20088 20058 20116 22200
rect 20258 20904 20314 20913
rect 20258 20839 20314 20848
rect 20168 20256 20220 20262
rect 20168 20198 20220 20204
rect 20076 20052 20128 20058
rect 20076 19994 20128 20000
rect 20076 19508 20128 19514
rect 19904 19468 20024 19496
rect 19892 19372 19944 19378
rect 19892 19314 19944 19320
rect 19798 19000 19854 19009
rect 19798 18935 19854 18944
rect 19904 18816 19932 19314
rect 19996 19145 20024 19468
rect 20076 19450 20128 19456
rect 20088 19417 20116 19450
rect 20180 19446 20208 20198
rect 20272 19922 20300 20839
rect 20352 20256 20404 20262
rect 20350 20224 20352 20233
rect 20404 20224 20406 20233
rect 20350 20159 20406 20168
rect 20260 19916 20312 19922
rect 20260 19858 20312 19864
rect 20456 19854 20484 22200
rect 20534 21448 20590 21457
rect 20534 21383 20590 21392
rect 20444 19848 20496 19854
rect 20444 19790 20496 19796
rect 20260 19780 20312 19786
rect 20260 19722 20312 19728
rect 20272 19446 20300 19722
rect 20168 19440 20220 19446
rect 20074 19408 20130 19417
rect 20168 19382 20220 19388
rect 20260 19440 20312 19446
rect 20260 19382 20312 19388
rect 20074 19343 20130 19352
rect 19982 19136 20038 19145
rect 19982 19071 20038 19080
rect 19812 18788 19932 18816
rect 19812 18714 19840 18788
rect 19984 18760 20036 18766
rect 19812 18686 19932 18714
rect 19984 18702 20036 18708
rect 19798 18456 19854 18465
rect 19904 18426 19932 18686
rect 19798 18391 19800 18400
rect 19852 18391 19854 18400
rect 19892 18420 19944 18426
rect 19800 18362 19852 18368
rect 19892 18362 19944 18368
rect 19798 18320 19854 18329
rect 19798 18255 19854 18264
rect 19708 17808 19760 17814
rect 19708 17750 19760 17756
rect 19708 17604 19760 17610
rect 19812 17592 19840 18255
rect 19996 17746 20024 18702
rect 19984 17740 20036 17746
rect 19984 17682 20036 17688
rect 19760 17564 19840 17592
rect 19708 17546 19760 17552
rect 19616 17332 19668 17338
rect 19616 17274 19668 17280
rect 18972 17196 19024 17202
rect 18972 17138 19024 17144
rect 18984 16046 19012 17138
rect 19616 16992 19668 16998
rect 19616 16934 19668 16940
rect 19143 16892 19451 16901
rect 19143 16890 19149 16892
rect 19205 16890 19229 16892
rect 19285 16890 19309 16892
rect 19365 16890 19389 16892
rect 19445 16890 19451 16892
rect 19205 16838 19207 16890
rect 19387 16838 19389 16890
rect 19143 16836 19149 16838
rect 19205 16836 19229 16838
rect 19285 16836 19309 16838
rect 19365 16836 19389 16838
rect 19445 16836 19451 16838
rect 19143 16827 19451 16836
rect 19524 16788 19576 16794
rect 19524 16730 19576 16736
rect 18972 16040 19024 16046
rect 18972 15982 19024 15988
rect 19064 16040 19116 16046
rect 19064 15982 19116 15988
rect 18880 15904 18932 15910
rect 18880 15846 18932 15852
rect 18892 15366 18920 15846
rect 18880 15360 18932 15366
rect 19076 15337 19104 15982
rect 19143 15804 19451 15813
rect 19143 15802 19149 15804
rect 19205 15802 19229 15804
rect 19285 15802 19309 15804
rect 19365 15802 19389 15804
rect 19445 15802 19451 15804
rect 19205 15750 19207 15802
rect 19387 15750 19389 15802
rect 19143 15748 19149 15750
rect 19205 15748 19229 15750
rect 19285 15748 19309 15750
rect 19365 15748 19389 15750
rect 19445 15748 19451 15750
rect 19143 15739 19451 15748
rect 19536 15638 19564 16730
rect 19628 16017 19656 16934
rect 19720 16538 19748 17546
rect 19996 16794 20024 17682
rect 20088 17678 20116 19343
rect 20180 18290 20208 19382
rect 20456 19378 20484 19790
rect 20548 19514 20576 21383
rect 20720 20460 20772 20466
rect 20720 20402 20772 20408
rect 20536 19508 20588 19514
rect 20536 19450 20588 19456
rect 20444 19372 20496 19378
rect 20496 19320 20576 19334
rect 20444 19314 20576 19320
rect 20456 19306 20576 19314
rect 20260 19236 20312 19242
rect 20260 19178 20312 19184
rect 20272 18340 20300 19178
rect 20548 18834 20576 19306
rect 20628 19304 20680 19310
rect 20628 19246 20680 19252
rect 20536 18828 20588 18834
rect 20456 18788 20536 18816
rect 20272 18312 20392 18340
rect 20168 18284 20220 18290
rect 20220 18244 20300 18272
rect 20168 18226 20220 18232
rect 20168 18148 20220 18154
rect 20168 18090 20220 18096
rect 20076 17672 20128 17678
rect 20076 17614 20128 17620
rect 20180 17542 20208 18090
rect 20272 17678 20300 18244
rect 20260 17672 20312 17678
rect 20260 17614 20312 17620
rect 20168 17536 20220 17542
rect 20168 17478 20220 17484
rect 19984 16788 20036 16794
rect 19984 16730 20036 16736
rect 19800 16652 19852 16658
rect 20260 16652 20312 16658
rect 19852 16612 20024 16640
rect 19800 16594 19852 16600
rect 19720 16510 19932 16538
rect 19708 16176 19760 16182
rect 19706 16144 19708 16153
rect 19760 16144 19762 16153
rect 19706 16079 19762 16088
rect 19800 16108 19852 16114
rect 19800 16050 19852 16056
rect 19614 16008 19670 16017
rect 19614 15943 19670 15952
rect 19812 15910 19840 16050
rect 19616 15904 19668 15910
rect 19616 15846 19668 15852
rect 19800 15904 19852 15910
rect 19800 15846 19852 15852
rect 19628 15706 19656 15846
rect 19616 15700 19668 15706
rect 19616 15642 19668 15648
rect 19524 15632 19576 15638
rect 19524 15574 19576 15580
rect 18880 15302 18932 15308
rect 19062 15328 19118 15337
rect 18788 14544 18840 14550
rect 18788 14486 18840 14492
rect 18800 14278 18828 14486
rect 18788 14272 18840 14278
rect 18788 14214 18840 14220
rect 18892 13433 18920 15302
rect 19062 15263 19118 15272
rect 19536 15094 19564 15574
rect 19628 15366 19656 15642
rect 19708 15496 19760 15502
rect 19708 15438 19760 15444
rect 19616 15360 19668 15366
rect 19616 15302 19668 15308
rect 19524 15088 19576 15094
rect 19524 15030 19576 15036
rect 19064 15020 19116 15026
rect 19064 14962 19116 14968
rect 19076 14929 19104 14962
rect 19062 14920 19118 14929
rect 19062 14855 19118 14864
rect 19524 14816 19576 14822
rect 19524 14758 19576 14764
rect 19143 14716 19451 14725
rect 19143 14714 19149 14716
rect 19205 14714 19229 14716
rect 19285 14714 19309 14716
rect 19365 14714 19389 14716
rect 19445 14714 19451 14716
rect 19205 14662 19207 14714
rect 19387 14662 19389 14714
rect 19143 14660 19149 14662
rect 19205 14660 19229 14662
rect 19285 14660 19309 14662
rect 19365 14660 19389 14662
rect 19445 14660 19451 14662
rect 19143 14651 19451 14660
rect 19536 14482 19564 14758
rect 19524 14476 19576 14482
rect 19524 14418 19576 14424
rect 19536 14006 19564 14418
rect 19628 14346 19656 15302
rect 19616 14340 19668 14346
rect 19616 14282 19668 14288
rect 19524 14000 19576 14006
rect 19524 13942 19576 13948
rect 19143 13628 19451 13637
rect 19143 13626 19149 13628
rect 19205 13626 19229 13628
rect 19285 13626 19309 13628
rect 19365 13626 19389 13628
rect 19445 13626 19451 13628
rect 19205 13574 19207 13626
rect 19387 13574 19389 13626
rect 19143 13572 19149 13574
rect 19205 13572 19229 13574
rect 19285 13572 19309 13574
rect 19365 13572 19389 13574
rect 19445 13572 19451 13574
rect 19143 13563 19451 13572
rect 18878 13424 18934 13433
rect 18788 13388 18840 13394
rect 19536 13394 19564 13942
rect 19720 13530 19748 15438
rect 19904 14618 19932 16510
rect 19892 14612 19944 14618
rect 19892 14554 19944 14560
rect 19800 14544 19852 14550
rect 19800 14486 19852 14492
rect 19812 14414 19840 14486
rect 19800 14408 19852 14414
rect 19800 14350 19852 14356
rect 19812 13938 19840 14350
rect 19800 13932 19852 13938
rect 19800 13874 19852 13880
rect 19708 13524 19760 13530
rect 19708 13466 19760 13472
rect 18878 13359 18934 13368
rect 19524 13388 19576 13394
rect 18788 13330 18840 13336
rect 19524 13330 19576 13336
rect 18694 13288 18750 13297
rect 18694 13223 18750 13232
rect 18696 13184 18748 13190
rect 18696 13126 18748 13132
rect 18708 12442 18736 13126
rect 18800 12782 18828 13330
rect 19892 13320 19944 13326
rect 19892 13262 19944 13268
rect 19064 13252 19116 13258
rect 19064 13194 19116 13200
rect 18788 12776 18840 12782
rect 18788 12718 18840 12724
rect 18328 12378 18380 12384
rect 18432 12406 18644 12434
rect 18696 12436 18748 12442
rect 18236 12300 18288 12306
rect 18236 12242 18288 12248
rect 18052 12164 18104 12170
rect 18052 12106 18104 12112
rect 18064 11898 18092 12106
rect 18144 12096 18196 12102
rect 18144 12038 18196 12044
rect 18052 11892 18104 11898
rect 18052 11834 18104 11840
rect 18050 11656 18106 11665
rect 18050 11591 18052 11600
rect 18104 11591 18106 11600
rect 18052 11562 18104 11568
rect 18052 11008 18104 11014
rect 18052 10950 18104 10956
rect 18064 9926 18092 10950
rect 18156 10577 18184 12038
rect 18328 11892 18380 11898
rect 18328 11834 18380 11840
rect 18340 11762 18368 11834
rect 18328 11756 18380 11762
rect 18328 11698 18380 11704
rect 18236 11552 18288 11558
rect 18236 11494 18288 11500
rect 18248 10606 18276 11494
rect 18328 10668 18380 10674
rect 18328 10610 18380 10616
rect 18236 10600 18288 10606
rect 18142 10568 18198 10577
rect 18236 10542 18288 10548
rect 18142 10503 18198 10512
rect 18144 10464 18196 10470
rect 18144 10406 18196 10412
rect 18052 9920 18104 9926
rect 18052 9862 18104 9868
rect 17972 9710 18092 9738
rect 18064 9625 18092 9710
rect 18050 9616 18106 9625
rect 17960 9580 18012 9586
rect 18156 9602 18184 10406
rect 18248 9722 18276 10542
rect 18340 9722 18368 10610
rect 18432 10305 18460 12406
rect 18696 12378 18748 12384
rect 18604 12232 18656 12238
rect 18604 12174 18656 12180
rect 18616 11014 18644 12174
rect 18972 12164 19024 12170
rect 19076 12152 19104 13194
rect 19904 12986 19932 13262
rect 19892 12980 19944 12986
rect 19892 12922 19944 12928
rect 19432 12776 19484 12782
rect 19432 12718 19484 12724
rect 19616 12776 19668 12782
rect 19616 12718 19668 12724
rect 19444 12646 19472 12718
rect 19432 12640 19484 12646
rect 19432 12582 19484 12588
rect 19143 12540 19451 12549
rect 19143 12538 19149 12540
rect 19205 12538 19229 12540
rect 19285 12538 19309 12540
rect 19365 12538 19389 12540
rect 19445 12538 19451 12540
rect 19205 12486 19207 12538
rect 19387 12486 19389 12538
rect 19143 12484 19149 12486
rect 19205 12484 19229 12486
rect 19285 12484 19309 12486
rect 19365 12484 19389 12486
rect 19445 12484 19451 12486
rect 19143 12475 19451 12484
rect 19246 12336 19302 12345
rect 19246 12271 19302 12280
rect 19076 12124 19196 12152
rect 18972 12106 19024 12112
rect 18880 12096 18932 12102
rect 18880 12038 18932 12044
rect 18696 11892 18748 11898
rect 18696 11834 18748 11840
rect 18708 11082 18736 11834
rect 18788 11756 18840 11762
rect 18788 11698 18840 11704
rect 18696 11076 18748 11082
rect 18696 11018 18748 11024
rect 18604 11008 18656 11014
rect 18604 10950 18656 10956
rect 18512 10600 18564 10606
rect 18708 10554 18736 11018
rect 18800 10810 18828 11698
rect 18788 10804 18840 10810
rect 18788 10746 18840 10752
rect 18788 10668 18840 10674
rect 18788 10610 18840 10616
rect 18564 10548 18736 10554
rect 18512 10542 18736 10548
rect 18524 10526 18736 10542
rect 18418 10296 18474 10305
rect 18524 10266 18552 10526
rect 18604 10464 18656 10470
rect 18604 10406 18656 10412
rect 18418 10231 18474 10240
rect 18512 10260 18564 10266
rect 18512 10202 18564 10208
rect 18418 10160 18474 10169
rect 18418 10095 18474 10104
rect 18236 9716 18288 9722
rect 18236 9658 18288 9664
rect 18328 9716 18380 9722
rect 18328 9658 18380 9664
rect 18156 9574 18276 9602
rect 18050 9551 18106 9560
rect 17960 9522 18012 9528
rect 17972 8090 18000 9522
rect 18052 9512 18104 9518
rect 18052 9454 18104 9460
rect 18144 9512 18196 9518
rect 18144 9454 18196 9460
rect 18064 8634 18092 9454
rect 18156 9042 18184 9454
rect 18144 9036 18196 9042
rect 18144 8978 18196 8984
rect 18144 8900 18196 8906
rect 18144 8842 18196 8848
rect 18052 8628 18104 8634
rect 18052 8570 18104 8576
rect 18156 8294 18184 8842
rect 18248 8514 18276 9574
rect 18340 9382 18368 9658
rect 18328 9376 18380 9382
rect 18328 9318 18380 9324
rect 18326 9208 18382 9217
rect 18326 9143 18382 9152
rect 18340 8945 18368 9143
rect 18326 8936 18382 8945
rect 18326 8871 18382 8880
rect 18328 8832 18380 8838
rect 18328 8774 18380 8780
rect 18340 8634 18368 8774
rect 18432 8634 18460 10095
rect 18512 9920 18564 9926
rect 18512 9862 18564 9868
rect 18328 8628 18380 8634
rect 18328 8570 18380 8576
rect 18420 8628 18472 8634
rect 18420 8570 18472 8576
rect 18248 8486 18368 8514
rect 18236 8356 18288 8362
rect 18236 8298 18288 8304
rect 18144 8288 18196 8294
rect 18144 8230 18196 8236
rect 17960 8084 18012 8090
rect 17960 8026 18012 8032
rect 18142 7984 18198 7993
rect 18142 7919 18198 7928
rect 17880 7806 18092 7834
rect 17960 7744 18012 7750
rect 17880 7704 17960 7732
rect 17776 7268 17828 7274
rect 17776 7210 17828 7216
rect 17684 7200 17736 7206
rect 17684 7142 17736 7148
rect 17604 6412 17724 6440
rect 17592 6316 17644 6322
rect 17592 6258 17644 6264
rect 17604 5846 17632 6258
rect 17592 5840 17644 5846
rect 17592 5782 17644 5788
rect 17500 5364 17552 5370
rect 17500 5306 17552 5312
rect 17592 5228 17644 5234
rect 17592 5170 17644 5176
rect 17500 3392 17552 3398
rect 17500 3334 17552 3340
rect 17406 2408 17462 2417
rect 17406 2343 17462 2352
rect 17512 2038 17540 3334
rect 17604 3194 17632 5170
rect 17696 4826 17724 6412
rect 17684 4820 17736 4826
rect 17684 4762 17736 4768
rect 17696 4690 17724 4762
rect 17684 4684 17736 4690
rect 17684 4626 17736 4632
rect 17696 4282 17724 4626
rect 17788 4554 17816 7210
rect 17880 5710 17908 7704
rect 17960 7686 18012 7692
rect 18064 7585 18092 7806
rect 18050 7576 18106 7585
rect 18156 7546 18184 7919
rect 18050 7511 18106 7520
rect 18144 7540 18196 7546
rect 18144 7482 18196 7488
rect 18144 7336 18196 7342
rect 18144 7278 18196 7284
rect 18050 7032 18106 7041
rect 18050 6967 18106 6976
rect 17958 6896 18014 6905
rect 17958 6831 18014 6840
rect 17972 6662 18000 6831
rect 17960 6656 18012 6662
rect 17960 6598 18012 6604
rect 17958 6488 18014 6497
rect 17958 6423 18014 6432
rect 17972 5817 18000 6423
rect 17958 5808 18014 5817
rect 17958 5743 18014 5752
rect 17868 5704 17920 5710
rect 17868 5646 17920 5652
rect 17868 5568 17920 5574
rect 17866 5536 17868 5545
rect 17920 5536 17922 5545
rect 17866 5471 17922 5480
rect 18064 4690 18092 6967
rect 18156 6730 18184 7278
rect 18144 6724 18196 6730
rect 18144 6666 18196 6672
rect 18156 5642 18184 6666
rect 18144 5636 18196 5642
rect 18144 5578 18196 5584
rect 18248 5234 18276 8298
rect 18340 7002 18368 8486
rect 18420 8492 18472 8498
rect 18420 8434 18472 8440
rect 18432 8090 18460 8434
rect 18524 8430 18552 9862
rect 18616 8974 18644 10406
rect 18694 10296 18750 10305
rect 18694 10231 18750 10240
rect 18708 10062 18736 10231
rect 18696 10056 18748 10062
rect 18696 9998 18748 10004
rect 18800 9926 18828 10610
rect 18696 9920 18748 9926
rect 18694 9888 18696 9897
rect 18788 9920 18840 9926
rect 18748 9888 18750 9897
rect 18788 9862 18840 9868
rect 18694 9823 18750 9832
rect 18708 9382 18736 9823
rect 18892 9738 18920 12038
rect 18984 10577 19012 12106
rect 19168 11694 19196 12124
rect 19260 11830 19288 12271
rect 19340 12096 19392 12102
rect 19340 12038 19392 12044
rect 19248 11824 19300 11830
rect 19352 11801 19380 12038
rect 19628 11937 19656 12718
rect 19800 12232 19852 12238
rect 19800 12174 19852 12180
rect 19614 11928 19670 11937
rect 19614 11863 19670 11872
rect 19524 11824 19576 11830
rect 19248 11766 19300 11772
rect 19338 11792 19394 11801
rect 19524 11766 19576 11772
rect 19338 11727 19394 11736
rect 19156 11688 19208 11694
rect 19156 11630 19208 11636
rect 19536 11558 19564 11766
rect 19524 11552 19576 11558
rect 19524 11494 19576 11500
rect 19143 11452 19451 11461
rect 19143 11450 19149 11452
rect 19205 11450 19229 11452
rect 19285 11450 19309 11452
rect 19365 11450 19389 11452
rect 19445 11450 19451 11452
rect 19205 11398 19207 11450
rect 19387 11398 19389 11450
rect 19143 11396 19149 11398
rect 19205 11396 19229 11398
rect 19285 11396 19309 11398
rect 19365 11396 19389 11398
rect 19445 11396 19451 11398
rect 19143 11387 19451 11396
rect 19248 11280 19300 11286
rect 19246 11248 19248 11257
rect 19300 11248 19302 11257
rect 19246 11183 19302 11192
rect 19156 11144 19208 11150
rect 19156 11086 19208 11092
rect 18970 10568 19026 10577
rect 18970 10503 19026 10512
rect 19168 10452 19196 11086
rect 19628 10810 19656 11863
rect 19812 11830 19840 12174
rect 19800 11824 19852 11830
rect 19800 11766 19852 11772
rect 19812 11014 19840 11766
rect 19892 11348 19944 11354
rect 19892 11290 19944 11296
rect 19904 11082 19932 11290
rect 19892 11076 19944 11082
rect 19892 11018 19944 11024
rect 19800 11008 19852 11014
rect 19800 10950 19852 10956
rect 19616 10804 19668 10810
rect 19616 10746 19668 10752
rect 19524 10668 19576 10674
rect 19524 10610 19576 10616
rect 18984 10424 19196 10452
rect 18984 9874 19012 10424
rect 19143 10364 19451 10373
rect 19143 10362 19149 10364
rect 19205 10362 19229 10364
rect 19285 10362 19309 10364
rect 19365 10362 19389 10364
rect 19445 10362 19451 10364
rect 19205 10310 19207 10362
rect 19387 10310 19389 10362
rect 19143 10308 19149 10310
rect 19205 10308 19229 10310
rect 19285 10308 19309 10310
rect 19365 10308 19389 10310
rect 19445 10308 19451 10310
rect 19143 10299 19451 10308
rect 18984 9846 19288 9874
rect 18892 9710 19012 9738
rect 18984 9674 19012 9710
rect 18984 9646 19104 9674
rect 18878 9616 18934 9625
rect 18788 9580 18840 9586
rect 18878 9551 18934 9560
rect 18788 9522 18840 9528
rect 18696 9376 18748 9382
rect 18694 9344 18696 9353
rect 18748 9344 18750 9353
rect 18694 9279 18750 9288
rect 18800 9178 18828 9522
rect 18892 9217 18920 9551
rect 18878 9208 18934 9217
rect 18696 9172 18748 9178
rect 18696 9114 18748 9120
rect 18788 9172 18840 9178
rect 18878 9143 18934 9152
rect 18788 9114 18840 9120
rect 18604 8968 18656 8974
rect 18604 8910 18656 8916
rect 18512 8424 18564 8430
rect 18512 8366 18564 8372
rect 18510 8256 18566 8265
rect 18510 8191 18566 8200
rect 18420 8084 18472 8090
rect 18420 8026 18472 8032
rect 18328 6996 18380 7002
rect 18328 6938 18380 6944
rect 18328 6860 18380 6866
rect 18432 6848 18460 8026
rect 18380 6820 18460 6848
rect 18328 6802 18380 6808
rect 18328 6656 18380 6662
rect 18328 6598 18380 6604
rect 18340 5914 18368 6598
rect 18432 6390 18460 6820
rect 18420 6384 18472 6390
rect 18420 6326 18472 6332
rect 18432 5914 18460 6326
rect 18328 5908 18380 5914
rect 18328 5850 18380 5856
rect 18420 5908 18472 5914
rect 18420 5850 18472 5856
rect 18524 5273 18552 8191
rect 18616 7954 18644 8910
rect 18708 8537 18736 9114
rect 18788 9036 18840 9042
rect 18788 8978 18840 8984
rect 18800 8945 18828 8978
rect 18786 8936 18842 8945
rect 18786 8871 18842 8880
rect 18788 8832 18840 8838
rect 18788 8774 18840 8780
rect 18800 8634 18828 8774
rect 18892 8634 18920 9143
rect 19076 8974 19104 9646
rect 19260 9602 19288 9846
rect 19536 9722 19564 10610
rect 19812 10606 19840 10950
rect 19616 10600 19668 10606
rect 19616 10542 19668 10548
rect 19800 10600 19852 10606
rect 19800 10542 19852 10548
rect 19628 10266 19656 10542
rect 19708 10464 19760 10470
rect 19708 10406 19760 10412
rect 19616 10260 19668 10266
rect 19616 10202 19668 10208
rect 19720 10130 19748 10406
rect 19708 10124 19760 10130
rect 19708 10066 19760 10072
rect 19800 10124 19852 10130
rect 19904 10112 19932 11018
rect 19852 10084 19932 10112
rect 19800 10066 19852 10072
rect 19812 10010 19840 10066
rect 19720 9982 19840 10010
rect 19524 9716 19576 9722
rect 19524 9658 19576 9664
rect 19260 9574 19564 9602
rect 19143 9276 19451 9285
rect 19143 9274 19149 9276
rect 19205 9274 19229 9276
rect 19285 9274 19309 9276
rect 19365 9274 19389 9276
rect 19445 9274 19451 9276
rect 19205 9222 19207 9274
rect 19387 9222 19389 9274
rect 19143 9220 19149 9222
rect 19205 9220 19229 9222
rect 19285 9220 19309 9222
rect 19365 9220 19389 9222
rect 19445 9220 19451 9222
rect 19143 9211 19451 9220
rect 19064 8968 19116 8974
rect 18970 8936 19026 8945
rect 19064 8910 19116 8916
rect 18970 8871 18972 8880
rect 19024 8871 19026 8880
rect 18972 8842 19024 8848
rect 18788 8628 18840 8634
rect 18788 8570 18840 8576
rect 18880 8628 18932 8634
rect 18880 8570 18932 8576
rect 18984 8566 19012 8842
rect 18972 8560 19024 8566
rect 18694 8528 18750 8537
rect 18972 8502 19024 8508
rect 18694 8463 18750 8472
rect 18880 8492 18932 8498
rect 18880 8434 18932 8440
rect 18696 8288 18748 8294
rect 18696 8230 18748 8236
rect 18604 7948 18656 7954
rect 18604 7890 18656 7896
rect 18708 7546 18736 8230
rect 18892 8129 18920 8434
rect 19076 8294 19104 8910
rect 19248 8832 19300 8838
rect 19248 8774 19300 8780
rect 19260 8498 19288 8774
rect 19340 8628 19392 8634
rect 19340 8570 19392 8576
rect 19248 8492 19300 8498
rect 19248 8434 19300 8440
rect 19352 8401 19380 8570
rect 19338 8392 19394 8401
rect 19338 8327 19394 8336
rect 19064 8288 19116 8294
rect 19064 8230 19116 8236
rect 18878 8120 18934 8129
rect 18878 8055 18934 8064
rect 18696 7540 18748 7546
rect 18696 7482 18748 7488
rect 18604 7472 18656 7478
rect 18604 7414 18656 7420
rect 18616 6458 18644 7414
rect 18788 6860 18840 6866
rect 18788 6802 18840 6808
rect 18696 6792 18748 6798
rect 18696 6734 18748 6740
rect 18604 6452 18656 6458
rect 18604 6394 18656 6400
rect 18616 6254 18644 6394
rect 18604 6248 18656 6254
rect 18604 6190 18656 6196
rect 18510 5264 18566 5273
rect 18236 5228 18288 5234
rect 18236 5170 18288 5176
rect 18420 5228 18472 5234
rect 18510 5199 18566 5208
rect 18420 5170 18472 5176
rect 18248 4826 18276 5170
rect 18236 4820 18288 4826
rect 18236 4762 18288 4768
rect 18052 4684 18104 4690
rect 18052 4626 18104 4632
rect 17776 4548 17828 4554
rect 17776 4490 17828 4496
rect 17960 4480 18012 4486
rect 17774 4448 17830 4457
rect 17960 4422 18012 4428
rect 17774 4383 17830 4392
rect 17684 4276 17736 4282
rect 17684 4218 17736 4224
rect 17682 3768 17738 3777
rect 17682 3703 17738 3712
rect 17696 3398 17724 3703
rect 17684 3392 17736 3398
rect 17684 3334 17736 3340
rect 17592 3188 17644 3194
rect 17592 3130 17644 3136
rect 17788 2961 17816 4383
rect 17868 3460 17920 3466
rect 17868 3402 17920 3408
rect 17880 3058 17908 3402
rect 17972 3233 18000 4422
rect 18248 4214 18276 4762
rect 18328 4480 18380 4486
rect 18328 4422 18380 4428
rect 18236 4208 18288 4214
rect 18236 4150 18288 4156
rect 18340 3602 18368 4422
rect 18432 4282 18460 5170
rect 18524 5114 18552 5199
rect 18524 5086 18644 5114
rect 18512 5024 18564 5030
rect 18512 4966 18564 4972
rect 18420 4276 18472 4282
rect 18420 4218 18472 4224
rect 18432 4078 18460 4218
rect 18420 4072 18472 4078
rect 18420 4014 18472 4020
rect 18432 3670 18460 4014
rect 18420 3664 18472 3670
rect 18420 3606 18472 3612
rect 18328 3596 18380 3602
rect 18328 3538 18380 3544
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 18144 3392 18196 3398
rect 18144 3334 18196 3340
rect 17958 3224 18014 3233
rect 18156 3194 18184 3334
rect 17958 3159 18014 3168
rect 18144 3188 18196 3194
rect 18144 3130 18196 3136
rect 17960 3120 18012 3126
rect 17960 3062 18012 3068
rect 17868 3052 17920 3058
rect 17868 2994 17920 3000
rect 17774 2952 17830 2961
rect 17774 2887 17830 2896
rect 17684 2644 17736 2650
rect 17684 2586 17736 2592
rect 17500 2032 17552 2038
rect 17500 1974 17552 1980
rect 17696 800 17724 2586
rect 17972 2446 18000 3062
rect 18052 2848 18104 2854
rect 18052 2790 18104 2796
rect 17960 2440 18012 2446
rect 17960 2382 18012 2388
rect 18064 800 18092 2790
rect 18248 2530 18276 3470
rect 18156 2514 18276 2530
rect 18420 2576 18472 2582
rect 18420 2518 18472 2524
rect 18144 2508 18276 2514
rect 18196 2502 18276 2508
rect 18144 2450 18196 2456
rect 18328 2440 18380 2446
rect 18328 2382 18380 2388
rect 18340 2106 18368 2382
rect 18328 2100 18380 2106
rect 18328 2042 18380 2048
rect 18432 800 18460 2518
rect 18524 2446 18552 4966
rect 18616 4486 18644 5086
rect 18604 4480 18656 4486
rect 18604 4422 18656 4428
rect 18708 4298 18736 6734
rect 18800 6322 18828 6802
rect 18892 6780 18920 8055
rect 19076 7886 19104 8230
rect 19143 8188 19451 8197
rect 19143 8186 19149 8188
rect 19205 8186 19229 8188
rect 19285 8186 19309 8188
rect 19365 8186 19389 8188
rect 19445 8186 19451 8188
rect 19205 8134 19207 8186
rect 19387 8134 19389 8186
rect 19143 8132 19149 8134
rect 19205 8132 19229 8134
rect 19285 8132 19309 8134
rect 19365 8132 19389 8134
rect 19445 8132 19451 8134
rect 19143 8123 19451 8132
rect 18972 7880 19024 7886
rect 18972 7822 19024 7828
rect 19064 7880 19116 7886
rect 19064 7822 19116 7828
rect 18984 6934 19012 7822
rect 19340 7744 19392 7750
rect 19340 7686 19392 7692
rect 19352 7342 19380 7686
rect 19536 7528 19564 9574
rect 19616 9580 19668 9586
rect 19616 9522 19668 9528
rect 19628 9450 19656 9522
rect 19616 9444 19668 9450
rect 19616 9386 19668 9392
rect 19720 9382 19748 9982
rect 19892 9920 19944 9926
rect 19892 9862 19944 9868
rect 19800 9716 19852 9722
rect 19800 9658 19852 9664
rect 19708 9376 19760 9382
rect 19708 9318 19760 9324
rect 19812 8838 19840 9658
rect 19904 9382 19932 9862
rect 19892 9376 19944 9382
rect 19892 9318 19944 9324
rect 19892 8900 19944 8906
rect 19892 8842 19944 8848
rect 19800 8832 19852 8838
rect 19800 8774 19852 8780
rect 19904 8634 19932 8842
rect 19892 8628 19944 8634
rect 19892 8570 19944 8576
rect 19800 8492 19852 8498
rect 19800 8434 19852 8440
rect 19812 7546 19840 8434
rect 19904 7886 19932 8570
rect 19892 7880 19944 7886
rect 19892 7822 19944 7828
rect 19996 7546 20024 16612
rect 20260 16594 20312 16600
rect 20076 16448 20128 16454
rect 20076 16390 20128 16396
rect 20168 16448 20220 16454
rect 20168 16390 20220 16396
rect 20088 14793 20116 16390
rect 20180 16250 20208 16390
rect 20168 16244 20220 16250
rect 20168 16186 20220 16192
rect 20168 15360 20220 15366
rect 20168 15302 20220 15308
rect 20180 15162 20208 15302
rect 20168 15156 20220 15162
rect 20168 15098 20220 15104
rect 20074 14784 20130 14793
rect 20074 14719 20130 14728
rect 20076 14272 20128 14278
rect 20076 14214 20128 14220
rect 20088 13326 20116 14214
rect 20168 14068 20220 14074
rect 20168 14010 20220 14016
rect 20180 13394 20208 14010
rect 20168 13388 20220 13394
rect 20168 13330 20220 13336
rect 20076 13320 20128 13326
rect 20272 13274 20300 16594
rect 20364 14550 20392 18312
rect 20456 17882 20484 18788
rect 20536 18770 20588 18776
rect 20536 18692 20588 18698
rect 20536 18634 20588 18640
rect 20444 17876 20496 17882
rect 20444 17818 20496 17824
rect 20548 17762 20576 18634
rect 20640 18630 20668 19246
rect 20732 18902 20760 20402
rect 20824 19938 20852 22200
rect 21192 20602 21220 22200
rect 21180 20596 21232 20602
rect 21180 20538 21232 20544
rect 21364 20460 21416 20466
rect 21364 20402 21416 20408
rect 21088 20256 21140 20262
rect 21088 20198 21140 20204
rect 20824 19910 21036 19938
rect 20812 19780 20864 19786
rect 20812 19722 20864 19728
rect 20720 18896 20772 18902
rect 20720 18838 20772 18844
rect 20628 18624 20680 18630
rect 20824 18601 20852 19722
rect 21008 19530 21036 19910
rect 21100 19825 21128 20198
rect 21180 19848 21232 19854
rect 21086 19816 21142 19825
rect 21180 19790 21232 19796
rect 21086 19751 21142 19760
rect 21008 19502 21128 19530
rect 20996 19372 21048 19378
rect 20996 19314 21048 19320
rect 21008 18873 21036 19314
rect 20994 18864 21050 18873
rect 20994 18799 21050 18808
rect 20904 18692 20956 18698
rect 20904 18634 20956 18640
rect 20628 18566 20680 18572
rect 20810 18592 20866 18601
rect 20810 18527 20866 18536
rect 20628 18420 20680 18426
rect 20628 18362 20680 18368
rect 20640 18329 20668 18362
rect 20626 18320 20682 18329
rect 20626 18255 20682 18264
rect 20812 18284 20864 18290
rect 20812 18226 20864 18232
rect 20628 18148 20680 18154
rect 20628 18090 20680 18096
rect 20640 18057 20668 18090
rect 20626 18048 20682 18057
rect 20626 17983 20682 17992
rect 20548 17734 20668 17762
rect 20536 17604 20588 17610
rect 20536 17546 20588 17552
rect 20548 16794 20576 17546
rect 20640 17134 20668 17734
rect 20720 17672 20772 17678
rect 20720 17614 20772 17620
rect 20732 17542 20760 17614
rect 20720 17536 20772 17542
rect 20720 17478 20772 17484
rect 20628 17128 20680 17134
rect 20628 17070 20680 17076
rect 20824 16998 20852 18226
rect 20916 18193 20944 18634
rect 21100 18290 21128 19502
rect 20996 18284 21048 18290
rect 20996 18226 21048 18232
rect 21088 18284 21140 18290
rect 21088 18226 21140 18232
rect 20902 18184 20958 18193
rect 20902 18119 20958 18128
rect 21008 17882 21036 18226
rect 21086 18184 21142 18193
rect 21086 18119 21088 18128
rect 21140 18119 21142 18128
rect 21088 18090 21140 18096
rect 21192 18057 21220 19790
rect 21272 19372 21324 19378
rect 21272 19314 21324 19320
rect 21284 18426 21312 19314
rect 21272 18420 21324 18426
rect 21272 18362 21324 18368
rect 21272 18284 21324 18290
rect 21272 18226 21324 18232
rect 21178 18048 21234 18057
rect 21178 17983 21234 17992
rect 20996 17876 21048 17882
rect 20996 17818 21048 17824
rect 21180 17672 21232 17678
rect 21180 17614 21232 17620
rect 21192 17066 21220 17614
rect 21284 17338 21312 18226
rect 21376 17814 21404 20402
rect 21560 20330 21588 22200
rect 21548 20324 21600 20330
rect 21548 20266 21600 20272
rect 21548 19712 21600 19718
rect 21548 19654 21600 19660
rect 21456 19508 21508 19514
rect 21456 19450 21508 19456
rect 21468 19009 21496 19450
rect 21560 19417 21588 19654
rect 21546 19408 21602 19417
rect 21546 19343 21602 19352
rect 21454 19000 21510 19009
rect 21454 18935 21510 18944
rect 21652 18873 21680 22222
rect 21836 22114 21864 22222
rect 21914 22200 21970 23000
rect 22282 22200 22338 23000
rect 21928 22114 21956 22200
rect 21836 22086 21956 22114
rect 21742 20700 22050 20709
rect 21742 20698 21748 20700
rect 21804 20698 21828 20700
rect 21884 20698 21908 20700
rect 21964 20698 21988 20700
rect 22044 20698 22050 20700
rect 21804 20646 21806 20698
rect 21986 20646 21988 20698
rect 21742 20644 21748 20646
rect 21804 20644 21828 20646
rect 21884 20644 21908 20646
rect 21964 20644 21988 20646
rect 22044 20644 22050 20646
rect 21742 20635 22050 20644
rect 22006 19952 22062 19961
rect 22062 19910 22232 19938
rect 22006 19887 22062 19896
rect 21742 19612 22050 19621
rect 21742 19610 21748 19612
rect 21804 19610 21828 19612
rect 21884 19610 21908 19612
rect 21964 19610 21988 19612
rect 22044 19610 22050 19612
rect 21804 19558 21806 19610
rect 21986 19558 21988 19610
rect 21742 19556 21748 19558
rect 21804 19556 21828 19558
rect 21884 19556 21908 19558
rect 21964 19556 21988 19558
rect 22044 19556 22050 19558
rect 21742 19547 22050 19556
rect 21638 18864 21694 18873
rect 21638 18799 21694 18808
rect 21454 18728 21510 18737
rect 21454 18663 21510 18672
rect 21468 18630 21496 18663
rect 21456 18624 21508 18630
rect 21456 18566 21508 18572
rect 21742 18524 22050 18533
rect 21742 18522 21748 18524
rect 21804 18522 21828 18524
rect 21884 18522 21908 18524
rect 21964 18522 21988 18524
rect 22044 18522 22050 18524
rect 21804 18470 21806 18522
rect 21986 18470 21988 18522
rect 21742 18468 21748 18470
rect 21804 18468 21828 18470
rect 21884 18468 21908 18470
rect 21964 18468 21988 18470
rect 22044 18468 22050 18470
rect 21742 18459 22050 18468
rect 22204 18272 22232 19910
rect 22296 18970 22324 22200
rect 22284 18964 22336 18970
rect 22284 18906 22336 18912
rect 22204 18244 22600 18272
rect 22192 18148 22244 18154
rect 22192 18090 22244 18096
rect 21456 18080 21508 18086
rect 21456 18022 21508 18028
rect 21364 17808 21416 17814
rect 21468 17785 21496 18022
rect 21548 17808 21600 17814
rect 21364 17750 21416 17756
rect 21454 17776 21510 17785
rect 21548 17750 21600 17756
rect 21454 17711 21510 17720
rect 21272 17332 21324 17338
rect 21272 17274 21324 17280
rect 21560 17241 21588 17750
rect 21742 17436 22050 17445
rect 21742 17434 21748 17436
rect 21804 17434 21828 17436
rect 21884 17434 21908 17436
rect 21964 17434 21988 17436
rect 22044 17434 22050 17436
rect 21804 17382 21806 17434
rect 21986 17382 21988 17434
rect 21742 17380 21748 17382
rect 21804 17380 21828 17382
rect 21884 17380 21908 17382
rect 21964 17380 21988 17382
rect 22044 17380 22050 17382
rect 21742 17371 22050 17380
rect 21546 17232 21602 17241
rect 21272 17196 21324 17202
rect 21546 17167 21602 17176
rect 21272 17138 21324 17144
rect 21180 17060 21232 17066
rect 21180 17002 21232 17008
rect 20812 16992 20864 16998
rect 20812 16934 20864 16940
rect 21284 16794 21312 17138
rect 21456 16992 21508 16998
rect 21454 16960 21456 16969
rect 21508 16960 21510 16969
rect 21454 16895 21510 16904
rect 20536 16788 20588 16794
rect 20536 16730 20588 16736
rect 21272 16788 21324 16794
rect 21272 16730 21324 16736
rect 20812 16652 20864 16658
rect 20812 16594 20864 16600
rect 20628 16584 20680 16590
rect 20628 16526 20680 16532
rect 20444 16516 20496 16522
rect 20444 16458 20496 16464
rect 20456 16114 20484 16458
rect 20534 16144 20590 16153
rect 20444 16108 20496 16114
rect 20534 16079 20536 16088
rect 20444 16050 20496 16056
rect 20588 16079 20590 16088
rect 20536 16050 20588 16056
rect 20536 15904 20588 15910
rect 20536 15846 20588 15852
rect 20548 15502 20576 15846
rect 20640 15638 20668 16526
rect 20824 16232 20852 16594
rect 21088 16584 21140 16590
rect 21086 16552 21088 16561
rect 21140 16552 21142 16561
rect 21086 16487 21142 16496
rect 21456 16448 21508 16454
rect 21456 16390 21508 16396
rect 20996 16244 21048 16250
rect 20824 16204 20944 16232
rect 20812 16108 20864 16114
rect 20812 16050 20864 16056
rect 20824 15706 20852 16050
rect 20812 15700 20864 15706
rect 20812 15642 20864 15648
rect 20628 15632 20680 15638
rect 20628 15574 20680 15580
rect 20720 15564 20772 15570
rect 20720 15506 20772 15512
rect 20536 15496 20588 15502
rect 20536 15438 20588 15444
rect 20444 14816 20496 14822
rect 20444 14758 20496 14764
rect 20352 14544 20404 14550
rect 20352 14486 20404 14492
rect 20456 14414 20484 14758
rect 20628 14476 20680 14482
rect 20628 14418 20680 14424
rect 20444 14408 20496 14414
rect 20444 14350 20496 14356
rect 20640 14006 20668 14418
rect 20628 14000 20680 14006
rect 20628 13942 20680 13948
rect 20352 13932 20404 13938
rect 20352 13874 20404 13880
rect 20364 13462 20392 13874
rect 20352 13456 20404 13462
rect 20352 13398 20404 13404
rect 20732 13326 20760 15506
rect 20812 15360 20864 15366
rect 20812 15302 20864 15308
rect 20824 15026 20852 15302
rect 20812 15020 20864 15026
rect 20812 14962 20864 14968
rect 20812 14272 20864 14278
rect 20812 14214 20864 14220
rect 20076 13262 20128 13268
rect 20180 13246 20300 13274
rect 20536 13320 20588 13326
rect 20536 13262 20588 13268
rect 20720 13320 20772 13326
rect 20720 13262 20772 13268
rect 20076 11552 20128 11558
rect 20076 11494 20128 11500
rect 19800 7540 19852 7546
rect 19536 7500 19748 7528
rect 19614 7440 19670 7449
rect 19614 7375 19670 7384
rect 19340 7336 19392 7342
rect 19340 7278 19392 7284
rect 19143 7100 19451 7109
rect 19143 7098 19149 7100
rect 19205 7098 19229 7100
rect 19285 7098 19309 7100
rect 19365 7098 19389 7100
rect 19445 7098 19451 7100
rect 19205 7046 19207 7098
rect 19387 7046 19389 7098
rect 19143 7044 19149 7046
rect 19205 7044 19229 7046
rect 19285 7044 19309 7046
rect 19365 7044 19389 7046
rect 19445 7044 19451 7046
rect 19143 7035 19451 7044
rect 18972 6928 19024 6934
rect 18972 6870 19024 6876
rect 19260 6888 19564 6916
rect 19156 6860 19208 6866
rect 19260 6848 19288 6888
rect 19208 6820 19288 6848
rect 19156 6802 19208 6808
rect 18892 6752 19012 6780
rect 19536 6769 19564 6888
rect 18984 6662 19012 6752
rect 19522 6760 19578 6769
rect 19522 6695 19578 6704
rect 18972 6656 19024 6662
rect 18878 6624 18934 6633
rect 18972 6598 19024 6604
rect 19248 6656 19300 6662
rect 19248 6598 19300 6604
rect 18878 6559 18934 6568
rect 18788 6316 18840 6322
rect 18788 6258 18840 6264
rect 18800 5778 18828 6258
rect 18892 5817 18920 6559
rect 19260 6458 19288 6598
rect 19248 6452 19300 6458
rect 19248 6394 19300 6400
rect 19628 6338 19656 7375
rect 19720 7177 19748 7500
rect 19800 7482 19852 7488
rect 19984 7540 20036 7546
rect 19984 7482 20036 7488
rect 19706 7168 19762 7177
rect 19706 7103 19762 7112
rect 19812 6866 19840 7482
rect 19984 7404 20036 7410
rect 19984 7346 20036 7352
rect 19996 7002 20024 7346
rect 19984 6996 20036 7002
rect 19984 6938 20036 6944
rect 19800 6860 19852 6866
rect 19800 6802 19852 6808
rect 19800 6724 19852 6730
rect 19800 6666 19852 6672
rect 19708 6656 19760 6662
rect 19708 6598 19760 6604
rect 19720 6458 19748 6598
rect 19812 6458 19840 6666
rect 19892 6656 19944 6662
rect 19892 6598 19944 6604
rect 19708 6452 19760 6458
rect 19708 6394 19760 6400
rect 19800 6452 19852 6458
rect 19800 6394 19852 6400
rect 19524 6316 19576 6322
rect 19628 6310 19840 6338
rect 19524 6258 19576 6264
rect 18972 6112 19024 6118
rect 18972 6054 19024 6060
rect 18878 5808 18934 5817
rect 18788 5772 18840 5778
rect 18878 5743 18934 5752
rect 18788 5714 18840 5720
rect 18892 5710 18920 5743
rect 18880 5704 18932 5710
rect 18786 5672 18842 5681
rect 18880 5646 18932 5652
rect 18786 5607 18788 5616
rect 18840 5607 18842 5616
rect 18788 5578 18840 5584
rect 18880 5024 18932 5030
rect 18880 4966 18932 4972
rect 18892 4826 18920 4966
rect 18880 4820 18932 4826
rect 18880 4762 18932 4768
rect 18880 4684 18932 4690
rect 18880 4626 18932 4632
rect 18616 4270 18736 4298
rect 18616 3369 18644 4270
rect 18892 4146 18920 4626
rect 18880 4140 18932 4146
rect 18880 4082 18932 4088
rect 18696 4072 18748 4078
rect 18696 4014 18748 4020
rect 18708 3738 18736 4014
rect 18696 3732 18748 3738
rect 18696 3674 18748 3680
rect 18788 3664 18840 3670
rect 18788 3606 18840 3612
rect 18696 3460 18748 3466
rect 18696 3402 18748 3408
rect 18602 3360 18658 3369
rect 18602 3295 18658 3304
rect 18708 2990 18736 3402
rect 18604 2984 18656 2990
rect 18604 2926 18656 2932
rect 18696 2984 18748 2990
rect 18696 2926 18748 2932
rect 18616 2582 18644 2926
rect 18696 2848 18748 2854
rect 18696 2790 18748 2796
rect 18604 2576 18656 2582
rect 18708 2553 18736 2790
rect 18604 2518 18656 2524
rect 18694 2544 18750 2553
rect 18694 2479 18750 2488
rect 18512 2440 18564 2446
rect 18512 2382 18564 2388
rect 18800 800 18828 3606
rect 18892 3534 18920 4082
rect 18880 3528 18932 3534
rect 18880 3470 18932 3476
rect 18880 3392 18932 3398
rect 18880 3334 18932 3340
rect 18892 3126 18920 3334
rect 18880 3120 18932 3126
rect 18880 3062 18932 3068
rect 18984 2972 19012 6054
rect 19143 6012 19451 6021
rect 19143 6010 19149 6012
rect 19205 6010 19229 6012
rect 19285 6010 19309 6012
rect 19365 6010 19389 6012
rect 19445 6010 19451 6012
rect 19205 5958 19207 6010
rect 19387 5958 19389 6010
rect 19143 5956 19149 5958
rect 19205 5956 19229 5958
rect 19285 5956 19309 5958
rect 19365 5956 19389 5958
rect 19445 5956 19451 5958
rect 19143 5947 19451 5956
rect 19536 5914 19564 6258
rect 19706 6216 19762 6225
rect 19706 6151 19762 6160
rect 19524 5908 19576 5914
rect 19524 5850 19576 5856
rect 19064 5704 19116 5710
rect 19064 5646 19116 5652
rect 19076 4078 19104 5646
rect 19720 5642 19748 6151
rect 19708 5636 19760 5642
rect 19708 5578 19760 5584
rect 19444 5370 19748 5386
rect 19432 5364 19748 5370
rect 19484 5358 19748 5364
rect 19432 5306 19484 5312
rect 19616 5296 19668 5302
rect 19616 5238 19668 5244
rect 19143 4924 19451 4933
rect 19143 4922 19149 4924
rect 19205 4922 19229 4924
rect 19285 4922 19309 4924
rect 19365 4922 19389 4924
rect 19445 4922 19451 4924
rect 19205 4870 19207 4922
rect 19387 4870 19389 4922
rect 19143 4868 19149 4870
rect 19205 4868 19229 4870
rect 19285 4868 19309 4870
rect 19365 4868 19389 4870
rect 19445 4868 19451 4870
rect 19143 4859 19451 4868
rect 19628 4690 19656 5238
rect 19616 4684 19668 4690
rect 19616 4626 19668 4632
rect 19524 4480 19576 4486
rect 19524 4422 19576 4428
rect 19616 4480 19668 4486
rect 19616 4422 19668 4428
rect 19154 4176 19210 4185
rect 19154 4111 19210 4120
rect 19064 4072 19116 4078
rect 19064 4014 19116 4020
rect 19168 3924 19196 4111
rect 19076 3896 19196 3924
rect 19076 3534 19104 3896
rect 19143 3836 19451 3845
rect 19143 3834 19149 3836
rect 19205 3834 19229 3836
rect 19285 3834 19309 3836
rect 19365 3834 19389 3836
rect 19445 3834 19451 3836
rect 19205 3782 19207 3834
rect 19387 3782 19389 3834
rect 19143 3780 19149 3782
rect 19205 3780 19229 3782
rect 19285 3780 19309 3782
rect 19365 3780 19389 3782
rect 19445 3780 19451 3782
rect 19143 3771 19451 3780
rect 19064 3528 19116 3534
rect 19536 3482 19564 4422
rect 19628 4010 19656 4422
rect 19616 4004 19668 4010
rect 19616 3946 19668 3952
rect 19064 3470 19116 3476
rect 19444 3466 19564 3482
rect 19432 3460 19564 3466
rect 19484 3454 19564 3460
rect 19432 3402 19484 3408
rect 19524 3120 19576 3126
rect 19524 3062 19576 3068
rect 18892 2944 19012 2972
rect 18892 2854 18920 2944
rect 18880 2848 18932 2854
rect 18880 2790 18932 2796
rect 18972 2848 19024 2854
rect 18972 2790 19024 2796
rect 19064 2848 19116 2854
rect 19064 2790 19116 2796
rect 18984 2446 19012 2790
rect 18972 2440 19024 2446
rect 18972 2382 19024 2388
rect 19076 1306 19104 2790
rect 19143 2748 19451 2757
rect 19143 2746 19149 2748
rect 19205 2746 19229 2748
rect 19285 2746 19309 2748
rect 19365 2746 19389 2748
rect 19445 2746 19451 2748
rect 19205 2694 19207 2746
rect 19387 2694 19389 2746
rect 19143 2692 19149 2694
rect 19205 2692 19229 2694
rect 19285 2692 19309 2694
rect 19365 2692 19389 2694
rect 19445 2692 19451 2694
rect 19143 2683 19451 2692
rect 19248 1964 19300 1970
rect 19248 1906 19300 1912
rect 19156 1896 19208 1902
rect 19260 1873 19288 1906
rect 19156 1838 19208 1844
rect 19246 1864 19302 1873
rect 19168 1465 19196 1838
rect 19246 1799 19302 1808
rect 19536 1578 19564 3062
rect 19616 2916 19668 2922
rect 19616 2858 19668 2864
rect 19444 1550 19564 1578
rect 19154 1456 19210 1465
rect 19154 1391 19210 1400
rect 19076 1278 19196 1306
rect 19168 800 19196 1278
rect 19444 921 19472 1550
rect 19628 1442 19656 2858
rect 19720 2446 19748 5358
rect 19812 4214 19840 6310
rect 19904 5710 19932 6598
rect 19892 5704 19944 5710
rect 19892 5646 19944 5652
rect 20088 5556 20116 11494
rect 20180 6440 20208 13246
rect 20260 12912 20312 12918
rect 20260 12854 20312 12860
rect 20272 9353 20300 12854
rect 20352 12640 20404 12646
rect 20352 12582 20404 12588
rect 20258 9344 20314 9353
rect 20258 9279 20314 9288
rect 20258 9208 20314 9217
rect 20258 9143 20260 9152
rect 20312 9143 20314 9152
rect 20260 9114 20312 9120
rect 20272 8634 20300 9114
rect 20260 8628 20312 8634
rect 20260 8570 20312 8576
rect 20260 7472 20312 7478
rect 20258 7440 20260 7449
rect 20312 7440 20314 7449
rect 20258 7375 20314 7384
rect 20260 7200 20312 7206
rect 20260 7142 20312 7148
rect 20272 6905 20300 7142
rect 20258 6896 20314 6905
rect 20258 6831 20314 6840
rect 20260 6724 20312 6730
rect 20260 6666 20312 6672
rect 20272 6633 20300 6666
rect 20258 6624 20314 6633
rect 20258 6559 20314 6568
rect 20180 6412 20300 6440
rect 20272 6361 20300 6412
rect 20258 6352 20314 6361
rect 20168 6316 20220 6322
rect 20258 6287 20314 6296
rect 20168 6258 20220 6264
rect 20180 5914 20208 6258
rect 20260 6248 20312 6254
rect 20260 6190 20312 6196
rect 20168 5908 20220 5914
rect 20168 5850 20220 5856
rect 20166 5808 20222 5817
rect 20166 5743 20222 5752
rect 19904 5528 20116 5556
rect 19800 4208 19852 4214
rect 19800 4150 19852 4156
rect 19904 3534 19932 5528
rect 19984 4480 20036 4486
rect 19984 4422 20036 4428
rect 20076 4480 20128 4486
rect 20076 4422 20128 4428
rect 19996 4146 20024 4422
rect 20088 4282 20116 4422
rect 20076 4276 20128 4282
rect 20076 4218 20128 4224
rect 19984 4140 20036 4146
rect 19984 4082 20036 4088
rect 19984 4004 20036 4010
rect 19984 3946 20036 3952
rect 19892 3528 19944 3534
rect 19892 3470 19944 3476
rect 19892 3392 19944 3398
rect 19892 3334 19944 3340
rect 19800 2984 19852 2990
rect 19800 2926 19852 2932
rect 19812 2514 19840 2926
rect 19800 2508 19852 2514
rect 19800 2450 19852 2456
rect 19708 2440 19760 2446
rect 19708 2382 19760 2388
rect 19904 2106 19932 3334
rect 19892 2100 19944 2106
rect 19892 2042 19944 2048
rect 19800 2032 19852 2038
rect 19852 1980 19932 1986
rect 19800 1974 19932 1980
rect 19812 1958 19932 1974
rect 19536 1414 19656 1442
rect 19430 912 19486 921
rect 19430 847 19486 856
rect 19536 800 19564 1414
rect 19904 800 19932 1958
rect 19996 1834 20024 3946
rect 20076 3052 20128 3058
rect 20076 2994 20128 3000
rect 20088 2650 20116 2994
rect 20076 2644 20128 2650
rect 20076 2586 20128 2592
rect 20180 2378 20208 5743
rect 20272 5234 20300 6190
rect 20260 5228 20312 5234
rect 20260 5170 20312 5176
rect 20364 4146 20392 12582
rect 20548 12434 20576 13262
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 20548 12406 20668 12434
rect 20444 11756 20496 11762
rect 20444 11698 20496 11704
rect 20456 10713 20484 11698
rect 20536 11552 20588 11558
rect 20536 11494 20588 11500
rect 20548 11257 20576 11494
rect 20534 11248 20590 11257
rect 20534 11183 20590 11192
rect 20442 10704 20498 10713
rect 20442 10639 20498 10648
rect 20456 9382 20484 10639
rect 20536 9988 20588 9994
rect 20536 9930 20588 9936
rect 20548 9518 20576 9930
rect 20640 9722 20668 12406
rect 20732 12322 20760 12582
rect 20824 12434 20852 14214
rect 20916 12646 20944 16204
rect 20996 16186 21048 16192
rect 21008 15502 21036 16186
rect 21468 16153 21496 16390
rect 21742 16348 22050 16357
rect 21742 16346 21748 16348
rect 21804 16346 21828 16348
rect 21884 16346 21908 16348
rect 21964 16346 21988 16348
rect 22044 16346 22050 16348
rect 21804 16294 21806 16346
rect 21986 16294 21988 16346
rect 21742 16292 21748 16294
rect 21804 16292 21828 16294
rect 21884 16292 21908 16294
rect 21964 16292 21988 16294
rect 22044 16292 22050 16294
rect 21742 16283 22050 16292
rect 21454 16144 21510 16153
rect 21454 16079 21510 16088
rect 22100 16040 22152 16046
rect 22100 15982 22152 15988
rect 21456 15904 21508 15910
rect 21456 15846 21508 15852
rect 21468 15745 21496 15846
rect 21454 15736 21510 15745
rect 21454 15671 21510 15680
rect 21638 15600 21694 15609
rect 21638 15535 21694 15544
rect 20996 15496 21048 15502
rect 20996 15438 21048 15444
rect 21454 15464 21510 15473
rect 21454 15399 21510 15408
rect 21468 15366 21496 15399
rect 20996 15360 21048 15366
rect 20996 15302 21048 15308
rect 21456 15360 21508 15366
rect 21456 15302 21508 15308
rect 21546 15328 21602 15337
rect 21008 15026 21036 15302
rect 21546 15263 21602 15272
rect 20996 15020 21048 15026
rect 20996 14962 21048 14968
rect 21364 14952 21416 14958
rect 21086 14920 21142 14929
rect 21364 14894 21416 14900
rect 21086 14855 21088 14864
rect 21140 14855 21142 14864
rect 21088 14826 21140 14832
rect 21272 14408 21324 14414
rect 21272 14350 21324 14356
rect 21180 13728 21232 13734
rect 21180 13670 21232 13676
rect 21192 13394 21220 13670
rect 21284 13530 21312 14350
rect 21272 13524 21324 13530
rect 21272 13466 21324 13472
rect 21180 13388 21232 13394
rect 21180 13330 21232 13336
rect 21088 13184 21140 13190
rect 21088 13126 21140 13132
rect 21100 12889 21128 13126
rect 21192 12918 21220 13330
rect 21272 13320 21324 13326
rect 21272 13262 21324 13268
rect 21284 12986 21312 13262
rect 21376 13002 21404 14894
rect 21456 14816 21508 14822
rect 21456 14758 21508 14764
rect 21468 14521 21496 14758
rect 21454 14512 21510 14521
rect 21454 14447 21510 14456
rect 21456 14272 21508 14278
rect 21456 14214 21508 14220
rect 21468 13977 21496 14214
rect 21454 13968 21510 13977
rect 21560 13938 21588 15263
rect 21454 13903 21510 13912
rect 21548 13932 21600 13938
rect 21548 13874 21600 13880
rect 21456 13728 21508 13734
rect 21454 13696 21456 13705
rect 21508 13696 21510 13705
rect 21454 13631 21510 13640
rect 21454 13288 21510 13297
rect 21454 13223 21510 13232
rect 21468 13190 21496 13223
rect 21456 13184 21508 13190
rect 21456 13126 21508 13132
rect 21272 12980 21324 12986
rect 21376 12974 21588 13002
rect 21272 12922 21324 12928
rect 21180 12912 21232 12918
rect 21086 12880 21142 12889
rect 21180 12854 21232 12860
rect 21086 12815 21142 12824
rect 20904 12640 20956 12646
rect 20904 12582 20956 12588
rect 20824 12406 20944 12434
rect 20732 12294 20852 12322
rect 20916 12306 20944 12406
rect 20718 12200 20774 12209
rect 20718 12135 20720 12144
rect 20772 12135 20774 12144
rect 20720 12106 20772 12112
rect 20824 11762 20852 12294
rect 20904 12300 20956 12306
rect 20904 12242 20956 12248
rect 20720 11756 20772 11762
rect 20720 11698 20772 11704
rect 20812 11756 20864 11762
rect 20812 11698 20864 11704
rect 20732 11665 20760 11698
rect 20718 11656 20774 11665
rect 20916 11626 20944 12242
rect 20996 12232 21048 12238
rect 20996 12174 21048 12180
rect 20718 11591 20774 11600
rect 20904 11620 20956 11626
rect 20904 11562 20956 11568
rect 20916 11150 20944 11562
rect 20904 11144 20956 11150
rect 20904 11086 20956 11092
rect 20812 11008 20864 11014
rect 20812 10950 20864 10956
rect 20720 10736 20772 10742
rect 20720 10678 20772 10684
rect 20732 10062 20760 10678
rect 20824 10130 20852 10950
rect 20916 10674 20944 11086
rect 20904 10668 20956 10674
rect 20904 10610 20956 10616
rect 20904 10192 20956 10198
rect 20904 10134 20956 10140
rect 20812 10124 20864 10130
rect 20812 10066 20864 10072
rect 20720 10056 20772 10062
rect 20718 10024 20720 10033
rect 20772 10024 20774 10033
rect 20718 9959 20774 9968
rect 20812 9920 20864 9926
rect 20812 9862 20864 9868
rect 20628 9716 20680 9722
rect 20628 9658 20680 9664
rect 20720 9648 20772 9654
rect 20720 9590 20772 9596
rect 20536 9512 20588 9518
rect 20588 9460 20668 9466
rect 20536 9454 20668 9460
rect 20548 9438 20668 9454
rect 20444 9376 20496 9382
rect 20444 9318 20496 9324
rect 20640 8838 20668 9438
rect 20732 9178 20760 9590
rect 20720 9172 20772 9178
rect 20720 9114 20772 9120
rect 20628 8832 20680 8838
rect 20442 8800 20498 8809
rect 20628 8774 20680 8780
rect 20442 8735 20498 8744
rect 20456 8634 20484 8735
rect 20444 8628 20496 8634
rect 20444 8570 20496 8576
rect 20444 8016 20496 8022
rect 20444 7958 20496 7964
rect 20536 8016 20588 8022
rect 20536 7958 20588 7964
rect 20456 5778 20484 7958
rect 20444 5772 20496 5778
rect 20444 5714 20496 5720
rect 20352 4140 20404 4146
rect 20352 4082 20404 4088
rect 20444 3936 20496 3942
rect 20444 3878 20496 3884
rect 20350 3768 20406 3777
rect 20350 3703 20406 3712
rect 20260 3664 20312 3670
rect 20260 3606 20312 3612
rect 20272 2961 20300 3606
rect 20364 3534 20392 3703
rect 20352 3528 20404 3534
rect 20352 3470 20404 3476
rect 20456 3058 20484 3878
rect 20444 3052 20496 3058
rect 20444 2994 20496 3000
rect 20258 2952 20314 2961
rect 20258 2887 20314 2896
rect 20352 2848 20404 2854
rect 20352 2790 20404 2796
rect 20168 2372 20220 2378
rect 20168 2314 20220 2320
rect 19984 1828 20036 1834
rect 19984 1770 20036 1776
rect 20364 1442 20392 2790
rect 20548 2774 20576 7958
rect 20640 7954 20668 8774
rect 20718 8528 20774 8537
rect 20718 8463 20720 8472
rect 20772 8463 20774 8472
rect 20720 8434 20772 8440
rect 20718 8392 20774 8401
rect 20718 8327 20720 8336
rect 20772 8327 20774 8336
rect 20720 8298 20772 8304
rect 20824 7954 20852 9862
rect 20916 9654 20944 10134
rect 21008 9722 21036 12174
rect 21088 12164 21140 12170
rect 21088 12106 21140 12112
rect 21100 11830 21128 12106
rect 21088 11824 21140 11830
rect 21088 11766 21140 11772
rect 21100 11257 21128 11766
rect 21086 11248 21142 11257
rect 21086 11183 21142 11192
rect 21088 11076 21140 11082
rect 21088 11018 21140 11024
rect 20996 9716 21048 9722
rect 20996 9658 21048 9664
rect 20904 9648 20956 9654
rect 20904 9590 20956 9596
rect 20996 9580 21048 9586
rect 20996 9522 21048 9528
rect 20902 9072 20958 9081
rect 20902 9007 20958 9016
rect 20916 7970 20944 9007
rect 21008 8090 21036 9522
rect 21100 8090 21128 11018
rect 21192 10742 21220 12854
rect 21272 12844 21324 12850
rect 21272 12786 21324 12792
rect 21284 12374 21312 12786
rect 21456 12640 21508 12646
rect 21456 12582 21508 12588
rect 21468 12481 21496 12582
rect 21454 12472 21510 12481
rect 21454 12407 21510 12416
rect 21272 12368 21324 12374
rect 21272 12310 21324 12316
rect 21362 12336 21418 12345
rect 21362 12271 21418 12280
rect 21272 11892 21324 11898
rect 21272 11834 21324 11840
rect 21284 11218 21312 11834
rect 21272 11212 21324 11218
rect 21376 11200 21404 12271
rect 21454 12200 21510 12209
rect 21454 12135 21510 12144
rect 21468 12102 21496 12135
rect 21456 12096 21508 12102
rect 21456 12038 21508 12044
rect 21376 11172 21496 11200
rect 21272 11154 21324 11160
rect 21180 10736 21232 10742
rect 21180 10678 21232 10684
rect 21180 9716 21232 9722
rect 21180 9658 21232 9664
rect 21192 8922 21220 9658
rect 21284 9518 21312 11154
rect 21364 11076 21416 11082
rect 21364 11018 21416 11024
rect 21272 9512 21324 9518
rect 21272 9454 21324 9460
rect 21284 9042 21312 9454
rect 21272 9036 21324 9042
rect 21272 8978 21324 8984
rect 21192 8894 21312 8922
rect 21180 8832 21232 8838
rect 21180 8774 21232 8780
rect 20996 8084 21048 8090
rect 20996 8026 21048 8032
rect 21088 8084 21140 8090
rect 21088 8026 21140 8032
rect 20628 7948 20680 7954
rect 20628 7890 20680 7896
rect 20812 7948 20864 7954
rect 20916 7942 21036 7970
rect 20812 7890 20864 7896
rect 20720 7744 20772 7750
rect 20720 7686 20772 7692
rect 20628 6792 20680 6798
rect 20626 6760 20628 6769
rect 20680 6760 20682 6769
rect 20626 6695 20682 6704
rect 20732 6458 20760 7686
rect 20824 7274 20852 7890
rect 20904 7336 20956 7342
rect 20902 7304 20904 7313
rect 20956 7304 20958 7313
rect 20812 7268 20864 7274
rect 20902 7239 20958 7248
rect 20812 7210 20864 7216
rect 20720 6452 20772 6458
rect 20720 6394 20772 6400
rect 20720 6316 20772 6322
rect 20720 6258 20772 6264
rect 20732 6225 20760 6258
rect 20824 6254 20852 7210
rect 20904 6860 20956 6866
rect 20904 6802 20956 6808
rect 20812 6248 20864 6254
rect 20718 6216 20774 6225
rect 20812 6190 20864 6196
rect 20718 6151 20774 6160
rect 20732 5658 20760 6151
rect 20732 5630 20852 5658
rect 20720 5568 20772 5574
rect 20720 5510 20772 5516
rect 20732 3738 20760 5510
rect 20824 5166 20852 5630
rect 20916 5370 20944 6802
rect 21008 5914 21036 7942
rect 21088 7948 21140 7954
rect 21088 7890 21140 7896
rect 21100 7857 21128 7890
rect 21086 7848 21142 7857
rect 21086 7783 21142 7792
rect 21088 7744 21140 7750
rect 21086 7712 21088 7721
rect 21140 7712 21142 7721
rect 21086 7647 21142 7656
rect 21192 7546 21220 8774
rect 21180 7540 21232 7546
rect 21180 7482 21232 7488
rect 21088 7404 21140 7410
rect 21088 7346 21140 7352
rect 20996 5908 21048 5914
rect 20996 5850 21048 5856
rect 20994 5808 21050 5817
rect 20994 5743 21050 5752
rect 20904 5364 20956 5370
rect 20904 5306 20956 5312
rect 20812 5160 20864 5166
rect 20812 5102 20864 5108
rect 20810 4176 20866 4185
rect 20810 4111 20866 4120
rect 20824 4078 20852 4111
rect 20812 4072 20864 4078
rect 20812 4014 20864 4020
rect 20824 3913 20852 4014
rect 20810 3904 20866 3913
rect 20810 3839 20866 3848
rect 20720 3732 20772 3738
rect 20720 3674 20772 3680
rect 20916 3602 20944 5306
rect 21008 5273 21036 5743
rect 20994 5264 21050 5273
rect 20994 5199 21050 5208
rect 20994 4720 21050 4729
rect 20994 4655 21050 4664
rect 21008 4622 21036 4655
rect 20996 4616 21048 4622
rect 20996 4558 21048 4564
rect 20994 4040 21050 4049
rect 20994 3975 21050 3984
rect 20904 3596 20956 3602
rect 20904 3538 20956 3544
rect 20810 3496 20866 3505
rect 20810 3431 20812 3440
rect 20864 3431 20866 3440
rect 20812 3402 20864 3408
rect 20720 3392 20772 3398
rect 20720 3334 20772 3340
rect 20732 3233 20760 3334
rect 20718 3224 20774 3233
rect 20718 3159 20774 3168
rect 20628 2916 20680 2922
rect 20628 2858 20680 2864
rect 20272 1414 20392 1442
rect 20456 2746 20576 2774
rect 20272 800 20300 1414
rect 16684 734 16896 762
rect 16946 0 17002 800
rect 17314 0 17370 800
rect 17682 0 17738 800
rect 18050 0 18106 800
rect 18418 0 18474 800
rect 18786 0 18842 800
rect 19154 0 19210 800
rect 19522 0 19578 800
rect 19890 0 19946 800
rect 20258 0 20314 800
rect 20456 66 20484 2746
rect 20534 2680 20590 2689
rect 20534 2615 20590 2624
rect 20548 2446 20576 2615
rect 20536 2440 20588 2446
rect 20536 2382 20588 2388
rect 20640 800 20668 2858
rect 20720 2440 20772 2446
rect 20720 2382 20772 2388
rect 20732 1057 20760 2382
rect 20718 1048 20774 1057
rect 20718 983 20774 992
rect 21008 800 21036 3975
rect 21100 3466 21128 7346
rect 21180 7336 21232 7342
rect 21180 7278 21232 7284
rect 21088 3460 21140 3466
rect 21088 3402 21140 3408
rect 21192 2990 21220 7278
rect 21284 5846 21312 8894
rect 21376 6458 21404 11018
rect 21468 8022 21496 11172
rect 21560 10130 21588 12974
rect 21548 10124 21600 10130
rect 21548 10066 21600 10072
rect 21548 9580 21600 9586
rect 21548 9522 21600 9528
rect 21560 8906 21588 9522
rect 21548 8900 21600 8906
rect 21548 8842 21600 8848
rect 21546 8664 21602 8673
rect 21546 8599 21602 8608
rect 21456 8016 21508 8022
rect 21456 7958 21508 7964
rect 21454 7576 21510 7585
rect 21454 7511 21510 7520
rect 21468 7478 21496 7511
rect 21456 7472 21508 7478
rect 21456 7414 21508 7420
rect 21454 7168 21510 7177
rect 21454 7103 21510 7112
rect 21468 6458 21496 7103
rect 21364 6452 21416 6458
rect 21364 6394 21416 6400
rect 21456 6452 21508 6458
rect 21456 6394 21508 6400
rect 21560 6338 21588 8599
rect 21376 6310 21588 6338
rect 21272 5840 21324 5846
rect 21272 5782 21324 5788
rect 21272 5704 21324 5710
rect 21270 5672 21272 5681
rect 21324 5672 21326 5681
rect 21270 5607 21326 5616
rect 21376 5370 21404 6310
rect 21454 6216 21510 6225
rect 21454 6151 21510 6160
rect 21364 5364 21416 5370
rect 21364 5306 21416 5312
rect 21468 5302 21496 6151
rect 21548 6112 21600 6118
rect 21548 6054 21600 6060
rect 21456 5296 21508 5302
rect 21456 5238 21508 5244
rect 21364 5228 21416 5234
rect 21364 5170 21416 5176
rect 21270 3904 21326 3913
rect 21270 3839 21326 3848
rect 21284 3369 21312 3839
rect 21376 3670 21404 5170
rect 21456 5160 21508 5166
rect 21456 5102 21508 5108
rect 21364 3664 21416 3670
rect 21364 3606 21416 3612
rect 21270 3360 21326 3369
rect 21270 3295 21326 3304
rect 21468 3210 21496 5102
rect 21284 3182 21496 3210
rect 21180 2984 21232 2990
rect 21180 2926 21232 2932
rect 21284 2310 21312 3182
rect 21560 3097 21588 6054
rect 21546 3088 21602 3097
rect 21546 3023 21602 3032
rect 21364 2848 21416 2854
rect 21364 2790 21416 2796
rect 21272 2304 21324 2310
rect 21272 2246 21324 2252
rect 21376 800 21404 2790
rect 21652 2774 21680 15535
rect 21742 15260 22050 15269
rect 21742 15258 21748 15260
rect 21804 15258 21828 15260
rect 21884 15258 21908 15260
rect 21964 15258 21988 15260
rect 22044 15258 22050 15260
rect 21804 15206 21806 15258
rect 21986 15206 21988 15258
rect 21742 15204 21748 15206
rect 21804 15204 21828 15206
rect 21884 15204 21908 15206
rect 21964 15204 21988 15206
rect 22044 15204 22050 15206
rect 21742 15195 22050 15204
rect 21742 14172 22050 14181
rect 21742 14170 21748 14172
rect 21804 14170 21828 14172
rect 21884 14170 21908 14172
rect 21964 14170 21988 14172
rect 22044 14170 22050 14172
rect 21804 14118 21806 14170
rect 21986 14118 21988 14170
rect 21742 14116 21748 14118
rect 21804 14116 21828 14118
rect 21884 14116 21908 14118
rect 21964 14116 21988 14118
rect 22044 14116 22050 14118
rect 21742 14107 22050 14116
rect 22006 13832 22062 13841
rect 22006 13767 22062 13776
rect 22020 13190 22048 13767
rect 22008 13184 22060 13190
rect 22008 13126 22060 13132
rect 21742 13084 22050 13093
rect 21742 13082 21748 13084
rect 21804 13082 21828 13084
rect 21884 13082 21908 13084
rect 21964 13082 21988 13084
rect 22044 13082 22050 13084
rect 21804 13030 21806 13082
rect 21986 13030 21988 13082
rect 21742 13028 21748 13030
rect 21804 13028 21828 13030
rect 21884 13028 21908 13030
rect 21964 13028 21988 13030
rect 22044 13028 22050 13030
rect 21742 13019 22050 13028
rect 21730 12336 21786 12345
rect 21730 12271 21786 12280
rect 21744 12102 21772 12271
rect 21732 12096 21784 12102
rect 21732 12038 21784 12044
rect 21742 11996 22050 12005
rect 21742 11994 21748 11996
rect 21804 11994 21828 11996
rect 21884 11994 21908 11996
rect 21964 11994 21988 11996
rect 22044 11994 22050 11996
rect 21804 11942 21806 11994
rect 21986 11942 21988 11994
rect 21742 11940 21748 11942
rect 21804 11940 21828 11942
rect 21884 11940 21908 11942
rect 21964 11940 21988 11942
rect 22044 11940 22050 11942
rect 21742 11931 22050 11940
rect 21742 10908 22050 10917
rect 21742 10906 21748 10908
rect 21804 10906 21828 10908
rect 21884 10906 21908 10908
rect 21964 10906 21988 10908
rect 22044 10906 22050 10908
rect 21804 10854 21806 10906
rect 21986 10854 21988 10906
rect 21742 10852 21748 10854
rect 21804 10852 21828 10854
rect 21884 10852 21908 10854
rect 21964 10852 21988 10854
rect 22044 10852 22050 10854
rect 21742 10843 22050 10852
rect 21742 9820 22050 9829
rect 21742 9818 21748 9820
rect 21804 9818 21828 9820
rect 21884 9818 21908 9820
rect 21964 9818 21988 9820
rect 22044 9818 22050 9820
rect 21804 9766 21806 9818
rect 21986 9766 21988 9818
rect 21742 9764 21748 9766
rect 21804 9764 21828 9766
rect 21884 9764 21908 9766
rect 21964 9764 21988 9766
rect 22044 9764 22050 9766
rect 21742 9755 22050 9764
rect 21742 8732 22050 8741
rect 21742 8730 21748 8732
rect 21804 8730 21828 8732
rect 21884 8730 21908 8732
rect 21964 8730 21988 8732
rect 22044 8730 22050 8732
rect 21804 8678 21806 8730
rect 21986 8678 21988 8730
rect 21742 8676 21748 8678
rect 21804 8676 21828 8678
rect 21884 8676 21908 8678
rect 21964 8676 21988 8678
rect 22044 8676 22050 8678
rect 21742 8667 22050 8676
rect 21732 8356 21784 8362
rect 21732 8298 21784 8304
rect 21744 8129 21772 8298
rect 21730 8120 21786 8129
rect 21730 8055 21786 8064
rect 21742 7644 22050 7653
rect 21742 7642 21748 7644
rect 21804 7642 21828 7644
rect 21884 7642 21908 7644
rect 21964 7642 21988 7644
rect 22044 7642 22050 7644
rect 21804 7590 21806 7642
rect 21986 7590 21988 7642
rect 21742 7588 21748 7590
rect 21804 7588 21828 7590
rect 21884 7588 21908 7590
rect 21964 7588 21988 7590
rect 22044 7588 22050 7590
rect 21742 7579 22050 7588
rect 21742 6556 22050 6565
rect 21742 6554 21748 6556
rect 21804 6554 21828 6556
rect 21884 6554 21908 6556
rect 21964 6554 21988 6556
rect 22044 6554 22050 6556
rect 21804 6502 21806 6554
rect 21986 6502 21988 6554
rect 21742 6500 21748 6502
rect 21804 6500 21828 6502
rect 21884 6500 21908 6502
rect 21964 6500 21988 6502
rect 22044 6500 22050 6502
rect 21742 6491 22050 6500
rect 21732 6452 21784 6458
rect 21732 6394 21784 6400
rect 21744 5642 21772 6394
rect 21732 5636 21784 5642
rect 21732 5578 21784 5584
rect 21742 5468 22050 5477
rect 21742 5466 21748 5468
rect 21804 5466 21828 5468
rect 21884 5466 21908 5468
rect 21964 5466 21988 5468
rect 22044 5466 22050 5468
rect 21804 5414 21806 5466
rect 21986 5414 21988 5466
rect 21742 5412 21748 5414
rect 21804 5412 21828 5414
rect 21884 5412 21908 5414
rect 21964 5412 21988 5414
rect 22044 5412 22050 5414
rect 21742 5403 22050 5412
rect 21732 5364 21784 5370
rect 21732 5306 21784 5312
rect 21744 5137 21772 5306
rect 21730 5128 21786 5137
rect 22006 5128 22062 5137
rect 21730 5063 21786 5072
rect 21928 5086 22006 5114
rect 21928 4690 21956 5086
rect 22112 5114 22140 15982
rect 22062 5086 22140 5114
rect 22006 5063 22062 5072
rect 22008 4752 22060 4758
rect 22006 4720 22008 4729
rect 22060 4720 22062 4729
rect 21916 4684 21968 4690
rect 22062 4678 22140 4706
rect 22006 4655 22062 4664
rect 21916 4626 21968 4632
rect 21742 4380 22050 4389
rect 21742 4378 21748 4380
rect 21804 4378 21828 4380
rect 21884 4378 21908 4380
rect 21964 4378 21988 4380
rect 22044 4378 22050 4380
rect 21804 4326 21806 4378
rect 21986 4326 21988 4378
rect 21742 4324 21748 4326
rect 21804 4324 21828 4326
rect 21884 4324 21908 4326
rect 21964 4324 21988 4326
rect 22044 4324 22050 4326
rect 21742 4315 22050 4324
rect 22112 3534 22140 4678
rect 22100 3528 22152 3534
rect 22100 3470 22152 3476
rect 21742 3292 22050 3301
rect 21742 3290 21748 3292
rect 21804 3290 21828 3292
rect 21884 3290 21908 3292
rect 21964 3290 21988 3292
rect 22044 3290 22050 3292
rect 21804 3238 21806 3290
rect 21986 3238 21988 3290
rect 21742 3236 21748 3238
rect 21804 3236 21828 3238
rect 21884 3236 21908 3238
rect 21964 3236 21988 3238
rect 22044 3236 22050 3238
rect 21742 3227 22050 3236
rect 22204 3194 22232 18090
rect 22284 17740 22336 17746
rect 22284 17682 22336 17688
rect 22192 3188 22244 3194
rect 22192 3130 22244 3136
rect 22296 3126 22324 17682
rect 22376 17604 22428 17610
rect 22376 17546 22428 17552
rect 22284 3120 22336 3126
rect 22284 3062 22336 3068
rect 22388 3058 22416 17546
rect 22468 11756 22520 11762
rect 22468 11698 22520 11704
rect 22480 5370 22508 11698
rect 22572 5710 22600 18244
rect 22928 17060 22980 17066
rect 22928 17002 22980 17008
rect 22652 13932 22704 13938
rect 22652 13874 22704 13880
rect 22560 5704 22612 5710
rect 22560 5646 22612 5652
rect 22468 5364 22520 5370
rect 22468 5306 22520 5312
rect 22664 4758 22692 13874
rect 22836 13184 22888 13190
rect 22836 13126 22888 13132
rect 22744 12096 22796 12102
rect 22744 12038 22796 12044
rect 22756 5234 22784 12038
rect 22744 5228 22796 5234
rect 22744 5170 22796 5176
rect 22652 4752 22704 4758
rect 22652 4694 22704 4700
rect 22376 3052 22428 3058
rect 22376 2994 22428 3000
rect 21560 2746 21680 2774
rect 21560 2446 21588 2746
rect 21548 2440 21600 2446
rect 21548 2382 21600 2388
rect 21742 2204 22050 2213
rect 21742 2202 21748 2204
rect 21804 2202 21828 2204
rect 21884 2202 21908 2204
rect 21964 2202 21988 2204
rect 22044 2202 22050 2204
rect 21804 2150 21806 2202
rect 21986 2150 21988 2202
rect 21742 2148 21748 2150
rect 21804 2148 21828 2150
rect 21884 2148 21908 2150
rect 21964 2148 21988 2150
rect 22044 2148 22050 2150
rect 21742 2139 22050 2148
rect 20444 60 20496 66
rect 20444 2 20496 8
rect 20626 0 20682 800
rect 20994 0 21050 800
rect 21362 0 21418 800
rect 22848 134 22876 13126
rect 22940 9586 22968 17002
rect 22928 9580 22980 9586
rect 22928 9522 22980 9528
rect 22928 9444 22980 9450
rect 22928 9386 22980 9392
rect 22940 8362 22968 9386
rect 22928 8356 22980 8362
rect 22928 8298 22980 8304
rect 22940 2514 22968 8298
rect 22928 2508 22980 2514
rect 22928 2450 22980 2456
rect 22836 128 22888 134
rect 22836 70 22888 76
<< via2 >>
rect 2318 22208 2374 22264
rect 1122 21256 1178 21312
rect 938 16260 940 16280
rect 940 16260 992 16280
rect 992 16260 994 16280
rect 938 16224 994 16260
rect 938 14184 994 14240
rect 938 13912 994 13968
rect 1030 13368 1086 13424
rect 938 13096 994 13152
rect 938 6296 994 6352
rect 938 5500 994 5536
rect 938 5480 940 5500
rect 940 5480 992 5500
rect 992 5480 994 5500
rect 1030 4664 1086 4720
rect 938 3304 994 3360
rect 1490 20204 1492 20224
rect 1492 20204 1544 20224
rect 1544 20204 1546 20224
rect 1490 20168 1546 20204
rect 1490 19352 1546 19408
rect 1306 17448 1362 17504
rect 1490 18944 1546 19000
rect 1490 18572 1492 18592
rect 1492 18572 1544 18592
rect 1544 18572 1546 18592
rect 1490 18536 1546 18572
rect 1766 21392 1822 21448
rect 2226 20984 2282 21040
rect 1858 20596 1914 20632
rect 1858 20576 1860 20596
rect 1860 20576 1912 20596
rect 1912 20576 1914 20596
rect 2134 20848 2190 20904
rect 2134 20204 2136 20224
rect 2136 20204 2188 20224
rect 2188 20204 2190 20224
rect 2134 20168 2190 20204
rect 1858 19760 1914 19816
rect 1490 17720 1546 17776
rect 1490 16904 1546 16960
rect 1582 16088 1638 16144
rect 1490 15680 1546 15736
rect 1490 15308 1492 15328
rect 1492 15308 1544 15328
rect 1544 15308 1546 15328
rect 1490 15272 1546 15308
rect 1858 18148 1914 18184
rect 1858 18128 1860 18148
rect 1860 18128 1912 18148
rect 1912 18128 1914 18148
rect 1858 17312 1914 17368
rect 1858 16496 1914 16552
rect 2042 19760 2098 19816
rect 2226 17040 2282 17096
rect 2042 16632 2098 16688
rect 1950 15952 2006 16008
rect 1858 14884 1914 14920
rect 1858 14864 1860 14884
rect 1860 14864 1912 14884
rect 1912 14864 1914 14884
rect 1490 14456 1546 14512
rect 1490 14048 1546 14104
rect 2502 19080 2558 19136
rect 2594 18808 2650 18864
rect 2686 18672 2742 18728
rect 2594 17720 2650 17776
rect 2686 16632 2742 16688
rect 2318 15544 2374 15600
rect 2594 16088 2650 16144
rect 1490 13676 1492 13696
rect 1492 13676 1544 13696
rect 1544 13676 1546 13696
rect 1490 13640 1546 13676
rect 1490 13232 1546 13288
rect 1490 12824 1546 12880
rect 1490 12708 1546 12744
rect 1490 12688 1492 12708
rect 1492 12688 1544 12708
rect 1544 12688 1546 12708
rect 1766 13252 1822 13288
rect 1766 13232 1768 13252
rect 1768 13232 1820 13252
rect 1820 13232 1822 13252
rect 1858 12416 1914 12472
rect 2042 12144 2098 12200
rect 1490 12008 1546 12064
rect 1950 11756 2006 11792
rect 1950 11736 1952 11756
rect 1952 11736 2004 11756
rect 2004 11736 2006 11756
rect 1858 11192 1914 11248
rect 1490 10784 1546 10840
rect 1490 10376 1546 10432
rect 1490 9596 1492 9616
rect 1492 9596 1544 9616
rect 1544 9596 1546 9616
rect 1490 9560 1546 9596
rect 1398 8744 1454 8800
rect 1582 8200 1638 8256
rect 1490 7112 1546 7168
rect 1398 4256 1454 4312
rect 1858 10512 1914 10568
rect 1858 10140 1860 10160
rect 1860 10140 1912 10160
rect 1912 10140 1914 10160
rect 1858 10104 1914 10140
rect 2870 20476 2872 20496
rect 2872 20476 2924 20496
rect 2924 20476 2926 20496
rect 2870 20440 2926 20476
rect 2870 19080 2926 19136
rect 2410 13812 2412 13832
rect 2412 13812 2464 13832
rect 2464 13812 2466 13832
rect 2410 13776 2466 13812
rect 2226 11600 2282 11656
rect 2042 9696 2098 9752
rect 1858 8880 1914 8936
rect 1766 7656 1822 7712
rect 2134 8628 2190 8664
rect 3146 19896 3202 19952
rect 2962 18672 3018 18728
rect 4066 21800 4122 21856
rect 3514 20304 3570 20360
rect 3555 20154 3611 20156
rect 3635 20154 3691 20156
rect 3715 20154 3771 20156
rect 3795 20154 3851 20156
rect 3555 20102 3601 20154
rect 3601 20102 3611 20154
rect 3635 20102 3665 20154
rect 3665 20102 3677 20154
rect 3677 20102 3691 20154
rect 3715 20102 3729 20154
rect 3729 20102 3741 20154
rect 3741 20102 3771 20154
rect 3795 20102 3805 20154
rect 3805 20102 3851 20154
rect 3555 20100 3611 20102
rect 3635 20100 3691 20102
rect 3715 20100 3771 20102
rect 3795 20100 3851 20102
rect 3422 19352 3478 19408
rect 3330 19216 3386 19272
rect 3555 19066 3611 19068
rect 3635 19066 3691 19068
rect 3715 19066 3771 19068
rect 3795 19066 3851 19068
rect 3555 19014 3601 19066
rect 3601 19014 3611 19066
rect 3635 19014 3665 19066
rect 3665 19014 3677 19066
rect 3677 19014 3691 19066
rect 3715 19014 3729 19066
rect 3729 19014 3741 19066
rect 3741 19014 3771 19066
rect 3795 19014 3805 19066
rect 3805 19014 3851 19066
rect 3555 19012 3611 19014
rect 3635 19012 3691 19014
rect 3715 19012 3771 19014
rect 3795 19012 3851 19014
rect 4158 20032 4214 20088
rect 4066 18420 4122 18456
rect 4066 18400 4068 18420
rect 4068 18400 4120 18420
rect 4120 18400 4122 18420
rect 3555 17978 3611 17980
rect 3635 17978 3691 17980
rect 3715 17978 3771 17980
rect 3795 17978 3851 17980
rect 3555 17926 3601 17978
rect 3601 17926 3611 17978
rect 3635 17926 3665 17978
rect 3665 17926 3677 17978
rect 3677 17926 3691 17978
rect 3715 17926 3729 17978
rect 3729 17926 3741 17978
rect 3741 17926 3771 17978
rect 3795 17926 3805 17978
rect 3805 17926 3851 17978
rect 3555 17924 3611 17926
rect 3635 17924 3691 17926
rect 3715 17924 3771 17926
rect 3795 17924 3851 17926
rect 2686 11872 2742 11928
rect 3238 15000 3294 15056
rect 3790 17176 3846 17232
rect 3555 16890 3611 16892
rect 3635 16890 3691 16892
rect 3715 16890 3771 16892
rect 3795 16890 3851 16892
rect 3555 16838 3601 16890
rect 3601 16838 3611 16890
rect 3635 16838 3665 16890
rect 3665 16838 3677 16890
rect 3677 16838 3691 16890
rect 3715 16838 3729 16890
rect 3729 16838 3741 16890
rect 3741 16838 3771 16890
rect 3795 16838 3805 16890
rect 3805 16838 3851 16890
rect 3555 16836 3611 16838
rect 3635 16836 3691 16838
rect 3715 16836 3771 16838
rect 3795 16836 3851 16838
rect 4066 16904 4122 16960
rect 4618 20304 4674 20360
rect 4526 19488 4582 19544
rect 4434 18264 4490 18320
rect 4342 16632 4398 16688
rect 3422 15952 3478 16008
rect 3555 15802 3611 15804
rect 3635 15802 3691 15804
rect 3715 15802 3771 15804
rect 3795 15802 3851 15804
rect 3555 15750 3601 15802
rect 3601 15750 3611 15802
rect 3635 15750 3665 15802
rect 3665 15750 3677 15802
rect 3677 15750 3691 15802
rect 3715 15750 3729 15802
rect 3729 15750 3741 15802
rect 3741 15750 3771 15802
rect 3795 15750 3805 15802
rect 3805 15750 3851 15802
rect 3555 15748 3611 15750
rect 3635 15748 3691 15750
rect 3715 15748 3771 15750
rect 3795 15748 3851 15750
rect 3790 15444 3792 15464
rect 3792 15444 3844 15464
rect 3844 15444 3846 15464
rect 3790 15408 3846 15444
rect 3555 14714 3611 14716
rect 3635 14714 3691 14716
rect 3715 14714 3771 14716
rect 3795 14714 3851 14716
rect 3555 14662 3601 14714
rect 3601 14662 3611 14714
rect 3635 14662 3665 14714
rect 3665 14662 3677 14714
rect 3677 14662 3691 14714
rect 3715 14662 3729 14714
rect 3729 14662 3741 14714
rect 3741 14662 3771 14714
rect 3795 14662 3805 14714
rect 3805 14662 3851 14714
rect 3555 14660 3611 14662
rect 3635 14660 3691 14662
rect 3715 14660 3771 14662
rect 3795 14660 3851 14662
rect 4342 16224 4398 16280
rect 4066 15544 4122 15600
rect 4710 18400 4766 18456
rect 4618 17584 4674 17640
rect 5354 20440 5410 20496
rect 4894 19080 4950 19136
rect 4526 16632 4582 16688
rect 4802 16768 4858 16824
rect 4342 15544 4398 15600
rect 4250 15444 4252 15464
rect 4252 15444 4304 15464
rect 4304 15444 4306 15464
rect 4250 15408 4306 15444
rect 4250 14592 4306 14648
rect 3330 13640 3386 13696
rect 2502 10648 2558 10704
rect 2502 9968 2558 10024
rect 2134 8608 2136 8628
rect 2136 8608 2188 8628
rect 2188 8608 2190 8628
rect 2042 7384 2098 7440
rect 2134 6740 2136 6760
rect 2136 6740 2188 6760
rect 2188 6740 2190 6760
rect 2134 6704 2190 6740
rect 1766 5108 1768 5128
rect 1768 5108 1820 5128
rect 1820 5108 1822 5128
rect 1766 5072 1822 5108
rect 1950 5072 2006 5128
rect 1766 4256 1822 4312
rect 1950 3612 1952 3632
rect 1952 3612 2004 3632
rect 2004 3612 2006 3632
rect 1950 3576 2006 3612
rect 2778 8472 2834 8528
rect 2502 7248 2558 7304
rect 2594 6724 2650 6760
rect 2594 6704 2596 6724
rect 2596 6704 2648 6724
rect 2648 6704 2650 6724
rect 3555 13626 3611 13628
rect 3635 13626 3691 13628
rect 3715 13626 3771 13628
rect 3795 13626 3851 13628
rect 3555 13574 3601 13626
rect 3601 13574 3611 13626
rect 3635 13574 3665 13626
rect 3665 13574 3677 13626
rect 3677 13574 3691 13626
rect 3715 13574 3729 13626
rect 3729 13574 3741 13626
rect 3741 13574 3771 13626
rect 3795 13574 3805 13626
rect 3805 13574 3851 13626
rect 3555 13572 3611 13574
rect 3635 13572 3691 13574
rect 3715 13572 3771 13574
rect 3795 13572 3851 13574
rect 4066 12960 4122 13016
rect 3555 12538 3611 12540
rect 3635 12538 3691 12540
rect 3715 12538 3771 12540
rect 3795 12538 3851 12540
rect 3555 12486 3601 12538
rect 3601 12486 3611 12538
rect 3635 12486 3665 12538
rect 3665 12486 3677 12538
rect 3677 12486 3691 12538
rect 3715 12486 3729 12538
rect 3729 12486 3741 12538
rect 3741 12486 3771 12538
rect 3795 12486 3805 12538
rect 3805 12486 3851 12538
rect 3555 12484 3611 12486
rect 3635 12484 3691 12486
rect 3715 12484 3771 12486
rect 3795 12484 3851 12486
rect 3054 9716 3110 9752
rect 3054 9696 3056 9716
rect 3056 9696 3108 9716
rect 3108 9696 3110 9716
rect 3974 12316 3976 12336
rect 3976 12316 4028 12336
rect 4028 12316 4030 12336
rect 3974 12280 4030 12316
rect 3555 11450 3611 11452
rect 3635 11450 3691 11452
rect 3715 11450 3771 11452
rect 3795 11450 3851 11452
rect 3555 11398 3601 11450
rect 3601 11398 3611 11450
rect 3635 11398 3665 11450
rect 3665 11398 3677 11450
rect 3677 11398 3691 11450
rect 3715 11398 3729 11450
rect 3729 11398 3741 11450
rect 3741 11398 3771 11450
rect 3795 11398 3805 11450
rect 3805 11398 3851 11450
rect 3555 11396 3611 11398
rect 3635 11396 3691 11398
rect 3715 11396 3771 11398
rect 3795 11396 3851 11398
rect 3882 10648 3938 10704
rect 3555 10362 3611 10364
rect 3635 10362 3691 10364
rect 3715 10362 3771 10364
rect 3795 10362 3851 10364
rect 3555 10310 3601 10362
rect 3601 10310 3611 10362
rect 3635 10310 3665 10362
rect 3665 10310 3677 10362
rect 3677 10310 3691 10362
rect 3715 10310 3729 10362
rect 3729 10310 3741 10362
rect 3741 10310 3771 10362
rect 3795 10310 3805 10362
rect 3805 10310 3851 10362
rect 3555 10308 3611 10310
rect 3635 10308 3691 10310
rect 3715 10308 3771 10310
rect 3795 10308 3851 10310
rect 3422 9596 3424 9616
rect 3424 9596 3476 9616
rect 3476 9596 3478 9616
rect 3422 9560 3478 9596
rect 3606 9696 3662 9752
rect 3790 9696 3846 9752
rect 3330 9424 3386 9480
rect 2870 6840 2926 6896
rect 2778 5888 2834 5944
rect 2502 5616 2558 5672
rect 2502 4664 2558 4720
rect 1766 2352 1822 2408
rect 1582 1264 1638 1320
rect 1030 584 1086 640
rect 2226 2488 2282 2544
rect 2870 4392 2926 4448
rect 2686 2896 2742 2952
rect 2778 2644 2834 2680
rect 2778 2624 2780 2644
rect 2780 2624 2832 2644
rect 2832 2624 2834 2644
rect 2686 2488 2742 2544
rect 3146 6740 3148 6760
rect 3148 6740 3200 6760
rect 3200 6740 3202 6760
rect 3146 6704 3202 6740
rect 3146 6432 3202 6488
rect 3146 6180 3202 6216
rect 3146 6160 3148 6180
rect 3148 6160 3200 6180
rect 3200 6160 3202 6180
rect 3054 5208 3110 5264
rect 3698 9424 3754 9480
rect 3555 9274 3611 9276
rect 3635 9274 3691 9276
rect 3715 9274 3771 9276
rect 3795 9274 3851 9276
rect 3555 9222 3601 9274
rect 3601 9222 3611 9274
rect 3635 9222 3665 9274
rect 3665 9222 3677 9274
rect 3677 9222 3691 9274
rect 3715 9222 3729 9274
rect 3729 9222 3741 9274
rect 3741 9222 3771 9274
rect 3795 9222 3805 9274
rect 3805 9222 3851 9274
rect 3555 9220 3611 9222
rect 3635 9220 3691 9222
rect 3715 9220 3771 9222
rect 3795 9220 3851 9222
rect 3606 9016 3662 9072
rect 4342 13776 4398 13832
rect 4342 11892 4398 11928
rect 4342 11872 4344 11892
rect 4344 11872 4396 11892
rect 4396 11872 4398 11892
rect 4434 11328 4490 11384
rect 4158 9968 4214 10024
rect 4066 9560 4122 9616
rect 4066 9444 4122 9480
rect 4066 9424 4068 9444
rect 4068 9424 4120 9444
rect 4120 9424 4122 9444
rect 4066 9288 4122 9344
rect 3422 8336 3478 8392
rect 3555 8186 3611 8188
rect 3635 8186 3691 8188
rect 3715 8186 3771 8188
rect 3795 8186 3851 8188
rect 3555 8134 3601 8186
rect 3601 8134 3611 8186
rect 3635 8134 3665 8186
rect 3665 8134 3677 8186
rect 3677 8134 3691 8186
rect 3715 8134 3729 8186
rect 3729 8134 3741 8186
rect 3741 8134 3771 8186
rect 3795 8134 3805 8186
rect 3805 8134 3851 8186
rect 3555 8132 3611 8134
rect 3635 8132 3691 8134
rect 3715 8132 3771 8134
rect 3795 8132 3851 8134
rect 3974 8064 4030 8120
rect 3882 7928 3938 7984
rect 3790 7812 3846 7848
rect 3790 7792 3792 7812
rect 3792 7792 3844 7812
rect 3844 7792 3846 7812
rect 3514 7520 3570 7576
rect 3555 7098 3611 7100
rect 3635 7098 3691 7100
rect 3715 7098 3771 7100
rect 3795 7098 3851 7100
rect 3555 7046 3601 7098
rect 3601 7046 3611 7098
rect 3635 7046 3665 7098
rect 3665 7046 3677 7098
rect 3677 7046 3691 7098
rect 3715 7046 3729 7098
rect 3729 7046 3741 7098
rect 3741 7046 3771 7098
rect 3795 7046 3805 7098
rect 3805 7046 3851 7098
rect 3555 7044 3611 7046
rect 3635 7044 3691 7046
rect 3715 7044 3771 7046
rect 3795 7044 3851 7046
rect 4250 9424 4306 9480
rect 5630 20032 5686 20088
rect 5354 18944 5410 19000
rect 5262 18284 5318 18320
rect 5262 18264 5264 18284
rect 5264 18264 5316 18284
rect 5316 18264 5318 18284
rect 5170 18128 5226 18184
rect 5078 17040 5134 17096
rect 5538 18400 5594 18456
rect 5446 17856 5502 17912
rect 5538 17332 5594 17368
rect 5538 17312 5540 17332
rect 5540 17312 5592 17332
rect 5592 17312 5594 17332
rect 5538 17176 5594 17232
rect 5170 15952 5226 16008
rect 5262 15544 5318 15600
rect 5446 15544 5502 15600
rect 4710 11600 4766 11656
rect 4802 11500 4804 11520
rect 4804 11500 4856 11520
rect 4856 11500 4858 11520
rect 4802 11464 4858 11500
rect 4618 11192 4674 11248
rect 4710 10648 4766 10704
rect 3555 6010 3611 6012
rect 3635 6010 3691 6012
rect 3715 6010 3771 6012
rect 3795 6010 3851 6012
rect 3555 5958 3601 6010
rect 3601 5958 3611 6010
rect 3635 5958 3665 6010
rect 3665 5958 3677 6010
rect 3677 5958 3691 6010
rect 3715 5958 3729 6010
rect 3729 5958 3741 6010
rect 3741 5958 3771 6010
rect 3795 5958 3805 6010
rect 3805 5958 3851 6010
rect 3555 5956 3611 5958
rect 3635 5956 3691 5958
rect 3715 5956 3771 5958
rect 3795 5956 3851 5958
rect 3882 5616 3938 5672
rect 3330 5228 3386 5264
rect 3330 5208 3332 5228
rect 3332 5208 3384 5228
rect 3384 5208 3386 5228
rect 2962 1536 3018 1592
rect 2778 992 2834 1048
rect 3555 4922 3611 4924
rect 3635 4922 3691 4924
rect 3715 4922 3771 4924
rect 3795 4922 3851 4924
rect 3555 4870 3601 4922
rect 3601 4870 3611 4922
rect 3635 4870 3665 4922
rect 3665 4870 3677 4922
rect 3677 4870 3691 4922
rect 3715 4870 3729 4922
rect 3729 4870 3741 4922
rect 3741 4870 3771 4922
rect 3795 4870 3805 4922
rect 3805 4870 3851 4922
rect 3555 4868 3611 4870
rect 3635 4868 3691 4870
rect 3715 4868 3771 4870
rect 3795 4868 3851 4870
rect 3882 4528 3938 4584
rect 3555 3834 3611 3836
rect 3635 3834 3691 3836
rect 3715 3834 3771 3836
rect 3795 3834 3851 3836
rect 3555 3782 3601 3834
rect 3601 3782 3611 3834
rect 3635 3782 3665 3834
rect 3665 3782 3677 3834
rect 3677 3782 3691 3834
rect 3715 3782 3729 3834
rect 3729 3782 3741 3834
rect 3741 3782 3771 3834
rect 3795 3782 3805 3834
rect 3805 3782 3851 3834
rect 3555 3780 3611 3782
rect 3635 3780 3691 3782
rect 3715 3780 3771 3782
rect 3795 3780 3851 3782
rect 3422 3576 3478 3632
rect 3422 3032 3478 3088
rect 3790 3612 3792 3632
rect 3792 3612 3844 3632
rect 3844 3612 3846 3632
rect 3790 3576 3846 3612
rect 3555 2746 3611 2748
rect 3635 2746 3691 2748
rect 3715 2746 3771 2748
rect 3795 2746 3851 2748
rect 3555 2694 3601 2746
rect 3601 2694 3611 2746
rect 3635 2694 3665 2746
rect 3665 2694 3677 2746
rect 3677 2694 3691 2746
rect 3715 2694 3729 2746
rect 3729 2694 3741 2746
rect 3741 2694 3771 2746
rect 3795 2694 3805 2746
rect 3805 2694 3851 2746
rect 3555 2692 3611 2694
rect 3635 2692 3691 2694
rect 3715 2692 3771 2694
rect 3795 2692 3851 2694
rect 3606 2524 3608 2544
rect 3608 2524 3660 2544
rect 3660 2524 3662 2544
rect 3606 2488 3662 2524
rect 3330 1944 3386 2000
rect 3146 1128 3202 1184
rect 3422 1128 3478 1184
rect 3422 856 3478 912
rect 3790 2216 3846 2272
rect 4710 9868 4712 9888
rect 4712 9868 4764 9888
rect 4764 9868 4766 9888
rect 4710 9832 4766 9868
rect 4618 9016 4674 9072
rect 4802 8608 4858 8664
rect 4618 8372 4620 8392
rect 4620 8372 4672 8392
rect 4672 8372 4674 8392
rect 4618 8336 4674 8372
rect 4710 7928 4766 7984
rect 5630 14048 5686 14104
rect 5262 8608 5318 8664
rect 5262 8472 5318 8528
rect 5906 18808 5962 18864
rect 5814 18672 5870 18728
rect 5814 18284 5870 18320
rect 5814 18264 5816 18284
rect 5816 18264 5868 18284
rect 5868 18264 5870 18284
rect 6154 20698 6210 20700
rect 6234 20698 6290 20700
rect 6314 20698 6370 20700
rect 6394 20698 6450 20700
rect 6154 20646 6200 20698
rect 6200 20646 6210 20698
rect 6234 20646 6264 20698
rect 6264 20646 6276 20698
rect 6276 20646 6290 20698
rect 6314 20646 6328 20698
rect 6328 20646 6340 20698
rect 6340 20646 6370 20698
rect 6394 20646 6404 20698
rect 6404 20646 6450 20698
rect 6154 20644 6210 20646
rect 6234 20644 6290 20646
rect 6314 20644 6370 20646
rect 6394 20644 6450 20646
rect 6154 19610 6210 19612
rect 6234 19610 6290 19612
rect 6314 19610 6370 19612
rect 6394 19610 6450 19612
rect 6154 19558 6200 19610
rect 6200 19558 6210 19610
rect 6234 19558 6264 19610
rect 6264 19558 6276 19610
rect 6276 19558 6290 19610
rect 6314 19558 6328 19610
rect 6328 19558 6340 19610
rect 6340 19558 6370 19610
rect 6394 19558 6404 19610
rect 6404 19558 6450 19610
rect 6154 19556 6210 19558
rect 6234 19556 6290 19558
rect 6314 19556 6370 19558
rect 6394 19556 6450 19558
rect 7102 21392 7158 21448
rect 7102 21120 7158 21176
rect 6458 19216 6514 19272
rect 6458 18672 6514 18728
rect 6154 18522 6210 18524
rect 6234 18522 6290 18524
rect 6314 18522 6370 18524
rect 6394 18522 6450 18524
rect 6154 18470 6200 18522
rect 6200 18470 6210 18522
rect 6234 18470 6264 18522
rect 6264 18470 6276 18522
rect 6276 18470 6290 18522
rect 6314 18470 6328 18522
rect 6328 18470 6340 18522
rect 6340 18470 6370 18522
rect 6394 18470 6404 18522
rect 6404 18470 6450 18522
rect 6154 18468 6210 18470
rect 6234 18468 6290 18470
rect 6314 18468 6370 18470
rect 6394 18468 6450 18470
rect 5906 17856 5962 17912
rect 5906 17448 5962 17504
rect 6154 17434 6210 17436
rect 6234 17434 6290 17436
rect 6314 17434 6370 17436
rect 6394 17434 6450 17436
rect 6154 17382 6200 17434
rect 6200 17382 6210 17434
rect 6234 17382 6264 17434
rect 6264 17382 6276 17434
rect 6276 17382 6290 17434
rect 6314 17382 6328 17434
rect 6328 17382 6340 17434
rect 6340 17382 6370 17434
rect 6394 17382 6404 17434
rect 6404 17382 6450 17434
rect 6154 17380 6210 17382
rect 6234 17380 6290 17382
rect 6314 17380 6370 17382
rect 6394 17380 6450 17382
rect 5814 16904 5870 16960
rect 6154 16346 6210 16348
rect 6234 16346 6290 16348
rect 6314 16346 6370 16348
rect 6394 16346 6450 16348
rect 6154 16294 6200 16346
rect 6200 16294 6210 16346
rect 6234 16294 6264 16346
rect 6264 16294 6276 16346
rect 6276 16294 6290 16346
rect 6314 16294 6328 16346
rect 6328 16294 6340 16346
rect 6340 16294 6370 16346
rect 6394 16294 6404 16346
rect 6404 16294 6450 16346
rect 6154 16292 6210 16294
rect 6234 16292 6290 16294
rect 6314 16292 6370 16294
rect 6394 16292 6450 16294
rect 5906 15308 5908 15328
rect 5908 15308 5960 15328
rect 5960 15308 5962 15328
rect 5906 15272 5962 15308
rect 6642 17076 6644 17096
rect 6644 17076 6696 17096
rect 6696 17076 6698 17096
rect 6642 17040 6698 17076
rect 6642 16088 6698 16144
rect 6642 15308 6644 15328
rect 6644 15308 6696 15328
rect 6696 15308 6698 15328
rect 6642 15272 6698 15308
rect 6154 15258 6210 15260
rect 6234 15258 6290 15260
rect 6314 15258 6370 15260
rect 6394 15258 6450 15260
rect 6154 15206 6200 15258
rect 6200 15206 6210 15258
rect 6234 15206 6264 15258
rect 6264 15206 6276 15258
rect 6276 15206 6290 15258
rect 6314 15206 6328 15258
rect 6328 15206 6340 15258
rect 6340 15206 6370 15258
rect 6394 15206 6404 15258
rect 6404 15206 6450 15258
rect 6154 15204 6210 15206
rect 6234 15204 6290 15206
rect 6314 15204 6370 15206
rect 6394 15204 6450 15206
rect 6090 14864 6146 14920
rect 6154 14170 6210 14172
rect 6234 14170 6290 14172
rect 6314 14170 6370 14172
rect 6394 14170 6450 14172
rect 6154 14118 6200 14170
rect 6200 14118 6210 14170
rect 6234 14118 6264 14170
rect 6264 14118 6276 14170
rect 6276 14118 6290 14170
rect 6314 14118 6328 14170
rect 6328 14118 6340 14170
rect 6340 14118 6370 14170
rect 6394 14118 6404 14170
rect 6404 14118 6450 14170
rect 6154 14116 6210 14118
rect 6234 14116 6290 14118
rect 6314 14116 6370 14118
rect 6394 14116 6450 14118
rect 6826 18808 6882 18864
rect 6918 18536 6974 18592
rect 6826 18400 6882 18456
rect 6918 17312 6974 17368
rect 7286 20460 7342 20496
rect 7286 20440 7288 20460
rect 7288 20440 7340 20460
rect 7340 20440 7342 20460
rect 7010 16632 7066 16688
rect 6918 16496 6974 16552
rect 6826 14048 6882 14104
rect 6826 13640 6882 13696
rect 6154 13082 6210 13084
rect 6234 13082 6290 13084
rect 6314 13082 6370 13084
rect 6394 13082 6450 13084
rect 6154 13030 6200 13082
rect 6200 13030 6210 13082
rect 6234 13030 6264 13082
rect 6264 13030 6276 13082
rect 6276 13030 6290 13082
rect 6314 13030 6328 13082
rect 6328 13030 6340 13082
rect 6340 13030 6370 13082
rect 6394 13030 6404 13082
rect 6404 13030 6450 13082
rect 6154 13028 6210 13030
rect 6234 13028 6290 13030
rect 6314 13028 6370 13030
rect 6394 13028 6450 13030
rect 5906 12416 5962 12472
rect 6154 11994 6210 11996
rect 6234 11994 6290 11996
rect 6314 11994 6370 11996
rect 6394 11994 6450 11996
rect 6154 11942 6200 11994
rect 6200 11942 6210 11994
rect 6234 11942 6264 11994
rect 6264 11942 6276 11994
rect 6276 11942 6290 11994
rect 6314 11942 6328 11994
rect 6328 11942 6340 11994
rect 6340 11942 6370 11994
rect 6394 11942 6404 11994
rect 6404 11942 6450 11994
rect 6154 11940 6210 11942
rect 6234 11940 6290 11942
rect 6314 11940 6370 11942
rect 6394 11940 6450 11942
rect 5722 11736 5778 11792
rect 6154 10906 6210 10908
rect 6234 10906 6290 10908
rect 6314 10906 6370 10908
rect 6394 10906 6450 10908
rect 6154 10854 6200 10906
rect 6200 10854 6210 10906
rect 6234 10854 6264 10906
rect 6264 10854 6276 10906
rect 6276 10854 6290 10906
rect 6314 10854 6328 10906
rect 6328 10854 6340 10906
rect 6340 10854 6370 10906
rect 6394 10854 6404 10906
rect 6404 10854 6450 10906
rect 6154 10852 6210 10854
rect 6234 10852 6290 10854
rect 6314 10852 6370 10854
rect 6394 10852 6450 10854
rect 6550 10240 6606 10296
rect 6154 9818 6210 9820
rect 6234 9818 6290 9820
rect 6314 9818 6370 9820
rect 6394 9818 6450 9820
rect 6154 9766 6200 9818
rect 6200 9766 6210 9818
rect 6234 9766 6264 9818
rect 6264 9766 6276 9818
rect 6276 9766 6290 9818
rect 6314 9766 6328 9818
rect 6328 9766 6340 9818
rect 6340 9766 6370 9818
rect 6394 9766 6404 9818
rect 6404 9766 6450 9818
rect 6154 9764 6210 9766
rect 6234 9764 6290 9766
rect 6314 9764 6370 9766
rect 6394 9764 6450 9766
rect 5078 8200 5134 8256
rect 4710 7384 4766 7440
rect 4434 6976 4490 7032
rect 4158 5888 4214 5944
rect 4066 5364 4122 5400
rect 4066 5344 4068 5364
rect 4068 5344 4120 5364
rect 4120 5344 4122 5364
rect 4250 5344 4306 5400
rect 4250 3576 4306 3632
rect 3974 3168 4030 3224
rect 3974 2760 4030 2816
rect 3882 1128 3938 1184
rect 4158 2624 4214 2680
rect 4618 5616 4674 5672
rect 4802 5888 4858 5944
rect 4434 2896 4490 2952
rect 5078 4936 5134 4992
rect 4986 4800 5042 4856
rect 5078 4428 5080 4448
rect 5080 4428 5132 4448
rect 5132 4428 5134 4448
rect 5078 4392 5134 4428
rect 4710 3712 4766 3768
rect 4802 3576 4858 3632
rect 4618 2760 4674 2816
rect 4986 2352 5042 2408
rect 4986 1400 5042 1456
rect 5630 9016 5686 9072
rect 5446 7520 5502 7576
rect 5354 6840 5410 6896
rect 5446 6568 5502 6624
rect 5354 6160 5410 6216
rect 5446 5752 5502 5808
rect 5630 8200 5686 8256
rect 5814 8608 5870 8664
rect 5814 8200 5870 8256
rect 6182 9288 6238 9344
rect 6154 8730 6210 8732
rect 6234 8730 6290 8732
rect 6314 8730 6370 8732
rect 6394 8730 6450 8732
rect 6154 8678 6200 8730
rect 6200 8678 6210 8730
rect 6234 8678 6264 8730
rect 6264 8678 6276 8730
rect 6276 8678 6290 8730
rect 6314 8678 6328 8730
rect 6328 8678 6340 8730
rect 6340 8678 6370 8730
rect 6394 8678 6404 8730
rect 6404 8678 6450 8730
rect 6154 8676 6210 8678
rect 6234 8676 6290 8678
rect 6314 8676 6370 8678
rect 6394 8676 6450 8678
rect 6642 8900 6698 8936
rect 6642 8880 6644 8900
rect 6644 8880 6696 8900
rect 6696 8880 6698 8900
rect 6090 7928 6146 7984
rect 5630 7656 5686 7712
rect 6918 9696 6974 9752
rect 7838 20304 7894 20360
rect 7746 20032 7802 20088
rect 8753 20154 8809 20156
rect 8833 20154 8889 20156
rect 8913 20154 8969 20156
rect 8993 20154 9049 20156
rect 8753 20102 8799 20154
rect 8799 20102 8809 20154
rect 8833 20102 8863 20154
rect 8863 20102 8875 20154
rect 8875 20102 8889 20154
rect 8913 20102 8927 20154
rect 8927 20102 8939 20154
rect 8939 20102 8969 20154
rect 8993 20102 9003 20154
rect 9003 20102 9049 20154
rect 8753 20100 8809 20102
rect 8833 20100 8889 20102
rect 8913 20100 8969 20102
rect 8993 20100 9049 20102
rect 8206 19508 8262 19544
rect 8206 19488 8208 19508
rect 8208 19488 8260 19508
rect 8260 19488 8262 19508
rect 8206 18944 8262 19000
rect 7838 17992 7894 18048
rect 7562 17484 7564 17504
rect 7564 17484 7616 17504
rect 7616 17484 7618 17504
rect 7562 17448 7618 17484
rect 7746 17448 7802 17504
rect 7470 16088 7526 16144
rect 7654 17312 7710 17368
rect 7746 17176 7802 17232
rect 7746 17040 7802 17096
rect 7654 16632 7710 16688
rect 7746 16532 7748 16552
rect 7748 16532 7800 16552
rect 7800 16532 7802 16552
rect 7746 16496 7802 16532
rect 7930 16652 7986 16688
rect 8753 19066 8809 19068
rect 8833 19066 8889 19068
rect 8913 19066 8969 19068
rect 8993 19066 9049 19068
rect 8753 19014 8799 19066
rect 8799 19014 8809 19066
rect 8833 19014 8863 19066
rect 8863 19014 8875 19066
rect 8875 19014 8889 19066
rect 8913 19014 8927 19066
rect 8927 19014 8939 19066
rect 8939 19014 8969 19066
rect 8993 19014 9003 19066
rect 9003 19014 9049 19066
rect 8753 19012 8809 19014
rect 8833 19012 8889 19014
rect 8913 19012 8969 19014
rect 8993 19012 9049 19014
rect 8482 17992 8538 18048
rect 8482 17856 8538 17912
rect 8753 17978 8809 17980
rect 8833 17978 8889 17980
rect 8913 17978 8969 17980
rect 8993 17978 9049 17980
rect 8753 17926 8799 17978
rect 8799 17926 8809 17978
rect 8833 17926 8863 17978
rect 8863 17926 8875 17978
rect 8875 17926 8889 17978
rect 8913 17926 8927 17978
rect 8927 17926 8939 17978
rect 8939 17926 8969 17978
rect 8993 17926 9003 17978
rect 9003 17926 9049 17978
rect 8753 17924 8809 17926
rect 8833 17924 8889 17926
rect 8913 17924 8969 17926
rect 8993 17924 9049 17926
rect 8850 17720 8906 17776
rect 9034 17720 9090 17776
rect 8206 16904 8262 16960
rect 7930 16632 7932 16652
rect 7932 16632 7984 16652
rect 7984 16632 7986 16652
rect 7654 15544 7710 15600
rect 7838 15564 7894 15600
rect 7838 15544 7840 15564
rect 7840 15544 7892 15564
rect 7892 15544 7894 15564
rect 7654 15272 7710 15328
rect 7378 12044 7380 12064
rect 7380 12044 7432 12064
rect 7432 12044 7434 12064
rect 7378 12008 7434 12044
rect 7378 11736 7434 11792
rect 7286 10376 7342 10432
rect 6642 8064 6698 8120
rect 6274 7964 6276 7984
rect 6276 7964 6328 7984
rect 6328 7964 6330 7984
rect 6274 7928 6330 7964
rect 6154 7642 6210 7644
rect 6234 7642 6290 7644
rect 6314 7642 6370 7644
rect 6394 7642 6450 7644
rect 6154 7590 6200 7642
rect 6200 7590 6210 7642
rect 6234 7590 6264 7642
rect 6264 7590 6276 7642
rect 6276 7590 6290 7642
rect 6314 7590 6328 7642
rect 6328 7590 6340 7642
rect 6340 7590 6370 7642
rect 6394 7590 6404 7642
rect 6404 7590 6450 7642
rect 6154 7588 6210 7590
rect 6234 7588 6290 7590
rect 6314 7588 6370 7590
rect 6394 7588 6450 7590
rect 5722 5652 5724 5672
rect 5724 5652 5776 5672
rect 5776 5652 5778 5672
rect 5722 5616 5778 5652
rect 5630 5344 5686 5400
rect 5906 5908 5962 5944
rect 5906 5888 5908 5908
rect 5908 5888 5960 5908
rect 5960 5888 5962 5908
rect 5906 5480 5962 5536
rect 5814 5072 5870 5128
rect 5630 4528 5686 4584
rect 5814 4528 5870 4584
rect 5906 4392 5962 4448
rect 6458 6840 6514 6896
rect 6642 7692 6644 7712
rect 6644 7692 6696 7712
rect 6696 7692 6698 7712
rect 6642 7656 6698 7692
rect 6642 7248 6698 7304
rect 6642 6840 6698 6896
rect 6154 6554 6210 6556
rect 6234 6554 6290 6556
rect 6314 6554 6370 6556
rect 6394 6554 6450 6556
rect 6154 6502 6200 6554
rect 6200 6502 6210 6554
rect 6234 6502 6264 6554
rect 6264 6502 6276 6554
rect 6276 6502 6290 6554
rect 6314 6502 6328 6554
rect 6328 6502 6340 6554
rect 6340 6502 6370 6554
rect 6394 6502 6404 6554
rect 6404 6502 6450 6554
rect 6154 6500 6210 6502
rect 6234 6500 6290 6502
rect 6314 6500 6370 6502
rect 6394 6500 6450 6502
rect 6642 6296 6698 6352
rect 6366 6160 6422 6216
rect 6274 5616 6330 5672
rect 6458 5752 6514 5808
rect 6154 5466 6210 5468
rect 6234 5466 6290 5468
rect 6314 5466 6370 5468
rect 6394 5466 6450 5468
rect 6154 5414 6200 5466
rect 6200 5414 6210 5466
rect 6234 5414 6264 5466
rect 6264 5414 6276 5466
rect 6276 5414 6290 5466
rect 6314 5414 6328 5466
rect 6328 5414 6340 5466
rect 6340 5414 6370 5466
rect 6394 5414 6404 5466
rect 6404 5414 6450 5466
rect 6154 5412 6210 5414
rect 6234 5412 6290 5414
rect 6314 5412 6370 5414
rect 6394 5412 6450 5414
rect 6182 5208 6238 5264
rect 6274 4936 6330 4992
rect 6274 4820 6330 4856
rect 6274 4800 6276 4820
rect 6276 4800 6328 4820
rect 6328 4800 6330 4820
rect 6154 4378 6210 4380
rect 6234 4378 6290 4380
rect 6314 4378 6370 4380
rect 6394 4378 6450 4380
rect 6154 4326 6200 4378
rect 6200 4326 6210 4378
rect 6234 4326 6264 4378
rect 6264 4326 6276 4378
rect 6276 4326 6290 4378
rect 6314 4326 6328 4378
rect 6328 4326 6340 4378
rect 6340 4326 6370 4378
rect 6394 4326 6404 4378
rect 6404 4326 6450 4378
rect 6154 4324 6210 4326
rect 6234 4324 6290 4326
rect 6314 4324 6370 4326
rect 6394 4324 6450 4326
rect 5354 3304 5410 3360
rect 5538 3032 5594 3088
rect 5446 2624 5502 2680
rect 5998 3848 6054 3904
rect 6366 3984 6422 4040
rect 7010 8744 7066 8800
rect 6918 8472 6974 8528
rect 7010 8064 7066 8120
rect 7010 6432 7066 6488
rect 6826 5072 6882 5128
rect 6550 3712 6606 3768
rect 5538 2352 5594 2408
rect 5538 1808 5594 1864
rect 6154 3290 6210 3292
rect 6234 3290 6290 3292
rect 6314 3290 6370 3292
rect 6394 3290 6450 3292
rect 6154 3238 6200 3290
rect 6200 3238 6210 3290
rect 6234 3238 6264 3290
rect 6264 3238 6276 3290
rect 6276 3238 6290 3290
rect 6314 3238 6328 3290
rect 6328 3238 6340 3290
rect 6340 3238 6370 3290
rect 6394 3238 6404 3290
rect 6404 3238 6450 3290
rect 6154 3236 6210 3238
rect 6234 3236 6290 3238
rect 6314 3236 6370 3238
rect 6394 3236 6450 3238
rect 7010 5344 7066 5400
rect 7654 9696 7710 9752
rect 7470 9152 7526 9208
rect 7562 8492 7618 8528
rect 7562 8472 7564 8492
rect 7564 8472 7616 8492
rect 7616 8472 7618 8492
rect 7470 7248 7526 7304
rect 7286 5480 7342 5536
rect 7286 5344 7342 5400
rect 6918 3304 6974 3360
rect 6826 3188 6882 3224
rect 6826 3168 6828 3188
rect 6828 3168 6880 3188
rect 6880 3168 6882 3188
rect 7102 3848 7158 3904
rect 7010 3032 7066 3088
rect 6550 2760 6606 2816
rect 5906 2352 5962 2408
rect 5906 2216 5962 2272
rect 6154 2202 6210 2204
rect 6234 2202 6290 2204
rect 6314 2202 6370 2204
rect 6394 2202 6450 2204
rect 6154 2150 6200 2202
rect 6200 2150 6210 2202
rect 6234 2150 6264 2202
rect 6264 2150 6276 2202
rect 6276 2150 6290 2202
rect 6314 2150 6328 2202
rect 6328 2150 6340 2202
rect 6340 2150 6370 2202
rect 6394 2150 6404 2202
rect 6404 2150 6450 2202
rect 6154 2148 6210 2150
rect 6234 2148 6290 2150
rect 6314 2148 6370 2150
rect 6394 2148 6450 2150
rect 4618 40 4674 96
rect 6826 2760 6882 2816
rect 6734 1808 6790 1864
rect 7838 11076 7894 11112
rect 7838 11056 7840 11076
rect 7840 11056 7892 11076
rect 7892 11056 7894 11076
rect 8022 10376 8078 10432
rect 8390 16496 8446 16552
rect 8850 17176 8906 17232
rect 9034 17448 9090 17504
rect 8753 16890 8809 16892
rect 8833 16890 8889 16892
rect 8913 16890 8969 16892
rect 8993 16890 9049 16892
rect 8753 16838 8799 16890
rect 8799 16838 8809 16890
rect 8833 16838 8863 16890
rect 8863 16838 8875 16890
rect 8875 16838 8889 16890
rect 8913 16838 8927 16890
rect 8927 16838 8939 16890
rect 8939 16838 8969 16890
rect 8993 16838 9003 16890
rect 9003 16838 9049 16890
rect 8753 16836 8809 16838
rect 8833 16836 8889 16838
rect 8913 16836 8969 16838
rect 8993 16836 9049 16838
rect 8758 16632 8814 16688
rect 9126 16632 9182 16688
rect 8753 15802 8809 15804
rect 8833 15802 8889 15804
rect 8913 15802 8969 15804
rect 8993 15802 9049 15804
rect 8753 15750 8799 15802
rect 8799 15750 8809 15802
rect 8833 15750 8863 15802
rect 8863 15750 8875 15802
rect 8875 15750 8889 15802
rect 8913 15750 8927 15802
rect 8927 15750 8939 15802
rect 8939 15750 8969 15802
rect 8993 15750 9003 15802
rect 9003 15750 9049 15802
rect 8753 15748 8809 15750
rect 8833 15748 8889 15750
rect 8913 15748 8969 15750
rect 8993 15748 9049 15750
rect 8666 15408 8722 15464
rect 8390 15272 8446 15328
rect 8574 15308 8576 15328
rect 8576 15308 8628 15328
rect 8628 15308 8630 15328
rect 8574 15272 8630 15308
rect 9494 19352 9550 19408
rect 9770 18400 9826 18456
rect 10230 19352 10286 19408
rect 10230 18536 10286 18592
rect 9586 17312 9642 17368
rect 9954 17448 10010 17504
rect 9678 16224 9734 16280
rect 9310 15816 9366 15872
rect 9126 15020 9182 15056
rect 9126 15000 9128 15020
rect 9128 15000 9180 15020
rect 9180 15000 9182 15020
rect 8390 14728 8446 14784
rect 8753 14714 8809 14716
rect 8833 14714 8889 14716
rect 8913 14714 8969 14716
rect 8993 14714 9049 14716
rect 8753 14662 8799 14714
rect 8799 14662 8809 14714
rect 8833 14662 8863 14714
rect 8863 14662 8875 14714
rect 8875 14662 8889 14714
rect 8913 14662 8927 14714
rect 8927 14662 8939 14714
rect 8939 14662 8969 14714
rect 8993 14662 9003 14714
rect 9003 14662 9049 14714
rect 8753 14660 8809 14662
rect 8833 14660 8889 14662
rect 8913 14660 8969 14662
rect 8993 14660 9049 14662
rect 8482 14592 8538 14648
rect 8206 13096 8262 13152
rect 8758 14220 8760 14240
rect 8760 14220 8812 14240
rect 8812 14220 8814 14240
rect 8758 14184 8814 14220
rect 9494 14220 9496 14240
rect 9496 14220 9548 14240
rect 9548 14220 9550 14240
rect 9494 14184 9550 14220
rect 8574 13524 8630 13560
rect 8574 13504 8576 13524
rect 8576 13504 8628 13524
rect 8628 13504 8630 13524
rect 8753 13626 8809 13628
rect 8833 13626 8889 13628
rect 8913 13626 8969 13628
rect 8993 13626 9049 13628
rect 8753 13574 8799 13626
rect 8799 13574 8809 13626
rect 8833 13574 8863 13626
rect 8863 13574 8875 13626
rect 8875 13574 8889 13626
rect 8913 13574 8927 13626
rect 8927 13574 8939 13626
rect 8939 13574 8969 13626
rect 8993 13574 9003 13626
rect 9003 13574 9049 13626
rect 8753 13572 8809 13574
rect 8833 13572 8889 13574
rect 8913 13572 8969 13574
rect 8993 13572 9049 13574
rect 8298 12416 8354 12472
rect 8390 12300 8446 12336
rect 8390 12280 8392 12300
rect 8392 12280 8444 12300
rect 8444 12280 8446 12300
rect 8298 11464 8354 11520
rect 8390 11328 8446 11384
rect 8114 10104 8170 10160
rect 8114 9832 8170 9888
rect 7838 9696 7894 9752
rect 7838 9152 7894 9208
rect 7838 8200 7894 8256
rect 8206 9696 8262 9752
rect 8114 9152 8170 9208
rect 8206 8472 8262 8528
rect 8022 6976 8078 7032
rect 8298 8200 8354 8256
rect 8298 6568 8354 6624
rect 8022 6024 8078 6080
rect 7838 5480 7894 5536
rect 7562 4392 7618 4448
rect 7470 2760 7526 2816
rect 8753 12538 8809 12540
rect 8833 12538 8889 12540
rect 8913 12538 8969 12540
rect 8993 12538 9049 12540
rect 8753 12486 8799 12538
rect 8799 12486 8809 12538
rect 8833 12486 8863 12538
rect 8863 12486 8875 12538
rect 8875 12486 8889 12538
rect 8913 12486 8927 12538
rect 8927 12486 8939 12538
rect 8939 12486 8969 12538
rect 8993 12486 9003 12538
rect 9003 12486 9049 12538
rect 8753 12484 8809 12486
rect 8833 12484 8889 12486
rect 8913 12484 8969 12486
rect 8993 12484 9049 12486
rect 9586 12552 9642 12608
rect 8753 11450 8809 11452
rect 8833 11450 8889 11452
rect 8913 11450 8969 11452
rect 8993 11450 9049 11452
rect 8753 11398 8799 11450
rect 8799 11398 8809 11450
rect 8833 11398 8863 11450
rect 8863 11398 8875 11450
rect 8875 11398 8889 11450
rect 8913 11398 8927 11450
rect 8927 11398 8939 11450
rect 8939 11398 8969 11450
rect 8993 11398 9003 11450
rect 9003 11398 9049 11450
rect 8753 11396 8809 11398
rect 8833 11396 8889 11398
rect 8913 11396 8969 11398
rect 8993 11396 9049 11398
rect 9218 11500 9220 11520
rect 9220 11500 9272 11520
rect 9272 11500 9274 11520
rect 9218 11464 9274 11500
rect 9034 11192 9090 11248
rect 9126 10920 9182 10976
rect 9586 11872 9642 11928
rect 10046 15136 10102 15192
rect 9954 13640 10010 13696
rect 9770 13504 9826 13560
rect 10322 17448 10378 17504
rect 10598 18536 10654 18592
rect 10782 20340 10784 20360
rect 10784 20340 10836 20360
rect 10836 20340 10838 20360
rect 10782 20304 10838 20340
rect 10782 19352 10838 19408
rect 10874 19216 10930 19272
rect 10598 17448 10654 17504
rect 10506 16224 10562 16280
rect 10322 14356 10324 14376
rect 10324 14356 10376 14376
rect 10376 14356 10378 14376
rect 10322 14320 10378 14356
rect 10230 14048 10286 14104
rect 10138 13912 10194 13968
rect 10138 13640 10194 13696
rect 9770 12552 9826 12608
rect 10230 13504 10286 13560
rect 9862 12008 9918 12064
rect 9770 11872 9826 11928
rect 9586 10920 9642 10976
rect 8753 10362 8809 10364
rect 8833 10362 8889 10364
rect 8913 10362 8969 10364
rect 8993 10362 9049 10364
rect 8753 10310 8799 10362
rect 8799 10310 8809 10362
rect 8833 10310 8863 10362
rect 8863 10310 8875 10362
rect 8875 10310 8889 10362
rect 8913 10310 8927 10362
rect 8927 10310 8939 10362
rect 8939 10310 8969 10362
rect 8993 10310 9003 10362
rect 9003 10310 9049 10362
rect 8753 10308 8809 10310
rect 8833 10308 8889 10310
rect 8913 10308 8969 10310
rect 8993 10308 9049 10310
rect 9310 10376 9366 10432
rect 8942 9868 8944 9888
rect 8944 9868 8996 9888
rect 8996 9868 8998 9888
rect 8942 9832 8998 9868
rect 9126 9696 9182 9752
rect 8758 9560 8814 9616
rect 8753 9274 8809 9276
rect 8833 9274 8889 9276
rect 8913 9274 8969 9276
rect 8993 9274 9049 9276
rect 8753 9222 8799 9274
rect 8799 9222 8809 9274
rect 8833 9222 8863 9274
rect 8863 9222 8875 9274
rect 8875 9222 8889 9274
rect 8913 9222 8927 9274
rect 8927 9222 8939 9274
rect 8939 9222 8969 9274
rect 8993 9222 9003 9274
rect 9003 9222 9049 9274
rect 8753 9220 8809 9222
rect 8833 9220 8889 9222
rect 8913 9220 8969 9222
rect 8993 9220 9049 9222
rect 9310 10104 9366 10160
rect 9310 8608 9366 8664
rect 8753 8186 8809 8188
rect 8833 8186 8889 8188
rect 8913 8186 8969 8188
rect 8993 8186 9049 8188
rect 8753 8134 8799 8186
rect 8799 8134 8809 8186
rect 8833 8134 8863 8186
rect 8863 8134 8875 8186
rect 8875 8134 8889 8186
rect 8913 8134 8927 8186
rect 8927 8134 8939 8186
rect 8939 8134 8969 8186
rect 8993 8134 9003 8186
rect 9003 8134 9049 8186
rect 8753 8132 8809 8134
rect 8833 8132 8889 8134
rect 8913 8132 8969 8134
rect 8993 8132 9049 8134
rect 8574 8064 8630 8120
rect 8753 7098 8809 7100
rect 8833 7098 8889 7100
rect 8913 7098 8969 7100
rect 8993 7098 9049 7100
rect 8753 7046 8799 7098
rect 8799 7046 8809 7098
rect 8833 7046 8863 7098
rect 8863 7046 8875 7098
rect 8875 7046 8889 7098
rect 8913 7046 8927 7098
rect 8927 7046 8939 7098
rect 8939 7046 8969 7098
rect 8993 7046 9003 7098
rect 9003 7046 9049 7098
rect 8753 7044 8809 7046
rect 8833 7044 8889 7046
rect 8913 7044 8969 7046
rect 8993 7044 9049 7046
rect 8850 6296 8906 6352
rect 8753 6010 8809 6012
rect 8833 6010 8889 6012
rect 8913 6010 8969 6012
rect 8993 6010 9049 6012
rect 8753 5958 8799 6010
rect 8799 5958 8809 6010
rect 8833 5958 8863 6010
rect 8863 5958 8875 6010
rect 8875 5958 8889 6010
rect 8913 5958 8927 6010
rect 8927 5958 8939 6010
rect 8939 5958 8969 6010
rect 8993 5958 9003 6010
rect 9003 5958 9049 6010
rect 8753 5956 8809 5958
rect 8833 5956 8889 5958
rect 8913 5956 8969 5958
rect 8993 5956 9049 5958
rect 8482 4256 8538 4312
rect 8942 5616 8998 5672
rect 8753 4922 8809 4924
rect 8833 4922 8889 4924
rect 8913 4922 8969 4924
rect 8993 4922 9049 4924
rect 8753 4870 8799 4922
rect 8799 4870 8809 4922
rect 8833 4870 8863 4922
rect 8863 4870 8875 4922
rect 8875 4870 8889 4922
rect 8913 4870 8927 4922
rect 8927 4870 8939 4922
rect 8939 4870 8969 4922
rect 8993 4870 9003 4922
rect 9003 4870 9049 4922
rect 8753 4868 8809 4870
rect 8833 4868 8889 4870
rect 8913 4868 8969 4870
rect 8993 4868 9049 4870
rect 7746 2896 7802 2952
rect 7654 2644 7710 2680
rect 7654 2624 7656 2644
rect 7656 2624 7708 2644
rect 7708 2624 7710 2644
rect 7654 2372 7710 2408
rect 7654 2352 7656 2372
rect 7656 2352 7708 2372
rect 7708 2352 7710 2372
rect 8114 3304 8170 3360
rect 9034 4392 9090 4448
rect 9034 4256 9090 4312
rect 9034 3984 9090 4040
rect 8753 3834 8809 3836
rect 8833 3834 8889 3836
rect 8913 3834 8969 3836
rect 8993 3834 9049 3836
rect 8753 3782 8799 3834
rect 8799 3782 8809 3834
rect 8833 3782 8863 3834
rect 8863 3782 8875 3834
rect 8875 3782 8889 3834
rect 8913 3782 8927 3834
rect 8927 3782 8939 3834
rect 8939 3782 8969 3834
rect 8993 3782 9003 3834
rect 9003 3782 9049 3834
rect 8753 3780 8809 3782
rect 8833 3780 8889 3782
rect 8913 3780 8969 3782
rect 8993 3780 9049 3782
rect 8114 2080 8170 2136
rect 9218 5344 9274 5400
rect 9678 10548 9680 10568
rect 9680 10548 9732 10568
rect 9732 10548 9734 10568
rect 9678 10512 9734 10548
rect 9586 9696 9642 9752
rect 9678 8200 9734 8256
rect 9954 7656 10010 7712
rect 10138 9580 10194 9616
rect 10138 9560 10140 9580
rect 10140 9560 10192 9580
rect 10192 9560 10194 9580
rect 10138 9016 10194 9072
rect 10230 8356 10286 8392
rect 10230 8336 10232 8356
rect 10232 8336 10284 8356
rect 10284 8336 10286 8356
rect 10046 7384 10102 7440
rect 10598 15444 10600 15464
rect 10600 15444 10652 15464
rect 10652 15444 10654 15464
rect 10598 15408 10654 15444
rect 10598 14728 10654 14784
rect 10506 14048 10562 14104
rect 10598 13912 10654 13968
rect 10598 13812 10600 13832
rect 10600 13812 10652 13832
rect 10652 13812 10654 13832
rect 10598 13776 10654 13812
rect 10598 12552 10654 12608
rect 10782 16224 10838 16280
rect 10966 17312 11022 17368
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11398 20698
rect 11398 20646 11408 20698
rect 11432 20646 11462 20698
rect 11462 20646 11474 20698
rect 11474 20646 11488 20698
rect 11512 20646 11526 20698
rect 11526 20646 11538 20698
rect 11538 20646 11568 20698
rect 11592 20646 11602 20698
rect 11602 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 13634 20440 13690 20496
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11398 19610
rect 11398 19558 11408 19610
rect 11432 19558 11462 19610
rect 11462 19558 11474 19610
rect 11474 19558 11488 19610
rect 11512 19558 11526 19610
rect 11526 19558 11538 19610
rect 11538 19558 11568 19610
rect 11592 19558 11602 19610
rect 11602 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11398 18522
rect 11398 18470 11408 18522
rect 11432 18470 11462 18522
rect 11462 18470 11474 18522
rect 11474 18470 11488 18522
rect 11512 18470 11526 18522
rect 11526 18470 11538 18522
rect 11538 18470 11568 18522
rect 11592 18470 11602 18522
rect 11602 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11398 17434
rect 11398 17382 11408 17434
rect 11432 17382 11462 17434
rect 11462 17382 11474 17434
rect 11474 17382 11488 17434
rect 11512 17382 11526 17434
rect 11526 17382 11538 17434
rect 11538 17382 11568 17434
rect 11592 17382 11602 17434
rect 11602 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11978 18264 12034 18320
rect 11886 18028 11888 18048
rect 11888 18028 11940 18048
rect 11940 18028 11942 18048
rect 11886 17992 11942 18028
rect 10782 14864 10838 14920
rect 10782 13504 10838 13560
rect 10690 10804 10746 10840
rect 10690 10784 10692 10804
rect 10692 10784 10744 10804
rect 10744 10784 10746 10804
rect 10598 9968 10654 10024
rect 11058 14456 11114 14512
rect 10966 14048 11022 14104
rect 11058 12980 11114 13016
rect 11058 12960 11060 12980
rect 11060 12960 11112 12980
rect 11112 12960 11114 12980
rect 11794 16360 11850 16416
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11398 16346
rect 11398 16294 11408 16346
rect 11432 16294 11462 16346
rect 11462 16294 11474 16346
rect 11474 16294 11488 16346
rect 11512 16294 11526 16346
rect 11526 16294 11538 16346
rect 11538 16294 11568 16346
rect 11592 16294 11602 16346
rect 11602 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11610 16108 11666 16144
rect 11610 16088 11612 16108
rect 11612 16088 11664 16108
rect 11664 16088 11666 16108
rect 11334 15952 11390 16008
rect 11518 15988 11520 16008
rect 11520 15988 11572 16008
rect 11572 15988 11574 16008
rect 11518 15952 11574 15988
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11398 15258
rect 11398 15206 11408 15258
rect 11432 15206 11462 15258
rect 11462 15206 11474 15258
rect 11474 15206 11488 15258
rect 11512 15206 11526 15258
rect 11526 15206 11538 15258
rect 11538 15206 11568 15258
rect 11592 15206 11602 15258
rect 11602 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11398 14170
rect 11398 14118 11408 14170
rect 11432 14118 11462 14170
rect 11462 14118 11474 14170
rect 11474 14118 11488 14170
rect 11512 14118 11526 14170
rect 11526 14118 11538 14170
rect 11538 14118 11568 14170
rect 11592 14118 11602 14170
rect 11602 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11886 16088 11942 16144
rect 12070 16224 12126 16280
rect 12254 16768 12310 16824
rect 12898 18264 12954 18320
rect 13082 17992 13138 18048
rect 13082 17720 13138 17776
rect 12438 16668 12440 16688
rect 12440 16668 12492 16688
rect 12492 16668 12494 16688
rect 12438 16632 12494 16668
rect 12438 16496 12494 16552
rect 12346 16360 12402 16416
rect 12254 16088 12310 16144
rect 12254 15816 12310 15872
rect 11978 15308 11980 15328
rect 11980 15308 12032 15328
rect 12032 15308 12034 15328
rect 11978 15272 12034 15308
rect 12070 14864 12126 14920
rect 11518 13812 11520 13832
rect 11520 13812 11572 13832
rect 11572 13812 11574 13832
rect 11518 13776 11574 13812
rect 11426 13640 11482 13696
rect 11978 13524 12034 13560
rect 11978 13504 11980 13524
rect 11980 13504 12032 13524
rect 12032 13504 12034 13524
rect 11702 13368 11758 13424
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11398 13082
rect 11398 13030 11408 13082
rect 11432 13030 11462 13082
rect 11462 13030 11474 13082
rect 11474 13030 11488 13082
rect 11512 13030 11526 13082
rect 11526 13030 11538 13082
rect 11538 13030 11568 13082
rect 11592 13030 11602 13082
rect 11602 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11398 11994
rect 11398 11942 11408 11994
rect 11432 11942 11462 11994
rect 11462 11942 11474 11994
rect 11474 11942 11488 11994
rect 11512 11942 11526 11994
rect 11526 11942 11538 11994
rect 11538 11942 11568 11994
rect 11592 11942 11602 11994
rect 11602 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11518 11192 11574 11248
rect 11794 11636 11796 11656
rect 11796 11636 11848 11656
rect 11848 11636 11850 11656
rect 10966 9968 11022 10024
rect 10414 7928 10470 7984
rect 10414 6976 10470 7032
rect 10322 6840 10378 6896
rect 9586 4936 9642 4992
rect 9862 4936 9918 4992
rect 10322 6160 10378 6216
rect 10230 5480 10286 5536
rect 10138 5208 10194 5264
rect 9586 4256 9642 4312
rect 9494 3576 9550 3632
rect 9494 3168 9550 3224
rect 8753 2746 8809 2748
rect 8833 2746 8889 2748
rect 8913 2746 8969 2748
rect 8993 2746 9049 2748
rect 8753 2694 8799 2746
rect 8799 2694 8809 2746
rect 8833 2694 8863 2746
rect 8863 2694 8875 2746
rect 8875 2694 8889 2746
rect 8913 2694 8927 2746
rect 8927 2694 8939 2746
rect 8939 2694 8969 2746
rect 8993 2694 9003 2746
rect 9003 2694 9049 2746
rect 8753 2692 8809 2694
rect 8833 2692 8889 2694
rect 8913 2692 8969 2694
rect 8993 2692 9049 2694
rect 9310 2624 9366 2680
rect 9402 2488 9458 2544
rect 9494 1536 9550 1592
rect 9310 1400 9366 1456
rect 9954 4392 10010 4448
rect 9862 3576 9918 3632
rect 9862 3304 9918 3360
rect 10322 3732 10378 3768
rect 10322 3712 10324 3732
rect 10324 3712 10376 3732
rect 10376 3712 10378 3732
rect 10322 2760 10378 2816
rect 11150 10920 11206 10976
rect 10874 9424 10930 9480
rect 10966 9288 11022 9344
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11398 10906
rect 11398 10854 11408 10906
rect 11432 10854 11462 10906
rect 11462 10854 11474 10906
rect 11474 10854 11488 10906
rect 11512 10854 11526 10906
rect 11526 10854 11538 10906
rect 11538 10854 11568 10906
rect 11592 10854 11602 10906
rect 11602 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11242 10668 11298 10704
rect 11242 10648 11244 10668
rect 11244 10648 11296 10668
rect 11296 10648 11298 10668
rect 11794 11600 11850 11636
rect 11518 10104 11574 10160
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11398 9818
rect 11398 9766 11408 9818
rect 11432 9766 11462 9818
rect 11462 9766 11474 9818
rect 11474 9766 11488 9818
rect 11512 9766 11526 9818
rect 11526 9766 11538 9818
rect 11538 9766 11568 9818
rect 11592 9766 11602 9818
rect 11602 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11794 9560 11850 9616
rect 11610 9152 11666 9208
rect 11794 9152 11850 9208
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11398 8730
rect 11398 8678 11408 8730
rect 11432 8678 11462 8730
rect 11462 8678 11474 8730
rect 11474 8678 11488 8730
rect 11512 8678 11526 8730
rect 11526 8678 11538 8730
rect 11538 8678 11568 8730
rect 11592 8678 11602 8730
rect 11602 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 10782 7520 10838 7576
rect 10690 7384 10746 7440
rect 10782 7112 10838 7168
rect 10506 6296 10562 6352
rect 10966 6568 11022 6624
rect 10874 6432 10930 6488
rect 10966 5888 11022 5944
rect 10138 2352 10194 2408
rect 11610 7928 11666 7984
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11398 7642
rect 11398 7590 11408 7642
rect 11432 7590 11462 7642
rect 11462 7590 11474 7642
rect 11474 7590 11488 7642
rect 11512 7590 11526 7642
rect 11526 7590 11538 7642
rect 11538 7590 11568 7642
rect 11592 7590 11602 7642
rect 11602 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11334 6704 11390 6760
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11398 6554
rect 11398 6502 11408 6554
rect 11432 6502 11462 6554
rect 11462 6502 11474 6554
rect 11474 6502 11488 6554
rect 11512 6502 11526 6554
rect 11526 6502 11538 6554
rect 11538 6502 11568 6554
rect 11592 6502 11602 6554
rect 11602 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 11150 6160 11206 6216
rect 11242 6060 11244 6080
rect 11244 6060 11296 6080
rect 11296 6060 11298 6080
rect 11242 6024 11298 6060
rect 11610 6180 11666 6216
rect 11610 6160 11612 6180
rect 11612 6160 11664 6180
rect 11664 6160 11666 6180
rect 11610 6024 11666 6080
rect 11334 5888 11390 5944
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11398 5466
rect 11398 5414 11408 5466
rect 11432 5414 11462 5466
rect 11462 5414 11474 5466
rect 11474 5414 11488 5466
rect 11512 5414 11526 5466
rect 11526 5414 11538 5466
rect 11538 5414 11568 5466
rect 11592 5414 11602 5466
rect 11602 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 11058 3168 11114 3224
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11398 4378
rect 11398 4326 11408 4378
rect 11432 4326 11462 4378
rect 11462 4326 11474 4378
rect 11474 4326 11488 4378
rect 11512 4326 11526 4378
rect 11526 4326 11538 4378
rect 11538 4326 11568 4378
rect 11592 4326 11602 4378
rect 11602 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11398 3290
rect 11398 3238 11408 3290
rect 11432 3238 11462 3290
rect 11462 3238 11474 3290
rect 11474 3238 11488 3290
rect 11512 3238 11526 3290
rect 11526 3238 11538 3290
rect 11538 3238 11568 3290
rect 11592 3238 11602 3290
rect 11602 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 12438 15680 12494 15736
rect 12346 14864 12402 14920
rect 12714 16668 12716 16688
rect 12716 16668 12768 16688
rect 12768 16668 12770 16688
rect 12714 16632 12770 16668
rect 12622 16088 12678 16144
rect 12530 14864 12586 14920
rect 12898 15136 12954 15192
rect 13174 16632 13230 16688
rect 14462 21392 14518 21448
rect 13951 20154 14007 20156
rect 14031 20154 14087 20156
rect 14111 20154 14167 20156
rect 14191 20154 14247 20156
rect 13951 20102 13997 20154
rect 13997 20102 14007 20154
rect 14031 20102 14061 20154
rect 14061 20102 14073 20154
rect 14073 20102 14087 20154
rect 14111 20102 14125 20154
rect 14125 20102 14137 20154
rect 14137 20102 14167 20154
rect 14191 20102 14201 20154
rect 14201 20102 14247 20154
rect 13951 20100 14007 20102
rect 14031 20100 14087 20102
rect 14111 20100 14167 20102
rect 14191 20100 14247 20102
rect 13726 17856 13782 17912
rect 13951 19066 14007 19068
rect 14031 19066 14087 19068
rect 14111 19066 14167 19068
rect 14191 19066 14247 19068
rect 13951 19014 13997 19066
rect 13997 19014 14007 19066
rect 14031 19014 14061 19066
rect 14061 19014 14073 19066
rect 14073 19014 14087 19066
rect 14111 19014 14125 19066
rect 14125 19014 14137 19066
rect 14137 19014 14167 19066
rect 14191 19014 14201 19066
rect 14201 19014 14247 19066
rect 13951 19012 14007 19014
rect 14031 19012 14087 19014
rect 14111 19012 14167 19014
rect 14191 19012 14247 19014
rect 13951 17978 14007 17980
rect 14031 17978 14087 17980
rect 14111 17978 14167 17980
rect 14191 17978 14247 17980
rect 13951 17926 13997 17978
rect 13997 17926 14007 17978
rect 14031 17926 14061 17978
rect 14061 17926 14073 17978
rect 14073 17926 14087 17978
rect 14111 17926 14125 17978
rect 14125 17926 14137 17978
rect 14137 17926 14167 17978
rect 14191 17926 14201 17978
rect 14201 17926 14247 17978
rect 13951 17924 14007 17926
rect 14031 17924 14087 17926
rect 14111 17924 14167 17926
rect 14191 17924 14247 17926
rect 13818 17604 13874 17640
rect 13818 17584 13820 17604
rect 13820 17584 13872 17604
rect 13872 17584 13874 17604
rect 12898 14864 12954 14920
rect 12162 11872 12218 11928
rect 12438 11872 12494 11928
rect 12070 11192 12126 11248
rect 11978 9696 12034 9752
rect 11978 9560 12034 9616
rect 12622 13388 12678 13424
rect 12622 13368 12624 13388
rect 12624 13368 12676 13388
rect 12676 13368 12678 13388
rect 12622 12552 12678 12608
rect 12806 12824 12862 12880
rect 12714 12144 12770 12200
rect 12714 11756 12770 11792
rect 12714 11736 12716 11756
rect 12716 11736 12768 11756
rect 12768 11736 12770 11756
rect 13174 14864 13230 14920
rect 13450 13776 13506 13832
rect 13542 13676 13544 13696
rect 13544 13676 13596 13696
rect 13596 13676 13598 13696
rect 13542 13640 13598 13676
rect 13726 16940 13728 16960
rect 13728 16940 13780 16960
rect 13780 16940 13782 16960
rect 13726 16904 13782 16940
rect 13951 16890 14007 16892
rect 14031 16890 14087 16892
rect 14111 16890 14167 16892
rect 14191 16890 14247 16892
rect 13951 16838 13997 16890
rect 13997 16838 14007 16890
rect 14031 16838 14061 16890
rect 14061 16838 14073 16890
rect 14073 16838 14087 16890
rect 14111 16838 14125 16890
rect 14125 16838 14137 16890
rect 14137 16838 14167 16890
rect 14191 16838 14201 16890
rect 14201 16838 14247 16890
rect 13951 16836 14007 16838
rect 14031 16836 14087 16838
rect 14111 16836 14167 16838
rect 14191 16836 14247 16838
rect 13951 15802 14007 15804
rect 14031 15802 14087 15804
rect 14111 15802 14167 15804
rect 14191 15802 14247 15804
rect 13951 15750 13997 15802
rect 13997 15750 14007 15802
rect 14031 15750 14061 15802
rect 14061 15750 14073 15802
rect 14073 15750 14087 15802
rect 14111 15750 14125 15802
rect 14125 15750 14137 15802
rect 14137 15750 14167 15802
rect 14191 15750 14201 15802
rect 14201 15750 14247 15802
rect 13951 15748 14007 15750
rect 14031 15748 14087 15750
rect 14111 15748 14167 15750
rect 14191 15748 14247 15750
rect 14186 15136 14242 15192
rect 13726 14592 13782 14648
rect 13951 14714 14007 14716
rect 14031 14714 14087 14716
rect 14111 14714 14167 14716
rect 14191 14714 14247 14716
rect 13951 14662 13997 14714
rect 13997 14662 14007 14714
rect 14031 14662 14061 14714
rect 14061 14662 14073 14714
rect 14073 14662 14087 14714
rect 14111 14662 14125 14714
rect 14125 14662 14137 14714
rect 14137 14662 14167 14714
rect 14191 14662 14201 14714
rect 14201 14662 14247 14714
rect 13951 14660 14007 14662
rect 14031 14660 14087 14662
rect 14111 14660 14167 14662
rect 14191 14660 14247 14662
rect 14002 14456 14058 14512
rect 14278 13912 14334 13968
rect 13726 13776 13782 13832
rect 13951 13626 14007 13628
rect 14031 13626 14087 13628
rect 14111 13626 14167 13628
rect 14191 13626 14247 13628
rect 13951 13574 13997 13626
rect 13997 13574 14007 13626
rect 14031 13574 14061 13626
rect 14061 13574 14073 13626
rect 14073 13574 14087 13626
rect 14111 13574 14125 13626
rect 14125 13574 14137 13626
rect 14137 13574 14167 13626
rect 14191 13574 14201 13626
rect 14201 13574 14247 13626
rect 13951 13572 14007 13574
rect 14031 13572 14087 13574
rect 14111 13572 14167 13574
rect 14191 13572 14247 13574
rect 15106 17856 15162 17912
rect 15566 18708 15568 18728
rect 15568 18708 15620 18728
rect 15620 18708 15622 18728
rect 15566 18672 15622 18708
rect 15382 18420 15438 18456
rect 15382 18400 15384 18420
rect 15384 18400 15436 18420
rect 15436 18400 15438 18420
rect 15290 17720 15346 17776
rect 15198 17176 15254 17232
rect 13358 12824 13414 12880
rect 13266 12392 13322 12448
rect 13634 12960 13690 13016
rect 13542 12688 13598 12744
rect 15566 18028 15568 18048
rect 15568 18028 15620 18048
rect 15620 18028 15622 18048
rect 15566 17992 15622 18028
rect 14094 13096 14150 13152
rect 14186 12824 14242 12880
rect 13450 12280 13506 12336
rect 12530 9560 12586 9616
rect 12438 9424 12494 9480
rect 12530 9016 12586 9072
rect 12254 7928 12310 7984
rect 12990 10512 13046 10568
rect 12714 8472 12770 8528
rect 12714 8064 12770 8120
rect 11978 6976 12034 7032
rect 11886 6160 11942 6216
rect 11886 5888 11942 5944
rect 11978 5752 12034 5808
rect 11978 4428 11980 4448
rect 11980 4428 12032 4448
rect 12032 4428 12034 4448
rect 11978 4392 12034 4428
rect 11978 4276 12034 4312
rect 11978 4256 11980 4276
rect 11980 4256 12032 4276
rect 12032 4256 12034 4276
rect 11886 4120 11942 4176
rect 12162 7248 12218 7304
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11398 2202
rect 11398 2150 11408 2202
rect 11432 2150 11462 2202
rect 11462 2150 11474 2202
rect 11474 2150 11488 2202
rect 11512 2150 11526 2202
rect 11526 2150 11538 2202
rect 11538 2150 11568 2202
rect 11592 2150 11602 2202
rect 11602 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 10966 1944 11022 2000
rect 11242 1128 11298 1184
rect 11242 856 11298 912
rect 12070 1672 12126 1728
rect 12806 7112 12862 7168
rect 12806 6996 12862 7032
rect 12806 6976 12808 6996
rect 12808 6976 12860 6996
rect 12860 6976 12862 6996
rect 12438 4664 12494 4720
rect 13358 9288 13414 9344
rect 13358 9152 13414 9208
rect 13358 8472 13414 8528
rect 12990 6568 13046 6624
rect 12898 6024 12954 6080
rect 12530 3712 12586 3768
rect 12346 3304 12402 3360
rect 12438 3168 12494 3224
rect 12530 2896 12586 2952
rect 12346 2760 12402 2816
rect 12346 2524 12348 2544
rect 12348 2524 12400 2544
rect 12400 2524 12402 2544
rect 12346 2488 12402 2524
rect 12714 4684 12770 4720
rect 12714 4664 12716 4684
rect 12716 4664 12768 4684
rect 12768 4664 12770 4684
rect 12714 3032 12770 3088
rect 13082 5752 13138 5808
rect 12990 5208 13046 5264
rect 12990 4820 13046 4856
rect 12990 4800 12992 4820
rect 12992 4800 13044 4820
rect 13044 4800 13046 4820
rect 13358 5480 13414 5536
rect 13951 12538 14007 12540
rect 14031 12538 14087 12540
rect 14111 12538 14167 12540
rect 14191 12538 14247 12540
rect 13951 12486 13997 12538
rect 13997 12486 14007 12538
rect 14031 12486 14061 12538
rect 14061 12486 14073 12538
rect 14073 12486 14087 12538
rect 14111 12486 14125 12538
rect 14125 12486 14137 12538
rect 14137 12486 14167 12538
rect 14191 12486 14201 12538
rect 14201 12486 14247 12538
rect 13951 12484 14007 12486
rect 14031 12484 14087 12486
rect 14111 12484 14167 12486
rect 14191 12484 14247 12486
rect 13910 12044 13912 12064
rect 13912 12044 13964 12064
rect 13964 12044 13966 12064
rect 13910 12008 13966 12044
rect 14094 11736 14150 11792
rect 13951 11450 14007 11452
rect 14031 11450 14087 11452
rect 14111 11450 14167 11452
rect 14191 11450 14247 11452
rect 13951 11398 13997 11450
rect 13997 11398 14007 11450
rect 14031 11398 14061 11450
rect 14061 11398 14073 11450
rect 14073 11398 14087 11450
rect 14111 11398 14125 11450
rect 14125 11398 14137 11450
rect 14137 11398 14167 11450
rect 14191 11398 14201 11450
rect 14201 11398 14247 11450
rect 13951 11396 14007 11398
rect 14031 11396 14087 11398
rect 14111 11396 14167 11398
rect 14191 11396 14247 11398
rect 14370 12688 14426 12744
rect 15106 14184 15162 14240
rect 14646 12144 14702 12200
rect 14554 11872 14610 11928
rect 14186 10784 14242 10840
rect 13951 10362 14007 10364
rect 14031 10362 14087 10364
rect 14111 10362 14167 10364
rect 14191 10362 14247 10364
rect 13951 10310 13997 10362
rect 13997 10310 14007 10362
rect 14031 10310 14061 10362
rect 14061 10310 14073 10362
rect 14073 10310 14087 10362
rect 14111 10310 14125 10362
rect 14125 10310 14137 10362
rect 14137 10310 14167 10362
rect 14191 10310 14201 10362
rect 14201 10310 14247 10362
rect 13951 10308 14007 10310
rect 14031 10308 14087 10310
rect 14111 10308 14167 10310
rect 14191 10308 14247 10310
rect 13818 10104 13874 10160
rect 14002 10140 14004 10160
rect 14004 10140 14056 10160
rect 14056 10140 14058 10160
rect 14002 10104 14058 10140
rect 13634 9832 13690 9888
rect 13726 9696 13782 9752
rect 13951 9274 14007 9276
rect 14031 9274 14087 9276
rect 14111 9274 14167 9276
rect 14191 9274 14247 9276
rect 13951 9222 13997 9274
rect 13997 9222 14007 9274
rect 14031 9222 14061 9274
rect 14061 9222 14073 9274
rect 14073 9222 14087 9274
rect 14111 9222 14125 9274
rect 14125 9222 14137 9274
rect 14137 9222 14167 9274
rect 14191 9222 14201 9274
rect 14201 9222 14247 9274
rect 13951 9220 14007 9222
rect 14031 9220 14087 9222
rect 14111 9220 14167 9222
rect 14191 9220 14247 9222
rect 14094 8492 14150 8528
rect 14094 8472 14096 8492
rect 14096 8472 14148 8492
rect 14148 8472 14150 8492
rect 14186 8356 14242 8392
rect 14186 8336 14188 8356
rect 14188 8336 14240 8356
rect 14240 8336 14242 8356
rect 13634 7248 13690 7304
rect 13951 8186 14007 8188
rect 14031 8186 14087 8188
rect 14111 8186 14167 8188
rect 14191 8186 14247 8188
rect 13951 8134 13997 8186
rect 13997 8134 14007 8186
rect 14031 8134 14061 8186
rect 14061 8134 14073 8186
rect 14073 8134 14087 8186
rect 14111 8134 14125 8186
rect 14125 8134 14137 8186
rect 14137 8134 14167 8186
rect 14191 8134 14201 8186
rect 14201 8134 14247 8186
rect 13951 8132 14007 8134
rect 14031 8132 14087 8134
rect 14111 8132 14167 8134
rect 14191 8132 14247 8134
rect 13818 7520 13874 7576
rect 13951 7098 14007 7100
rect 14031 7098 14087 7100
rect 14111 7098 14167 7100
rect 14191 7098 14247 7100
rect 13951 7046 13997 7098
rect 13997 7046 14007 7098
rect 14031 7046 14061 7098
rect 14061 7046 14073 7098
rect 14073 7046 14087 7098
rect 14111 7046 14125 7098
rect 14125 7046 14137 7098
rect 14137 7046 14167 7098
rect 14191 7046 14201 7098
rect 14201 7046 14247 7098
rect 13951 7044 14007 7046
rect 14031 7044 14087 7046
rect 14111 7044 14167 7046
rect 14191 7044 14247 7046
rect 13818 6976 13874 7032
rect 14646 11192 14702 11248
rect 14554 9832 14610 9888
rect 14462 7928 14518 7984
rect 14646 9324 14648 9344
rect 14648 9324 14700 9344
rect 14700 9324 14702 9344
rect 14646 9288 14702 9324
rect 14830 9560 14886 9616
rect 14738 8608 14794 8664
rect 15106 12008 15162 12064
rect 15198 11736 15254 11792
rect 15198 11500 15200 11520
rect 15200 11500 15252 11520
rect 15252 11500 15254 11520
rect 15198 11464 15254 11500
rect 15014 8880 15070 8936
rect 14738 8200 14794 8256
rect 14646 8064 14702 8120
rect 13542 5072 13598 5128
rect 13266 3032 13322 3088
rect 13951 6010 14007 6012
rect 14031 6010 14087 6012
rect 14111 6010 14167 6012
rect 14191 6010 14247 6012
rect 13951 5958 13997 6010
rect 13997 5958 14007 6010
rect 14031 5958 14061 6010
rect 14061 5958 14073 6010
rect 14073 5958 14087 6010
rect 14111 5958 14125 6010
rect 14125 5958 14137 6010
rect 14137 5958 14167 6010
rect 14191 5958 14201 6010
rect 14201 5958 14247 6010
rect 13951 5956 14007 5958
rect 14031 5956 14087 5958
rect 14111 5956 14167 5958
rect 14191 5956 14247 5958
rect 14186 5752 14242 5808
rect 14462 5344 14518 5400
rect 13818 4936 13874 4992
rect 13951 4922 14007 4924
rect 14031 4922 14087 4924
rect 14111 4922 14167 4924
rect 14191 4922 14247 4924
rect 13951 4870 13997 4922
rect 13997 4870 14007 4922
rect 14031 4870 14061 4922
rect 14061 4870 14073 4922
rect 14073 4870 14087 4922
rect 14111 4870 14125 4922
rect 14125 4870 14137 4922
rect 14137 4870 14167 4922
rect 14191 4870 14201 4922
rect 14201 4870 14247 4922
rect 13951 4868 14007 4870
rect 14031 4868 14087 4870
rect 14111 4868 14167 4870
rect 14191 4868 14247 4870
rect 13726 4684 13782 4720
rect 13726 4664 13728 4684
rect 13728 4664 13780 4684
rect 13780 4664 13782 4684
rect 13634 4392 13690 4448
rect 13542 4120 13598 4176
rect 12990 1264 13046 1320
rect 13951 3834 14007 3836
rect 14031 3834 14087 3836
rect 14111 3834 14167 3836
rect 14191 3834 14247 3836
rect 13951 3782 13997 3834
rect 13997 3782 14007 3834
rect 14031 3782 14061 3834
rect 14061 3782 14073 3834
rect 14073 3782 14087 3834
rect 14111 3782 14125 3834
rect 14125 3782 14137 3834
rect 14137 3782 14167 3834
rect 14191 3782 14201 3834
rect 14201 3782 14247 3834
rect 13951 3780 14007 3782
rect 14031 3780 14087 3782
rect 14111 3780 14167 3782
rect 14191 3780 14247 3782
rect 13818 3576 13874 3632
rect 14462 4684 14518 4720
rect 14462 4664 14464 4684
rect 14464 4664 14516 4684
rect 14516 4664 14518 4684
rect 14554 4428 14556 4448
rect 14556 4428 14608 4448
rect 14608 4428 14610 4448
rect 14554 4392 14610 4428
rect 15474 14320 15530 14376
rect 16550 20698 16606 20700
rect 16630 20698 16686 20700
rect 16710 20698 16766 20700
rect 16790 20698 16846 20700
rect 16550 20646 16596 20698
rect 16596 20646 16606 20698
rect 16630 20646 16660 20698
rect 16660 20646 16672 20698
rect 16672 20646 16686 20698
rect 16710 20646 16724 20698
rect 16724 20646 16736 20698
rect 16736 20646 16766 20698
rect 16790 20646 16800 20698
rect 16800 20646 16846 20698
rect 16550 20644 16606 20646
rect 16630 20644 16686 20646
rect 16710 20644 16766 20646
rect 16790 20644 16846 20646
rect 17774 20984 17830 21040
rect 16394 20032 16450 20088
rect 15566 11056 15622 11112
rect 15474 10648 15530 10704
rect 15290 9560 15346 9616
rect 15474 9288 15530 9344
rect 15474 9152 15530 9208
rect 14922 7792 14978 7848
rect 14738 3576 14794 3632
rect 14738 3168 14794 3224
rect 14830 3068 14832 3088
rect 14832 3068 14884 3088
rect 14884 3068 14886 3088
rect 13951 2746 14007 2748
rect 14031 2746 14087 2748
rect 14111 2746 14167 2748
rect 14191 2746 14247 2748
rect 13951 2694 13997 2746
rect 13997 2694 14007 2746
rect 14031 2694 14061 2746
rect 14061 2694 14073 2746
rect 14073 2694 14087 2746
rect 14111 2694 14125 2746
rect 14125 2694 14137 2746
rect 14137 2694 14167 2746
rect 14191 2694 14201 2746
rect 14201 2694 14247 2746
rect 13951 2692 14007 2694
rect 14031 2692 14087 2694
rect 14111 2692 14167 2694
rect 14191 2692 14247 2694
rect 14830 3032 14886 3068
rect 15566 8064 15622 8120
rect 15474 7520 15530 7576
rect 15106 6840 15162 6896
rect 15382 7248 15438 7304
rect 15014 4256 15070 4312
rect 15566 6976 15622 7032
rect 15290 4120 15346 4176
rect 15198 3984 15254 4040
rect 15014 3712 15070 3768
rect 16550 19610 16606 19612
rect 16630 19610 16686 19612
rect 16710 19610 16766 19612
rect 16790 19610 16846 19612
rect 16550 19558 16596 19610
rect 16596 19558 16606 19610
rect 16630 19558 16660 19610
rect 16660 19558 16672 19610
rect 16672 19558 16686 19610
rect 16710 19558 16724 19610
rect 16724 19558 16736 19610
rect 16736 19558 16766 19610
rect 16790 19558 16800 19610
rect 16800 19558 16846 19610
rect 16550 19556 16606 19558
rect 16630 19556 16686 19558
rect 16710 19556 16766 19558
rect 16790 19556 16846 19558
rect 16854 19372 16910 19408
rect 16854 19352 16856 19372
rect 16856 19352 16908 19372
rect 16908 19352 16910 19372
rect 16550 18522 16606 18524
rect 16630 18522 16686 18524
rect 16710 18522 16766 18524
rect 16790 18522 16846 18524
rect 16550 18470 16596 18522
rect 16596 18470 16606 18522
rect 16630 18470 16660 18522
rect 16660 18470 16672 18522
rect 16672 18470 16686 18522
rect 16710 18470 16724 18522
rect 16724 18470 16736 18522
rect 16736 18470 16766 18522
rect 16790 18470 16800 18522
rect 16800 18470 16846 18522
rect 16550 18468 16606 18470
rect 16630 18468 16686 18470
rect 16710 18468 16766 18470
rect 16790 18468 16846 18470
rect 17222 17992 17278 18048
rect 16550 17434 16606 17436
rect 16630 17434 16686 17436
rect 16710 17434 16766 17436
rect 16790 17434 16846 17436
rect 16550 17382 16596 17434
rect 16596 17382 16606 17434
rect 16630 17382 16660 17434
rect 16660 17382 16672 17434
rect 16672 17382 16686 17434
rect 16710 17382 16724 17434
rect 16724 17382 16736 17434
rect 16736 17382 16766 17434
rect 16790 17382 16800 17434
rect 16800 17382 16846 17434
rect 16550 17380 16606 17382
rect 16630 17380 16686 17382
rect 16710 17380 16766 17382
rect 16790 17380 16846 17382
rect 16210 16652 16266 16688
rect 16210 16632 16212 16652
rect 16212 16632 16264 16652
rect 16264 16632 16266 16652
rect 16118 16224 16174 16280
rect 16550 16346 16606 16348
rect 16630 16346 16686 16348
rect 16710 16346 16766 16348
rect 16790 16346 16846 16348
rect 16550 16294 16596 16346
rect 16596 16294 16606 16346
rect 16630 16294 16660 16346
rect 16660 16294 16672 16346
rect 16672 16294 16686 16346
rect 16710 16294 16724 16346
rect 16724 16294 16736 16346
rect 16736 16294 16766 16346
rect 16790 16294 16800 16346
rect 16800 16294 16846 16346
rect 16550 16292 16606 16294
rect 16630 16292 16686 16294
rect 16710 16292 16766 16294
rect 16790 16292 16846 16294
rect 16550 15258 16606 15260
rect 16630 15258 16686 15260
rect 16710 15258 16766 15260
rect 16790 15258 16846 15260
rect 16550 15206 16596 15258
rect 16596 15206 16606 15258
rect 16630 15206 16660 15258
rect 16660 15206 16672 15258
rect 16672 15206 16686 15258
rect 16710 15206 16724 15258
rect 16724 15206 16736 15258
rect 16736 15206 16766 15258
rect 16790 15206 16800 15258
rect 16800 15206 16846 15258
rect 16550 15204 16606 15206
rect 16630 15204 16686 15206
rect 16710 15204 16766 15206
rect 16790 15204 16846 15206
rect 16550 14170 16606 14172
rect 16630 14170 16686 14172
rect 16710 14170 16766 14172
rect 16790 14170 16846 14172
rect 16550 14118 16596 14170
rect 16596 14118 16606 14170
rect 16630 14118 16660 14170
rect 16660 14118 16672 14170
rect 16672 14118 16686 14170
rect 16710 14118 16724 14170
rect 16724 14118 16736 14170
rect 16736 14118 16766 14170
rect 16790 14118 16800 14170
rect 16800 14118 16846 14170
rect 16550 14116 16606 14118
rect 16630 14116 16686 14118
rect 16710 14116 16766 14118
rect 16790 14116 16846 14118
rect 17038 15408 17094 15464
rect 16550 13082 16606 13084
rect 16630 13082 16686 13084
rect 16710 13082 16766 13084
rect 16790 13082 16846 13084
rect 16550 13030 16596 13082
rect 16596 13030 16606 13082
rect 16630 13030 16660 13082
rect 16660 13030 16672 13082
rect 16672 13030 16686 13082
rect 16710 13030 16724 13082
rect 16724 13030 16736 13082
rect 16736 13030 16766 13082
rect 16790 13030 16800 13082
rect 16800 13030 16846 13082
rect 16550 13028 16606 13030
rect 16630 13028 16686 13030
rect 16710 13028 16766 13030
rect 16790 13028 16846 13030
rect 17958 19932 17960 19952
rect 17960 19932 18012 19952
rect 18012 19932 18014 19952
rect 17958 19896 18014 19932
rect 17682 19116 17684 19136
rect 17684 19116 17736 19136
rect 17736 19116 17738 19136
rect 17682 19080 17738 19116
rect 18510 21800 18566 21856
rect 18234 19760 18290 19816
rect 18050 18808 18106 18864
rect 18786 22072 18842 22128
rect 18786 19216 18842 19272
rect 19522 20984 19578 21040
rect 19149 20154 19205 20156
rect 19229 20154 19285 20156
rect 19309 20154 19365 20156
rect 19389 20154 19445 20156
rect 19149 20102 19195 20154
rect 19195 20102 19205 20154
rect 19229 20102 19259 20154
rect 19259 20102 19271 20154
rect 19271 20102 19285 20154
rect 19309 20102 19323 20154
rect 19323 20102 19335 20154
rect 19335 20102 19365 20154
rect 19389 20102 19399 20154
rect 19399 20102 19445 20154
rect 19149 20100 19205 20102
rect 19229 20100 19285 20102
rect 19309 20100 19365 20102
rect 19389 20100 19445 20102
rect 19154 19760 19210 19816
rect 19614 19916 19670 19952
rect 19614 19896 19616 19916
rect 19616 19896 19668 19916
rect 19668 19896 19670 19916
rect 19614 19216 19670 19272
rect 19149 19066 19205 19068
rect 19229 19066 19285 19068
rect 19309 19066 19365 19068
rect 19389 19066 19445 19068
rect 19149 19014 19195 19066
rect 19195 19014 19205 19066
rect 19229 19014 19259 19066
rect 19259 19014 19271 19066
rect 19271 19014 19285 19066
rect 19309 19014 19323 19066
rect 19323 19014 19335 19066
rect 19335 19014 19365 19066
rect 19389 19014 19399 19066
rect 19399 19014 19445 19066
rect 19149 19012 19205 19014
rect 19229 19012 19285 19014
rect 19309 19012 19365 19014
rect 19389 19012 19445 19014
rect 19614 19080 19670 19136
rect 19292 18672 19348 18728
rect 19430 18672 19486 18728
rect 17774 16652 17830 16688
rect 17774 16632 17776 16652
rect 17776 16632 17828 16652
rect 17828 16632 17830 16652
rect 17038 13132 17040 13152
rect 17040 13132 17092 13152
rect 17092 13132 17094 13152
rect 17038 13096 17094 13132
rect 16210 12008 16266 12064
rect 16210 11872 16266 11928
rect 16550 11994 16606 11996
rect 16630 11994 16686 11996
rect 16710 11994 16766 11996
rect 16790 11994 16846 11996
rect 16550 11942 16596 11994
rect 16596 11942 16606 11994
rect 16630 11942 16660 11994
rect 16660 11942 16672 11994
rect 16672 11942 16686 11994
rect 16710 11942 16724 11994
rect 16724 11942 16736 11994
rect 16736 11942 16766 11994
rect 16790 11942 16800 11994
rect 16800 11942 16846 11994
rect 16550 11940 16606 11942
rect 16630 11940 16686 11942
rect 16710 11940 16766 11942
rect 16790 11940 16846 11942
rect 16946 11892 17002 11928
rect 16946 11872 16948 11892
rect 16948 11872 17000 11892
rect 17000 11872 17002 11892
rect 16854 11600 16910 11656
rect 16210 10240 16266 10296
rect 16118 9968 16174 10024
rect 16118 9868 16120 9888
rect 16120 9868 16172 9888
rect 16172 9868 16174 9888
rect 16118 9832 16174 9868
rect 16118 7792 16174 7848
rect 16026 7284 16028 7304
rect 16028 7284 16080 7304
rect 16080 7284 16082 7304
rect 16026 7248 16082 7284
rect 15934 6432 15990 6488
rect 15658 3848 15714 3904
rect 16210 7148 16212 7168
rect 16212 7148 16264 7168
rect 16264 7148 16266 7168
rect 16210 7112 16266 7148
rect 16550 10906 16606 10908
rect 16630 10906 16686 10908
rect 16710 10906 16766 10908
rect 16790 10906 16846 10908
rect 16550 10854 16596 10906
rect 16596 10854 16606 10906
rect 16630 10854 16660 10906
rect 16660 10854 16672 10906
rect 16672 10854 16686 10906
rect 16710 10854 16724 10906
rect 16724 10854 16736 10906
rect 16736 10854 16766 10906
rect 16790 10854 16800 10906
rect 16800 10854 16846 10906
rect 16550 10852 16606 10854
rect 16630 10852 16686 10854
rect 16710 10852 16766 10854
rect 16790 10852 16846 10854
rect 16762 10512 16818 10568
rect 16550 9818 16606 9820
rect 16630 9818 16686 9820
rect 16710 9818 16766 9820
rect 16790 9818 16846 9820
rect 16550 9766 16596 9818
rect 16596 9766 16606 9818
rect 16630 9766 16660 9818
rect 16660 9766 16672 9818
rect 16672 9766 16686 9818
rect 16710 9766 16724 9818
rect 16724 9766 16736 9818
rect 16736 9766 16766 9818
rect 16790 9766 16800 9818
rect 16800 9766 16846 9818
rect 16550 9764 16606 9766
rect 16630 9764 16686 9766
rect 16710 9764 16766 9766
rect 16790 9764 16846 9766
rect 16550 8730 16606 8732
rect 16630 8730 16686 8732
rect 16710 8730 16766 8732
rect 16790 8730 16846 8732
rect 16550 8678 16596 8730
rect 16596 8678 16606 8730
rect 16630 8678 16660 8730
rect 16660 8678 16672 8730
rect 16672 8678 16686 8730
rect 16710 8678 16724 8730
rect 16724 8678 16736 8730
rect 16736 8678 16766 8730
rect 16790 8678 16800 8730
rect 16800 8678 16846 8730
rect 16550 8676 16606 8678
rect 16630 8676 16686 8678
rect 16710 8676 16766 8678
rect 16790 8676 16846 8678
rect 16394 8200 16450 8256
rect 16394 7656 16450 7712
rect 16550 7642 16606 7644
rect 16630 7642 16686 7644
rect 16710 7642 16766 7644
rect 16790 7642 16846 7644
rect 16550 7590 16596 7642
rect 16596 7590 16606 7642
rect 16630 7590 16660 7642
rect 16660 7590 16672 7642
rect 16672 7590 16686 7642
rect 16710 7590 16724 7642
rect 16724 7590 16736 7642
rect 16736 7590 16766 7642
rect 16790 7590 16800 7642
rect 16800 7590 16846 7642
rect 16550 7588 16606 7590
rect 16630 7588 16686 7590
rect 16710 7588 16766 7590
rect 16790 7588 16846 7590
rect 16210 5480 16266 5536
rect 16118 4664 16174 4720
rect 16026 4120 16082 4176
rect 15842 3304 15898 3360
rect 17130 10512 17186 10568
rect 17590 15544 17646 15600
rect 17590 12436 17646 12472
rect 17590 12416 17592 12436
rect 17592 12416 17644 12436
rect 17644 12416 17646 12436
rect 17498 9696 17554 9752
rect 17314 7656 17370 7712
rect 17130 7248 17186 7304
rect 16550 6554 16606 6556
rect 16630 6554 16686 6556
rect 16710 6554 16766 6556
rect 16790 6554 16846 6556
rect 16550 6502 16596 6554
rect 16596 6502 16606 6554
rect 16630 6502 16660 6554
rect 16660 6502 16672 6554
rect 16672 6502 16686 6554
rect 16710 6502 16724 6554
rect 16724 6502 16736 6554
rect 16736 6502 16766 6554
rect 16790 6502 16800 6554
rect 16800 6502 16846 6554
rect 16550 6500 16606 6502
rect 16630 6500 16686 6502
rect 16710 6500 16766 6502
rect 16790 6500 16846 6502
rect 16550 5466 16606 5468
rect 16630 5466 16686 5468
rect 16710 5466 16766 5468
rect 16790 5466 16846 5468
rect 16550 5414 16596 5466
rect 16596 5414 16606 5466
rect 16630 5414 16660 5466
rect 16660 5414 16672 5466
rect 16672 5414 16686 5466
rect 16710 5414 16724 5466
rect 16724 5414 16736 5466
rect 16736 5414 16766 5466
rect 16790 5414 16800 5466
rect 16800 5414 16846 5466
rect 16550 5412 16606 5414
rect 16630 5412 16686 5414
rect 16710 5412 16766 5414
rect 16790 5412 16846 5414
rect 17038 6568 17094 6624
rect 16578 5208 16634 5264
rect 16486 5108 16488 5128
rect 16488 5108 16540 5128
rect 16540 5108 16542 5128
rect 16486 5072 16542 5108
rect 16762 4528 16818 4584
rect 16302 4392 16358 4448
rect 16550 4378 16606 4380
rect 16630 4378 16686 4380
rect 16710 4378 16766 4380
rect 16790 4378 16846 4380
rect 16550 4326 16596 4378
rect 16596 4326 16606 4378
rect 16630 4326 16660 4378
rect 16660 4326 16672 4378
rect 16672 4326 16686 4378
rect 16710 4326 16724 4378
rect 16724 4326 16736 4378
rect 16736 4326 16766 4378
rect 16790 4326 16800 4378
rect 16800 4326 16846 4378
rect 16550 4324 16606 4326
rect 16630 4324 16686 4326
rect 16710 4324 16766 4326
rect 16790 4324 16846 4326
rect 16550 3290 16606 3292
rect 16630 3290 16686 3292
rect 16710 3290 16766 3292
rect 16790 3290 16846 3292
rect 16550 3238 16596 3290
rect 16596 3238 16606 3290
rect 16630 3238 16660 3290
rect 16660 3238 16672 3290
rect 16672 3238 16686 3290
rect 16710 3238 16724 3290
rect 16724 3238 16736 3290
rect 16736 3238 16766 3290
rect 16790 3238 16800 3290
rect 16800 3238 16846 3290
rect 16550 3236 16606 3238
rect 16630 3236 16686 3238
rect 16710 3236 16766 3238
rect 16790 3236 16846 3238
rect 17222 4548 17278 4584
rect 17222 4528 17224 4548
rect 17224 4528 17276 4548
rect 17276 4528 17278 4548
rect 17314 3576 17370 3632
rect 17314 3304 17370 3360
rect 16762 3032 16818 3088
rect 16946 3052 17002 3088
rect 16946 3032 16948 3052
rect 16948 3032 17000 3052
rect 17000 3032 17002 3052
rect 16118 2760 16174 2816
rect 16550 2202 16606 2204
rect 16630 2202 16686 2204
rect 16710 2202 16766 2204
rect 16790 2202 16846 2204
rect 16550 2150 16596 2202
rect 16596 2150 16606 2202
rect 16630 2150 16660 2202
rect 16660 2150 16672 2202
rect 16672 2150 16686 2202
rect 16710 2150 16724 2202
rect 16724 2150 16736 2202
rect 16736 2150 16766 2202
rect 16790 2150 16800 2202
rect 16800 2150 16846 2202
rect 16550 2148 16606 2150
rect 16630 2148 16686 2150
rect 16710 2148 16766 2150
rect 16790 2148 16846 2150
rect 19149 17978 19205 17980
rect 19229 17978 19285 17980
rect 19309 17978 19365 17980
rect 19389 17978 19445 17980
rect 19149 17926 19195 17978
rect 19195 17926 19205 17978
rect 19229 17926 19259 17978
rect 19259 17926 19271 17978
rect 19271 17926 19285 17978
rect 19309 17926 19323 17978
rect 19323 17926 19335 17978
rect 19335 17926 19365 17978
rect 19389 17926 19399 17978
rect 19399 17926 19445 17978
rect 19149 17924 19205 17926
rect 19229 17924 19285 17926
rect 19309 17924 19365 17926
rect 19389 17924 19445 17926
rect 19614 18420 19670 18456
rect 19614 18400 19616 18420
rect 19616 18400 19668 18420
rect 19668 18400 19670 18420
rect 18142 15580 18144 15600
rect 18144 15580 18196 15600
rect 18196 15580 18198 15600
rect 18142 15544 18198 15580
rect 18326 15408 18382 15464
rect 18050 15000 18106 15056
rect 18142 12688 18198 12744
rect 17866 12144 17922 12200
rect 17866 11600 17922 11656
rect 17866 10648 17922 10704
rect 17774 9968 17830 10024
rect 17774 9460 17776 9480
rect 17776 9460 17828 9480
rect 17828 9460 17830 9480
rect 17774 9424 17830 9460
rect 17590 7792 17646 7848
rect 19982 20440 20038 20496
rect 20258 20848 20314 20904
rect 19798 18944 19854 19000
rect 20350 20204 20352 20224
rect 20352 20204 20404 20224
rect 20404 20204 20406 20224
rect 20350 20168 20406 20204
rect 20534 21392 20590 21448
rect 20074 19352 20130 19408
rect 19982 19080 20038 19136
rect 19798 18420 19854 18456
rect 19798 18400 19800 18420
rect 19800 18400 19852 18420
rect 19852 18400 19854 18420
rect 19798 18264 19854 18320
rect 19149 16890 19205 16892
rect 19229 16890 19285 16892
rect 19309 16890 19365 16892
rect 19389 16890 19445 16892
rect 19149 16838 19195 16890
rect 19195 16838 19205 16890
rect 19229 16838 19259 16890
rect 19259 16838 19271 16890
rect 19271 16838 19285 16890
rect 19309 16838 19323 16890
rect 19323 16838 19335 16890
rect 19335 16838 19365 16890
rect 19389 16838 19399 16890
rect 19399 16838 19445 16890
rect 19149 16836 19205 16838
rect 19229 16836 19285 16838
rect 19309 16836 19365 16838
rect 19389 16836 19445 16838
rect 19149 15802 19205 15804
rect 19229 15802 19285 15804
rect 19309 15802 19365 15804
rect 19389 15802 19445 15804
rect 19149 15750 19195 15802
rect 19195 15750 19205 15802
rect 19229 15750 19259 15802
rect 19259 15750 19271 15802
rect 19271 15750 19285 15802
rect 19309 15750 19323 15802
rect 19323 15750 19335 15802
rect 19335 15750 19365 15802
rect 19389 15750 19399 15802
rect 19399 15750 19445 15802
rect 19149 15748 19205 15750
rect 19229 15748 19285 15750
rect 19309 15748 19365 15750
rect 19389 15748 19445 15750
rect 19706 16124 19708 16144
rect 19708 16124 19760 16144
rect 19760 16124 19762 16144
rect 19706 16088 19762 16124
rect 19614 15952 19670 16008
rect 19062 15272 19118 15328
rect 19062 14864 19118 14920
rect 19149 14714 19205 14716
rect 19229 14714 19285 14716
rect 19309 14714 19365 14716
rect 19389 14714 19445 14716
rect 19149 14662 19195 14714
rect 19195 14662 19205 14714
rect 19229 14662 19259 14714
rect 19259 14662 19271 14714
rect 19271 14662 19285 14714
rect 19309 14662 19323 14714
rect 19323 14662 19335 14714
rect 19335 14662 19365 14714
rect 19389 14662 19399 14714
rect 19399 14662 19445 14714
rect 19149 14660 19205 14662
rect 19229 14660 19285 14662
rect 19309 14660 19365 14662
rect 19389 14660 19445 14662
rect 19149 13626 19205 13628
rect 19229 13626 19285 13628
rect 19309 13626 19365 13628
rect 19389 13626 19445 13628
rect 19149 13574 19195 13626
rect 19195 13574 19205 13626
rect 19229 13574 19259 13626
rect 19259 13574 19271 13626
rect 19271 13574 19285 13626
rect 19309 13574 19323 13626
rect 19323 13574 19335 13626
rect 19335 13574 19365 13626
rect 19389 13574 19399 13626
rect 19399 13574 19445 13626
rect 19149 13572 19205 13574
rect 19229 13572 19285 13574
rect 19309 13572 19365 13574
rect 19389 13572 19445 13574
rect 18878 13368 18934 13424
rect 18694 13232 18750 13288
rect 18050 11620 18106 11656
rect 18050 11600 18052 11620
rect 18052 11600 18104 11620
rect 18104 11600 18106 11620
rect 18142 10512 18198 10568
rect 18050 9560 18106 9616
rect 19149 12538 19205 12540
rect 19229 12538 19285 12540
rect 19309 12538 19365 12540
rect 19389 12538 19445 12540
rect 19149 12486 19195 12538
rect 19195 12486 19205 12538
rect 19229 12486 19259 12538
rect 19259 12486 19271 12538
rect 19271 12486 19285 12538
rect 19309 12486 19323 12538
rect 19323 12486 19335 12538
rect 19335 12486 19365 12538
rect 19389 12486 19399 12538
rect 19399 12486 19445 12538
rect 19149 12484 19205 12486
rect 19229 12484 19285 12486
rect 19309 12484 19365 12486
rect 19389 12484 19445 12486
rect 19246 12280 19302 12336
rect 18418 10240 18474 10296
rect 18418 10104 18474 10160
rect 18326 9152 18382 9208
rect 18326 8880 18382 8936
rect 18142 7928 18198 7984
rect 17406 2352 17462 2408
rect 18050 7520 18106 7576
rect 18050 6976 18106 7032
rect 17958 6840 18014 6896
rect 17958 6432 18014 6488
rect 17958 5752 18014 5808
rect 17866 5516 17868 5536
rect 17868 5516 17920 5536
rect 17920 5516 17922 5536
rect 17866 5480 17922 5516
rect 18694 10240 18750 10296
rect 18694 9868 18696 9888
rect 18696 9868 18748 9888
rect 18748 9868 18750 9888
rect 18694 9832 18750 9868
rect 19614 11872 19670 11928
rect 19338 11736 19394 11792
rect 19149 11450 19205 11452
rect 19229 11450 19285 11452
rect 19309 11450 19365 11452
rect 19389 11450 19445 11452
rect 19149 11398 19195 11450
rect 19195 11398 19205 11450
rect 19229 11398 19259 11450
rect 19259 11398 19271 11450
rect 19271 11398 19285 11450
rect 19309 11398 19323 11450
rect 19323 11398 19335 11450
rect 19335 11398 19365 11450
rect 19389 11398 19399 11450
rect 19399 11398 19445 11450
rect 19149 11396 19205 11398
rect 19229 11396 19285 11398
rect 19309 11396 19365 11398
rect 19389 11396 19445 11398
rect 19246 11228 19248 11248
rect 19248 11228 19300 11248
rect 19300 11228 19302 11248
rect 19246 11192 19302 11228
rect 18970 10512 19026 10568
rect 19149 10362 19205 10364
rect 19229 10362 19285 10364
rect 19309 10362 19365 10364
rect 19389 10362 19445 10364
rect 19149 10310 19195 10362
rect 19195 10310 19205 10362
rect 19229 10310 19259 10362
rect 19259 10310 19271 10362
rect 19271 10310 19285 10362
rect 19309 10310 19323 10362
rect 19323 10310 19335 10362
rect 19335 10310 19365 10362
rect 19389 10310 19399 10362
rect 19399 10310 19445 10362
rect 19149 10308 19205 10310
rect 19229 10308 19285 10310
rect 19309 10308 19365 10310
rect 19389 10308 19445 10310
rect 18878 9560 18934 9616
rect 18694 9324 18696 9344
rect 18696 9324 18748 9344
rect 18748 9324 18750 9344
rect 18694 9288 18750 9324
rect 18878 9152 18934 9208
rect 18510 8200 18566 8256
rect 18786 8880 18842 8936
rect 19149 9274 19205 9276
rect 19229 9274 19285 9276
rect 19309 9274 19365 9276
rect 19389 9274 19445 9276
rect 19149 9222 19195 9274
rect 19195 9222 19205 9274
rect 19229 9222 19259 9274
rect 19259 9222 19271 9274
rect 19271 9222 19285 9274
rect 19309 9222 19323 9274
rect 19323 9222 19335 9274
rect 19335 9222 19365 9274
rect 19389 9222 19399 9274
rect 19399 9222 19445 9274
rect 19149 9220 19205 9222
rect 19229 9220 19285 9222
rect 19309 9220 19365 9222
rect 19389 9220 19445 9222
rect 18970 8900 19026 8936
rect 18970 8880 18972 8900
rect 18972 8880 19024 8900
rect 19024 8880 19026 8900
rect 18694 8472 18750 8528
rect 19338 8336 19394 8392
rect 18878 8064 18934 8120
rect 18510 5208 18566 5264
rect 17774 4392 17830 4448
rect 17682 3712 17738 3768
rect 17958 3168 18014 3224
rect 17774 2896 17830 2952
rect 19149 8186 19205 8188
rect 19229 8186 19285 8188
rect 19309 8186 19365 8188
rect 19389 8186 19445 8188
rect 19149 8134 19195 8186
rect 19195 8134 19205 8186
rect 19229 8134 19259 8186
rect 19259 8134 19271 8186
rect 19271 8134 19285 8186
rect 19309 8134 19323 8186
rect 19323 8134 19335 8186
rect 19335 8134 19365 8186
rect 19389 8134 19399 8186
rect 19399 8134 19445 8186
rect 19149 8132 19205 8134
rect 19229 8132 19285 8134
rect 19309 8132 19365 8134
rect 19389 8132 19445 8134
rect 20074 14728 20130 14784
rect 21086 19760 21142 19816
rect 20994 18808 21050 18864
rect 20810 18536 20866 18592
rect 20626 18264 20682 18320
rect 20626 17992 20682 18048
rect 20902 18128 20958 18184
rect 21086 18148 21142 18184
rect 21086 18128 21088 18148
rect 21088 18128 21140 18148
rect 21140 18128 21142 18148
rect 21178 17992 21234 18048
rect 21546 19352 21602 19408
rect 21454 18944 21510 19000
rect 21748 20698 21804 20700
rect 21828 20698 21884 20700
rect 21908 20698 21964 20700
rect 21988 20698 22044 20700
rect 21748 20646 21794 20698
rect 21794 20646 21804 20698
rect 21828 20646 21858 20698
rect 21858 20646 21870 20698
rect 21870 20646 21884 20698
rect 21908 20646 21922 20698
rect 21922 20646 21934 20698
rect 21934 20646 21964 20698
rect 21988 20646 21998 20698
rect 21998 20646 22044 20698
rect 21748 20644 21804 20646
rect 21828 20644 21884 20646
rect 21908 20644 21964 20646
rect 21988 20644 22044 20646
rect 22006 19896 22062 19952
rect 21748 19610 21804 19612
rect 21828 19610 21884 19612
rect 21908 19610 21964 19612
rect 21988 19610 22044 19612
rect 21748 19558 21794 19610
rect 21794 19558 21804 19610
rect 21828 19558 21858 19610
rect 21858 19558 21870 19610
rect 21870 19558 21884 19610
rect 21908 19558 21922 19610
rect 21922 19558 21934 19610
rect 21934 19558 21964 19610
rect 21988 19558 21998 19610
rect 21998 19558 22044 19610
rect 21748 19556 21804 19558
rect 21828 19556 21884 19558
rect 21908 19556 21964 19558
rect 21988 19556 22044 19558
rect 21638 18808 21694 18864
rect 21454 18672 21510 18728
rect 21748 18522 21804 18524
rect 21828 18522 21884 18524
rect 21908 18522 21964 18524
rect 21988 18522 22044 18524
rect 21748 18470 21794 18522
rect 21794 18470 21804 18522
rect 21828 18470 21858 18522
rect 21858 18470 21870 18522
rect 21870 18470 21884 18522
rect 21908 18470 21922 18522
rect 21922 18470 21934 18522
rect 21934 18470 21964 18522
rect 21988 18470 21998 18522
rect 21998 18470 22044 18522
rect 21748 18468 21804 18470
rect 21828 18468 21884 18470
rect 21908 18468 21964 18470
rect 21988 18468 22044 18470
rect 21454 17720 21510 17776
rect 21748 17434 21804 17436
rect 21828 17434 21884 17436
rect 21908 17434 21964 17436
rect 21988 17434 22044 17436
rect 21748 17382 21794 17434
rect 21794 17382 21804 17434
rect 21828 17382 21858 17434
rect 21858 17382 21870 17434
rect 21870 17382 21884 17434
rect 21908 17382 21922 17434
rect 21922 17382 21934 17434
rect 21934 17382 21964 17434
rect 21988 17382 21998 17434
rect 21998 17382 22044 17434
rect 21748 17380 21804 17382
rect 21828 17380 21884 17382
rect 21908 17380 21964 17382
rect 21988 17380 22044 17382
rect 21546 17176 21602 17232
rect 21454 16940 21456 16960
rect 21456 16940 21508 16960
rect 21508 16940 21510 16960
rect 21454 16904 21510 16940
rect 20534 16108 20590 16144
rect 20534 16088 20536 16108
rect 20536 16088 20588 16108
rect 20588 16088 20590 16108
rect 21086 16532 21088 16552
rect 21088 16532 21140 16552
rect 21140 16532 21142 16552
rect 21086 16496 21142 16532
rect 19614 7384 19670 7440
rect 19149 7098 19205 7100
rect 19229 7098 19285 7100
rect 19309 7098 19365 7100
rect 19389 7098 19445 7100
rect 19149 7046 19195 7098
rect 19195 7046 19205 7098
rect 19229 7046 19259 7098
rect 19259 7046 19271 7098
rect 19271 7046 19285 7098
rect 19309 7046 19323 7098
rect 19323 7046 19335 7098
rect 19335 7046 19365 7098
rect 19389 7046 19399 7098
rect 19399 7046 19445 7098
rect 19149 7044 19205 7046
rect 19229 7044 19285 7046
rect 19309 7044 19365 7046
rect 19389 7044 19445 7046
rect 19522 6704 19578 6760
rect 18878 6568 18934 6624
rect 19706 7112 19762 7168
rect 18878 5752 18934 5808
rect 18786 5636 18842 5672
rect 18786 5616 18788 5636
rect 18788 5616 18840 5636
rect 18840 5616 18842 5636
rect 18602 3304 18658 3360
rect 18694 2488 18750 2544
rect 19149 6010 19205 6012
rect 19229 6010 19285 6012
rect 19309 6010 19365 6012
rect 19389 6010 19445 6012
rect 19149 5958 19195 6010
rect 19195 5958 19205 6010
rect 19229 5958 19259 6010
rect 19259 5958 19271 6010
rect 19271 5958 19285 6010
rect 19309 5958 19323 6010
rect 19323 5958 19335 6010
rect 19335 5958 19365 6010
rect 19389 5958 19399 6010
rect 19399 5958 19445 6010
rect 19149 5956 19205 5958
rect 19229 5956 19285 5958
rect 19309 5956 19365 5958
rect 19389 5956 19445 5958
rect 19706 6160 19762 6216
rect 19149 4922 19205 4924
rect 19229 4922 19285 4924
rect 19309 4922 19365 4924
rect 19389 4922 19445 4924
rect 19149 4870 19195 4922
rect 19195 4870 19205 4922
rect 19229 4870 19259 4922
rect 19259 4870 19271 4922
rect 19271 4870 19285 4922
rect 19309 4870 19323 4922
rect 19323 4870 19335 4922
rect 19335 4870 19365 4922
rect 19389 4870 19399 4922
rect 19399 4870 19445 4922
rect 19149 4868 19205 4870
rect 19229 4868 19285 4870
rect 19309 4868 19365 4870
rect 19389 4868 19445 4870
rect 19154 4120 19210 4176
rect 19149 3834 19205 3836
rect 19229 3834 19285 3836
rect 19309 3834 19365 3836
rect 19389 3834 19445 3836
rect 19149 3782 19195 3834
rect 19195 3782 19205 3834
rect 19229 3782 19259 3834
rect 19259 3782 19271 3834
rect 19271 3782 19285 3834
rect 19309 3782 19323 3834
rect 19323 3782 19335 3834
rect 19335 3782 19365 3834
rect 19389 3782 19399 3834
rect 19399 3782 19445 3834
rect 19149 3780 19205 3782
rect 19229 3780 19285 3782
rect 19309 3780 19365 3782
rect 19389 3780 19445 3782
rect 19149 2746 19205 2748
rect 19229 2746 19285 2748
rect 19309 2746 19365 2748
rect 19389 2746 19445 2748
rect 19149 2694 19195 2746
rect 19195 2694 19205 2746
rect 19229 2694 19259 2746
rect 19259 2694 19271 2746
rect 19271 2694 19285 2746
rect 19309 2694 19323 2746
rect 19323 2694 19335 2746
rect 19335 2694 19365 2746
rect 19389 2694 19399 2746
rect 19399 2694 19445 2746
rect 19149 2692 19205 2694
rect 19229 2692 19285 2694
rect 19309 2692 19365 2694
rect 19389 2692 19445 2694
rect 19246 1808 19302 1864
rect 19154 1400 19210 1456
rect 20258 9288 20314 9344
rect 20258 9172 20314 9208
rect 20258 9152 20260 9172
rect 20260 9152 20312 9172
rect 20312 9152 20314 9172
rect 20258 7420 20260 7440
rect 20260 7420 20312 7440
rect 20312 7420 20314 7440
rect 20258 7384 20314 7420
rect 20258 6840 20314 6896
rect 20258 6568 20314 6624
rect 20258 6296 20314 6352
rect 20166 5752 20222 5808
rect 19430 856 19486 912
rect 20534 11192 20590 11248
rect 20442 10648 20498 10704
rect 21748 16346 21804 16348
rect 21828 16346 21884 16348
rect 21908 16346 21964 16348
rect 21988 16346 22044 16348
rect 21748 16294 21794 16346
rect 21794 16294 21804 16346
rect 21828 16294 21858 16346
rect 21858 16294 21870 16346
rect 21870 16294 21884 16346
rect 21908 16294 21922 16346
rect 21922 16294 21934 16346
rect 21934 16294 21964 16346
rect 21988 16294 21998 16346
rect 21998 16294 22044 16346
rect 21748 16292 21804 16294
rect 21828 16292 21884 16294
rect 21908 16292 21964 16294
rect 21988 16292 22044 16294
rect 21454 16088 21510 16144
rect 21454 15680 21510 15736
rect 21638 15544 21694 15600
rect 21454 15408 21510 15464
rect 21546 15272 21602 15328
rect 21086 14884 21142 14920
rect 21086 14864 21088 14884
rect 21088 14864 21140 14884
rect 21140 14864 21142 14884
rect 21454 14456 21510 14512
rect 21454 13912 21510 13968
rect 21454 13676 21456 13696
rect 21456 13676 21508 13696
rect 21508 13676 21510 13696
rect 21454 13640 21510 13676
rect 21454 13232 21510 13288
rect 21086 12824 21142 12880
rect 20718 12164 20774 12200
rect 20718 12144 20720 12164
rect 20720 12144 20772 12164
rect 20772 12144 20774 12164
rect 20718 11600 20774 11656
rect 20718 10004 20720 10024
rect 20720 10004 20772 10024
rect 20772 10004 20774 10024
rect 20718 9968 20774 10004
rect 20442 8744 20498 8800
rect 20350 3712 20406 3768
rect 20258 2896 20314 2952
rect 20718 8492 20774 8528
rect 20718 8472 20720 8492
rect 20720 8472 20772 8492
rect 20772 8472 20774 8492
rect 20718 8356 20774 8392
rect 20718 8336 20720 8356
rect 20720 8336 20772 8356
rect 20772 8336 20774 8356
rect 21086 11192 21142 11248
rect 20902 9016 20958 9072
rect 21454 12416 21510 12472
rect 21362 12280 21418 12336
rect 21454 12144 21510 12200
rect 20626 6740 20628 6760
rect 20628 6740 20680 6760
rect 20680 6740 20682 6760
rect 20626 6704 20682 6740
rect 20902 7284 20904 7304
rect 20904 7284 20956 7304
rect 20956 7284 20958 7304
rect 20902 7248 20958 7284
rect 20718 6160 20774 6216
rect 21086 7792 21142 7848
rect 21086 7692 21088 7712
rect 21088 7692 21140 7712
rect 21140 7692 21142 7712
rect 21086 7656 21142 7692
rect 20994 5752 21050 5808
rect 20810 4120 20866 4176
rect 20810 3848 20866 3904
rect 20994 5208 21050 5264
rect 20994 4664 21050 4720
rect 20994 3984 21050 4040
rect 20810 3460 20866 3496
rect 20810 3440 20812 3460
rect 20812 3440 20864 3460
rect 20864 3440 20866 3460
rect 20718 3168 20774 3224
rect 20534 2624 20590 2680
rect 20718 992 20774 1048
rect 21546 8608 21602 8664
rect 21454 7520 21510 7576
rect 21454 7112 21510 7168
rect 21270 5652 21272 5672
rect 21272 5652 21324 5672
rect 21324 5652 21326 5672
rect 21270 5616 21326 5652
rect 21454 6160 21510 6216
rect 21270 3848 21326 3904
rect 21270 3304 21326 3360
rect 21546 3032 21602 3088
rect 21748 15258 21804 15260
rect 21828 15258 21884 15260
rect 21908 15258 21964 15260
rect 21988 15258 22044 15260
rect 21748 15206 21794 15258
rect 21794 15206 21804 15258
rect 21828 15206 21858 15258
rect 21858 15206 21870 15258
rect 21870 15206 21884 15258
rect 21908 15206 21922 15258
rect 21922 15206 21934 15258
rect 21934 15206 21964 15258
rect 21988 15206 21998 15258
rect 21998 15206 22044 15258
rect 21748 15204 21804 15206
rect 21828 15204 21884 15206
rect 21908 15204 21964 15206
rect 21988 15204 22044 15206
rect 21748 14170 21804 14172
rect 21828 14170 21884 14172
rect 21908 14170 21964 14172
rect 21988 14170 22044 14172
rect 21748 14118 21794 14170
rect 21794 14118 21804 14170
rect 21828 14118 21858 14170
rect 21858 14118 21870 14170
rect 21870 14118 21884 14170
rect 21908 14118 21922 14170
rect 21922 14118 21934 14170
rect 21934 14118 21964 14170
rect 21988 14118 21998 14170
rect 21998 14118 22044 14170
rect 21748 14116 21804 14118
rect 21828 14116 21884 14118
rect 21908 14116 21964 14118
rect 21988 14116 22044 14118
rect 22006 13776 22062 13832
rect 21748 13082 21804 13084
rect 21828 13082 21884 13084
rect 21908 13082 21964 13084
rect 21988 13082 22044 13084
rect 21748 13030 21794 13082
rect 21794 13030 21804 13082
rect 21828 13030 21858 13082
rect 21858 13030 21870 13082
rect 21870 13030 21884 13082
rect 21908 13030 21922 13082
rect 21922 13030 21934 13082
rect 21934 13030 21964 13082
rect 21988 13030 21998 13082
rect 21998 13030 22044 13082
rect 21748 13028 21804 13030
rect 21828 13028 21884 13030
rect 21908 13028 21964 13030
rect 21988 13028 22044 13030
rect 21730 12280 21786 12336
rect 21748 11994 21804 11996
rect 21828 11994 21884 11996
rect 21908 11994 21964 11996
rect 21988 11994 22044 11996
rect 21748 11942 21794 11994
rect 21794 11942 21804 11994
rect 21828 11942 21858 11994
rect 21858 11942 21870 11994
rect 21870 11942 21884 11994
rect 21908 11942 21922 11994
rect 21922 11942 21934 11994
rect 21934 11942 21964 11994
rect 21988 11942 21998 11994
rect 21998 11942 22044 11994
rect 21748 11940 21804 11942
rect 21828 11940 21884 11942
rect 21908 11940 21964 11942
rect 21988 11940 22044 11942
rect 21748 10906 21804 10908
rect 21828 10906 21884 10908
rect 21908 10906 21964 10908
rect 21988 10906 22044 10908
rect 21748 10854 21794 10906
rect 21794 10854 21804 10906
rect 21828 10854 21858 10906
rect 21858 10854 21870 10906
rect 21870 10854 21884 10906
rect 21908 10854 21922 10906
rect 21922 10854 21934 10906
rect 21934 10854 21964 10906
rect 21988 10854 21998 10906
rect 21998 10854 22044 10906
rect 21748 10852 21804 10854
rect 21828 10852 21884 10854
rect 21908 10852 21964 10854
rect 21988 10852 22044 10854
rect 21748 9818 21804 9820
rect 21828 9818 21884 9820
rect 21908 9818 21964 9820
rect 21988 9818 22044 9820
rect 21748 9766 21794 9818
rect 21794 9766 21804 9818
rect 21828 9766 21858 9818
rect 21858 9766 21870 9818
rect 21870 9766 21884 9818
rect 21908 9766 21922 9818
rect 21922 9766 21934 9818
rect 21934 9766 21964 9818
rect 21988 9766 21998 9818
rect 21998 9766 22044 9818
rect 21748 9764 21804 9766
rect 21828 9764 21884 9766
rect 21908 9764 21964 9766
rect 21988 9764 22044 9766
rect 21748 8730 21804 8732
rect 21828 8730 21884 8732
rect 21908 8730 21964 8732
rect 21988 8730 22044 8732
rect 21748 8678 21794 8730
rect 21794 8678 21804 8730
rect 21828 8678 21858 8730
rect 21858 8678 21870 8730
rect 21870 8678 21884 8730
rect 21908 8678 21922 8730
rect 21922 8678 21934 8730
rect 21934 8678 21964 8730
rect 21988 8678 21998 8730
rect 21998 8678 22044 8730
rect 21748 8676 21804 8678
rect 21828 8676 21884 8678
rect 21908 8676 21964 8678
rect 21988 8676 22044 8678
rect 21730 8064 21786 8120
rect 21748 7642 21804 7644
rect 21828 7642 21884 7644
rect 21908 7642 21964 7644
rect 21988 7642 22044 7644
rect 21748 7590 21794 7642
rect 21794 7590 21804 7642
rect 21828 7590 21858 7642
rect 21858 7590 21870 7642
rect 21870 7590 21884 7642
rect 21908 7590 21922 7642
rect 21922 7590 21934 7642
rect 21934 7590 21964 7642
rect 21988 7590 21998 7642
rect 21998 7590 22044 7642
rect 21748 7588 21804 7590
rect 21828 7588 21884 7590
rect 21908 7588 21964 7590
rect 21988 7588 22044 7590
rect 21748 6554 21804 6556
rect 21828 6554 21884 6556
rect 21908 6554 21964 6556
rect 21988 6554 22044 6556
rect 21748 6502 21794 6554
rect 21794 6502 21804 6554
rect 21828 6502 21858 6554
rect 21858 6502 21870 6554
rect 21870 6502 21884 6554
rect 21908 6502 21922 6554
rect 21922 6502 21934 6554
rect 21934 6502 21964 6554
rect 21988 6502 21998 6554
rect 21998 6502 22044 6554
rect 21748 6500 21804 6502
rect 21828 6500 21884 6502
rect 21908 6500 21964 6502
rect 21988 6500 22044 6502
rect 21748 5466 21804 5468
rect 21828 5466 21884 5468
rect 21908 5466 21964 5468
rect 21988 5466 22044 5468
rect 21748 5414 21794 5466
rect 21794 5414 21804 5466
rect 21828 5414 21858 5466
rect 21858 5414 21870 5466
rect 21870 5414 21884 5466
rect 21908 5414 21922 5466
rect 21922 5414 21934 5466
rect 21934 5414 21964 5466
rect 21988 5414 21998 5466
rect 21998 5414 22044 5466
rect 21748 5412 21804 5414
rect 21828 5412 21884 5414
rect 21908 5412 21964 5414
rect 21988 5412 22044 5414
rect 21730 5072 21786 5128
rect 22006 5072 22062 5128
rect 22006 4700 22008 4720
rect 22008 4700 22060 4720
rect 22060 4700 22062 4720
rect 22006 4664 22062 4700
rect 21748 4378 21804 4380
rect 21828 4378 21884 4380
rect 21908 4378 21964 4380
rect 21988 4378 22044 4380
rect 21748 4326 21794 4378
rect 21794 4326 21804 4378
rect 21828 4326 21858 4378
rect 21858 4326 21870 4378
rect 21870 4326 21884 4378
rect 21908 4326 21922 4378
rect 21922 4326 21934 4378
rect 21934 4326 21964 4378
rect 21988 4326 21998 4378
rect 21998 4326 22044 4378
rect 21748 4324 21804 4326
rect 21828 4324 21884 4326
rect 21908 4324 21964 4326
rect 21988 4324 22044 4326
rect 21748 3290 21804 3292
rect 21828 3290 21884 3292
rect 21908 3290 21964 3292
rect 21988 3290 22044 3292
rect 21748 3238 21794 3290
rect 21794 3238 21804 3290
rect 21828 3238 21858 3290
rect 21858 3238 21870 3290
rect 21870 3238 21884 3290
rect 21908 3238 21922 3290
rect 21922 3238 21934 3290
rect 21934 3238 21964 3290
rect 21988 3238 21998 3290
rect 21998 3238 22044 3290
rect 21748 3236 21804 3238
rect 21828 3236 21884 3238
rect 21908 3236 21964 3238
rect 21988 3236 22044 3238
rect 21748 2202 21804 2204
rect 21828 2202 21884 2204
rect 21908 2202 21964 2204
rect 21988 2202 22044 2204
rect 21748 2150 21794 2202
rect 21794 2150 21804 2202
rect 21828 2150 21858 2202
rect 21858 2150 21870 2202
rect 21870 2150 21884 2202
rect 21908 2150 21922 2202
rect 21922 2150 21934 2202
rect 21934 2150 21964 2202
rect 21988 2150 21998 2202
rect 21998 2150 22044 2202
rect 21748 2148 21804 2150
rect 21828 2148 21884 2150
rect 21908 2148 21964 2150
rect 21988 2148 22044 2150
<< metal3 >>
rect 54 22476 60 22540
rect 124 22538 130 22540
rect 14406 22538 14412 22540
rect 124 22478 14412 22538
rect 124 22476 130 22478
rect 14406 22476 14412 22478
rect 14476 22476 14482 22540
rect 0 22266 800 22296
rect 2313 22266 2379 22269
rect 22200 22266 23000 22296
rect 0 22264 2379 22266
rect 0 22208 2318 22264
rect 2374 22208 2379 22264
rect 0 22206 2379 22208
rect 0 22176 800 22206
rect 2313 22203 2379 22206
rect 19014 22206 23000 22266
rect 18781 22130 18847 22133
rect 19014 22130 19074 22206
rect 22200 22176 23000 22206
rect 18781 22128 19074 22130
rect 18781 22072 18786 22128
rect 18842 22072 19074 22128
rect 18781 22070 19074 22072
rect 18781 22067 18847 22070
rect 0 21858 800 21888
rect 4061 21858 4127 21861
rect 0 21856 4127 21858
rect 0 21800 4066 21856
rect 4122 21800 4127 21856
rect 0 21798 4127 21800
rect 0 21768 800 21798
rect 4061 21795 4127 21798
rect 18505 21858 18571 21861
rect 22200 21858 23000 21888
rect 18505 21856 23000 21858
rect 18505 21800 18510 21856
rect 18566 21800 23000 21856
rect 18505 21798 23000 21800
rect 18505 21795 18571 21798
rect 22200 21768 23000 21798
rect 0 21450 800 21480
rect 1761 21450 1827 21453
rect 0 21448 1827 21450
rect 0 21392 1766 21448
rect 1822 21392 1827 21448
rect 0 21390 1827 21392
rect 0 21360 800 21390
rect 1761 21387 1827 21390
rect 7097 21450 7163 21453
rect 14457 21450 14523 21453
rect 7097 21448 14523 21450
rect 7097 21392 7102 21448
rect 7158 21392 14462 21448
rect 14518 21392 14523 21448
rect 7097 21390 14523 21392
rect 7097 21387 7163 21390
rect 14457 21387 14523 21390
rect 20529 21450 20595 21453
rect 22200 21450 23000 21480
rect 20529 21448 23000 21450
rect 20529 21392 20534 21448
rect 20590 21392 23000 21448
rect 20529 21390 23000 21392
rect 20529 21387 20595 21390
rect 22200 21360 23000 21390
rect 1117 21314 1183 21317
rect 12750 21314 12756 21316
rect 1117 21312 12756 21314
rect 1117 21256 1122 21312
rect 1178 21256 12756 21312
rect 1117 21254 12756 21256
rect 1117 21251 1183 21254
rect 12750 21252 12756 21254
rect 12820 21252 12826 21316
rect 1158 21116 1164 21180
rect 1228 21178 1234 21180
rect 7097 21178 7163 21181
rect 1228 21176 7163 21178
rect 1228 21120 7102 21176
rect 7158 21120 7163 21176
rect 1228 21118 7163 21120
rect 1228 21116 1234 21118
rect 7097 21115 7163 21118
rect 0 21042 800 21072
rect 2221 21042 2287 21045
rect 0 21040 2287 21042
rect 0 20984 2226 21040
rect 2282 20984 2287 21040
rect 0 20982 2287 20984
rect 0 20952 800 20982
rect 2221 20979 2287 20982
rect 4838 20980 4844 21044
rect 4908 21042 4914 21044
rect 17769 21042 17835 21045
rect 4908 21040 17835 21042
rect 4908 20984 17774 21040
rect 17830 20984 17835 21040
rect 4908 20982 17835 20984
rect 4908 20980 4914 20982
rect 17769 20979 17835 20982
rect 19517 21042 19583 21045
rect 22200 21042 23000 21072
rect 19517 21040 23000 21042
rect 19517 20984 19522 21040
rect 19578 20984 23000 21040
rect 19517 20982 23000 20984
rect 19517 20979 19583 20982
rect 22200 20952 23000 20982
rect 2129 20906 2195 20909
rect 2129 20904 8080 20906
rect 2129 20848 2134 20904
rect 2190 20848 8080 20904
rect 2129 20846 8080 20848
rect 2129 20843 2195 20846
rect 8020 20770 8080 20846
rect 8150 20844 8156 20908
rect 8220 20906 8226 20908
rect 20253 20906 20319 20909
rect 8220 20904 20319 20906
rect 8220 20848 20258 20904
rect 20314 20848 20319 20904
rect 8220 20846 20319 20848
rect 8220 20844 8226 20846
rect 20253 20843 20319 20846
rect 11094 20770 11100 20772
rect 8020 20710 11100 20770
rect 11094 20708 11100 20710
rect 11164 20708 11170 20772
rect 6144 20704 6460 20705
rect 0 20634 800 20664
rect 6144 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6460 20704
rect 6144 20639 6460 20640
rect 11342 20704 11658 20705
rect 11342 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11658 20704
rect 11342 20639 11658 20640
rect 16540 20704 16856 20705
rect 16540 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16856 20704
rect 16540 20639 16856 20640
rect 21738 20704 22054 20705
rect 21738 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22054 20704
rect 21738 20639 22054 20640
rect 1853 20634 1919 20637
rect 22200 20634 23000 20664
rect 0 20632 1919 20634
rect 0 20576 1858 20632
rect 1914 20576 1919 20632
rect 0 20574 1919 20576
rect 0 20544 800 20574
rect 1853 20571 1919 20574
rect 22142 20544 23000 20634
rect 2865 20498 2931 20501
rect 5349 20498 5415 20501
rect 7281 20498 7347 20501
rect 13629 20498 13695 20501
rect 2865 20496 5274 20498
rect 2865 20440 2870 20496
rect 2926 20440 5274 20496
rect 2865 20438 5274 20440
rect 2865 20435 2931 20438
rect 3509 20362 3575 20365
rect 4613 20362 4679 20365
rect 3509 20360 4679 20362
rect 3509 20304 3514 20360
rect 3570 20304 4618 20360
rect 4674 20304 4679 20360
rect 3509 20302 4679 20304
rect 5214 20362 5274 20438
rect 5349 20496 13695 20498
rect 5349 20440 5354 20496
rect 5410 20440 7286 20496
rect 7342 20440 13634 20496
rect 13690 20440 13695 20496
rect 5349 20438 13695 20440
rect 5349 20435 5415 20438
rect 7281 20435 7347 20438
rect 13629 20435 13695 20438
rect 19977 20498 20043 20501
rect 22142 20498 22202 20544
rect 19977 20496 22202 20498
rect 19977 20440 19982 20496
rect 20038 20440 22202 20496
rect 19977 20438 22202 20440
rect 19977 20435 20043 20438
rect 7833 20362 7899 20365
rect 5214 20360 7899 20362
rect 5214 20304 7838 20360
rect 7894 20304 7899 20360
rect 5214 20302 7899 20304
rect 3509 20299 3575 20302
rect 4613 20299 4679 20302
rect 7833 20299 7899 20302
rect 10777 20362 10843 20365
rect 14590 20362 14596 20364
rect 10777 20360 14596 20362
rect 10777 20304 10782 20360
rect 10838 20304 14596 20360
rect 10777 20302 14596 20304
rect 10777 20299 10843 20302
rect 14590 20300 14596 20302
rect 14660 20300 14666 20364
rect 0 20226 800 20256
rect 1485 20226 1551 20229
rect 0 20224 1551 20226
rect 0 20168 1490 20224
rect 1546 20168 1551 20224
rect 0 20166 1551 20168
rect 0 20136 800 20166
rect 1485 20163 1551 20166
rect 2129 20226 2195 20229
rect 2446 20226 2452 20228
rect 2129 20224 2452 20226
rect 2129 20168 2134 20224
rect 2190 20168 2452 20224
rect 2129 20166 2452 20168
rect 2129 20163 2195 20166
rect 2446 20164 2452 20166
rect 2516 20164 2522 20228
rect 20345 20226 20411 20229
rect 22200 20226 23000 20256
rect 20345 20224 23000 20226
rect 20345 20168 20350 20224
rect 20406 20168 23000 20224
rect 20345 20166 23000 20168
rect 20345 20163 20411 20166
rect 3545 20160 3861 20161
rect 3545 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3861 20160
rect 3545 20095 3861 20096
rect 8743 20160 9059 20161
rect 8743 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9059 20160
rect 8743 20095 9059 20096
rect 13941 20160 14257 20161
rect 13941 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14257 20160
rect 13941 20095 14257 20096
rect 19139 20160 19455 20161
rect 19139 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19455 20160
rect 22200 20136 23000 20166
rect 19139 20095 19455 20096
rect 4153 20090 4219 20093
rect 5625 20090 5691 20093
rect 4153 20088 5691 20090
rect 4153 20032 4158 20088
rect 4214 20032 5630 20088
rect 5686 20032 5691 20088
rect 4153 20030 5691 20032
rect 4153 20027 4219 20030
rect 5625 20027 5691 20030
rect 7741 20090 7807 20093
rect 8334 20090 8340 20092
rect 7741 20088 8340 20090
rect 7741 20032 7746 20088
rect 7802 20032 8340 20088
rect 7741 20030 8340 20032
rect 7741 20027 7807 20030
rect 8334 20028 8340 20030
rect 8404 20028 8410 20092
rect 16389 20090 16455 20093
rect 16389 20088 19074 20090
rect 16389 20032 16394 20088
rect 16450 20032 19074 20088
rect 16389 20030 19074 20032
rect 16389 20027 16455 20030
rect 3141 19954 3207 19957
rect 17953 19954 18019 19957
rect 3141 19952 18019 19954
rect 3141 19896 3146 19952
rect 3202 19896 17958 19952
rect 18014 19896 18019 19952
rect 3141 19894 18019 19896
rect 19014 19954 19074 20030
rect 19609 19954 19675 19957
rect 22001 19954 22067 19957
rect 19014 19952 19675 19954
rect 19014 19896 19614 19952
rect 19670 19896 19675 19952
rect 19014 19894 19675 19896
rect 3141 19891 3207 19894
rect 17953 19891 18019 19894
rect 19609 19891 19675 19894
rect 20854 19952 22067 19954
rect 20854 19896 22006 19952
rect 22062 19896 22067 19952
rect 20854 19894 22067 19896
rect 0 19818 800 19848
rect 1853 19818 1919 19821
rect 0 19816 1919 19818
rect 0 19760 1858 19816
rect 1914 19760 1919 19816
rect 0 19758 1919 19760
rect 0 19728 800 19758
rect 1853 19755 1919 19758
rect 2037 19818 2103 19821
rect 18229 19818 18295 19821
rect 2037 19816 18295 19818
rect 2037 19760 2042 19816
rect 2098 19760 18234 19816
rect 18290 19760 18295 19816
rect 2037 19758 18295 19760
rect 2037 19755 2103 19758
rect 18229 19755 18295 19758
rect 19149 19818 19215 19821
rect 20854 19818 20914 19894
rect 22001 19891 22067 19894
rect 19149 19816 20914 19818
rect 19149 19760 19154 19816
rect 19210 19760 20914 19816
rect 19149 19758 20914 19760
rect 21081 19818 21147 19821
rect 22200 19818 23000 19848
rect 21081 19816 23000 19818
rect 21081 19760 21086 19816
rect 21142 19760 23000 19816
rect 21081 19758 23000 19760
rect 19149 19755 19215 19758
rect 21081 19755 21147 19758
rect 22200 19728 23000 19758
rect 6144 19616 6460 19617
rect 6144 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6460 19616
rect 6144 19551 6460 19552
rect 11342 19616 11658 19617
rect 11342 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11658 19616
rect 11342 19551 11658 19552
rect 16540 19616 16856 19617
rect 16540 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16856 19616
rect 16540 19551 16856 19552
rect 21738 19616 22054 19617
rect 21738 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22054 19616
rect 21738 19551 22054 19552
rect 4521 19548 4587 19549
rect 4470 19546 4476 19548
rect 4430 19486 4476 19546
rect 4540 19544 4587 19548
rect 4582 19488 4587 19544
rect 4470 19484 4476 19486
rect 4540 19484 4587 19488
rect 4521 19483 4587 19484
rect 8201 19546 8267 19549
rect 8518 19546 8524 19548
rect 8201 19544 8524 19546
rect 8201 19488 8206 19544
rect 8262 19488 8524 19544
rect 8201 19486 8524 19488
rect 8201 19483 8267 19486
rect 8518 19484 8524 19486
rect 8588 19484 8594 19548
rect 0 19410 800 19440
rect 1485 19410 1551 19413
rect 0 19408 1551 19410
rect 0 19352 1490 19408
rect 1546 19352 1551 19408
rect 0 19350 1551 19352
rect 0 19320 800 19350
rect 1485 19347 1551 19350
rect 3417 19410 3483 19413
rect 7414 19410 7420 19412
rect 3417 19408 7420 19410
rect 3417 19352 3422 19408
rect 3478 19352 7420 19408
rect 3417 19350 7420 19352
rect 3417 19347 3483 19350
rect 7414 19348 7420 19350
rect 7484 19348 7490 19412
rect 7782 19348 7788 19412
rect 7852 19410 7858 19412
rect 9489 19410 9555 19413
rect 7852 19408 9555 19410
rect 7852 19352 9494 19408
rect 9550 19352 9555 19408
rect 7852 19350 9555 19352
rect 7852 19348 7858 19350
rect 9489 19347 9555 19350
rect 10225 19410 10291 19413
rect 10777 19410 10843 19413
rect 10225 19408 10843 19410
rect 10225 19352 10230 19408
rect 10286 19352 10782 19408
rect 10838 19352 10843 19408
rect 10225 19350 10843 19352
rect 10225 19347 10291 19350
rect 10777 19347 10843 19350
rect 16849 19410 16915 19413
rect 20069 19410 20135 19413
rect 16849 19408 20135 19410
rect 16849 19352 16854 19408
rect 16910 19352 20074 19408
rect 20130 19352 20135 19408
rect 16849 19350 20135 19352
rect 16849 19347 16915 19350
rect 3325 19274 3391 19277
rect 6453 19274 6519 19277
rect 10869 19274 10935 19277
rect 3325 19272 6519 19274
rect 3325 19216 3330 19272
rect 3386 19216 6458 19272
rect 6514 19216 6519 19272
rect 3325 19214 6519 19216
rect 3325 19211 3391 19214
rect 6453 19211 6519 19214
rect 6686 19272 10935 19274
rect 6686 19216 10874 19272
rect 10930 19216 10935 19272
rect 6686 19214 10935 19216
rect 18646 19274 18706 19350
rect 20069 19347 20135 19350
rect 21541 19410 21607 19413
rect 22200 19410 23000 19440
rect 21541 19408 23000 19410
rect 21541 19352 21546 19408
rect 21602 19352 23000 19408
rect 21541 19350 23000 19352
rect 21541 19347 21607 19350
rect 22200 19320 23000 19350
rect 18781 19274 18847 19277
rect 19609 19276 19675 19277
rect 19558 19274 19564 19276
rect 18646 19272 18847 19274
rect 18646 19216 18786 19272
rect 18842 19216 18847 19272
rect 18646 19214 18847 19216
rect 19518 19214 19564 19274
rect 19628 19272 19675 19276
rect 19670 19216 19675 19272
rect 2497 19138 2563 19141
rect 2865 19138 2931 19141
rect 4889 19138 4955 19141
rect 6686 19138 6746 19214
rect 10869 19211 10935 19214
rect 18781 19211 18847 19214
rect 19558 19212 19564 19214
rect 19628 19212 19675 19216
rect 19609 19211 19675 19212
rect 2497 19136 2931 19138
rect 2497 19080 2502 19136
rect 2558 19080 2870 19136
rect 2926 19080 2931 19136
rect 2497 19078 2931 19080
rect 2497 19075 2563 19078
rect 2865 19075 2931 19078
rect 3926 19136 6746 19138
rect 3926 19080 4894 19136
rect 4950 19080 6746 19136
rect 3926 19078 6746 19080
rect 17677 19138 17743 19141
rect 17902 19138 17908 19140
rect 17677 19136 17908 19138
rect 17677 19080 17682 19136
rect 17738 19080 17908 19136
rect 17677 19078 17908 19080
rect 3545 19072 3861 19073
rect 0 19002 800 19032
rect 3545 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3861 19072
rect 3545 19007 3861 19008
rect 1485 19002 1551 19005
rect 0 19000 1551 19002
rect 0 18944 1490 19000
rect 1546 18944 1551 19000
rect 0 18942 1551 18944
rect 0 18912 800 18942
rect 1485 18939 1551 18942
rect 2589 18866 2655 18869
rect 3926 18866 3986 19078
rect 4889 19075 4955 19078
rect 17677 19075 17743 19078
rect 17902 19076 17908 19078
rect 17972 19076 17978 19140
rect 19609 19138 19675 19141
rect 19977 19138 20043 19141
rect 19609 19136 20043 19138
rect 19609 19080 19614 19136
rect 19670 19080 19982 19136
rect 20038 19080 20043 19136
rect 19609 19078 20043 19080
rect 19609 19075 19675 19078
rect 19977 19075 20043 19078
rect 8743 19072 9059 19073
rect 8743 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9059 19072
rect 8743 19007 9059 19008
rect 13941 19072 14257 19073
rect 13941 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14257 19072
rect 13941 19007 14257 19008
rect 19139 19072 19455 19073
rect 19139 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19455 19072
rect 19139 19007 19455 19008
rect 5349 19002 5415 19005
rect 8201 19002 8267 19005
rect 5349 19000 8267 19002
rect 5349 18944 5354 19000
rect 5410 18944 8206 19000
rect 8262 18944 8267 19000
rect 5349 18942 8267 18944
rect 5349 18939 5415 18942
rect 8201 18939 8267 18942
rect 19793 19002 19859 19005
rect 19926 19002 19932 19004
rect 19793 19000 19932 19002
rect 19793 18944 19798 19000
rect 19854 18944 19932 19000
rect 19793 18942 19932 18944
rect 19793 18939 19859 18942
rect 19926 18940 19932 18942
rect 19996 18940 20002 19004
rect 21449 19002 21515 19005
rect 22200 19002 23000 19032
rect 21449 19000 23000 19002
rect 21449 18944 21454 19000
rect 21510 18944 23000 19000
rect 21449 18942 23000 18944
rect 21449 18939 21515 18942
rect 22200 18912 23000 18942
rect 2589 18864 3986 18866
rect 2589 18808 2594 18864
rect 2650 18808 3986 18864
rect 2589 18806 3986 18808
rect 2589 18803 2655 18806
rect 5758 18804 5764 18868
rect 5828 18866 5834 18868
rect 5901 18866 5967 18869
rect 5828 18864 5967 18866
rect 5828 18808 5906 18864
rect 5962 18808 5967 18864
rect 5828 18806 5967 18808
rect 5828 18804 5834 18806
rect 5901 18803 5967 18806
rect 6821 18866 6887 18869
rect 10726 18866 10732 18868
rect 6821 18864 10732 18866
rect 6821 18808 6826 18864
rect 6882 18808 10732 18864
rect 6821 18806 10732 18808
rect 6821 18803 6887 18806
rect 10726 18804 10732 18806
rect 10796 18804 10802 18868
rect 18045 18866 18111 18869
rect 20989 18866 21055 18869
rect 21633 18866 21699 18869
rect 18045 18864 21055 18866
rect 18045 18808 18050 18864
rect 18106 18808 20994 18864
rect 21050 18808 21055 18864
rect 18045 18806 21055 18808
rect 18045 18803 18111 18806
rect 20989 18803 21055 18806
rect 21222 18864 21699 18866
rect 21222 18808 21638 18864
rect 21694 18808 21699 18864
rect 21222 18806 21699 18808
rect 2681 18730 2747 18733
rect 2957 18730 3023 18733
rect 5809 18730 5875 18733
rect 6453 18730 6519 18733
rect 2681 18728 2790 18730
rect 2681 18672 2686 18728
rect 2742 18672 2790 18728
rect 2681 18667 2790 18672
rect 2957 18728 6010 18730
rect 2957 18672 2962 18728
rect 3018 18672 5814 18728
rect 5870 18672 6010 18728
rect 2957 18670 6010 18672
rect 2957 18667 3023 18670
rect 5809 18667 5875 18670
rect 0 18594 800 18624
rect 1485 18594 1551 18597
rect 0 18592 1551 18594
rect 0 18536 1490 18592
rect 1546 18536 1551 18592
rect 0 18534 1551 18536
rect 0 18504 800 18534
rect 1485 18531 1551 18534
rect 0 18186 800 18216
rect 1853 18186 1919 18189
rect 0 18184 1919 18186
rect 0 18128 1858 18184
rect 1914 18128 1919 18184
rect 0 18126 1919 18128
rect 2730 18186 2790 18667
rect 4061 18458 4127 18461
rect 4705 18458 4771 18461
rect 4061 18456 4771 18458
rect 4061 18400 4066 18456
rect 4122 18400 4710 18456
rect 4766 18400 4771 18456
rect 4061 18398 4771 18400
rect 4061 18395 4127 18398
rect 4705 18395 4771 18398
rect 5533 18460 5599 18461
rect 5533 18456 5580 18460
rect 5644 18458 5650 18460
rect 5533 18400 5538 18456
rect 5533 18396 5580 18400
rect 5644 18398 5690 18458
rect 5644 18396 5650 18398
rect 5533 18395 5599 18396
rect 4429 18322 4495 18325
rect 5257 18322 5323 18325
rect 5809 18324 5875 18325
rect 5758 18322 5764 18324
rect 4429 18320 5323 18322
rect 4429 18264 4434 18320
rect 4490 18264 5262 18320
rect 5318 18264 5323 18320
rect 4429 18262 5323 18264
rect 5718 18262 5764 18322
rect 5828 18320 5875 18324
rect 5870 18264 5875 18320
rect 4429 18259 4495 18262
rect 5257 18259 5323 18262
rect 5758 18260 5764 18262
rect 5828 18260 5875 18264
rect 5950 18322 6010 18670
rect 6453 18728 12450 18730
rect 6453 18672 6458 18728
rect 6514 18672 12450 18728
rect 6453 18670 12450 18672
rect 6453 18667 6519 18670
rect 6913 18594 6979 18597
rect 10225 18594 10291 18597
rect 10593 18596 10659 18597
rect 6913 18592 10291 18594
rect 6913 18536 6918 18592
rect 6974 18536 10230 18592
rect 10286 18536 10291 18592
rect 6913 18534 10291 18536
rect 6913 18531 6979 18534
rect 10225 18531 10291 18534
rect 10542 18532 10548 18596
rect 10612 18594 10659 18596
rect 10612 18592 10704 18594
rect 10654 18536 10704 18592
rect 10612 18534 10704 18536
rect 10612 18532 10659 18534
rect 10593 18531 10659 18532
rect 6144 18528 6460 18529
rect 6144 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6460 18528
rect 6144 18463 6460 18464
rect 11342 18528 11658 18529
rect 11342 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11658 18528
rect 11342 18463 11658 18464
rect 6821 18458 6887 18461
rect 9765 18458 9831 18461
rect 6821 18456 9831 18458
rect 6821 18400 6826 18456
rect 6882 18400 9770 18456
rect 9826 18400 9831 18456
rect 6821 18398 9831 18400
rect 12390 18458 12450 18670
rect 15326 18668 15332 18732
rect 15396 18730 15402 18732
rect 15561 18730 15627 18733
rect 15396 18728 15627 18730
rect 15396 18672 15566 18728
rect 15622 18672 15627 18728
rect 15396 18670 15627 18672
rect 15396 18668 15402 18670
rect 15561 18667 15627 18670
rect 19287 18728 19353 18733
rect 19287 18672 19292 18728
rect 19348 18672 19353 18728
rect 19287 18667 19353 18672
rect 19425 18730 19491 18733
rect 21222 18730 21282 18806
rect 21633 18803 21699 18806
rect 19425 18728 21282 18730
rect 19425 18672 19430 18728
rect 19486 18672 21282 18728
rect 19425 18670 21282 18672
rect 21449 18730 21515 18733
rect 21449 18728 22202 18730
rect 21449 18672 21454 18728
rect 21510 18672 22202 18728
rect 21449 18670 22202 18672
rect 19425 18667 19491 18670
rect 21449 18667 21515 18670
rect 19290 18594 19350 18667
rect 22142 18624 22202 18670
rect 20805 18594 20871 18597
rect 19290 18592 20871 18594
rect 19290 18536 20810 18592
rect 20866 18536 20871 18592
rect 19290 18534 20871 18536
rect 22142 18534 23000 18624
rect 20805 18531 20871 18534
rect 16540 18528 16856 18529
rect 16540 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16856 18528
rect 16540 18463 16856 18464
rect 21738 18528 22054 18529
rect 21738 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22054 18528
rect 22200 18504 23000 18534
rect 21738 18463 22054 18464
rect 15377 18458 15443 18461
rect 19609 18460 19675 18461
rect 12390 18456 15443 18458
rect 12390 18400 15382 18456
rect 15438 18400 15443 18456
rect 12390 18398 15443 18400
rect 6821 18395 6887 18398
rect 9765 18395 9831 18398
rect 15377 18395 15443 18398
rect 19558 18396 19564 18460
rect 19628 18458 19675 18460
rect 19793 18458 19859 18461
rect 19926 18458 19932 18460
rect 19628 18456 19720 18458
rect 19670 18400 19720 18456
rect 19628 18398 19720 18400
rect 19793 18456 19932 18458
rect 19793 18400 19798 18456
rect 19854 18400 19932 18456
rect 19793 18398 19932 18400
rect 19628 18396 19675 18398
rect 19609 18395 19675 18396
rect 19793 18395 19859 18398
rect 19926 18396 19932 18398
rect 19996 18396 20002 18460
rect 11973 18322 12039 18325
rect 5950 18320 12039 18322
rect 5950 18264 11978 18320
rect 12034 18264 12039 18320
rect 5950 18262 12039 18264
rect 5809 18259 5875 18260
rect 11973 18259 12039 18262
rect 12893 18322 12959 18325
rect 19793 18322 19859 18325
rect 20621 18322 20687 18325
rect 12893 18320 20687 18322
rect 12893 18264 12898 18320
rect 12954 18264 19798 18320
rect 19854 18264 20626 18320
rect 20682 18264 20687 18320
rect 12893 18262 20687 18264
rect 12893 18259 12959 18262
rect 19793 18259 19859 18262
rect 20621 18259 20687 18262
rect 5165 18186 5231 18189
rect 2730 18184 14474 18186
rect 2730 18128 5170 18184
rect 5226 18128 14474 18184
rect 2730 18126 14474 18128
rect 0 18096 800 18126
rect 1853 18123 1919 18126
rect 5165 18123 5231 18126
rect 4102 17988 4108 18052
rect 4172 18050 4178 18052
rect 7833 18050 7899 18053
rect 8477 18050 8543 18053
rect 4172 18048 8543 18050
rect 4172 17992 7838 18048
rect 7894 17992 8482 18048
rect 8538 17992 8543 18048
rect 4172 17990 8543 17992
rect 4172 17988 4178 17990
rect 7833 17987 7899 17990
rect 8477 17987 8543 17990
rect 11881 18050 11947 18053
rect 13077 18050 13143 18053
rect 11881 18048 13143 18050
rect 11881 17992 11886 18048
rect 11942 17992 13082 18048
rect 13138 17992 13143 18048
rect 11881 17990 13143 17992
rect 14414 18050 14474 18126
rect 14958 18124 14964 18188
rect 15028 18186 15034 18188
rect 20897 18186 20963 18189
rect 15028 18184 20963 18186
rect 15028 18128 20902 18184
rect 20958 18128 20963 18184
rect 15028 18126 20963 18128
rect 15028 18124 15034 18126
rect 20897 18123 20963 18126
rect 21081 18186 21147 18189
rect 22200 18186 23000 18216
rect 21081 18184 23000 18186
rect 21081 18128 21086 18184
rect 21142 18128 23000 18184
rect 21081 18126 23000 18128
rect 21081 18123 21147 18126
rect 22200 18096 23000 18126
rect 15561 18050 15627 18053
rect 14414 18048 15627 18050
rect 14414 17992 15566 18048
rect 15622 17992 15627 18048
rect 14414 17990 15627 17992
rect 11881 17987 11947 17990
rect 13077 17987 13143 17990
rect 15561 17987 15627 17990
rect 16246 17988 16252 18052
rect 16316 18050 16322 18052
rect 17217 18050 17283 18053
rect 16316 18048 17283 18050
rect 16316 17992 17222 18048
rect 17278 17992 17283 18048
rect 16316 17990 17283 17992
rect 16316 17988 16322 17990
rect 17217 17987 17283 17990
rect 20621 18050 20687 18053
rect 21173 18050 21239 18053
rect 20621 18048 21239 18050
rect 20621 17992 20626 18048
rect 20682 17992 21178 18048
rect 21234 17992 21239 18048
rect 20621 17990 21239 17992
rect 20621 17987 20687 17990
rect 21173 17987 21239 17990
rect 3545 17984 3861 17985
rect 3545 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3861 17984
rect 3545 17919 3861 17920
rect 8743 17984 9059 17985
rect 8743 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9059 17984
rect 8743 17919 9059 17920
rect 13941 17984 14257 17985
rect 13941 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14257 17984
rect 13941 17919 14257 17920
rect 19139 17984 19455 17985
rect 19139 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19455 17984
rect 19139 17919 19455 17920
rect 5441 17914 5507 17917
rect 5901 17914 5967 17917
rect 5441 17912 5967 17914
rect 5441 17856 5446 17912
rect 5502 17856 5906 17912
rect 5962 17856 5967 17912
rect 5441 17854 5967 17856
rect 5441 17851 5507 17854
rect 5901 17851 5967 17854
rect 7598 17852 7604 17916
rect 7668 17914 7674 17916
rect 8477 17914 8543 17917
rect 13721 17914 13787 17917
rect 7668 17912 8543 17914
rect 7668 17856 8482 17912
rect 8538 17856 8543 17912
rect 7668 17854 8543 17856
rect 7668 17852 7674 17854
rect 8477 17851 8543 17854
rect 9998 17912 13787 17914
rect 9998 17856 13726 17912
rect 13782 17856 13787 17912
rect 9998 17854 13787 17856
rect 0 17778 800 17808
rect 1485 17778 1551 17781
rect 0 17776 1551 17778
rect 0 17720 1490 17776
rect 1546 17720 1551 17776
rect 0 17718 1551 17720
rect 0 17688 800 17718
rect 1485 17715 1551 17718
rect 2589 17778 2655 17781
rect 8845 17778 8911 17781
rect 2589 17776 8911 17778
rect 2589 17720 2594 17776
rect 2650 17720 8850 17776
rect 8906 17720 8911 17776
rect 2589 17718 8911 17720
rect 2589 17715 2655 17718
rect 8845 17715 8911 17718
rect 9029 17778 9095 17781
rect 9998 17780 10058 17854
rect 13721 17851 13787 17854
rect 15101 17912 15167 17917
rect 15101 17856 15106 17912
rect 15162 17856 15167 17912
rect 15101 17851 15167 17856
rect 9990 17778 9996 17780
rect 9029 17776 9996 17778
rect 9029 17720 9034 17776
rect 9090 17720 9996 17776
rect 9029 17718 9996 17720
rect 9029 17715 9095 17718
rect 9990 17716 9996 17718
rect 10060 17716 10066 17780
rect 13077 17778 13143 17781
rect 15104 17778 15164 17851
rect 13077 17776 15164 17778
rect 13077 17720 13082 17776
rect 13138 17720 15164 17776
rect 13077 17718 15164 17720
rect 15285 17778 15351 17781
rect 20294 17778 20300 17780
rect 15285 17776 20300 17778
rect 15285 17720 15290 17776
rect 15346 17720 20300 17776
rect 15285 17718 20300 17720
rect 13077 17715 13143 17718
rect 15285 17715 15351 17718
rect 20294 17716 20300 17718
rect 20364 17716 20370 17780
rect 21449 17778 21515 17781
rect 22200 17778 23000 17808
rect 21449 17776 23000 17778
rect 21449 17720 21454 17776
rect 21510 17720 23000 17776
rect 21449 17718 23000 17720
rect 21449 17715 21515 17718
rect 22200 17688 23000 17718
rect 4613 17642 4679 17645
rect 13813 17642 13879 17645
rect 4613 17640 13879 17642
rect 4613 17584 4618 17640
rect 4674 17584 13818 17640
rect 13874 17584 13879 17640
rect 4613 17582 13879 17584
rect 4613 17579 4679 17582
rect 13813 17579 13879 17582
rect 1301 17506 1367 17509
rect 5901 17506 5967 17509
rect 1301 17504 5967 17506
rect 1301 17448 1306 17504
rect 1362 17448 5906 17504
rect 5962 17448 5967 17504
rect 1301 17446 5967 17448
rect 1301 17443 1367 17446
rect 5901 17443 5967 17446
rect 6678 17444 6684 17508
rect 6748 17506 6754 17508
rect 7557 17506 7623 17509
rect 6748 17504 7623 17506
rect 6748 17448 7562 17504
rect 7618 17448 7623 17504
rect 6748 17446 7623 17448
rect 6748 17444 6754 17446
rect 7557 17443 7623 17446
rect 7741 17506 7807 17509
rect 9029 17506 9095 17509
rect 7741 17504 9095 17506
rect 7741 17448 7746 17504
rect 7802 17448 9034 17504
rect 9090 17448 9095 17504
rect 7741 17446 9095 17448
rect 7741 17443 7807 17446
rect 9029 17443 9095 17446
rect 9949 17506 10015 17509
rect 10317 17506 10383 17509
rect 10593 17506 10659 17509
rect 9949 17504 10659 17506
rect 9949 17448 9954 17504
rect 10010 17448 10322 17504
rect 10378 17448 10598 17504
rect 10654 17448 10659 17504
rect 9949 17446 10659 17448
rect 9949 17443 10015 17446
rect 10317 17443 10383 17446
rect 10593 17443 10659 17446
rect 6144 17440 6460 17441
rect 0 17370 800 17400
rect 6144 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6460 17440
rect 6144 17375 6460 17376
rect 11342 17440 11658 17441
rect 11342 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11658 17440
rect 11342 17375 11658 17376
rect 16540 17440 16856 17441
rect 16540 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16856 17440
rect 16540 17375 16856 17376
rect 21738 17440 22054 17441
rect 21738 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22054 17440
rect 21738 17375 22054 17376
rect 1853 17370 1919 17373
rect 0 17368 1919 17370
rect 0 17312 1858 17368
rect 1914 17312 1919 17368
rect 0 17310 1919 17312
rect 0 17280 800 17310
rect 1853 17307 1919 17310
rect 3918 17308 3924 17372
rect 3988 17370 3994 17372
rect 5533 17370 5599 17373
rect 3988 17368 5599 17370
rect 3988 17312 5538 17368
rect 5594 17312 5599 17368
rect 3988 17310 5599 17312
rect 3988 17308 3994 17310
rect 5533 17307 5599 17310
rect 6913 17368 6979 17373
rect 6913 17312 6918 17368
rect 6974 17312 6979 17368
rect 6913 17307 6979 17312
rect 7649 17370 7715 17373
rect 9581 17370 9647 17373
rect 10961 17370 11027 17373
rect 22200 17370 23000 17400
rect 7649 17368 11027 17370
rect 7649 17312 7654 17368
rect 7710 17312 9586 17368
rect 9642 17312 10966 17368
rect 11022 17312 11027 17368
rect 7649 17310 11027 17312
rect 7649 17307 7715 17310
rect 9581 17307 9647 17310
rect 10961 17307 11027 17310
rect 3366 17172 3372 17236
rect 3436 17234 3442 17236
rect 3785 17234 3851 17237
rect 5533 17234 5599 17237
rect 6916 17234 6976 17307
rect 22142 17280 23000 17370
rect 7741 17234 7807 17237
rect 3436 17232 5274 17234
rect 3436 17176 3790 17232
rect 3846 17176 5274 17232
rect 3436 17174 5274 17176
rect 3436 17172 3442 17174
rect 3785 17171 3851 17174
rect 2221 17098 2287 17101
rect 5073 17098 5139 17101
rect 2221 17096 5139 17098
rect 2221 17040 2226 17096
rect 2282 17040 5078 17096
rect 5134 17040 5139 17096
rect 2221 17038 5139 17040
rect 5214 17098 5274 17174
rect 5533 17232 6976 17234
rect 5533 17176 5538 17232
rect 5594 17176 6976 17232
rect 5533 17174 6976 17176
rect 7054 17232 7807 17234
rect 7054 17176 7746 17232
rect 7802 17176 7807 17232
rect 7054 17174 7807 17176
rect 5533 17171 5599 17174
rect 6637 17098 6703 17101
rect 7054 17098 7114 17174
rect 7741 17171 7807 17174
rect 8845 17234 8911 17237
rect 15193 17234 15259 17237
rect 8845 17232 15259 17234
rect 8845 17176 8850 17232
rect 8906 17176 15198 17232
rect 15254 17176 15259 17232
rect 8845 17174 15259 17176
rect 8845 17171 8911 17174
rect 15193 17171 15259 17174
rect 21541 17234 21607 17237
rect 22142 17234 22202 17280
rect 21541 17232 22202 17234
rect 21541 17176 21546 17232
rect 21602 17176 22202 17232
rect 21541 17174 22202 17176
rect 21541 17171 21607 17174
rect 5214 17096 7114 17098
rect 5214 17040 6642 17096
rect 6698 17040 7114 17096
rect 5214 17038 7114 17040
rect 7741 17098 7807 17101
rect 15326 17098 15332 17100
rect 7741 17096 15332 17098
rect 7741 17040 7746 17096
rect 7802 17040 15332 17096
rect 7741 17038 15332 17040
rect 2221 17035 2287 17038
rect 5073 17035 5139 17038
rect 6637 17035 6703 17038
rect 7741 17035 7807 17038
rect 15326 17036 15332 17038
rect 15396 17036 15402 17100
rect 0 16962 800 16992
rect 1485 16962 1551 16965
rect 0 16960 1551 16962
rect 0 16904 1490 16960
rect 1546 16904 1551 16960
rect 0 16902 1551 16904
rect 0 16872 800 16902
rect 1485 16899 1551 16902
rect 4061 16962 4127 16965
rect 5809 16962 5875 16965
rect 8201 16962 8267 16965
rect 13721 16964 13787 16965
rect 13670 16962 13676 16964
rect 4061 16960 8267 16962
rect 4061 16904 4066 16960
rect 4122 16904 5814 16960
rect 5870 16904 8206 16960
rect 8262 16904 8267 16960
rect 4061 16902 8267 16904
rect 4061 16899 4127 16902
rect 5809 16899 5875 16902
rect 8201 16899 8267 16902
rect 9262 16902 13676 16962
rect 13740 16960 13787 16964
rect 13782 16904 13787 16960
rect 3545 16896 3861 16897
rect 3545 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3861 16896
rect 3545 16831 3861 16832
rect 8743 16896 9059 16897
rect 8743 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9059 16896
rect 8743 16831 9059 16832
rect 4797 16826 4863 16829
rect 4797 16824 8402 16826
rect 4797 16768 4802 16824
rect 4858 16768 8402 16824
rect 4797 16766 8402 16768
rect 4797 16763 4863 16766
rect 2037 16690 2103 16693
rect 2681 16690 2747 16693
rect 4337 16690 4403 16693
rect 2037 16688 2747 16690
rect 2037 16632 2042 16688
rect 2098 16632 2686 16688
rect 2742 16632 2747 16688
rect 2037 16630 2747 16632
rect 2037 16627 2103 16630
rect 2681 16627 2747 16630
rect 4294 16688 4403 16690
rect 4294 16632 4342 16688
rect 4398 16632 4403 16688
rect 4294 16627 4403 16632
rect 4521 16690 4587 16693
rect 7005 16690 7071 16693
rect 7649 16690 7715 16693
rect 7925 16692 7991 16693
rect 7925 16690 7972 16692
rect 4521 16688 7715 16690
rect 4521 16632 4526 16688
rect 4582 16632 7010 16688
rect 7066 16632 7654 16688
rect 7710 16632 7715 16688
rect 4521 16630 7715 16632
rect 7880 16688 7972 16690
rect 7880 16632 7930 16688
rect 7880 16630 7972 16632
rect 4521 16627 4587 16630
rect 7005 16627 7071 16630
rect 7649 16627 7715 16630
rect 7925 16628 7972 16630
rect 8036 16628 8042 16692
rect 7925 16627 7991 16628
rect 0 16554 800 16584
rect 1853 16554 1919 16557
rect 0 16552 1919 16554
rect 0 16496 1858 16552
rect 1914 16496 1919 16552
rect 0 16494 1919 16496
rect 4294 16554 4354 16627
rect 8342 16557 8402 16766
rect 8518 16628 8524 16692
rect 8588 16690 8594 16692
rect 8753 16690 8819 16693
rect 8588 16688 8819 16690
rect 8588 16632 8758 16688
rect 8814 16632 8819 16688
rect 8588 16630 8819 16632
rect 8588 16628 8594 16630
rect 8753 16627 8819 16630
rect 9121 16690 9187 16693
rect 9262 16690 9322 16902
rect 13670 16900 13676 16902
rect 13740 16900 13787 16904
rect 13721 16899 13787 16900
rect 21449 16962 21515 16965
rect 22200 16962 23000 16992
rect 21449 16960 23000 16962
rect 21449 16904 21454 16960
rect 21510 16904 23000 16960
rect 21449 16902 23000 16904
rect 21449 16899 21515 16902
rect 13941 16896 14257 16897
rect 13941 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14257 16896
rect 13941 16831 14257 16832
rect 19139 16896 19455 16897
rect 19139 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19455 16896
rect 22200 16872 23000 16902
rect 19139 16831 19455 16832
rect 12249 16826 12315 16829
rect 12249 16824 12634 16826
rect 12249 16768 12254 16824
rect 12310 16768 12634 16824
rect 12249 16766 12634 16768
rect 12249 16763 12315 16766
rect 9121 16688 9322 16690
rect 9121 16632 9126 16688
rect 9182 16632 9322 16688
rect 9121 16630 9322 16632
rect 9121 16627 9187 16630
rect 10910 16628 10916 16692
rect 10980 16690 10986 16692
rect 12433 16690 12499 16693
rect 10980 16688 12499 16690
rect 10980 16632 12438 16688
rect 12494 16632 12499 16688
rect 10980 16630 12499 16632
rect 10980 16628 10986 16630
rect 12433 16627 12499 16630
rect 4294 16494 6746 16554
rect 0 16464 800 16494
rect 1853 16491 1919 16494
rect 6144 16352 6460 16353
rect 6144 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6460 16352
rect 6144 16287 6460 16288
rect 933 16282 999 16285
rect 4337 16282 4403 16285
rect 933 16280 4403 16282
rect 933 16224 938 16280
rect 994 16224 4342 16280
rect 4398 16224 4403 16280
rect 933 16222 4403 16224
rect 6686 16282 6746 16494
rect 6913 16552 6979 16557
rect 6913 16496 6918 16552
rect 6974 16496 6979 16552
rect 6913 16491 6979 16496
rect 7741 16554 7807 16557
rect 8150 16554 8156 16556
rect 7741 16552 8156 16554
rect 7741 16496 7746 16552
rect 7802 16496 8156 16552
rect 7741 16494 8156 16496
rect 7741 16491 7807 16494
rect 8150 16492 8156 16494
rect 8220 16492 8226 16556
rect 8342 16552 8451 16557
rect 12433 16554 12499 16557
rect 8342 16496 8390 16552
rect 8446 16496 8451 16552
rect 8342 16494 8451 16496
rect 8385 16491 8451 16494
rect 8710 16552 12499 16554
rect 8710 16496 12438 16552
rect 12494 16496 12499 16552
rect 8710 16494 12499 16496
rect 6916 16418 6976 16491
rect 8518 16418 8524 16420
rect 6916 16358 8524 16418
rect 8518 16356 8524 16358
rect 8588 16356 8594 16420
rect 8710 16282 8770 16494
rect 12433 16491 12499 16494
rect 11789 16418 11855 16421
rect 12341 16418 12407 16421
rect 12574 16418 12634 16766
rect 12709 16690 12775 16693
rect 13169 16690 13235 16693
rect 15694 16690 15700 16692
rect 12709 16688 15700 16690
rect 12709 16632 12714 16688
rect 12770 16632 13174 16688
rect 13230 16632 15700 16688
rect 12709 16630 15700 16632
rect 12709 16627 12775 16630
rect 13169 16627 13235 16630
rect 15694 16628 15700 16630
rect 15764 16628 15770 16692
rect 16205 16690 16271 16693
rect 17769 16690 17835 16693
rect 16205 16688 17835 16690
rect 16205 16632 16210 16688
rect 16266 16632 17774 16688
rect 17830 16632 17835 16688
rect 16205 16630 17835 16632
rect 16205 16627 16271 16630
rect 17769 16627 17835 16630
rect 21081 16554 21147 16557
rect 22200 16554 23000 16584
rect 21081 16552 23000 16554
rect 21081 16496 21086 16552
rect 21142 16496 23000 16552
rect 21081 16494 23000 16496
rect 21081 16491 21147 16494
rect 22200 16464 23000 16494
rect 11789 16416 11898 16418
rect 11789 16360 11794 16416
rect 11850 16360 11898 16416
rect 11789 16355 11898 16360
rect 12341 16416 12634 16418
rect 12341 16360 12346 16416
rect 12402 16360 12634 16416
rect 12341 16358 12634 16360
rect 12341 16355 12407 16358
rect 11342 16352 11658 16353
rect 11342 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11658 16352
rect 11342 16287 11658 16288
rect 6686 16222 8770 16282
rect 9673 16282 9739 16285
rect 9806 16282 9812 16284
rect 9673 16280 9812 16282
rect 9673 16224 9678 16280
rect 9734 16224 9812 16280
rect 9673 16222 9812 16224
rect 933 16219 999 16222
rect 4337 16219 4403 16222
rect 9673 16219 9739 16222
rect 9806 16220 9812 16222
rect 9876 16220 9882 16284
rect 10501 16282 10567 16285
rect 10777 16282 10843 16285
rect 10501 16280 10843 16282
rect 10501 16224 10506 16280
rect 10562 16224 10782 16280
rect 10838 16224 10843 16280
rect 10501 16222 10843 16224
rect 10501 16219 10567 16222
rect 10777 16219 10843 16222
rect 0 16146 800 16176
rect 11838 16149 11898 16355
rect 16540 16352 16856 16353
rect 16540 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16856 16352
rect 16540 16287 16856 16288
rect 21738 16352 22054 16353
rect 21738 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22054 16352
rect 21738 16287 22054 16288
rect 12065 16282 12131 16285
rect 16113 16282 16179 16285
rect 12065 16280 16179 16282
rect 12065 16224 12070 16280
rect 12126 16224 16118 16280
rect 16174 16224 16179 16280
rect 12065 16222 16179 16224
rect 12065 16219 12131 16222
rect 16113 16219 16179 16222
rect 1577 16146 1643 16149
rect 0 16144 1643 16146
rect 0 16088 1582 16144
rect 1638 16088 1643 16144
rect 0 16086 1643 16088
rect 0 16056 800 16086
rect 1577 16083 1643 16086
rect 2589 16146 2655 16149
rect 6637 16146 6703 16149
rect 7465 16146 7531 16149
rect 10174 16146 10180 16148
rect 2589 16144 10180 16146
rect 2589 16088 2594 16144
rect 2650 16088 6642 16144
rect 6698 16088 7470 16144
rect 7526 16088 10180 16144
rect 2589 16086 10180 16088
rect 2589 16083 2655 16086
rect 6637 16083 6703 16086
rect 7465 16083 7531 16086
rect 10174 16084 10180 16086
rect 10244 16146 10250 16148
rect 11605 16146 11671 16149
rect 10244 16144 11671 16146
rect 10244 16088 11610 16144
rect 11666 16088 11671 16144
rect 10244 16086 11671 16088
rect 11838 16144 11947 16149
rect 11838 16088 11886 16144
rect 11942 16088 11947 16144
rect 11838 16086 11947 16088
rect 10244 16084 10250 16086
rect 11605 16083 11671 16086
rect 11881 16083 11947 16086
rect 12249 16146 12315 16149
rect 12617 16146 12683 16149
rect 12249 16144 12683 16146
rect 12249 16088 12254 16144
rect 12310 16088 12622 16144
rect 12678 16088 12683 16144
rect 12249 16086 12683 16088
rect 12249 16083 12315 16086
rect 12617 16083 12683 16086
rect 19701 16146 19767 16149
rect 20529 16146 20595 16149
rect 19701 16144 20595 16146
rect 19701 16088 19706 16144
rect 19762 16088 20534 16144
rect 20590 16088 20595 16144
rect 19701 16086 20595 16088
rect 19701 16083 19767 16086
rect 20529 16083 20595 16086
rect 21449 16146 21515 16149
rect 22200 16146 23000 16176
rect 21449 16144 23000 16146
rect 21449 16088 21454 16144
rect 21510 16088 23000 16144
rect 21449 16086 23000 16088
rect 21449 16083 21515 16086
rect 22200 16056 23000 16086
rect 1945 16010 2011 16013
rect 3417 16010 3483 16013
rect 1945 16008 3483 16010
rect 1945 15952 1950 16008
rect 2006 15952 3422 16008
rect 3478 15952 3483 16008
rect 1945 15950 3483 15952
rect 1945 15947 2011 15950
rect 3417 15947 3483 15950
rect 5165 16010 5231 16013
rect 11329 16010 11395 16013
rect 5165 16008 11395 16010
rect 5165 15952 5170 16008
rect 5226 15952 11334 16008
rect 11390 15952 11395 16008
rect 5165 15950 11395 15952
rect 5165 15947 5231 15950
rect 11329 15947 11395 15950
rect 11513 16010 11579 16013
rect 16246 16010 16252 16012
rect 11513 16008 16252 16010
rect 11513 15952 11518 16008
rect 11574 15952 16252 16008
rect 11513 15950 16252 15952
rect 11513 15947 11579 15950
rect 16246 15948 16252 15950
rect 16316 15948 16322 16012
rect 19609 16010 19675 16013
rect 17910 16008 19675 16010
rect 17910 15952 19614 16008
rect 19670 15952 19675 16008
rect 17910 15950 19675 15952
rect 9305 15874 9371 15877
rect 12249 15874 12315 15877
rect 9305 15872 12315 15874
rect 9305 15816 9310 15872
rect 9366 15816 12254 15872
rect 12310 15816 12315 15872
rect 9305 15814 12315 15816
rect 9305 15811 9371 15814
rect 12249 15811 12315 15814
rect 3545 15808 3861 15809
rect 0 15738 800 15768
rect 3545 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3861 15808
rect 3545 15743 3861 15744
rect 8743 15808 9059 15809
rect 8743 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9059 15808
rect 8743 15743 9059 15744
rect 13941 15808 14257 15809
rect 13941 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14257 15808
rect 13941 15743 14257 15744
rect 1485 15738 1551 15741
rect 12433 15738 12499 15741
rect 0 15736 1551 15738
rect 0 15680 1490 15736
rect 1546 15680 1551 15736
rect 0 15678 1551 15680
rect 0 15648 800 15678
rect 1485 15675 1551 15678
rect 9262 15736 12499 15738
rect 9262 15680 12438 15736
rect 12494 15680 12499 15736
rect 9262 15678 12499 15680
rect 2313 15602 2379 15605
rect 4061 15602 4127 15605
rect 2313 15600 4127 15602
rect 2313 15544 2318 15600
rect 2374 15544 4066 15600
rect 4122 15544 4127 15600
rect 2313 15542 4127 15544
rect 2313 15539 2379 15542
rect 4061 15539 4127 15542
rect 4337 15602 4403 15605
rect 5257 15602 5323 15605
rect 4337 15600 5323 15602
rect 4337 15544 4342 15600
rect 4398 15544 5262 15600
rect 5318 15544 5323 15600
rect 4337 15542 5323 15544
rect 4337 15539 4403 15542
rect 5257 15539 5323 15542
rect 5441 15602 5507 15605
rect 7649 15602 7715 15605
rect 5441 15600 7715 15602
rect 5441 15544 5446 15600
rect 5502 15544 7654 15600
rect 7710 15544 7715 15600
rect 5441 15542 7715 15544
rect 5441 15539 5507 15542
rect 7649 15539 7715 15542
rect 7833 15602 7899 15605
rect 9262 15602 9322 15678
rect 12433 15675 12499 15678
rect 7833 15600 9322 15602
rect 7833 15544 7838 15600
rect 7894 15544 9322 15600
rect 7833 15542 9322 15544
rect 7833 15539 7899 15542
rect 10726 15540 10732 15604
rect 10796 15602 10802 15604
rect 17585 15602 17651 15605
rect 10796 15600 17651 15602
rect 10796 15544 17590 15600
rect 17646 15544 17651 15600
rect 10796 15542 17651 15544
rect 10796 15540 10802 15542
rect 17585 15539 17651 15542
rect 3785 15466 3851 15469
rect 4245 15466 4311 15469
rect 3785 15464 4311 15466
rect 3785 15408 3790 15464
rect 3846 15408 4250 15464
rect 4306 15408 4311 15464
rect 3785 15406 4311 15408
rect 3785 15403 3851 15406
rect 4245 15403 4311 15406
rect 8150 15404 8156 15468
rect 8220 15466 8226 15468
rect 8661 15466 8727 15469
rect 8220 15464 8727 15466
rect 8220 15408 8666 15464
rect 8722 15408 8727 15464
rect 8220 15406 8727 15408
rect 8220 15404 8226 15406
rect 8661 15403 8727 15406
rect 10593 15466 10659 15469
rect 17033 15466 17099 15469
rect 17910 15466 17970 15950
rect 19609 15947 19675 15950
rect 19139 15808 19455 15809
rect 19139 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19455 15808
rect 19139 15743 19455 15744
rect 21449 15738 21515 15741
rect 22200 15738 23000 15768
rect 21449 15736 23000 15738
rect 21449 15680 21454 15736
rect 21510 15680 23000 15736
rect 21449 15678 23000 15680
rect 21449 15675 21515 15678
rect 22200 15648 23000 15678
rect 18137 15602 18203 15605
rect 21633 15602 21699 15605
rect 18137 15600 21699 15602
rect 18137 15544 18142 15600
rect 18198 15544 21638 15600
rect 21694 15544 21699 15600
rect 18137 15542 21699 15544
rect 18137 15539 18203 15542
rect 21633 15539 21699 15542
rect 10593 15464 17970 15466
rect 10593 15408 10598 15464
rect 10654 15408 17038 15464
rect 17094 15408 17970 15464
rect 10593 15406 17970 15408
rect 18321 15466 18387 15469
rect 21449 15466 21515 15469
rect 18321 15464 21282 15466
rect 18321 15408 18326 15464
rect 18382 15408 21282 15464
rect 18321 15406 21282 15408
rect 10593 15403 10659 15406
rect 17033 15403 17099 15406
rect 18321 15403 18387 15406
rect 0 15330 800 15360
rect 1485 15330 1551 15333
rect 5901 15332 5967 15333
rect 5901 15330 5948 15332
rect 0 15328 1551 15330
rect 0 15272 1490 15328
rect 1546 15272 1551 15328
rect 0 15270 1551 15272
rect 5856 15328 5948 15330
rect 5856 15272 5906 15328
rect 5856 15270 5948 15272
rect 0 15240 800 15270
rect 1485 15267 1551 15270
rect 5901 15268 5948 15270
rect 6012 15268 6018 15332
rect 6637 15330 6703 15333
rect 7649 15330 7715 15333
rect 8385 15330 8451 15333
rect 6637 15328 6930 15330
rect 6637 15272 6642 15328
rect 6698 15272 6930 15328
rect 6637 15270 6930 15272
rect 5901 15267 5967 15268
rect 6637 15267 6703 15270
rect 6144 15264 6460 15265
rect 6144 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6460 15264
rect 6144 15199 6460 15200
rect 6870 15194 6930 15270
rect 7649 15328 8451 15330
rect 7649 15272 7654 15328
rect 7710 15272 8390 15328
rect 8446 15272 8451 15328
rect 7649 15270 8451 15272
rect 7649 15267 7715 15270
rect 8385 15267 8451 15270
rect 8569 15330 8635 15333
rect 9438 15330 9444 15332
rect 8569 15328 9444 15330
rect 8569 15272 8574 15328
rect 8630 15272 9444 15328
rect 8569 15270 9444 15272
rect 8569 15267 8635 15270
rect 9438 15268 9444 15270
rect 9508 15268 9514 15332
rect 11973 15330 12039 15333
rect 19057 15330 19123 15333
rect 19926 15330 19932 15332
rect 11973 15328 12266 15330
rect 11973 15272 11978 15328
rect 12034 15272 12266 15328
rect 11973 15270 12266 15272
rect 11973 15267 12039 15270
rect 11342 15264 11658 15265
rect 11342 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11658 15264
rect 11342 15199 11658 15200
rect 10041 15194 10107 15197
rect 10542 15194 10548 15196
rect 6870 15192 10548 15194
rect 6870 15136 10046 15192
rect 10102 15136 10548 15192
rect 6870 15134 10548 15136
rect 10041 15131 10107 15134
rect 10542 15132 10548 15134
rect 10612 15132 10618 15196
rect 12206 15194 12266 15270
rect 19057 15328 19932 15330
rect 19057 15272 19062 15328
rect 19118 15272 19932 15328
rect 19057 15270 19932 15272
rect 19057 15267 19123 15270
rect 19926 15268 19932 15270
rect 19996 15268 20002 15332
rect 21222 15330 21282 15406
rect 21449 15464 22202 15466
rect 21449 15408 21454 15464
rect 21510 15408 22202 15464
rect 21449 15406 22202 15408
rect 21449 15403 21515 15406
rect 22142 15360 22202 15406
rect 21541 15330 21607 15333
rect 21222 15328 21607 15330
rect 21222 15272 21546 15328
rect 21602 15272 21607 15328
rect 21222 15270 21607 15272
rect 22142 15270 23000 15360
rect 21541 15267 21607 15270
rect 16540 15264 16856 15265
rect 16540 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16856 15264
rect 16540 15199 16856 15200
rect 21738 15264 22054 15265
rect 21738 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22054 15264
rect 22200 15240 23000 15270
rect 21738 15199 22054 15200
rect 12566 15194 12572 15196
rect 12206 15134 12572 15194
rect 12566 15132 12572 15134
rect 12636 15132 12642 15196
rect 12893 15194 12959 15197
rect 14181 15194 14247 15197
rect 12893 15192 14247 15194
rect 12893 15136 12898 15192
rect 12954 15136 14186 15192
rect 14242 15136 14247 15192
rect 12893 15134 14247 15136
rect 12893 15131 12959 15134
rect 14181 15131 14247 15134
rect 3233 15058 3299 15061
rect 9121 15058 9187 15061
rect 15510 15058 15516 15060
rect 3233 15056 15516 15058
rect 3233 15000 3238 15056
rect 3294 15000 9126 15056
rect 9182 15000 15516 15056
rect 3233 14998 15516 15000
rect 3233 14995 3299 14998
rect 9121 14995 9187 14998
rect 15510 14996 15516 14998
rect 15580 15058 15586 15060
rect 18045 15058 18111 15061
rect 15580 15056 18111 15058
rect 15580 15000 18050 15056
rect 18106 15000 18111 15056
rect 15580 14998 18111 15000
rect 15580 14996 15586 14998
rect 18045 14995 18111 14998
rect 0 14922 800 14952
rect 1853 14922 1919 14925
rect 0 14920 1919 14922
rect 0 14864 1858 14920
rect 1914 14864 1919 14920
rect 0 14862 1919 14864
rect 0 14832 800 14862
rect 1853 14859 1919 14862
rect 3918 14860 3924 14924
rect 3988 14860 3994 14924
rect 6085 14922 6151 14925
rect 10777 14922 10843 14925
rect 10910 14922 10916 14924
rect 6085 14920 10916 14922
rect 6085 14864 6090 14920
rect 6146 14864 10782 14920
rect 10838 14864 10916 14920
rect 6085 14862 10916 14864
rect 3926 14786 3986 14860
rect 6085 14859 6151 14862
rect 10777 14859 10843 14862
rect 10910 14860 10916 14862
rect 10980 14860 10986 14924
rect 12065 14922 12131 14925
rect 12341 14922 12407 14925
rect 12065 14920 12407 14922
rect 12065 14864 12070 14920
rect 12126 14864 12346 14920
rect 12402 14864 12407 14920
rect 12065 14862 12407 14864
rect 12065 14859 12131 14862
rect 12341 14859 12407 14862
rect 12525 14922 12591 14925
rect 12893 14922 12959 14925
rect 13169 14924 13235 14925
rect 13118 14922 13124 14924
rect 12525 14920 12959 14922
rect 12525 14864 12530 14920
rect 12586 14864 12898 14920
rect 12954 14864 12959 14920
rect 12525 14862 12959 14864
rect 13078 14862 13124 14922
rect 13188 14920 13235 14924
rect 19057 14922 19123 14925
rect 13230 14864 13235 14920
rect 12525 14859 12591 14862
rect 12893 14859 12959 14862
rect 13118 14860 13124 14862
rect 13188 14860 13235 14864
rect 13169 14859 13235 14860
rect 13816 14920 19123 14922
rect 13816 14864 19062 14920
rect 19118 14864 19123 14920
rect 13816 14862 19123 14864
rect 8385 14786 8451 14789
rect 10593 14788 10659 14789
rect 3926 14784 8451 14786
rect 3926 14728 8390 14784
rect 8446 14728 8451 14784
rect 3926 14726 8451 14728
rect 8385 14723 8451 14726
rect 10542 14724 10548 14788
rect 10612 14786 10659 14788
rect 12896 14786 12956 14859
rect 13816 14786 13876 14862
rect 19057 14859 19123 14862
rect 21081 14922 21147 14925
rect 22200 14922 23000 14952
rect 21081 14920 23000 14922
rect 21081 14864 21086 14920
rect 21142 14864 23000 14920
rect 21081 14862 23000 14864
rect 21081 14859 21147 14862
rect 22200 14832 23000 14862
rect 10612 14784 10704 14786
rect 10654 14728 10704 14784
rect 10612 14726 10704 14728
rect 12896 14726 13876 14786
rect 20069 14788 20135 14789
rect 20069 14784 20116 14788
rect 20180 14786 20186 14788
rect 20069 14728 20074 14784
rect 10612 14724 10659 14726
rect 10593 14723 10659 14724
rect 20069 14724 20116 14728
rect 20180 14726 20226 14786
rect 20180 14724 20186 14726
rect 20069 14723 20135 14724
rect 3545 14720 3861 14721
rect 3545 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3861 14720
rect 3545 14655 3861 14656
rect 8743 14720 9059 14721
rect 8743 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9059 14720
rect 8743 14655 9059 14656
rect 13941 14720 14257 14721
rect 13941 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14257 14720
rect 13941 14655 14257 14656
rect 19139 14720 19455 14721
rect 19139 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19455 14720
rect 19139 14655 19455 14656
rect 4245 14650 4311 14653
rect 8477 14650 8543 14653
rect 4245 14648 8543 14650
rect 4245 14592 4250 14648
rect 4306 14592 8482 14648
rect 8538 14592 8543 14648
rect 4245 14590 8543 14592
rect 4245 14587 4311 14590
rect 8477 14587 8543 14590
rect 11094 14588 11100 14652
rect 11164 14650 11170 14652
rect 11830 14650 11836 14652
rect 11164 14590 11836 14650
rect 11164 14588 11170 14590
rect 11830 14588 11836 14590
rect 11900 14588 11906 14652
rect 12014 14588 12020 14652
rect 12084 14650 12090 14652
rect 13721 14650 13787 14653
rect 12084 14648 13787 14650
rect 12084 14592 13726 14648
rect 13782 14592 13787 14648
rect 12084 14590 13787 14592
rect 12084 14588 12090 14590
rect 13721 14587 13787 14590
rect 0 14514 800 14544
rect 1485 14514 1551 14517
rect 11053 14514 11119 14517
rect 0 14512 1551 14514
rect 0 14456 1490 14512
rect 1546 14456 1551 14512
rect 0 14454 1551 14456
rect 0 14424 800 14454
rect 1485 14451 1551 14454
rect 1718 14512 11119 14514
rect 1718 14456 11058 14512
rect 11114 14456 11119 14512
rect 1718 14454 11119 14456
rect 1158 14316 1164 14380
rect 1228 14378 1234 14380
rect 1718 14378 1778 14454
rect 11053 14451 11119 14454
rect 13997 14514 14063 14517
rect 14406 14514 14412 14516
rect 13997 14512 14412 14514
rect 13997 14456 14002 14512
rect 14058 14456 14412 14512
rect 13997 14454 14412 14456
rect 13997 14451 14063 14454
rect 14406 14452 14412 14454
rect 14476 14452 14482 14516
rect 21449 14514 21515 14517
rect 22200 14514 23000 14544
rect 21449 14512 23000 14514
rect 21449 14456 21454 14512
rect 21510 14456 23000 14512
rect 21449 14454 23000 14456
rect 21449 14451 21515 14454
rect 22200 14424 23000 14454
rect 10317 14378 10383 14381
rect 15469 14378 15535 14381
rect 1228 14318 1778 14378
rect 2730 14376 10383 14378
rect 2730 14320 10322 14376
rect 10378 14320 10383 14376
rect 2730 14318 10383 14320
rect 1228 14316 1234 14318
rect 933 14242 999 14245
rect 2730 14242 2790 14318
rect 10317 14315 10383 14318
rect 10550 14376 15535 14378
rect 10550 14320 15474 14376
rect 15530 14320 15535 14376
rect 10550 14318 15535 14320
rect 933 14240 2790 14242
rect 933 14184 938 14240
rect 994 14184 2790 14240
rect 933 14182 2790 14184
rect 933 14179 999 14182
rect 8334 14180 8340 14244
rect 8404 14242 8410 14244
rect 8753 14242 8819 14245
rect 9254 14242 9260 14244
rect 8404 14240 9260 14242
rect 8404 14184 8758 14240
rect 8814 14184 9260 14240
rect 8404 14182 9260 14184
rect 8404 14180 8410 14182
rect 8753 14179 8819 14182
rect 9254 14180 9260 14182
rect 9324 14242 9330 14244
rect 9489 14242 9555 14245
rect 10550 14242 10610 14318
rect 15469 14315 15535 14318
rect 9324 14240 10610 14242
rect 9324 14184 9494 14240
rect 9550 14184 10610 14240
rect 9324 14182 10610 14184
rect 9324 14180 9330 14182
rect 9489 14179 9555 14182
rect 11830 14180 11836 14244
rect 11900 14242 11906 14244
rect 15101 14242 15167 14245
rect 11900 14240 15167 14242
rect 11900 14184 15106 14240
rect 15162 14184 15167 14240
rect 11900 14182 15167 14184
rect 11900 14180 11906 14182
rect 15101 14179 15167 14182
rect 6144 14176 6460 14177
rect 0 14106 800 14136
rect 6144 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6460 14176
rect 6144 14111 6460 14112
rect 11342 14176 11658 14177
rect 11342 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11658 14176
rect 11342 14111 11658 14112
rect 16540 14176 16856 14177
rect 16540 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16856 14176
rect 16540 14111 16856 14112
rect 21738 14176 22054 14177
rect 21738 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22054 14176
rect 21738 14111 22054 14112
rect 1485 14106 1551 14109
rect 5625 14108 5691 14109
rect 0 14104 1551 14106
rect 0 14048 1490 14104
rect 1546 14048 1551 14104
rect 0 14046 1551 14048
rect 0 14016 800 14046
rect 1485 14043 1551 14046
rect 5574 14044 5580 14108
rect 5644 14106 5691 14108
rect 6821 14106 6887 14109
rect 10225 14106 10291 14109
rect 5644 14104 5736 14106
rect 5686 14048 5736 14104
rect 5644 14046 5736 14048
rect 6821 14104 10291 14106
rect 6821 14048 6826 14104
rect 6882 14048 10230 14104
rect 10286 14048 10291 14104
rect 6821 14046 10291 14048
rect 5644 14044 5691 14046
rect 5625 14043 5691 14044
rect 6821 14043 6887 14046
rect 10225 14043 10291 14046
rect 10358 14044 10364 14108
rect 10428 14106 10434 14108
rect 10501 14106 10567 14109
rect 10961 14106 11027 14109
rect 22200 14106 23000 14136
rect 10428 14104 11027 14106
rect 10428 14048 10506 14104
rect 10562 14048 10966 14104
rect 11022 14048 11027 14104
rect 10428 14046 11027 14048
rect 10428 14044 10434 14046
rect 10501 14043 10567 14046
rect 10961 14043 11027 14046
rect 22142 14016 23000 14106
rect 933 13970 999 13973
rect 10133 13970 10199 13973
rect 933 13968 10199 13970
rect 933 13912 938 13968
rect 994 13912 10138 13968
rect 10194 13912 10199 13968
rect 933 13910 10199 13912
rect 933 13907 999 13910
rect 10133 13907 10199 13910
rect 10593 13970 10659 13973
rect 14273 13970 14339 13973
rect 10593 13968 14339 13970
rect 10593 13912 10598 13968
rect 10654 13912 14278 13968
rect 14334 13912 14339 13968
rect 10593 13910 14339 13912
rect 10593 13907 10659 13910
rect 14273 13907 14339 13910
rect 21449 13970 21515 13973
rect 22142 13970 22202 14016
rect 21449 13968 22202 13970
rect 21449 13912 21454 13968
rect 21510 13912 22202 13968
rect 21449 13910 22202 13912
rect 21449 13907 21515 13910
rect 2262 13772 2268 13836
rect 2332 13834 2338 13836
rect 2405 13834 2471 13837
rect 4337 13834 4403 13837
rect 2332 13832 4403 13834
rect 2332 13776 2410 13832
rect 2466 13776 4342 13832
rect 4398 13776 4403 13832
rect 2332 13774 4403 13776
rect 2332 13772 2338 13774
rect 2405 13771 2471 13774
rect 4337 13771 4403 13774
rect 5022 13772 5028 13836
rect 5092 13834 5098 13836
rect 10593 13834 10659 13837
rect 5092 13832 10659 13834
rect 5092 13776 10598 13832
rect 10654 13776 10659 13832
rect 5092 13774 10659 13776
rect 5092 13772 5098 13774
rect 10593 13771 10659 13774
rect 11094 13772 11100 13836
rect 11164 13834 11170 13836
rect 11513 13834 11579 13837
rect 13445 13836 13511 13837
rect 11830 13834 11836 13836
rect 11164 13832 11579 13834
rect 11164 13776 11518 13832
rect 11574 13776 11579 13832
rect 11164 13774 11579 13776
rect 11164 13772 11170 13774
rect 11513 13771 11579 13774
rect 11654 13774 11836 13834
rect 0 13698 800 13728
rect 1485 13698 1551 13701
rect 0 13696 1551 13698
rect 0 13640 1490 13696
rect 1546 13640 1551 13696
rect 0 13638 1551 13640
rect 0 13608 800 13638
rect 1485 13635 1551 13638
rect 2630 13636 2636 13700
rect 2700 13698 2706 13700
rect 3325 13698 3391 13701
rect 2700 13696 3391 13698
rect 2700 13640 3330 13696
rect 3386 13640 3391 13696
rect 2700 13638 3391 13640
rect 2700 13636 2706 13638
rect 3325 13635 3391 13638
rect 4470 13636 4476 13700
rect 4540 13698 4546 13700
rect 6821 13698 6887 13701
rect 4540 13696 6887 13698
rect 4540 13640 6826 13696
rect 6882 13640 6887 13696
rect 4540 13638 6887 13640
rect 4540 13636 4546 13638
rect 6821 13635 6887 13638
rect 9949 13698 10015 13701
rect 10133 13698 10199 13701
rect 9949 13696 10199 13698
rect 9949 13640 9954 13696
rect 10010 13640 10138 13696
rect 10194 13640 10199 13696
rect 9949 13638 10199 13640
rect 9949 13635 10015 13638
rect 10133 13635 10199 13638
rect 11421 13698 11487 13701
rect 11654 13698 11714 13774
rect 11830 13772 11836 13774
rect 11900 13772 11906 13836
rect 13445 13832 13492 13836
rect 13556 13834 13562 13836
rect 13721 13834 13787 13837
rect 22001 13834 22067 13837
rect 13445 13776 13450 13832
rect 13445 13772 13492 13776
rect 13556 13774 13602 13834
rect 13721 13832 22067 13834
rect 13721 13776 13726 13832
rect 13782 13776 22006 13832
rect 22062 13776 22067 13832
rect 13721 13774 22067 13776
rect 13556 13772 13562 13774
rect 13445 13771 13511 13772
rect 13721 13771 13787 13774
rect 22001 13771 22067 13774
rect 11421 13696 11714 13698
rect 11421 13640 11426 13696
rect 11482 13640 11714 13696
rect 11421 13638 11714 13640
rect 11421 13635 11487 13638
rect 12934 13636 12940 13700
rect 13004 13698 13010 13700
rect 13537 13698 13603 13701
rect 13004 13696 13603 13698
rect 13004 13640 13542 13696
rect 13598 13640 13603 13696
rect 13004 13638 13603 13640
rect 13004 13636 13010 13638
rect 13537 13635 13603 13638
rect 21449 13698 21515 13701
rect 22200 13698 23000 13728
rect 21449 13696 23000 13698
rect 21449 13640 21454 13696
rect 21510 13640 23000 13696
rect 21449 13638 23000 13640
rect 21449 13635 21515 13638
rect 3545 13632 3861 13633
rect 3545 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3861 13632
rect 3545 13567 3861 13568
rect 8743 13632 9059 13633
rect 8743 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9059 13632
rect 8743 13567 9059 13568
rect 13941 13632 14257 13633
rect 13941 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14257 13632
rect 13941 13567 14257 13568
rect 19139 13632 19455 13633
rect 19139 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19455 13632
rect 22200 13608 23000 13638
rect 19139 13567 19455 13568
rect 5574 13500 5580 13564
rect 5644 13562 5650 13564
rect 8569 13562 8635 13565
rect 5644 13560 8635 13562
rect 5644 13504 8574 13560
rect 8630 13504 8635 13560
rect 5644 13502 8635 13504
rect 5644 13500 5650 13502
rect 8569 13499 8635 13502
rect 9765 13562 9831 13565
rect 10225 13562 10291 13565
rect 10777 13564 10843 13565
rect 9765 13560 10291 13562
rect 9765 13504 9770 13560
rect 9826 13504 10230 13560
rect 10286 13504 10291 13560
rect 9765 13502 10291 13504
rect 9765 13499 9831 13502
rect 10225 13499 10291 13502
rect 10726 13500 10732 13564
rect 10796 13562 10843 13564
rect 11973 13562 12039 13565
rect 12750 13562 12756 13564
rect 10796 13560 10888 13562
rect 10838 13504 10888 13560
rect 10796 13502 10888 13504
rect 11973 13560 12756 13562
rect 11973 13504 11978 13560
rect 12034 13504 12756 13560
rect 11973 13502 12756 13504
rect 10796 13500 10843 13502
rect 10777 13499 10843 13500
rect 11973 13499 12039 13502
rect 12750 13500 12756 13502
rect 12820 13500 12826 13564
rect 1025 13426 1091 13429
rect 11697 13426 11763 13429
rect 12617 13426 12683 13429
rect 1025 13424 11763 13426
rect 1025 13368 1030 13424
rect 1086 13368 11702 13424
rect 11758 13368 11763 13424
rect 1025 13366 11763 13368
rect 1025 13363 1091 13366
rect 11697 13363 11763 13366
rect 12390 13424 12683 13426
rect 12390 13368 12622 13424
rect 12678 13368 12683 13424
rect 12390 13366 12683 13368
rect 0 13290 800 13320
rect 1485 13290 1551 13293
rect 0 13288 1551 13290
rect 0 13232 1490 13288
rect 1546 13232 1551 13288
rect 0 13230 1551 13232
rect 0 13200 800 13230
rect 1485 13227 1551 13230
rect 1761 13290 1827 13293
rect 12390 13290 12450 13366
rect 12617 13363 12683 13366
rect 18873 13426 18939 13429
rect 21582 13426 21588 13428
rect 18873 13424 21588 13426
rect 18873 13368 18878 13424
rect 18934 13368 21588 13424
rect 18873 13366 21588 13368
rect 18873 13363 18939 13366
rect 21582 13364 21588 13366
rect 21652 13364 21658 13428
rect 18689 13290 18755 13293
rect 1761 13288 12450 13290
rect 1761 13232 1766 13288
rect 1822 13232 12450 13288
rect 1761 13230 12450 13232
rect 18646 13288 18755 13290
rect 18646 13232 18694 13288
rect 18750 13232 18755 13288
rect 1761 13227 1827 13230
rect 18646 13227 18755 13232
rect 21449 13290 21515 13293
rect 22200 13290 23000 13320
rect 21449 13288 23000 13290
rect 21449 13232 21454 13288
rect 21510 13232 23000 13288
rect 21449 13230 23000 13232
rect 21449 13227 21515 13230
rect 933 13154 999 13157
rect 8201 13154 8267 13157
rect 10910 13154 10916 13156
rect 933 13152 6010 13154
rect 933 13096 938 13152
rect 994 13096 6010 13152
rect 933 13094 6010 13096
rect 933 13091 999 13094
rect 1710 12956 1716 13020
rect 1780 13018 1786 13020
rect 4061 13018 4127 13021
rect 1780 13016 4127 13018
rect 1780 12960 4066 13016
rect 4122 12960 4127 13016
rect 1780 12958 4127 12960
rect 1780 12956 1786 12958
rect 4061 12955 4127 12958
rect 0 12882 800 12912
rect 1485 12882 1551 12885
rect 0 12880 1551 12882
rect 0 12824 1490 12880
rect 1546 12824 1551 12880
rect 0 12822 1551 12824
rect 5950 12882 6010 13094
rect 8201 13152 10916 13154
rect 8201 13096 8206 13152
rect 8262 13096 10916 13152
rect 8201 13094 10916 13096
rect 8201 13091 8267 13094
rect 10910 13092 10916 13094
rect 10980 13092 10986 13156
rect 14089 13154 14155 13157
rect 14590 13154 14596 13156
rect 14089 13152 14596 13154
rect 14089 13096 14094 13152
rect 14150 13096 14596 13152
rect 14089 13094 14596 13096
rect 14089 13091 14155 13094
rect 14590 13092 14596 13094
rect 14660 13092 14666 13156
rect 17033 13154 17099 13157
rect 18646 13154 18706 13227
rect 22200 13200 23000 13230
rect 20478 13154 20484 13156
rect 17033 13152 20484 13154
rect 17033 13096 17038 13152
rect 17094 13096 20484 13152
rect 17033 13094 20484 13096
rect 17033 13091 17099 13094
rect 20478 13092 20484 13094
rect 20548 13092 20554 13156
rect 6144 13088 6460 13089
rect 6144 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6460 13088
rect 6144 13023 6460 13024
rect 11342 13088 11658 13089
rect 11342 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11658 13088
rect 11342 13023 11658 13024
rect 16540 13088 16856 13089
rect 16540 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16856 13088
rect 16540 13023 16856 13024
rect 21738 13088 22054 13089
rect 21738 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22054 13088
rect 21738 13023 22054 13024
rect 8334 12956 8340 13020
rect 8404 13018 8410 13020
rect 11053 13018 11119 13021
rect 8404 13016 11119 13018
rect 8404 12960 11058 13016
rect 11114 12960 11119 13016
rect 8404 12958 11119 12960
rect 8404 12956 8410 12958
rect 11053 12955 11119 12958
rect 13629 13018 13695 13021
rect 13629 13016 16360 13018
rect 13629 12960 13634 13016
rect 13690 12960 16360 13016
rect 13629 12958 16360 12960
rect 13629 12955 13695 12958
rect 12801 12882 12867 12885
rect 13353 12884 13419 12885
rect 13302 12882 13308 12884
rect 5950 12880 12867 12882
rect 5950 12824 12806 12880
rect 12862 12824 12867 12880
rect 5950 12822 12867 12824
rect 13262 12822 13308 12882
rect 13372 12880 13419 12884
rect 13414 12824 13419 12880
rect 0 12792 800 12822
rect 1485 12819 1551 12822
rect 12801 12819 12867 12822
rect 13302 12820 13308 12822
rect 13372 12820 13419 12824
rect 13353 12819 13419 12820
rect 14181 12882 14247 12885
rect 14774 12882 14780 12884
rect 14181 12880 14780 12882
rect 14181 12824 14186 12880
rect 14242 12824 14780 12880
rect 14181 12822 14780 12824
rect 14181 12819 14247 12822
rect 14774 12820 14780 12822
rect 14844 12820 14850 12884
rect 16300 12882 16360 12958
rect 21081 12882 21147 12885
rect 22200 12882 23000 12912
rect 16300 12822 20914 12882
rect 1485 12746 1551 12749
rect 13537 12746 13603 12749
rect 1485 12744 13603 12746
rect 1485 12688 1490 12744
rect 1546 12688 13542 12744
rect 13598 12688 13603 12744
rect 1485 12686 13603 12688
rect 1485 12683 1551 12686
rect 13537 12683 13603 12686
rect 14365 12746 14431 12749
rect 18137 12746 18203 12749
rect 14365 12744 18203 12746
rect 14365 12688 14370 12744
rect 14426 12688 18142 12744
rect 18198 12688 18203 12744
rect 14365 12686 18203 12688
rect 20854 12746 20914 12822
rect 21081 12880 23000 12882
rect 21081 12824 21086 12880
rect 21142 12824 23000 12880
rect 21081 12822 23000 12824
rect 21081 12819 21147 12822
rect 22200 12792 23000 12822
rect 21214 12746 21220 12748
rect 20854 12686 21220 12746
rect 14365 12683 14431 12686
rect 18137 12683 18203 12686
rect 21214 12684 21220 12686
rect 21284 12684 21290 12748
rect 9438 12548 9444 12612
rect 9508 12610 9514 12612
rect 9581 12610 9647 12613
rect 9508 12608 9647 12610
rect 9508 12552 9586 12608
rect 9642 12552 9647 12608
rect 9508 12550 9647 12552
rect 9508 12548 9514 12550
rect 9581 12547 9647 12550
rect 9765 12610 9831 12613
rect 10593 12610 10659 12613
rect 9765 12608 10659 12610
rect 9765 12552 9770 12608
rect 9826 12552 10598 12608
rect 10654 12552 10659 12608
rect 9765 12550 10659 12552
rect 9765 12547 9831 12550
rect 10593 12547 10659 12550
rect 12617 12610 12683 12613
rect 12617 12608 13186 12610
rect 12617 12552 12622 12608
rect 12678 12552 13186 12608
rect 12617 12550 13186 12552
rect 12617 12547 12683 12550
rect 3545 12544 3861 12545
rect 0 12474 800 12504
rect 3545 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3861 12544
rect 3545 12479 3861 12480
rect 8743 12544 9059 12545
rect 8743 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9059 12544
rect 8743 12479 9059 12480
rect 1853 12474 1919 12477
rect 0 12472 1919 12474
rect 0 12416 1858 12472
rect 1914 12416 1919 12472
rect 0 12414 1919 12416
rect 0 12384 800 12414
rect 1853 12411 1919 12414
rect 5901 12474 5967 12477
rect 8293 12474 8359 12477
rect 5901 12472 8359 12474
rect 5901 12416 5906 12472
rect 5962 12416 8298 12472
rect 8354 12416 8359 12472
rect 5901 12414 8359 12416
rect 5901 12411 5967 12414
rect 8293 12411 8359 12414
rect 9438 12412 9444 12476
rect 9508 12474 9514 12476
rect 10358 12474 10364 12476
rect 9508 12414 10364 12474
rect 9508 12412 9514 12414
rect 10358 12412 10364 12414
rect 10428 12412 10434 12476
rect 13126 12450 13186 12550
rect 13941 12544 14257 12545
rect 13941 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14257 12544
rect 13941 12479 14257 12480
rect 19139 12544 19455 12545
rect 19139 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19455 12544
rect 19139 12479 19455 12480
rect 17585 12474 17651 12477
rect 21449 12474 21515 12477
rect 22200 12474 23000 12504
rect 17585 12472 19028 12474
rect 13261 12450 13327 12453
rect 13126 12448 13327 12450
rect 13126 12392 13266 12448
rect 13322 12392 13327 12448
rect 17585 12416 17590 12472
rect 17646 12416 19028 12472
rect 17585 12414 19028 12416
rect 17585 12411 17651 12414
rect 13126 12390 13327 12392
rect 13261 12387 13327 12390
rect 3969 12338 4035 12341
rect 4102 12338 4108 12340
rect 3969 12336 4108 12338
rect 3969 12280 3974 12336
rect 4030 12280 4108 12336
rect 3969 12278 4108 12280
rect 3969 12275 4035 12278
rect 4102 12276 4108 12278
rect 4172 12276 4178 12340
rect 8385 12338 8451 12341
rect 8518 12338 8524 12340
rect 8385 12336 8524 12338
rect 8385 12280 8390 12336
rect 8446 12280 8524 12336
rect 8385 12278 8524 12280
rect 8385 12275 8451 12278
rect 8518 12276 8524 12278
rect 8588 12338 8594 12340
rect 12566 12338 12572 12340
rect 8588 12278 12572 12338
rect 8588 12276 8594 12278
rect 12566 12276 12572 12278
rect 12636 12338 12642 12340
rect 13445 12338 13511 12341
rect 17718 12338 17724 12340
rect 12636 12278 13002 12338
rect 12636 12276 12642 12278
rect 2037 12202 2103 12205
rect 12709 12202 12775 12205
rect 2037 12200 12775 12202
rect 2037 12144 2042 12200
rect 2098 12144 12714 12200
rect 12770 12144 12775 12200
rect 2037 12142 12775 12144
rect 12942 12202 13002 12278
rect 13445 12336 17724 12338
rect 13445 12280 13450 12336
rect 13506 12280 17724 12336
rect 13445 12278 17724 12280
rect 13445 12275 13511 12278
rect 17718 12276 17724 12278
rect 17788 12276 17794 12340
rect 18968 12338 19028 12414
rect 21449 12472 23000 12474
rect 21449 12416 21454 12472
rect 21510 12416 23000 12472
rect 21449 12414 23000 12416
rect 21449 12411 21515 12414
rect 22200 12384 23000 12414
rect 19241 12338 19307 12341
rect 18968 12336 19307 12338
rect 18968 12280 19246 12336
rect 19302 12280 19307 12336
rect 18968 12278 19307 12280
rect 19241 12275 19307 12278
rect 21214 12276 21220 12340
rect 21284 12338 21290 12340
rect 21357 12338 21423 12341
rect 21284 12336 21423 12338
rect 21284 12280 21362 12336
rect 21418 12280 21423 12336
rect 21284 12278 21423 12280
rect 21284 12276 21290 12278
rect 21357 12275 21423 12278
rect 21582 12276 21588 12340
rect 21652 12338 21658 12340
rect 21725 12338 21791 12341
rect 21652 12336 21791 12338
rect 21652 12280 21730 12336
rect 21786 12280 21791 12336
rect 21652 12278 21791 12280
rect 21652 12276 21658 12278
rect 21725 12275 21791 12278
rect 14641 12202 14707 12205
rect 17861 12202 17927 12205
rect 20713 12202 20779 12205
rect 12942 12142 14290 12202
rect 2037 12139 2103 12142
rect 12709 12139 12775 12142
rect 0 12066 800 12096
rect 1485 12066 1551 12069
rect 7373 12068 7439 12069
rect 7373 12066 7420 12068
rect 0 12064 1551 12066
rect 0 12008 1490 12064
rect 1546 12008 1551 12064
rect 0 12006 1551 12008
rect 7328 12064 7420 12066
rect 7328 12008 7378 12064
rect 7328 12006 7420 12008
rect 0 11976 800 12006
rect 1485 12003 1551 12006
rect 7373 12004 7420 12006
rect 7484 12004 7490 12068
rect 9857 12066 9923 12069
rect 10542 12066 10548 12068
rect 9857 12064 10548 12066
rect 9857 12008 9862 12064
rect 9918 12008 10548 12064
rect 9857 12006 10548 12008
rect 7373 12003 7439 12004
rect 9857 12003 9923 12006
rect 10542 12004 10548 12006
rect 10612 12004 10618 12068
rect 13905 12066 13971 12069
rect 12390 12064 13971 12066
rect 12390 12008 13910 12064
rect 13966 12008 13971 12064
rect 12390 12006 13971 12008
rect 6144 12000 6460 12001
rect 6144 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6460 12000
rect 6144 11935 6460 11936
rect 11342 12000 11658 12001
rect 11342 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11658 12000
rect 11342 11935 11658 11936
rect 12390 11933 12450 12006
rect 13905 12003 13971 12006
rect 2681 11930 2747 11933
rect 4337 11930 4403 11933
rect 9581 11930 9647 11933
rect 9765 11930 9831 11933
rect 2681 11928 6010 11930
rect 2681 11872 2686 11928
rect 2742 11872 4342 11928
rect 4398 11872 6010 11928
rect 2681 11870 6010 11872
rect 2681 11867 2747 11870
rect 4337 11867 4403 11870
rect 1945 11794 2011 11797
rect 5717 11796 5783 11797
rect 1945 11792 2790 11794
rect 1945 11736 1950 11792
rect 2006 11736 2790 11792
rect 1945 11734 2790 11736
rect 1945 11731 2011 11734
rect 0 11658 800 11688
rect 2221 11658 2287 11661
rect 0 11656 2287 11658
rect 0 11600 2226 11656
rect 2282 11600 2287 11656
rect 0 11598 2287 11600
rect 2730 11658 2790 11734
rect 5717 11792 5764 11796
rect 5828 11794 5834 11796
rect 5950 11794 6010 11870
rect 6640 11928 9831 11930
rect 6640 11872 9586 11928
rect 9642 11872 9770 11928
rect 9826 11872 9831 11928
rect 6640 11870 9831 11872
rect 6640 11794 6700 11870
rect 9581 11867 9647 11870
rect 9765 11867 9831 11870
rect 11830 11868 11836 11932
rect 11900 11930 11906 11932
rect 12157 11930 12223 11933
rect 11900 11928 12223 11930
rect 11900 11872 12162 11928
rect 12218 11872 12223 11928
rect 11900 11870 12223 11872
rect 11900 11868 11906 11870
rect 12157 11867 12223 11870
rect 12390 11928 12499 11933
rect 12390 11872 12438 11928
rect 12494 11872 12499 11928
rect 12390 11867 12499 11872
rect 5717 11736 5722 11792
rect 5717 11732 5764 11736
rect 5828 11734 5874 11794
rect 5950 11734 6700 11794
rect 7373 11794 7439 11797
rect 12390 11794 12450 11867
rect 7373 11792 12450 11794
rect 7373 11736 7378 11792
rect 7434 11736 12450 11792
rect 7373 11734 12450 11736
rect 12709 11794 12775 11797
rect 14089 11794 14155 11797
rect 12709 11792 14155 11794
rect 12709 11736 12714 11792
rect 12770 11736 14094 11792
rect 14150 11736 14155 11792
rect 12709 11734 14155 11736
rect 14230 11794 14290 12142
rect 14641 12200 20779 12202
rect 14641 12144 14646 12200
rect 14702 12144 17866 12200
rect 17922 12144 20718 12200
rect 20774 12144 20779 12200
rect 14641 12142 20779 12144
rect 14641 12139 14707 12142
rect 17861 12139 17927 12142
rect 20713 12139 20779 12142
rect 21449 12202 21515 12205
rect 21449 12200 22202 12202
rect 21449 12144 21454 12200
rect 21510 12144 22202 12200
rect 21449 12142 22202 12144
rect 21449 12139 21515 12142
rect 22142 12096 22202 12142
rect 15101 12066 15167 12069
rect 16205 12066 16271 12069
rect 15101 12064 16271 12066
rect 15101 12008 15106 12064
rect 15162 12008 16210 12064
rect 16266 12008 16271 12064
rect 15101 12006 16271 12008
rect 22142 12006 23000 12096
rect 15101 12003 15167 12006
rect 16205 12003 16271 12006
rect 16540 12000 16856 12001
rect 16540 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16856 12000
rect 16540 11935 16856 11936
rect 21738 12000 22054 12001
rect 21738 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22054 12000
rect 22200 11976 23000 12006
rect 21738 11935 22054 11936
rect 14549 11930 14615 11933
rect 16205 11930 16271 11933
rect 14549 11928 16271 11930
rect 14549 11872 14554 11928
rect 14610 11872 16210 11928
rect 16266 11872 16271 11928
rect 14549 11870 16271 11872
rect 14549 11867 14615 11870
rect 16205 11867 16271 11870
rect 16941 11930 17007 11933
rect 17166 11930 17172 11932
rect 16941 11928 17172 11930
rect 16941 11872 16946 11928
rect 17002 11872 17172 11928
rect 16941 11870 17172 11872
rect 16941 11867 17007 11870
rect 17166 11868 17172 11870
rect 17236 11930 17242 11932
rect 19609 11930 19675 11933
rect 17236 11928 19675 11930
rect 17236 11872 19614 11928
rect 19670 11872 19675 11928
rect 17236 11870 19675 11872
rect 17236 11868 17242 11870
rect 19609 11867 19675 11870
rect 15193 11794 15259 11797
rect 19333 11794 19399 11797
rect 14230 11792 19399 11794
rect 14230 11736 15198 11792
rect 15254 11736 19338 11792
rect 19394 11736 19399 11792
rect 14230 11734 19399 11736
rect 5828 11732 5834 11734
rect 5717 11731 5783 11732
rect 7373 11731 7439 11734
rect 12709 11731 12775 11734
rect 14089 11731 14155 11734
rect 15193 11731 15259 11734
rect 19333 11731 19399 11734
rect 4705 11658 4771 11661
rect 11789 11658 11855 11661
rect 16849 11658 16915 11661
rect 17861 11658 17927 11661
rect 2730 11656 11855 11658
rect 2730 11600 4710 11656
rect 4766 11600 11794 11656
rect 11850 11600 11855 11656
rect 2730 11598 11855 11600
rect 0 11568 800 11598
rect 2221 11595 2287 11598
rect 4705 11595 4771 11598
rect 11789 11595 11855 11598
rect 13816 11656 17927 11658
rect 13816 11600 16854 11656
rect 16910 11600 17866 11656
rect 17922 11600 17927 11656
rect 13816 11598 17927 11600
rect 4797 11524 4863 11525
rect 4797 11522 4844 11524
rect 4752 11520 4844 11522
rect 4752 11464 4802 11520
rect 4752 11462 4844 11464
rect 4797 11460 4844 11462
rect 4908 11460 4914 11524
rect 7598 11460 7604 11524
rect 7668 11522 7674 11524
rect 8293 11522 8359 11525
rect 7668 11520 8359 11522
rect 7668 11464 8298 11520
rect 8354 11464 8359 11520
rect 7668 11462 8359 11464
rect 7668 11460 7674 11462
rect 4797 11459 4863 11460
rect 8293 11459 8359 11462
rect 9213 11522 9279 11525
rect 9806 11522 9812 11524
rect 9213 11520 9812 11522
rect 9213 11464 9218 11520
rect 9274 11464 9812 11520
rect 9213 11462 9812 11464
rect 9213 11459 9279 11462
rect 9806 11460 9812 11462
rect 9876 11522 9882 11524
rect 10726 11522 10732 11524
rect 9876 11462 10732 11522
rect 9876 11460 9882 11462
rect 10726 11460 10732 11462
rect 10796 11522 10802 11524
rect 13816 11522 13876 11598
rect 16849 11595 16915 11598
rect 17861 11595 17927 11598
rect 18045 11658 18111 11661
rect 20713 11658 20779 11661
rect 22200 11658 23000 11688
rect 18045 11656 23000 11658
rect 18045 11600 18050 11656
rect 18106 11600 20718 11656
rect 20774 11600 23000 11656
rect 18045 11598 23000 11600
rect 18045 11595 18111 11598
rect 20713 11595 20779 11598
rect 22200 11568 23000 11598
rect 15193 11524 15259 11525
rect 10796 11462 13876 11522
rect 10796 11460 10802 11462
rect 15142 11460 15148 11524
rect 15212 11522 15259 11524
rect 15510 11522 15516 11524
rect 15212 11520 15516 11522
rect 15254 11464 15516 11520
rect 15212 11462 15516 11464
rect 15212 11460 15259 11462
rect 15510 11460 15516 11462
rect 15580 11460 15586 11524
rect 15193 11459 15259 11460
rect 3545 11456 3861 11457
rect 3545 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3861 11456
rect 3545 11391 3861 11392
rect 8743 11456 9059 11457
rect 8743 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9059 11456
rect 8743 11391 9059 11392
rect 13941 11456 14257 11457
rect 13941 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14257 11456
rect 13941 11391 14257 11392
rect 19139 11456 19455 11457
rect 19139 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19455 11456
rect 19139 11391 19455 11392
rect 4429 11386 4495 11389
rect 8385 11386 8451 11389
rect 4429 11384 8451 11386
rect 4429 11328 4434 11384
rect 4490 11328 8390 11384
rect 8446 11328 8451 11384
rect 4429 11326 8451 11328
rect 4429 11323 4495 11326
rect 8385 11323 8451 11326
rect 9308 11326 11208 11386
rect 0 11250 800 11280
rect 1853 11250 1919 11253
rect 0 11248 1919 11250
rect 0 11192 1858 11248
rect 1914 11192 1919 11248
rect 0 11190 1919 11192
rect 0 11160 800 11190
rect 1853 11187 1919 11190
rect 4613 11250 4679 11253
rect 9029 11250 9095 11253
rect 4613 11248 9095 11250
rect 4613 11192 4618 11248
rect 4674 11192 9034 11248
rect 9090 11192 9095 11248
rect 4613 11190 9095 11192
rect 4613 11187 4679 11190
rect 9029 11187 9095 11190
rect 5390 11052 5396 11116
rect 5460 11114 5466 11116
rect 7833 11114 7899 11117
rect 9308 11114 9368 11326
rect 5460 11112 9368 11114
rect 5460 11056 7838 11112
rect 7894 11056 9368 11112
rect 5460 11054 9368 11056
rect 5460 11052 5466 11054
rect 7833 11051 7899 11054
rect 9438 11052 9444 11116
rect 9508 11114 9514 11116
rect 11148 11114 11208 11326
rect 11513 11250 11579 11253
rect 12065 11250 12131 11253
rect 14641 11250 14707 11253
rect 11513 11248 14707 11250
rect 11513 11192 11518 11248
rect 11574 11192 12070 11248
rect 12126 11192 14646 11248
rect 14702 11192 14707 11248
rect 11513 11190 14707 11192
rect 11513 11187 11579 11190
rect 12065 11187 12131 11190
rect 14641 11187 14707 11190
rect 19241 11250 19307 11253
rect 20529 11250 20595 11253
rect 19241 11248 20595 11250
rect 19241 11192 19246 11248
rect 19302 11192 20534 11248
rect 20590 11192 20595 11248
rect 19241 11190 20595 11192
rect 19241 11187 19307 11190
rect 20529 11187 20595 11190
rect 21081 11250 21147 11253
rect 22200 11250 23000 11280
rect 21081 11248 23000 11250
rect 21081 11192 21086 11248
rect 21142 11192 23000 11248
rect 21081 11190 23000 11192
rect 21081 11187 21147 11190
rect 22200 11160 23000 11190
rect 15561 11114 15627 11117
rect 9508 11054 10426 11114
rect 11148 11112 15627 11114
rect 11148 11056 15566 11112
rect 15622 11056 15627 11112
rect 11148 11054 15627 11056
rect 9508 11052 9514 11054
rect 9121 10978 9187 10981
rect 9581 10978 9647 10981
rect 9121 10976 9647 10978
rect 9121 10920 9126 10976
rect 9182 10920 9586 10976
rect 9642 10920 9647 10976
rect 9121 10918 9647 10920
rect 10366 10978 10426 11054
rect 15561 11051 15627 11054
rect 11145 10978 11211 10981
rect 10366 10976 11211 10978
rect 10366 10920 11150 10976
rect 11206 10920 11211 10976
rect 10366 10918 11211 10920
rect 9121 10915 9187 10918
rect 9581 10915 9647 10918
rect 11145 10915 11211 10918
rect 6144 10912 6460 10913
rect 0 10842 800 10872
rect 6144 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6460 10912
rect 6144 10847 6460 10848
rect 11342 10912 11658 10913
rect 11342 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11658 10912
rect 11342 10847 11658 10848
rect 16540 10912 16856 10913
rect 16540 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16856 10912
rect 16540 10847 16856 10848
rect 21738 10912 22054 10913
rect 21738 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22054 10912
rect 21738 10847 22054 10848
rect 1485 10842 1551 10845
rect 9438 10842 9444 10844
rect 0 10840 1551 10842
rect 0 10784 1490 10840
rect 1546 10784 1551 10840
rect 0 10782 1551 10784
rect 0 10752 800 10782
rect 1485 10779 1551 10782
rect 6686 10782 9444 10842
rect 2497 10706 2563 10709
rect 3877 10706 3943 10709
rect 2497 10704 3943 10706
rect 2497 10648 2502 10704
rect 2558 10648 3882 10704
rect 3938 10648 3943 10704
rect 2497 10646 3943 10648
rect 2497 10643 2563 10646
rect 3877 10643 3943 10646
rect 4705 10706 4771 10709
rect 6686 10706 6746 10782
rect 9438 10780 9444 10782
rect 9508 10780 9514 10844
rect 10174 10780 10180 10844
rect 10244 10842 10250 10844
rect 10685 10842 10751 10845
rect 10244 10840 10751 10842
rect 10244 10784 10690 10840
rect 10746 10784 10751 10840
rect 10244 10782 10751 10784
rect 10244 10780 10250 10782
rect 10685 10779 10751 10782
rect 13118 10780 13124 10844
rect 13188 10842 13194 10844
rect 14181 10842 14247 10845
rect 22200 10842 23000 10872
rect 13188 10840 14247 10842
rect 13188 10784 14186 10840
rect 14242 10784 14247 10840
rect 13188 10782 14247 10784
rect 13188 10780 13194 10782
rect 14181 10779 14247 10782
rect 22142 10752 23000 10842
rect 4705 10704 6746 10706
rect 4705 10648 4710 10704
rect 4766 10648 6746 10704
rect 4705 10646 6746 10648
rect 4705 10643 4771 10646
rect 9990 10644 9996 10708
rect 10060 10706 10066 10708
rect 11237 10706 11303 10709
rect 10060 10704 11303 10706
rect 10060 10648 11242 10704
rect 11298 10648 11303 10704
rect 10060 10646 11303 10648
rect 10060 10644 10066 10646
rect 11237 10643 11303 10646
rect 15469 10706 15535 10709
rect 17861 10706 17927 10709
rect 15469 10704 17927 10706
rect 15469 10648 15474 10704
rect 15530 10648 17866 10704
rect 17922 10648 17927 10704
rect 15469 10646 17927 10648
rect 15469 10643 15535 10646
rect 17861 10643 17927 10646
rect 20437 10706 20503 10709
rect 22142 10706 22202 10752
rect 20437 10704 22202 10706
rect 20437 10648 20442 10704
rect 20498 10648 22202 10704
rect 20437 10646 22202 10648
rect 20437 10643 20503 10646
rect 1853 10570 1919 10573
rect 9673 10570 9739 10573
rect 1853 10568 9739 10570
rect 1853 10512 1858 10568
rect 1914 10512 9678 10568
rect 9734 10512 9739 10568
rect 1853 10510 9739 10512
rect 1853 10507 1919 10510
rect 9673 10507 9739 10510
rect 12985 10570 13051 10573
rect 16757 10570 16823 10573
rect 12985 10568 16823 10570
rect 12985 10512 12990 10568
rect 13046 10512 16762 10568
rect 16818 10512 16823 10568
rect 12985 10510 16823 10512
rect 12985 10507 13051 10510
rect 16757 10507 16823 10510
rect 17125 10570 17191 10573
rect 18137 10570 18203 10573
rect 17125 10568 18203 10570
rect 17125 10512 17130 10568
rect 17186 10512 18142 10568
rect 18198 10512 18203 10568
rect 17125 10510 18203 10512
rect 17125 10507 17191 10510
rect 18137 10507 18203 10510
rect 18965 10570 19031 10573
rect 18965 10568 19626 10570
rect 18965 10512 18970 10568
rect 19026 10512 19626 10568
rect 18965 10510 19626 10512
rect 18965 10507 19031 10510
rect 0 10434 800 10464
rect 1485 10434 1551 10437
rect 0 10432 1551 10434
rect 0 10376 1490 10432
rect 1546 10376 1551 10432
rect 0 10374 1551 10376
rect 0 10344 800 10374
rect 1485 10371 1551 10374
rect 7281 10434 7347 10437
rect 8017 10434 8083 10437
rect 7281 10432 8083 10434
rect 7281 10376 7286 10432
rect 7342 10376 8022 10432
rect 8078 10376 8083 10432
rect 7281 10374 8083 10376
rect 7281 10371 7347 10374
rect 8017 10371 8083 10374
rect 9305 10434 9371 10437
rect 9622 10434 9628 10436
rect 9305 10432 9628 10434
rect 9305 10376 9310 10432
rect 9366 10376 9628 10432
rect 9305 10374 9628 10376
rect 9305 10371 9371 10374
rect 9622 10372 9628 10374
rect 9692 10372 9698 10436
rect 19566 10434 19626 10510
rect 22200 10434 23000 10464
rect 19566 10374 23000 10434
rect 3545 10368 3861 10369
rect 3545 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3861 10368
rect 3545 10303 3861 10304
rect 8743 10368 9059 10369
rect 8743 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9059 10368
rect 8743 10303 9059 10304
rect 13941 10368 14257 10369
rect 13941 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14257 10368
rect 13941 10303 14257 10304
rect 19139 10368 19455 10369
rect 19139 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19455 10368
rect 22200 10344 23000 10374
rect 19139 10303 19455 10304
rect 4654 10236 4660 10300
rect 4724 10298 4730 10300
rect 6545 10298 6611 10301
rect 13118 10298 13124 10300
rect 4724 10296 8402 10298
rect 4724 10240 6550 10296
rect 6606 10240 8402 10296
rect 4724 10238 8402 10240
rect 4724 10236 4730 10238
rect 6545 10235 6611 10238
rect 1853 10162 1919 10165
rect 8109 10162 8175 10165
rect 1853 10160 8175 10162
rect 1853 10104 1858 10160
rect 1914 10104 8114 10160
rect 8170 10104 8175 10160
rect 1853 10102 8175 10104
rect 8342 10162 8402 10238
rect 9124 10238 13124 10298
rect 9124 10162 9184 10238
rect 13118 10236 13124 10238
rect 13188 10236 13194 10300
rect 16205 10298 16271 10301
rect 18413 10298 18479 10301
rect 18689 10298 18755 10301
rect 16205 10296 18755 10298
rect 16205 10240 16210 10296
rect 16266 10240 18418 10296
rect 18474 10240 18694 10296
rect 18750 10240 18755 10296
rect 16205 10238 18755 10240
rect 16205 10235 16271 10238
rect 18413 10235 18479 10238
rect 18689 10235 18755 10238
rect 8342 10102 9184 10162
rect 9305 10162 9371 10165
rect 11094 10162 11100 10164
rect 9305 10160 11100 10162
rect 9305 10104 9310 10160
rect 9366 10104 11100 10160
rect 9305 10102 11100 10104
rect 1853 10099 1919 10102
rect 8109 10099 8175 10102
rect 9305 10099 9371 10102
rect 11094 10100 11100 10102
rect 11164 10100 11170 10164
rect 11513 10162 11579 10165
rect 11830 10162 11836 10164
rect 11513 10160 11836 10162
rect 11513 10104 11518 10160
rect 11574 10104 11836 10160
rect 11513 10102 11836 10104
rect 11513 10099 11579 10102
rect 11830 10100 11836 10102
rect 11900 10100 11906 10164
rect 12934 10100 12940 10164
rect 13004 10162 13010 10164
rect 13813 10162 13879 10165
rect 13004 10160 13879 10162
rect 13004 10104 13818 10160
rect 13874 10104 13879 10160
rect 13004 10102 13879 10104
rect 13004 10100 13010 10102
rect 13813 10099 13879 10102
rect 13997 10162 14063 10165
rect 18413 10162 18479 10165
rect 13997 10160 18479 10162
rect 13997 10104 14002 10160
rect 14058 10104 18418 10160
rect 18474 10104 18479 10160
rect 13997 10102 18479 10104
rect 13997 10099 14063 10102
rect 18413 10099 18479 10102
rect 0 10026 800 10056
rect 2497 10026 2563 10029
rect 0 10024 2563 10026
rect 0 9968 2502 10024
rect 2558 9968 2563 10024
rect 0 9966 2563 9968
rect 0 9936 800 9966
rect 2497 9963 2563 9966
rect 4153 10026 4219 10029
rect 10593 10026 10659 10029
rect 10961 10026 11027 10029
rect 16113 10026 16179 10029
rect 4153 10024 11027 10026
rect 4153 9968 4158 10024
rect 4214 9968 10598 10024
rect 10654 9968 10966 10024
rect 11022 9968 11027 10024
rect 4153 9966 11027 9968
rect 4153 9963 4219 9966
rect 10593 9963 10659 9966
rect 10961 9963 11027 9966
rect 11148 10024 16179 10026
rect 11148 9968 16118 10024
rect 16174 9968 16179 10024
rect 11148 9966 16179 9968
rect 4705 9890 4771 9893
rect 2730 9888 4771 9890
rect 2730 9832 4710 9888
rect 4766 9832 4771 9888
rect 2730 9830 4771 9832
rect 2037 9754 2103 9757
rect 2730 9754 2790 9830
rect 4705 9827 4771 9830
rect 8109 9890 8175 9893
rect 8937 9890 9003 9893
rect 11148 9890 11208 9966
rect 16113 9963 16179 9966
rect 17769 10026 17835 10029
rect 19742 10026 19748 10028
rect 17769 10024 19748 10026
rect 17769 9968 17774 10024
rect 17830 9968 19748 10024
rect 17769 9966 19748 9968
rect 17769 9963 17835 9966
rect 19742 9964 19748 9966
rect 19812 10026 19818 10028
rect 20110 10026 20116 10028
rect 19812 9966 20116 10026
rect 19812 9964 19818 9966
rect 20110 9964 20116 9966
rect 20180 9964 20186 10028
rect 20713 10026 20779 10029
rect 22200 10026 23000 10056
rect 20713 10024 23000 10026
rect 20713 9968 20718 10024
rect 20774 9968 23000 10024
rect 20713 9966 23000 9968
rect 20713 9963 20779 9966
rect 22200 9936 23000 9966
rect 13629 9892 13695 9893
rect 13629 9890 13676 9892
rect 8109 9888 11208 9890
rect 8109 9832 8114 9888
rect 8170 9832 8942 9888
rect 8998 9832 11208 9888
rect 8109 9830 11208 9832
rect 13584 9888 13676 9890
rect 13584 9832 13634 9888
rect 13584 9830 13676 9832
rect 8109 9827 8175 9830
rect 8937 9827 9003 9830
rect 13629 9828 13676 9830
rect 13740 9828 13746 9892
rect 14549 9890 14615 9893
rect 15326 9890 15332 9892
rect 14549 9888 15332 9890
rect 14549 9832 14554 9888
rect 14610 9832 15332 9888
rect 14549 9830 15332 9832
rect 13629 9827 13695 9828
rect 14549 9827 14615 9830
rect 15326 9828 15332 9830
rect 15396 9828 15402 9892
rect 16113 9890 16179 9893
rect 16246 9890 16252 9892
rect 16113 9888 16252 9890
rect 16113 9832 16118 9888
rect 16174 9832 16252 9888
rect 16113 9830 16252 9832
rect 16113 9827 16179 9830
rect 16246 9828 16252 9830
rect 16316 9828 16322 9892
rect 17902 9828 17908 9892
rect 17972 9890 17978 9892
rect 18689 9890 18755 9893
rect 17972 9888 18755 9890
rect 17972 9832 18694 9888
rect 18750 9832 18755 9888
rect 17972 9830 18755 9832
rect 17972 9828 17978 9830
rect 18689 9827 18755 9830
rect 6144 9824 6460 9825
rect 6144 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6460 9824
rect 6144 9759 6460 9760
rect 11342 9824 11658 9825
rect 11342 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11658 9824
rect 11342 9759 11658 9760
rect 16540 9824 16856 9825
rect 16540 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16856 9824
rect 16540 9759 16856 9760
rect 21738 9824 22054 9825
rect 21738 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22054 9824
rect 21738 9759 22054 9760
rect 2037 9752 2790 9754
rect 2037 9696 2042 9752
rect 2098 9696 2790 9752
rect 2037 9694 2790 9696
rect 3049 9754 3115 9757
rect 3601 9754 3667 9757
rect 3049 9752 3667 9754
rect 3049 9696 3054 9752
rect 3110 9696 3606 9752
rect 3662 9696 3667 9752
rect 3049 9694 3667 9696
rect 2037 9691 2103 9694
rect 3049 9691 3115 9694
rect 3601 9691 3667 9694
rect 3785 9754 3851 9757
rect 6913 9754 6979 9757
rect 7649 9754 7715 9757
rect 3785 9752 5964 9754
rect 3785 9696 3790 9752
rect 3846 9696 5964 9752
rect 3785 9694 5964 9696
rect 3785 9691 3851 9694
rect 0 9618 800 9648
rect 1485 9618 1551 9621
rect 0 9616 1551 9618
rect 0 9560 1490 9616
rect 1546 9560 1551 9616
rect 0 9558 1551 9560
rect 0 9528 800 9558
rect 1485 9555 1551 9558
rect 3417 9618 3483 9621
rect 4061 9618 4127 9621
rect 3417 9616 4127 9618
rect 3417 9560 3422 9616
rect 3478 9560 4066 9616
rect 4122 9560 4127 9616
rect 3417 9558 4127 9560
rect 5904 9618 5964 9694
rect 6913 9752 7715 9754
rect 6913 9696 6918 9752
rect 6974 9696 7654 9752
rect 7710 9696 7715 9752
rect 6913 9694 7715 9696
rect 6913 9691 6979 9694
rect 7649 9691 7715 9694
rect 7833 9754 7899 9757
rect 8201 9756 8267 9757
rect 8150 9754 8156 9756
rect 7833 9752 8156 9754
rect 8220 9752 8267 9756
rect 7833 9696 7838 9752
rect 7894 9696 8156 9752
rect 8262 9696 8267 9752
rect 7833 9694 8156 9696
rect 7833 9691 7899 9694
rect 8150 9692 8156 9694
rect 8220 9692 8267 9696
rect 8334 9692 8340 9756
rect 8404 9754 8410 9756
rect 9121 9754 9187 9757
rect 8404 9752 9187 9754
rect 8404 9696 9126 9752
rect 9182 9696 9187 9752
rect 8404 9694 9187 9696
rect 8404 9692 8410 9694
rect 8201 9691 8267 9692
rect 9121 9691 9187 9694
rect 9254 9692 9260 9756
rect 9324 9754 9330 9756
rect 9581 9754 9647 9757
rect 9324 9752 9647 9754
rect 9324 9696 9586 9752
rect 9642 9696 9647 9752
rect 9324 9694 9647 9696
rect 9324 9692 9330 9694
rect 9581 9691 9647 9694
rect 11973 9754 12039 9757
rect 12198 9754 12204 9756
rect 11973 9752 12204 9754
rect 11973 9696 11978 9752
rect 12034 9696 12204 9752
rect 11973 9694 12204 9696
rect 11973 9691 12039 9694
rect 12198 9692 12204 9694
rect 12268 9692 12274 9756
rect 13721 9754 13787 9757
rect 17493 9756 17559 9757
rect 17493 9754 17540 9756
rect 13721 9752 16314 9754
rect 13721 9696 13726 9752
rect 13782 9696 16314 9752
rect 13721 9694 16314 9696
rect 17448 9752 17540 9754
rect 17448 9696 17498 9752
rect 17448 9694 17540 9696
rect 13721 9691 13787 9694
rect 8753 9618 8819 9621
rect 5904 9616 8819 9618
rect 5904 9560 8758 9616
rect 8814 9560 8819 9616
rect 5904 9558 8819 9560
rect 3417 9555 3483 9558
rect 4061 9555 4127 9558
rect 8753 9555 8819 9558
rect 9622 9556 9628 9620
rect 9692 9618 9698 9620
rect 10133 9618 10199 9621
rect 11789 9618 11855 9621
rect 9692 9616 10199 9618
rect 9692 9560 10138 9616
rect 10194 9560 10199 9616
rect 9692 9558 10199 9560
rect 9692 9556 9698 9558
rect 10133 9555 10199 9558
rect 10734 9616 11855 9618
rect 10734 9560 11794 9616
rect 11850 9560 11855 9616
rect 10734 9558 11855 9560
rect 3325 9482 3391 9485
rect 3693 9482 3759 9485
rect 3325 9480 3759 9482
rect 3325 9424 3330 9480
rect 3386 9424 3698 9480
rect 3754 9424 3759 9480
rect 3325 9422 3759 9424
rect 3325 9419 3391 9422
rect 3693 9419 3759 9422
rect 3918 9420 3924 9484
rect 3988 9482 3994 9484
rect 4061 9482 4127 9485
rect 3988 9480 4127 9482
rect 3988 9424 4066 9480
rect 4122 9424 4127 9480
rect 3988 9422 4127 9424
rect 3988 9420 3994 9422
rect 4061 9419 4127 9422
rect 4245 9484 4311 9485
rect 4245 9480 4292 9484
rect 4356 9482 4362 9484
rect 4245 9424 4250 9480
rect 4245 9420 4292 9424
rect 4356 9422 4402 9482
rect 4356 9420 4362 9422
rect 7782 9420 7788 9484
rect 7852 9482 7858 9484
rect 10734 9482 10794 9558
rect 11789 9555 11855 9558
rect 11973 9618 12039 9621
rect 12525 9618 12591 9621
rect 14825 9618 14891 9621
rect 15285 9618 15351 9621
rect 11973 9616 12718 9618
rect 11973 9560 11978 9616
rect 12034 9560 12530 9616
rect 12586 9560 12718 9616
rect 11973 9558 12718 9560
rect 14825 9616 15351 9618
rect 14825 9560 14830 9616
rect 14886 9560 15290 9616
rect 15346 9560 15351 9616
rect 14825 9558 15351 9560
rect 16254 9618 16314 9694
rect 17493 9692 17540 9694
rect 17604 9692 17610 9756
rect 17493 9691 17559 9692
rect 16982 9618 16988 9620
rect 16254 9558 16988 9618
rect 11973 9555 12039 9558
rect 12525 9555 12634 9558
rect 14825 9555 14891 9558
rect 15285 9555 15351 9558
rect 16982 9556 16988 9558
rect 17052 9556 17058 9620
rect 18045 9618 18111 9621
rect 18270 9618 18276 9620
rect 18045 9616 18276 9618
rect 18045 9560 18050 9616
rect 18106 9560 18276 9616
rect 18045 9558 18276 9560
rect 18045 9555 18111 9558
rect 18270 9556 18276 9558
rect 18340 9556 18346 9620
rect 18873 9618 18939 9621
rect 22200 9618 23000 9648
rect 18873 9616 23000 9618
rect 18873 9560 18878 9616
rect 18934 9560 23000 9616
rect 18873 9558 23000 9560
rect 18873 9555 18939 9558
rect 7852 9422 10794 9482
rect 10869 9482 10935 9485
rect 12433 9482 12499 9485
rect 10869 9480 12499 9482
rect 10869 9424 10874 9480
rect 10930 9424 12438 9480
rect 12494 9424 12499 9480
rect 10869 9422 12499 9424
rect 12574 9482 12634 9555
rect 22200 9528 23000 9558
rect 17769 9482 17835 9485
rect 12574 9480 17835 9482
rect 12574 9424 17774 9480
rect 17830 9424 17835 9480
rect 12574 9422 17835 9424
rect 7852 9420 7858 9422
rect 4245 9419 4311 9420
rect 10869 9419 10935 9422
rect 12433 9419 12499 9422
rect 17769 9419 17835 9422
rect 4061 9346 4127 9349
rect 6177 9346 6243 9349
rect 7966 9346 7972 9348
rect 4061 9344 6243 9346
rect 4061 9288 4066 9344
rect 4122 9288 6182 9344
rect 6238 9288 6243 9344
rect 4061 9286 6243 9288
rect 4061 9283 4127 9286
rect 6177 9283 6243 9286
rect 7468 9286 7972 9346
rect 3545 9280 3861 9281
rect 0 9210 800 9240
rect 3545 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3861 9280
rect 3545 9215 3861 9216
rect 7468 9213 7528 9286
rect 7966 9284 7972 9286
rect 8036 9284 8042 9348
rect 10961 9346 11027 9349
rect 13353 9346 13419 9349
rect 10961 9344 13419 9346
rect 10961 9288 10966 9344
rect 11022 9288 13358 9344
rect 13414 9288 13419 9344
rect 10961 9286 13419 9288
rect 10961 9283 11027 9286
rect 13353 9283 13419 9286
rect 14406 9284 14412 9348
rect 14476 9346 14482 9348
rect 14641 9346 14707 9349
rect 14476 9344 14707 9346
rect 14476 9288 14646 9344
rect 14702 9288 14707 9344
rect 14476 9286 14707 9288
rect 14476 9284 14482 9286
rect 14641 9283 14707 9286
rect 15469 9346 15535 9349
rect 18689 9348 18755 9349
rect 15469 9344 18568 9346
rect 15469 9288 15474 9344
rect 15530 9288 18568 9344
rect 15469 9286 18568 9288
rect 15469 9283 15535 9286
rect 8743 9280 9059 9281
rect 8743 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9059 9280
rect 8743 9215 9059 9216
rect 13941 9280 14257 9281
rect 13941 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14257 9280
rect 13941 9215 14257 9216
rect 7465 9210 7531 9213
rect 7833 9212 7899 9213
rect 0 9150 2790 9210
rect 0 9120 800 9150
rect 2730 9074 2790 9150
rect 4156 9208 7531 9210
rect 4156 9152 7470 9208
rect 7526 9152 7531 9208
rect 4156 9150 7531 9152
rect 3601 9074 3667 9077
rect 2730 9072 3667 9074
rect 2730 9016 3606 9072
rect 3662 9016 3667 9072
rect 2730 9014 3667 9016
rect 3601 9011 3667 9014
rect 1853 8938 1919 8941
rect 4156 8938 4216 9150
rect 7465 9147 7531 9150
rect 7782 9148 7788 9212
rect 7852 9210 7899 9212
rect 8109 9212 8175 9213
rect 7852 9208 7944 9210
rect 7894 9152 7944 9208
rect 7852 9150 7944 9152
rect 8109 9208 8156 9212
rect 8220 9210 8226 9212
rect 8109 9152 8114 9208
rect 7852 9148 7899 9150
rect 7833 9147 7899 9148
rect 8109 9148 8156 9152
rect 8220 9150 8266 9210
rect 8220 9148 8226 9150
rect 11094 9148 11100 9212
rect 11164 9210 11170 9212
rect 11605 9210 11671 9213
rect 11164 9208 11671 9210
rect 11164 9152 11610 9208
rect 11666 9152 11671 9208
rect 11164 9150 11671 9152
rect 11164 9148 11170 9150
rect 8109 9147 8175 9148
rect 11605 9147 11671 9150
rect 11789 9210 11855 9213
rect 13353 9210 13419 9213
rect 11789 9208 13419 9210
rect 11789 9152 11794 9208
rect 11850 9152 13358 9208
rect 13414 9152 13419 9208
rect 11789 9150 13419 9152
rect 11789 9147 11855 9150
rect 13353 9147 13419 9150
rect 15469 9210 15535 9213
rect 15694 9210 15700 9212
rect 15469 9208 15700 9210
rect 15469 9152 15474 9208
rect 15530 9152 15700 9208
rect 15469 9150 15700 9152
rect 15469 9147 15535 9150
rect 15694 9148 15700 9150
rect 15764 9210 15770 9212
rect 17902 9210 17908 9212
rect 15764 9150 17908 9210
rect 15764 9148 15770 9150
rect 17902 9148 17908 9150
rect 17972 9210 17978 9212
rect 18321 9210 18387 9213
rect 17972 9208 18387 9210
rect 17972 9152 18326 9208
rect 18382 9152 18387 9208
rect 17972 9150 18387 9152
rect 18508 9210 18568 9286
rect 18638 9284 18644 9348
rect 18708 9346 18755 9348
rect 20253 9346 20319 9349
rect 20662 9346 20668 9348
rect 18708 9344 18800 9346
rect 18750 9288 18800 9344
rect 18708 9286 18800 9288
rect 20253 9344 20668 9346
rect 20253 9288 20258 9344
rect 20314 9288 20668 9344
rect 20253 9286 20668 9288
rect 18708 9284 18755 9286
rect 18689 9283 18755 9284
rect 20253 9283 20319 9286
rect 20662 9284 20668 9286
rect 20732 9284 20738 9348
rect 19139 9280 19455 9281
rect 19139 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19455 9280
rect 19139 9215 19455 9216
rect 18873 9210 18939 9213
rect 18508 9208 18939 9210
rect 18508 9152 18878 9208
rect 18934 9152 18939 9208
rect 18508 9150 18939 9152
rect 17972 9148 17978 9150
rect 18321 9147 18387 9150
rect 18873 9147 18939 9150
rect 20253 9210 20319 9213
rect 22200 9210 23000 9240
rect 20253 9208 23000 9210
rect 20253 9152 20258 9208
rect 20314 9152 23000 9208
rect 20253 9150 23000 9152
rect 20253 9147 20319 9150
rect 22200 9120 23000 9150
rect 4286 9012 4292 9076
rect 4356 9074 4362 9076
rect 4613 9074 4679 9077
rect 4356 9072 4679 9074
rect 4356 9016 4618 9072
rect 4674 9016 4679 9072
rect 4356 9014 4679 9016
rect 4356 9012 4362 9014
rect 4613 9011 4679 9014
rect 5625 9074 5691 9077
rect 10133 9074 10199 9077
rect 12382 9074 12388 9076
rect 5625 9072 12388 9074
rect 5625 9016 5630 9072
rect 5686 9016 10138 9072
rect 10194 9016 12388 9072
rect 5625 9014 12388 9016
rect 5625 9011 5691 9014
rect 10133 9011 10199 9014
rect 12382 9012 12388 9014
rect 12452 9012 12458 9076
rect 12525 9074 12591 9077
rect 20897 9074 20963 9077
rect 12525 9072 20963 9074
rect 12525 9016 12530 9072
rect 12586 9016 20902 9072
rect 20958 9016 20963 9072
rect 12525 9014 20963 9016
rect 12525 9011 12591 9014
rect 20897 9011 20963 9014
rect 6637 8940 6703 8941
rect 1853 8936 4216 8938
rect 1853 8880 1858 8936
rect 1914 8880 4216 8936
rect 1853 8878 4216 8880
rect 1853 8875 1919 8878
rect 4286 8876 4292 8940
rect 4356 8938 4362 8940
rect 6637 8938 6684 8940
rect 4356 8878 6010 8938
rect 6556 8936 6684 8938
rect 6748 8938 6754 8940
rect 15009 8938 15075 8941
rect 18321 8938 18387 8941
rect 18781 8938 18847 8941
rect 6748 8936 15075 8938
rect 6556 8880 6642 8936
rect 6748 8880 15014 8936
rect 15070 8880 15075 8936
rect 6556 8878 6684 8880
rect 4356 8876 4362 8878
rect 0 8802 800 8832
rect 1393 8802 1459 8805
rect 5574 8802 5580 8804
rect 0 8800 5580 8802
rect 0 8744 1398 8800
rect 1454 8744 5580 8800
rect 0 8742 5580 8744
rect 0 8712 800 8742
rect 1393 8739 1459 8742
rect 5574 8740 5580 8742
rect 5644 8740 5650 8804
rect 2129 8666 2195 8669
rect 4797 8666 4863 8669
rect 2129 8664 4863 8666
rect 2129 8608 2134 8664
rect 2190 8608 4802 8664
rect 4858 8608 4863 8664
rect 2129 8606 4863 8608
rect 2129 8603 2195 8606
rect 4797 8603 4863 8606
rect 5257 8666 5323 8669
rect 5809 8666 5875 8669
rect 5257 8664 5875 8666
rect 5257 8608 5262 8664
rect 5318 8608 5814 8664
rect 5870 8608 5875 8664
rect 5257 8606 5875 8608
rect 5257 8603 5323 8606
rect 5809 8603 5875 8606
rect 2773 8530 2839 8533
rect 5257 8530 5323 8533
rect 2773 8528 5323 8530
rect 2773 8472 2778 8528
rect 2834 8472 5262 8528
rect 5318 8472 5323 8528
rect 2773 8470 5323 8472
rect 5950 8530 6010 8878
rect 6637 8876 6684 8878
rect 6748 8878 15075 8880
rect 6748 8876 6754 8878
rect 6637 8875 6703 8876
rect 15009 8875 15075 8878
rect 16254 8878 17970 8938
rect 6862 8740 6868 8804
rect 6932 8802 6938 8804
rect 7005 8802 7071 8805
rect 7598 8802 7604 8804
rect 6932 8800 7604 8802
rect 6932 8744 7010 8800
rect 7066 8744 7604 8800
rect 6932 8742 7604 8744
rect 6932 8740 6938 8742
rect 7005 8739 7071 8742
rect 7598 8740 7604 8742
rect 7668 8740 7674 8804
rect 7966 8740 7972 8804
rect 8036 8802 8042 8804
rect 10910 8802 10916 8804
rect 8036 8742 10916 8802
rect 8036 8740 8042 8742
rect 10910 8740 10916 8742
rect 10980 8740 10986 8804
rect 12566 8740 12572 8804
rect 12636 8802 12642 8804
rect 16254 8802 16314 8878
rect 12636 8742 16314 8802
rect 17910 8802 17970 8878
rect 18321 8936 18847 8938
rect 18321 8880 18326 8936
rect 18382 8880 18786 8936
rect 18842 8880 18847 8936
rect 18321 8878 18847 8880
rect 18321 8875 18387 8878
rect 18781 8875 18847 8878
rect 18965 8938 19031 8941
rect 18965 8936 22202 8938
rect 18965 8880 18970 8936
rect 19026 8880 22202 8936
rect 18965 8878 22202 8880
rect 18965 8875 19031 8878
rect 22142 8832 22202 8878
rect 20294 8802 20300 8804
rect 17910 8742 20300 8802
rect 12636 8740 12642 8742
rect 20294 8740 20300 8742
rect 20364 8802 20370 8804
rect 20437 8802 20503 8805
rect 20364 8800 20503 8802
rect 20364 8744 20442 8800
rect 20498 8744 20503 8800
rect 20364 8742 20503 8744
rect 22142 8742 23000 8832
rect 20364 8740 20370 8742
rect 20437 8739 20503 8742
rect 6144 8736 6460 8737
rect 6144 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6460 8736
rect 6144 8671 6460 8672
rect 11342 8736 11658 8737
rect 11342 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11658 8736
rect 11342 8671 11658 8672
rect 16540 8736 16856 8737
rect 16540 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16856 8736
rect 16540 8671 16856 8672
rect 21738 8736 22054 8737
rect 21738 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22054 8736
rect 22200 8712 23000 8742
rect 21738 8671 22054 8672
rect 9305 8666 9371 8669
rect 14406 8666 14412 8668
rect 6686 8664 9371 8666
rect 6686 8608 9310 8664
rect 9366 8608 9371 8664
rect 6686 8606 9371 8608
rect 6686 8530 6746 8606
rect 9305 8603 9371 8606
rect 12574 8606 14412 8666
rect 6913 8532 6979 8533
rect 5950 8470 6746 8530
rect 2773 8467 2839 8470
rect 5257 8467 5323 8470
rect 6862 8468 6868 8532
rect 6932 8530 6979 8532
rect 7557 8532 7623 8533
rect 7557 8530 7604 8532
rect 6932 8528 7024 8530
rect 6974 8472 7024 8528
rect 6932 8470 7024 8472
rect 7512 8528 7604 8530
rect 7512 8472 7562 8528
rect 7512 8470 7604 8472
rect 6932 8468 6979 8470
rect 6913 8467 6979 8468
rect 7557 8468 7604 8470
rect 7668 8468 7674 8532
rect 8201 8530 8267 8533
rect 12574 8530 12634 8606
rect 14406 8604 14412 8606
rect 14476 8604 14482 8668
rect 14733 8666 14799 8669
rect 15326 8666 15332 8668
rect 14733 8664 15332 8666
rect 14733 8608 14738 8664
rect 14794 8608 15332 8664
rect 14733 8606 15332 8608
rect 14733 8603 14799 8606
rect 15326 8604 15332 8606
rect 15396 8604 15402 8668
rect 21541 8666 21607 8669
rect 16990 8664 21607 8666
rect 16990 8608 21546 8664
rect 21602 8608 21607 8664
rect 16990 8606 21607 8608
rect 8201 8528 12634 8530
rect 8201 8472 8206 8528
rect 8262 8472 12634 8528
rect 8201 8470 12634 8472
rect 12709 8530 12775 8533
rect 13118 8530 13124 8532
rect 12709 8528 13124 8530
rect 12709 8472 12714 8528
rect 12770 8472 13124 8528
rect 12709 8470 13124 8472
rect 7557 8467 7623 8468
rect 8201 8467 8267 8470
rect 12709 8467 12775 8470
rect 13118 8468 13124 8470
rect 13188 8530 13194 8532
rect 13353 8530 13419 8533
rect 13188 8528 13419 8530
rect 13188 8472 13358 8528
rect 13414 8472 13419 8528
rect 13188 8470 13419 8472
rect 13188 8468 13194 8470
rect 13353 8467 13419 8470
rect 14089 8530 14155 8533
rect 16990 8530 17050 8606
rect 21541 8603 21607 8606
rect 14089 8528 17050 8530
rect 14089 8472 14094 8528
rect 14150 8472 17050 8528
rect 14089 8470 17050 8472
rect 18689 8530 18755 8533
rect 20713 8530 20779 8533
rect 18689 8528 20914 8530
rect 18689 8472 18694 8528
rect 18750 8472 20718 8528
rect 20774 8472 20914 8528
rect 18689 8470 20914 8472
rect 14089 8467 14155 8470
rect 18689 8467 18755 8470
rect 20713 8467 20779 8470
rect 0 8394 800 8424
rect 3417 8394 3483 8397
rect 0 8392 3483 8394
rect 0 8336 3422 8392
rect 3478 8336 3483 8392
rect 0 8334 3483 8336
rect 0 8304 800 8334
rect 3417 8331 3483 8334
rect 3918 8332 3924 8396
rect 3988 8332 3994 8396
rect 4613 8394 4679 8397
rect 10225 8394 10291 8397
rect 4613 8392 10291 8394
rect 4613 8336 4618 8392
rect 4674 8336 10230 8392
rect 10286 8336 10291 8392
rect 4613 8334 10291 8336
rect 1577 8258 1643 8261
rect 2630 8258 2636 8260
rect 1577 8256 2636 8258
rect 1577 8200 1582 8256
rect 1638 8200 2636 8256
rect 1577 8198 2636 8200
rect 1577 8195 1643 8198
rect 2630 8196 2636 8198
rect 2700 8196 2706 8260
rect 3926 8258 3986 8332
rect 4613 8331 4679 8334
rect 10225 8331 10291 8334
rect 10910 8332 10916 8396
rect 10980 8394 10986 8396
rect 14181 8394 14247 8397
rect 19333 8394 19399 8397
rect 10980 8392 19399 8394
rect 10980 8336 14186 8392
rect 14242 8336 19338 8392
rect 19394 8336 19399 8392
rect 10980 8334 19399 8336
rect 10980 8332 10986 8334
rect 14181 8331 14247 8334
rect 19333 8331 19399 8334
rect 19558 8332 19564 8396
rect 19628 8394 19634 8396
rect 20713 8394 20779 8397
rect 19628 8392 20779 8394
rect 19628 8336 20718 8392
rect 20774 8336 20779 8392
rect 19628 8334 20779 8336
rect 20854 8394 20914 8470
rect 22200 8394 23000 8424
rect 20854 8334 23000 8394
rect 19628 8332 19634 8334
rect 20713 8331 20779 8334
rect 22200 8304 23000 8334
rect 5073 8258 5139 8261
rect 5625 8258 5691 8261
rect 3926 8256 5691 8258
rect 3926 8200 5078 8256
rect 5134 8200 5630 8256
rect 5686 8200 5691 8256
rect 3926 8198 5691 8200
rect 5073 8195 5139 8198
rect 5625 8195 5691 8198
rect 5809 8258 5875 8261
rect 7414 8258 7420 8260
rect 5809 8256 7420 8258
rect 5809 8200 5814 8256
rect 5870 8200 7420 8256
rect 5809 8198 7420 8200
rect 5809 8195 5875 8198
rect 7414 8196 7420 8198
rect 7484 8196 7490 8260
rect 7833 8258 7899 8261
rect 8293 8258 8359 8261
rect 7833 8256 8359 8258
rect 7833 8200 7838 8256
rect 7894 8200 8298 8256
rect 8354 8200 8359 8256
rect 7833 8198 8359 8200
rect 7833 8195 7899 8198
rect 8293 8195 8359 8198
rect 9673 8258 9739 8261
rect 14733 8258 14799 8261
rect 15142 8258 15148 8260
rect 9673 8256 13002 8258
rect 9673 8200 9678 8256
rect 9734 8200 13002 8256
rect 9673 8198 13002 8200
rect 9673 8195 9739 8198
rect 3545 8192 3861 8193
rect 3545 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3861 8192
rect 3545 8127 3861 8128
rect 8743 8192 9059 8193
rect 8743 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9059 8192
rect 8743 8127 9059 8128
rect 3969 8122 4035 8125
rect 6637 8122 6703 8125
rect 3969 8120 6703 8122
rect 3969 8064 3974 8120
rect 4030 8064 6642 8120
rect 6698 8064 6703 8120
rect 3969 8062 6703 8064
rect 3969 8059 4035 8062
rect 6637 8059 6703 8062
rect 7005 8122 7071 8125
rect 8569 8122 8635 8125
rect 7005 8120 8635 8122
rect 7005 8064 7010 8120
rect 7066 8064 8574 8120
rect 8630 8064 8635 8120
rect 7005 8062 8635 8064
rect 7005 8059 7071 8062
rect 8569 8059 8635 8062
rect 10726 8060 10732 8124
rect 10796 8122 10802 8124
rect 12709 8122 12775 8125
rect 10796 8120 12775 8122
rect 10796 8064 12714 8120
rect 12770 8064 12775 8120
rect 10796 8062 12775 8064
rect 10796 8060 10802 8062
rect 12709 8059 12775 8062
rect 0 7986 800 8016
rect 3877 7986 3943 7989
rect 0 7984 3943 7986
rect 0 7928 3882 7984
rect 3938 7928 3943 7984
rect 0 7926 3943 7928
rect 0 7896 800 7926
rect 3877 7923 3943 7926
rect 4102 7924 4108 7988
rect 4172 7986 4178 7988
rect 4705 7986 4771 7989
rect 6085 7986 6151 7989
rect 4172 7984 6151 7986
rect 4172 7928 4710 7984
rect 4766 7928 6090 7984
rect 6146 7928 6151 7984
rect 4172 7926 6151 7928
rect 4172 7924 4178 7926
rect 4705 7923 4771 7926
rect 6085 7923 6151 7926
rect 6269 7986 6335 7989
rect 10409 7986 10475 7989
rect 6269 7984 10475 7986
rect 6269 7928 6274 7984
rect 6330 7928 10414 7984
rect 10470 7928 10475 7984
rect 6269 7926 10475 7928
rect 6269 7923 6335 7926
rect 10409 7923 10475 7926
rect 10910 7924 10916 7988
rect 10980 7986 10986 7988
rect 11605 7986 11671 7989
rect 12249 7986 12315 7989
rect 10980 7984 11671 7986
rect 10980 7928 11610 7984
rect 11666 7928 11671 7984
rect 10980 7926 11671 7928
rect 10980 7924 10986 7926
rect 11605 7923 11671 7926
rect 12022 7984 12315 7986
rect 12022 7928 12254 7984
rect 12310 7928 12315 7984
rect 12022 7926 12315 7928
rect 3785 7850 3851 7853
rect 12022 7850 12082 7926
rect 12249 7923 12315 7926
rect 3785 7848 12082 7850
rect 3785 7792 3790 7848
rect 3846 7792 12082 7848
rect 3785 7790 12082 7792
rect 3785 7787 3851 7790
rect 1761 7714 1827 7717
rect 5625 7714 5691 7717
rect 1761 7712 5691 7714
rect 1761 7656 1766 7712
rect 1822 7656 5630 7712
rect 5686 7656 5691 7712
rect 1761 7654 5691 7656
rect 1761 7651 1827 7654
rect 5625 7651 5691 7654
rect 6637 7714 6703 7717
rect 9949 7716 10015 7717
rect 9622 7714 9628 7716
rect 6637 7712 9628 7714
rect 6637 7656 6642 7712
rect 6698 7656 9628 7712
rect 6637 7654 9628 7656
rect 6637 7651 6703 7654
rect 9622 7652 9628 7654
rect 9692 7652 9698 7716
rect 9949 7714 9996 7716
rect 9904 7712 9996 7714
rect 9904 7656 9954 7712
rect 9904 7654 9996 7656
rect 9949 7652 9996 7654
rect 10060 7652 10066 7716
rect 12942 7714 13002 8198
rect 14733 8256 15148 8258
rect 14733 8200 14738 8256
rect 14794 8200 15148 8256
rect 14733 8198 15148 8200
rect 14733 8195 14799 8198
rect 15142 8196 15148 8198
rect 15212 8196 15218 8260
rect 16389 8258 16455 8261
rect 17350 8258 17356 8260
rect 16389 8256 17356 8258
rect 16389 8200 16394 8256
rect 16450 8200 17356 8256
rect 16389 8198 17356 8200
rect 16389 8195 16455 8198
rect 17350 8196 17356 8198
rect 17420 8196 17426 8260
rect 18270 8196 18276 8260
rect 18340 8258 18346 8260
rect 18505 8258 18571 8261
rect 18340 8256 18571 8258
rect 18340 8200 18510 8256
rect 18566 8200 18571 8256
rect 18340 8198 18571 8200
rect 18340 8196 18346 8198
rect 18505 8195 18571 8198
rect 13941 8192 14257 8193
rect 13941 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14257 8192
rect 13941 8127 14257 8128
rect 19139 8192 19455 8193
rect 19139 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19455 8192
rect 19139 8127 19455 8128
rect 14641 8122 14707 8125
rect 15561 8122 15627 8125
rect 18873 8122 18939 8125
rect 21725 8122 21791 8125
rect 14641 8120 15627 8122
rect 14641 8064 14646 8120
rect 14702 8064 15566 8120
rect 15622 8064 15627 8120
rect 14641 8062 15627 8064
rect 14641 8059 14707 8062
rect 15561 8059 15627 8062
rect 16806 8120 18939 8122
rect 16806 8064 18878 8120
rect 18934 8064 18939 8120
rect 16806 8062 18939 8064
rect 14457 7986 14523 7989
rect 16806 7986 16866 8062
rect 18873 8059 18939 8062
rect 19566 8120 21791 8122
rect 19566 8064 21730 8120
rect 21786 8064 21791 8120
rect 19566 8062 21791 8064
rect 14457 7984 16866 7986
rect 14457 7928 14462 7984
rect 14518 7928 16866 7984
rect 14457 7926 16866 7928
rect 14457 7923 14523 7926
rect 17534 7924 17540 7988
rect 17604 7986 17610 7988
rect 18137 7986 18203 7989
rect 19566 7986 19626 8062
rect 21725 8059 21791 8062
rect 22200 7986 23000 8016
rect 17604 7984 19626 7986
rect 17604 7928 18142 7984
rect 18198 7928 19626 7984
rect 17604 7926 19626 7928
rect 21452 7926 23000 7986
rect 17604 7924 17610 7926
rect 18137 7923 18203 7926
rect 14406 7788 14412 7852
rect 14476 7850 14482 7852
rect 14917 7850 14983 7853
rect 14476 7848 14983 7850
rect 14476 7792 14922 7848
rect 14978 7792 14983 7848
rect 14476 7790 14983 7792
rect 14476 7788 14482 7790
rect 14917 7787 14983 7790
rect 16113 7850 16179 7853
rect 17585 7850 17651 7853
rect 21081 7850 21147 7853
rect 16113 7848 21147 7850
rect 16113 7792 16118 7848
rect 16174 7792 17590 7848
rect 17646 7792 21086 7848
rect 21142 7792 21147 7848
rect 16113 7790 21147 7792
rect 16113 7787 16179 7790
rect 17585 7787 17651 7790
rect 21081 7787 21147 7790
rect 16389 7714 16455 7717
rect 12942 7712 16455 7714
rect 12942 7656 16394 7712
rect 16450 7656 16455 7712
rect 12942 7654 16455 7656
rect 9949 7651 10015 7652
rect 16389 7651 16455 7654
rect 17309 7714 17375 7717
rect 20110 7714 20116 7716
rect 17309 7712 20116 7714
rect 17309 7656 17314 7712
rect 17370 7656 20116 7712
rect 17309 7654 20116 7656
rect 17309 7651 17375 7654
rect 20110 7652 20116 7654
rect 20180 7714 20186 7716
rect 21081 7714 21147 7717
rect 20180 7712 21147 7714
rect 20180 7656 21086 7712
rect 21142 7656 21147 7712
rect 20180 7654 21147 7656
rect 20180 7652 20186 7654
rect 21081 7651 21147 7654
rect 6144 7648 6460 7649
rect 0 7578 800 7608
rect 6144 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6460 7648
rect 6144 7583 6460 7584
rect 11342 7648 11658 7649
rect 11342 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11658 7648
rect 11342 7583 11658 7584
rect 16540 7648 16856 7649
rect 16540 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16856 7648
rect 16540 7583 16856 7584
rect 21452 7581 21512 7926
rect 22200 7896 23000 7926
rect 21738 7648 22054 7649
rect 21738 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22054 7648
rect 21738 7583 22054 7584
rect 3509 7578 3575 7581
rect 5441 7578 5507 7581
rect 10777 7578 10843 7581
rect 0 7576 3575 7578
rect 0 7520 3514 7576
rect 3570 7520 3575 7576
rect 0 7518 3575 7520
rect 0 7488 800 7518
rect 3509 7515 3575 7518
rect 4340 7576 5507 7578
rect 4340 7520 5446 7576
rect 5502 7520 5507 7576
rect 4340 7518 5507 7520
rect 2037 7442 2103 7445
rect 4340 7442 4400 7518
rect 5441 7515 5507 7518
rect 6548 7576 10843 7578
rect 6548 7520 10782 7576
rect 10838 7520 10843 7576
rect 6548 7518 10843 7520
rect 2037 7440 4400 7442
rect 2037 7384 2042 7440
rect 2098 7384 4400 7440
rect 2037 7382 4400 7384
rect 4705 7442 4771 7445
rect 6548 7442 6608 7518
rect 10777 7515 10843 7518
rect 13813 7578 13879 7581
rect 15469 7578 15535 7581
rect 13813 7576 15535 7578
rect 13813 7520 13818 7576
rect 13874 7520 15474 7576
rect 15530 7520 15535 7576
rect 13813 7518 15535 7520
rect 13813 7515 13879 7518
rect 15469 7515 15535 7518
rect 18045 7578 18111 7581
rect 21449 7578 21515 7581
rect 22200 7578 23000 7608
rect 18045 7576 21515 7578
rect 18045 7520 18050 7576
rect 18106 7520 21454 7576
rect 21510 7520 21515 7576
rect 18045 7518 21515 7520
rect 18045 7515 18111 7518
rect 21449 7515 21515 7518
rect 22142 7488 23000 7578
rect 10041 7442 10107 7445
rect 4705 7440 6608 7442
rect 4705 7384 4710 7440
rect 4766 7384 6608 7440
rect 4705 7382 6608 7384
rect 6870 7440 10107 7442
rect 6870 7384 10046 7440
rect 10102 7384 10107 7440
rect 6870 7382 10107 7384
rect 2037 7379 2103 7382
rect 4705 7379 4771 7382
rect 2497 7306 2563 7309
rect 6637 7306 6703 7309
rect 2497 7304 6703 7306
rect 2497 7248 2502 7304
rect 2558 7248 6642 7304
rect 6698 7248 6703 7304
rect 2497 7246 6703 7248
rect 2497 7243 2563 7246
rect 6637 7243 6703 7246
rect 0 7170 800 7200
rect 1485 7170 1551 7173
rect 6870 7170 6930 7382
rect 10041 7379 10107 7382
rect 10685 7442 10751 7445
rect 19609 7442 19675 7445
rect 10685 7440 19675 7442
rect 10685 7384 10690 7440
rect 10746 7384 19614 7440
rect 19670 7384 19675 7440
rect 10685 7382 19675 7384
rect 10685 7379 10751 7382
rect 19609 7379 19675 7382
rect 20253 7442 20319 7445
rect 22142 7442 22202 7488
rect 20253 7440 22202 7442
rect 20253 7384 20258 7440
rect 20314 7384 22202 7440
rect 20253 7382 22202 7384
rect 20253 7379 20319 7382
rect 7465 7306 7531 7309
rect 12157 7306 12223 7309
rect 7465 7304 12223 7306
rect 7465 7248 7470 7304
rect 7526 7248 12162 7304
rect 12218 7248 12223 7304
rect 7465 7246 12223 7248
rect 7465 7243 7531 7246
rect 12157 7243 12223 7246
rect 13629 7306 13695 7309
rect 15377 7306 15443 7309
rect 13629 7304 15443 7306
rect 13629 7248 13634 7304
rect 13690 7248 15382 7304
rect 15438 7248 15443 7304
rect 13629 7246 15443 7248
rect 13629 7243 13695 7246
rect 15377 7243 15443 7246
rect 16021 7306 16087 7309
rect 17125 7306 17191 7309
rect 20897 7306 20963 7309
rect 16021 7304 16452 7306
rect 16021 7248 16026 7304
rect 16082 7248 16452 7304
rect 16021 7246 16452 7248
rect 16021 7243 16087 7246
rect 0 7168 1551 7170
rect 0 7112 1490 7168
rect 1546 7112 1551 7168
rect 0 7110 1551 7112
rect 0 7080 800 7110
rect 1485 7107 1551 7110
rect 5398 7110 6930 7170
rect 10777 7170 10843 7173
rect 12801 7170 12867 7173
rect 10777 7168 12867 7170
rect 10777 7112 10782 7168
rect 10838 7112 12806 7168
rect 12862 7112 12867 7168
rect 10777 7110 12867 7112
rect 3545 7104 3861 7105
rect 3545 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3861 7104
rect 3545 7039 3861 7040
rect 4429 7036 4495 7037
rect 4429 7034 4476 7036
rect 4384 7032 4476 7034
rect 4384 6976 4434 7032
rect 4384 6974 4476 6976
rect 4429 6972 4476 6974
rect 4540 6972 4546 7036
rect 4429 6971 4495 6972
rect 5398 6901 5458 7110
rect 10777 7107 10843 7110
rect 12801 7107 12867 7110
rect 16062 7108 16068 7172
rect 16132 7170 16138 7172
rect 16205 7170 16271 7173
rect 16132 7168 16271 7170
rect 16132 7112 16210 7168
rect 16266 7112 16271 7168
rect 16132 7110 16271 7112
rect 16392 7170 16452 7246
rect 17125 7304 20963 7306
rect 17125 7248 17130 7304
rect 17186 7248 20902 7304
rect 20958 7248 20963 7304
rect 17125 7246 20963 7248
rect 17125 7243 17191 7246
rect 20897 7243 20963 7246
rect 19701 7170 19767 7173
rect 21449 7170 21515 7173
rect 22200 7170 23000 7200
rect 16392 7110 19074 7170
rect 16132 7108 16138 7110
rect 16205 7107 16271 7110
rect 8743 7104 9059 7105
rect 8743 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9059 7104
rect 8743 7039 9059 7040
rect 13941 7104 14257 7105
rect 13941 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14257 7104
rect 13941 7039 14257 7040
rect 8017 7034 8083 7037
rect 8150 7034 8156 7036
rect 8017 7032 8156 7034
rect 8017 6976 8022 7032
rect 8078 6976 8156 7032
rect 8017 6974 8156 6976
rect 8017 6971 8083 6974
rect 8150 6972 8156 6974
rect 8220 6972 8226 7036
rect 10409 7034 10475 7037
rect 11973 7036 12039 7037
rect 11973 7034 12020 7036
rect 10409 7032 12020 7034
rect 10409 6976 10414 7032
rect 10470 6976 11978 7032
rect 10409 6974 12020 6976
rect 10409 6971 10475 6974
rect 11973 6972 12020 6974
rect 12084 6972 12090 7036
rect 12801 7034 12867 7037
rect 13813 7034 13879 7037
rect 12801 7032 13879 7034
rect 12801 6976 12806 7032
rect 12862 6976 13818 7032
rect 13874 6976 13879 7032
rect 12801 6974 13879 6976
rect 11973 6971 12039 6972
rect 12801 6971 12867 6974
rect 13813 6971 13879 6974
rect 15561 7034 15627 7037
rect 18045 7034 18111 7037
rect 15561 7032 18111 7034
rect 15561 6976 15566 7032
rect 15622 6976 18050 7032
rect 18106 6976 18111 7032
rect 15561 6974 18111 6976
rect 15561 6971 15627 6974
rect 18045 6971 18111 6974
rect 19014 6932 19074 7110
rect 19701 7168 23000 7170
rect 19701 7112 19706 7168
rect 19762 7112 21454 7168
rect 21510 7112 23000 7168
rect 19701 7110 23000 7112
rect 19701 7107 19767 7110
rect 21449 7107 21515 7110
rect 19139 7104 19455 7105
rect 19139 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19455 7104
rect 22200 7080 23000 7110
rect 19139 7039 19455 7040
rect 2865 6898 2931 6901
rect 4102 6898 4108 6900
rect 2865 6896 4108 6898
rect 2865 6840 2870 6896
rect 2926 6840 4108 6896
rect 2865 6838 4108 6840
rect 2865 6835 2931 6838
rect 4102 6836 4108 6838
rect 4172 6836 4178 6900
rect 5349 6896 5458 6901
rect 5349 6840 5354 6896
rect 5410 6840 5458 6896
rect 5349 6838 5458 6840
rect 5349 6835 5415 6838
rect 5574 6836 5580 6900
rect 5644 6898 5650 6900
rect 6453 6898 6519 6901
rect 5644 6896 6519 6898
rect 5644 6840 6458 6896
rect 6514 6840 6519 6896
rect 5644 6838 6519 6840
rect 5644 6836 5650 6838
rect 6453 6835 6519 6838
rect 6637 6898 6703 6901
rect 7782 6898 7788 6900
rect 6637 6896 7788 6898
rect 6637 6840 6642 6896
rect 6698 6840 7788 6896
rect 6637 6838 7788 6840
rect 6637 6835 6703 6838
rect 7782 6836 7788 6838
rect 7852 6836 7858 6900
rect 8150 6836 8156 6900
rect 8220 6898 8226 6900
rect 8518 6898 8524 6900
rect 8220 6838 8524 6898
rect 8220 6836 8226 6838
rect 8518 6836 8524 6838
rect 8588 6836 8594 6900
rect 10317 6898 10383 6901
rect 10317 6896 12450 6898
rect 10317 6840 10322 6896
rect 10378 6840 12450 6896
rect 10317 6838 12450 6840
rect 10317 6835 10383 6838
rect 0 6762 800 6792
rect 2129 6762 2195 6765
rect 0 6760 2195 6762
rect 0 6704 2134 6760
rect 2190 6704 2195 6760
rect 0 6702 2195 6704
rect 0 6672 800 6702
rect 2129 6699 2195 6702
rect 2589 6762 2655 6765
rect 3141 6762 3207 6765
rect 11329 6762 11395 6765
rect 12390 6762 12450 6838
rect 14958 6836 14964 6900
rect 15028 6898 15034 6900
rect 15101 6898 15167 6901
rect 15028 6896 15167 6898
rect 15028 6840 15106 6896
rect 15162 6840 15167 6896
rect 15028 6838 15167 6840
rect 15028 6836 15034 6838
rect 15101 6835 15167 6838
rect 17718 6836 17724 6900
rect 17788 6898 17794 6900
rect 17953 6898 18019 6901
rect 17788 6896 18019 6898
rect 17788 6840 17958 6896
rect 18014 6840 18019 6896
rect 19014 6898 19488 6932
rect 20253 6898 20319 6901
rect 19014 6896 20319 6898
rect 19014 6872 20258 6896
rect 17788 6838 18019 6840
rect 19428 6840 20258 6872
rect 20314 6840 20319 6896
rect 19428 6838 20319 6840
rect 17788 6836 17794 6838
rect 17953 6835 18019 6838
rect 20253 6835 20319 6838
rect 19517 6762 19583 6765
rect 20621 6762 20687 6765
rect 22200 6762 23000 6792
rect 2589 6760 2790 6762
rect 2589 6704 2594 6760
rect 2650 6704 2790 6760
rect 2589 6702 2790 6704
rect 2589 6699 2655 6702
rect 0 6354 800 6384
rect 933 6354 999 6357
rect 0 6352 999 6354
rect 0 6296 938 6352
rect 994 6296 999 6352
rect 0 6294 999 6296
rect 2730 6354 2790 6702
rect 3141 6760 11898 6762
rect 3141 6704 3146 6760
rect 3202 6704 11334 6760
rect 11390 6704 11898 6760
rect 3141 6702 11898 6704
rect 12390 6702 19350 6762
rect 3141 6699 3207 6702
rect 11329 6699 11395 6702
rect 3366 6564 3372 6628
rect 3436 6626 3442 6628
rect 5441 6626 5507 6629
rect 3436 6624 5507 6626
rect 3436 6568 5446 6624
rect 5502 6568 5507 6624
rect 3436 6566 5507 6568
rect 3436 6564 3442 6566
rect 5441 6563 5507 6566
rect 7598 6564 7604 6628
rect 7668 6626 7674 6628
rect 8293 6626 8359 6629
rect 10961 6626 11027 6629
rect 7668 6624 11027 6626
rect 7668 6568 8298 6624
rect 8354 6568 10966 6624
rect 11022 6568 11027 6624
rect 7668 6566 11027 6568
rect 7668 6564 7674 6566
rect 8293 6563 8359 6566
rect 10961 6563 11027 6566
rect 6144 6560 6460 6561
rect 6144 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6460 6560
rect 6144 6495 6460 6496
rect 11342 6560 11658 6561
rect 11342 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11658 6560
rect 11342 6495 11658 6496
rect 3141 6490 3207 6493
rect 5758 6490 5764 6492
rect 3141 6488 5764 6490
rect 3141 6432 3146 6488
rect 3202 6432 5764 6488
rect 3141 6430 5764 6432
rect 3141 6427 3207 6430
rect 5758 6428 5764 6430
rect 5828 6428 5834 6492
rect 7005 6490 7071 6493
rect 10869 6490 10935 6493
rect 7005 6488 10935 6490
rect 7005 6432 7010 6488
rect 7066 6432 10874 6488
rect 10930 6432 10935 6488
rect 7005 6430 10935 6432
rect 11838 6490 11898 6702
rect 12985 6626 13051 6629
rect 15878 6626 15884 6628
rect 12985 6624 15884 6626
rect 12985 6568 12990 6624
rect 13046 6568 15884 6624
rect 12985 6566 15884 6568
rect 12985 6563 13051 6566
rect 15878 6564 15884 6566
rect 15948 6564 15954 6628
rect 17033 6626 17099 6629
rect 18873 6626 18939 6629
rect 17033 6624 18939 6626
rect 17033 6568 17038 6624
rect 17094 6568 18878 6624
rect 18934 6568 18939 6624
rect 17033 6566 18939 6568
rect 19290 6626 19350 6702
rect 19517 6760 23000 6762
rect 19517 6704 19522 6760
rect 19578 6704 20626 6760
rect 20682 6704 23000 6760
rect 19517 6702 23000 6704
rect 19517 6699 19583 6702
rect 20621 6699 20687 6702
rect 22200 6672 23000 6702
rect 20253 6626 20319 6629
rect 19290 6624 20319 6626
rect 19290 6568 20258 6624
rect 20314 6568 20319 6624
rect 19290 6566 20319 6568
rect 17033 6563 17099 6566
rect 18873 6563 18939 6566
rect 20253 6563 20319 6566
rect 16540 6560 16856 6561
rect 16540 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16856 6560
rect 16540 6495 16856 6496
rect 21738 6560 22054 6561
rect 21738 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22054 6560
rect 21738 6495 22054 6496
rect 15929 6490 15995 6493
rect 11838 6488 15995 6490
rect 11838 6432 15934 6488
rect 15990 6432 15995 6488
rect 11838 6430 15995 6432
rect 7005 6427 7071 6430
rect 10869 6427 10935 6430
rect 15929 6427 15995 6430
rect 17953 6490 18019 6493
rect 20662 6490 20668 6492
rect 17953 6488 20668 6490
rect 17953 6432 17958 6488
rect 18014 6432 20668 6488
rect 17953 6430 20668 6432
rect 17953 6427 18019 6430
rect 20662 6428 20668 6430
rect 20732 6428 20738 6492
rect 6637 6354 6703 6357
rect 8518 6354 8524 6356
rect 2730 6294 6562 6354
rect 0 6264 800 6294
rect 933 6291 999 6294
rect 3141 6218 3207 6221
rect 3141 6216 4216 6218
rect 3141 6160 3146 6216
rect 3202 6160 4216 6216
rect 3141 6158 4216 6160
rect 3141 6155 3207 6158
rect 4156 6082 4216 6158
rect 4286 6156 4292 6220
rect 4356 6218 4362 6220
rect 5349 6218 5415 6221
rect 4356 6216 5415 6218
rect 4356 6160 5354 6216
rect 5410 6160 5415 6216
rect 4356 6158 5415 6160
rect 4356 6156 4362 6158
rect 5349 6155 5415 6158
rect 5758 6156 5764 6220
rect 5828 6218 5834 6220
rect 6361 6218 6427 6221
rect 5828 6216 6427 6218
rect 5828 6160 6366 6216
rect 6422 6160 6427 6216
rect 5828 6158 6427 6160
rect 6502 6218 6562 6294
rect 6637 6352 8524 6354
rect 6637 6296 6642 6352
rect 6698 6296 8524 6352
rect 6637 6294 8524 6296
rect 6637 6291 6703 6294
rect 8518 6292 8524 6294
rect 8588 6292 8594 6356
rect 8845 6354 8911 6357
rect 9254 6354 9260 6356
rect 8845 6352 9260 6354
rect 8845 6296 8850 6352
rect 8906 6296 9260 6352
rect 8845 6294 9260 6296
rect 8845 6291 8911 6294
rect 9254 6292 9260 6294
rect 9324 6292 9330 6356
rect 10501 6354 10567 6357
rect 9630 6352 10567 6354
rect 9630 6296 10506 6352
rect 10562 6296 10567 6352
rect 9630 6294 10567 6296
rect 9630 6218 9690 6294
rect 10501 6291 10567 6294
rect 12750 6292 12756 6356
rect 12820 6354 12826 6356
rect 13670 6354 13676 6356
rect 12820 6294 13676 6354
rect 12820 6292 12826 6294
rect 13670 6292 13676 6294
rect 13740 6354 13746 6356
rect 20253 6354 20319 6357
rect 22200 6354 23000 6384
rect 13740 6294 19810 6354
rect 13740 6292 13746 6294
rect 19750 6221 19810 6294
rect 20253 6352 23000 6354
rect 20253 6296 20258 6352
rect 20314 6296 23000 6352
rect 20253 6294 23000 6296
rect 20253 6291 20319 6294
rect 21452 6221 21512 6294
rect 22200 6264 23000 6294
rect 6502 6158 9690 6218
rect 10317 6218 10383 6221
rect 11145 6218 11211 6221
rect 11605 6218 11671 6221
rect 10317 6216 11671 6218
rect 10317 6160 10322 6216
rect 10378 6160 11150 6216
rect 11206 6160 11610 6216
rect 11666 6160 11671 6216
rect 10317 6158 11671 6160
rect 5828 6156 5834 6158
rect 6361 6155 6427 6158
rect 10317 6155 10383 6158
rect 11145 6155 11211 6158
rect 11605 6155 11671 6158
rect 11881 6218 11947 6221
rect 19558 6218 19564 6220
rect 11881 6216 19564 6218
rect 11881 6160 11886 6216
rect 11942 6160 19564 6216
rect 11881 6158 19564 6160
rect 11881 6155 11947 6158
rect 19558 6156 19564 6158
rect 19628 6156 19634 6220
rect 19701 6216 19810 6221
rect 20713 6220 20779 6221
rect 19701 6160 19706 6216
rect 19762 6160 19810 6216
rect 19701 6158 19810 6160
rect 19701 6155 19767 6158
rect 20662 6156 20668 6220
rect 20732 6218 20779 6220
rect 20732 6216 20824 6218
rect 20774 6160 20824 6216
rect 20732 6158 20824 6160
rect 21449 6216 21515 6221
rect 21449 6160 21454 6216
rect 21510 6160 21515 6216
rect 20732 6156 20779 6158
rect 20713 6155 20779 6156
rect 21449 6155 21515 6160
rect 8017 6082 8083 6085
rect 9990 6082 9996 6084
rect 4156 6080 8083 6082
rect 4156 6024 8022 6080
rect 8078 6024 8083 6080
rect 4156 6022 8083 6024
rect 8017 6019 8083 6022
rect 9630 6022 9996 6082
rect 3545 6016 3861 6017
rect 0 5946 800 5976
rect 3545 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3861 6016
rect 3545 5951 3861 5952
rect 8743 6016 9059 6017
rect 8743 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9059 6016
rect 8743 5951 9059 5952
rect 1158 5946 1164 5948
rect 0 5886 1164 5946
rect 0 5856 800 5886
rect 1158 5884 1164 5886
rect 1228 5946 1234 5948
rect 2773 5946 2839 5949
rect 1228 5944 2839 5946
rect 1228 5888 2778 5944
rect 2834 5888 2839 5944
rect 1228 5886 2839 5888
rect 1228 5884 1234 5886
rect 2773 5883 2839 5886
rect 4153 5946 4219 5949
rect 4797 5946 4863 5949
rect 4153 5944 4863 5946
rect 4153 5888 4158 5944
rect 4214 5888 4802 5944
rect 4858 5888 4863 5944
rect 4153 5886 4863 5888
rect 4153 5883 4219 5886
rect 4797 5883 4863 5886
rect 5901 5946 5967 5949
rect 6678 5946 6684 5948
rect 5901 5944 6684 5946
rect 5901 5888 5906 5944
rect 5962 5888 6684 5944
rect 5901 5886 6684 5888
rect 5901 5883 5967 5886
rect 6678 5884 6684 5886
rect 6748 5884 6754 5948
rect 5441 5810 5507 5813
rect 2730 5808 5507 5810
rect 2730 5752 5446 5808
rect 5502 5752 5507 5808
rect 2730 5750 5507 5752
rect 2497 5674 2563 5677
rect 2730 5674 2790 5750
rect 5441 5747 5507 5750
rect 6453 5810 6519 5813
rect 9630 5810 9690 6022
rect 9990 6020 9996 6022
rect 10060 6082 10066 6084
rect 11237 6082 11303 6085
rect 10060 6080 11303 6082
rect 10060 6024 11242 6080
rect 11298 6024 11303 6080
rect 10060 6022 11303 6024
rect 10060 6020 10066 6022
rect 11237 6019 11303 6022
rect 11605 6082 11671 6085
rect 12566 6082 12572 6084
rect 11605 6080 12572 6082
rect 11605 6024 11610 6080
rect 11666 6024 12572 6080
rect 11605 6022 12572 6024
rect 11605 6019 11671 6022
rect 12566 6020 12572 6022
rect 12636 6082 12642 6084
rect 12893 6082 12959 6085
rect 12636 6080 12959 6082
rect 12636 6024 12898 6080
rect 12954 6024 12959 6080
rect 12636 6022 12959 6024
rect 12636 6020 12642 6022
rect 12893 6019 12959 6022
rect 13941 6016 14257 6017
rect 13941 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14257 6016
rect 13941 5951 14257 5952
rect 19139 6016 19455 6017
rect 19139 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19455 6016
rect 19139 5951 19455 5952
rect 10961 5946 11027 5949
rect 11329 5946 11395 5949
rect 11881 5946 11947 5949
rect 22200 5946 23000 5976
rect 10961 5944 11162 5946
rect 10961 5888 10966 5944
rect 11022 5888 11162 5944
rect 10961 5886 11162 5888
rect 10961 5883 11027 5886
rect 6453 5808 9690 5810
rect 6453 5752 6458 5808
rect 6514 5752 9690 5808
rect 6453 5750 9690 5752
rect 6453 5747 6519 5750
rect 2497 5672 2790 5674
rect 2497 5616 2502 5672
rect 2558 5616 2790 5672
rect 2497 5614 2790 5616
rect 3877 5674 3943 5677
rect 4613 5674 4679 5677
rect 3877 5672 4679 5674
rect 3877 5616 3882 5672
rect 3938 5616 4618 5672
rect 4674 5616 4679 5672
rect 3877 5614 4679 5616
rect 2497 5611 2563 5614
rect 3877 5611 3943 5614
rect 4613 5611 4679 5614
rect 5574 5612 5580 5676
rect 5644 5674 5650 5676
rect 5717 5674 5783 5677
rect 5644 5672 5783 5674
rect 5644 5616 5722 5672
rect 5778 5616 5783 5672
rect 5644 5614 5783 5616
rect 5644 5612 5650 5614
rect 5717 5611 5783 5614
rect 6269 5674 6335 5677
rect 6862 5674 6868 5676
rect 6269 5672 6868 5674
rect 6269 5616 6274 5672
rect 6330 5616 6868 5672
rect 6269 5614 6868 5616
rect 6269 5611 6335 5614
rect 6862 5612 6868 5614
rect 6932 5612 6938 5676
rect 8937 5674 9003 5677
rect 7054 5672 9003 5674
rect 7054 5616 8942 5672
rect 8998 5616 9003 5672
rect 7054 5614 9003 5616
rect 11102 5674 11162 5886
rect 11329 5944 11947 5946
rect 11329 5888 11334 5944
rect 11390 5888 11886 5944
rect 11942 5888 11947 5944
rect 11329 5886 11947 5888
rect 11329 5883 11395 5886
rect 11881 5883 11947 5886
rect 19934 5886 23000 5946
rect 11973 5810 12039 5813
rect 12750 5810 12756 5812
rect 11973 5808 12756 5810
rect 11973 5752 11978 5808
rect 12034 5752 12756 5808
rect 11973 5750 12756 5752
rect 11973 5747 12039 5750
rect 12750 5748 12756 5750
rect 12820 5748 12826 5812
rect 12934 5748 12940 5812
rect 13004 5810 13010 5812
rect 13077 5810 13143 5813
rect 13004 5808 13143 5810
rect 13004 5752 13082 5808
rect 13138 5752 13143 5808
rect 13004 5750 13143 5752
rect 13004 5748 13010 5750
rect 13077 5747 13143 5750
rect 14181 5810 14247 5813
rect 17953 5810 18019 5813
rect 14181 5808 18019 5810
rect 14181 5752 14186 5808
rect 14242 5752 17958 5808
rect 18014 5752 18019 5808
rect 14181 5750 18019 5752
rect 14181 5747 14247 5750
rect 17953 5747 18019 5750
rect 18873 5810 18939 5813
rect 19934 5810 19994 5886
rect 22200 5856 23000 5886
rect 20161 5812 20227 5813
rect 20110 5810 20116 5812
rect 18873 5808 19994 5810
rect 18873 5752 18878 5808
rect 18934 5752 19994 5808
rect 18873 5750 19994 5752
rect 20070 5750 20116 5810
rect 20180 5808 20227 5812
rect 20222 5752 20227 5808
rect 18873 5747 18939 5750
rect 20110 5748 20116 5750
rect 20180 5748 20227 5752
rect 20161 5747 20227 5748
rect 20989 5810 21055 5813
rect 20989 5808 22064 5810
rect 20989 5752 20994 5808
rect 21050 5752 22064 5808
rect 20989 5750 22064 5752
rect 20989 5747 21055 5750
rect 18781 5674 18847 5677
rect 21265 5674 21331 5677
rect 11102 5672 18847 5674
rect 11102 5616 18786 5672
rect 18842 5616 18847 5672
rect 11102 5614 18847 5616
rect 0 5538 800 5568
rect 933 5538 999 5541
rect 0 5536 999 5538
rect 0 5480 938 5536
rect 994 5480 999 5536
rect 0 5478 999 5480
rect 0 5448 800 5478
rect 933 5475 999 5478
rect 2998 5476 3004 5540
rect 3068 5538 3074 5540
rect 5901 5538 5967 5541
rect 3068 5536 5967 5538
rect 3068 5480 5906 5536
rect 5962 5480 5967 5536
rect 3068 5478 5967 5480
rect 3068 5476 3074 5478
rect 5901 5475 5967 5478
rect 6144 5472 6460 5473
rect 6144 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6460 5472
rect 6144 5407 6460 5408
rect 7054 5405 7114 5614
rect 8937 5611 9003 5614
rect 18781 5611 18847 5614
rect 19014 5672 21331 5674
rect 19014 5616 21270 5672
rect 21326 5616 21331 5672
rect 19014 5614 21331 5616
rect 22004 5674 22064 5750
rect 22004 5614 22202 5674
rect 7281 5540 7347 5541
rect 7230 5538 7236 5540
rect 7190 5478 7236 5538
rect 7300 5536 7347 5540
rect 7342 5480 7347 5536
rect 7230 5476 7236 5478
rect 7300 5476 7347 5480
rect 7281 5475 7347 5476
rect 7833 5538 7899 5541
rect 7833 5536 9506 5538
rect 7833 5480 7838 5536
rect 7894 5480 9506 5536
rect 7833 5478 9506 5480
rect 7833 5475 7899 5478
rect 2814 5340 2820 5404
rect 2884 5402 2890 5404
rect 4061 5402 4127 5405
rect 2884 5400 4127 5402
rect 2884 5344 4066 5400
rect 4122 5344 4127 5400
rect 2884 5342 4127 5344
rect 2884 5340 2890 5342
rect 4061 5339 4127 5342
rect 4245 5402 4311 5405
rect 5625 5402 5691 5405
rect 7005 5404 7114 5405
rect 7005 5402 7052 5404
rect 4245 5400 5691 5402
rect 4245 5344 4250 5400
rect 4306 5344 5630 5400
rect 5686 5344 5691 5400
rect 4245 5342 5691 5344
rect 6960 5400 7052 5402
rect 6960 5344 7010 5400
rect 6960 5342 7052 5344
rect 4245 5339 4311 5342
rect 5625 5339 5691 5342
rect 7005 5340 7052 5342
rect 7116 5340 7122 5404
rect 7281 5402 7347 5405
rect 9213 5402 9279 5405
rect 7281 5400 9279 5402
rect 7281 5344 7286 5400
rect 7342 5344 9218 5400
rect 9274 5344 9279 5400
rect 7281 5342 9279 5344
rect 9446 5402 9506 5478
rect 9622 5476 9628 5540
rect 9692 5538 9698 5540
rect 10225 5538 10291 5541
rect 9692 5536 10291 5538
rect 9692 5480 10230 5536
rect 10286 5480 10291 5536
rect 9692 5478 10291 5480
rect 9692 5476 9698 5478
rect 10225 5475 10291 5478
rect 13353 5538 13419 5541
rect 16205 5538 16271 5541
rect 13353 5536 16271 5538
rect 13353 5480 13358 5536
rect 13414 5480 16210 5536
rect 16266 5480 16271 5536
rect 13353 5478 16271 5480
rect 13353 5475 13419 5478
rect 16205 5475 16271 5478
rect 17861 5538 17927 5541
rect 19014 5538 19074 5614
rect 21265 5611 21331 5614
rect 17861 5536 19074 5538
rect 17861 5480 17866 5536
rect 17922 5480 19074 5536
rect 17861 5478 19074 5480
rect 22142 5568 22202 5614
rect 22142 5478 23000 5568
rect 17861 5475 17927 5478
rect 11342 5472 11658 5473
rect 11342 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11658 5472
rect 11342 5407 11658 5408
rect 16540 5472 16856 5473
rect 16540 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16856 5472
rect 16540 5407 16856 5408
rect 21738 5472 22054 5473
rect 21738 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22054 5472
rect 22200 5448 23000 5478
rect 21738 5407 22054 5408
rect 10910 5402 10916 5404
rect 9446 5342 10916 5402
rect 7005 5339 7071 5340
rect 7281 5339 7347 5342
rect 9213 5339 9279 5342
rect 10910 5340 10916 5342
rect 10980 5340 10986 5404
rect 14457 5402 14523 5405
rect 12804 5400 14523 5402
rect 12804 5344 14462 5400
rect 14518 5344 14523 5400
rect 12804 5342 14523 5344
rect 3049 5266 3115 5269
rect 3182 5266 3188 5268
rect 3049 5264 3188 5266
rect 3049 5208 3054 5264
rect 3110 5208 3188 5264
rect 3049 5206 3188 5208
rect 3049 5203 3115 5206
rect 3182 5204 3188 5206
rect 3252 5204 3258 5268
rect 3325 5266 3391 5269
rect 6177 5266 6243 5269
rect 8150 5266 8156 5268
rect 3325 5264 6056 5266
rect 3325 5208 3330 5264
rect 3386 5208 6056 5264
rect 3325 5206 6056 5208
rect 3325 5203 3391 5206
rect 0 5130 800 5160
rect 1761 5130 1827 5133
rect 0 5128 1827 5130
rect 0 5072 1766 5128
rect 1822 5072 1827 5128
rect 0 5070 1827 5072
rect 0 5040 800 5070
rect 1761 5067 1827 5070
rect 1945 5130 2011 5133
rect 5809 5130 5875 5133
rect 1945 5128 5875 5130
rect 1945 5072 1950 5128
rect 2006 5072 5814 5128
rect 5870 5072 5875 5128
rect 1945 5070 5875 5072
rect 5996 5130 6056 5206
rect 6177 5264 8156 5266
rect 6177 5208 6182 5264
rect 6238 5208 8156 5264
rect 6177 5206 8156 5208
rect 6177 5203 6243 5206
rect 8150 5204 8156 5206
rect 8220 5204 8226 5268
rect 10133 5266 10199 5269
rect 12804 5266 12864 5342
rect 14457 5339 14523 5342
rect 10133 5264 12864 5266
rect 10133 5208 10138 5264
rect 10194 5208 12864 5264
rect 10133 5206 12864 5208
rect 12985 5266 13051 5269
rect 16573 5266 16639 5269
rect 12985 5264 16639 5266
rect 12985 5208 12990 5264
rect 13046 5208 16578 5264
rect 16634 5208 16639 5264
rect 12985 5206 16639 5208
rect 10133 5203 10199 5206
rect 12985 5203 13051 5206
rect 16573 5203 16639 5206
rect 18505 5266 18571 5269
rect 20989 5266 21055 5269
rect 18505 5264 21055 5266
rect 18505 5208 18510 5264
rect 18566 5208 20994 5264
rect 21050 5208 21055 5264
rect 18505 5206 21055 5208
rect 18505 5203 18571 5206
rect 20989 5203 21055 5206
rect 6821 5130 6887 5133
rect 13537 5130 13603 5133
rect 5996 5128 6887 5130
rect 5996 5072 6826 5128
rect 6882 5072 6887 5128
rect 5996 5070 6887 5072
rect 1945 5067 2011 5070
rect 5809 5067 5875 5070
rect 6821 5067 6887 5070
rect 7054 5128 13603 5130
rect 7054 5072 13542 5128
rect 13598 5072 13603 5128
rect 7054 5070 13603 5072
rect 5073 4996 5139 4997
rect 5022 4932 5028 4996
rect 5092 4994 5139 4996
rect 6269 4994 6335 4997
rect 7054 4994 7114 5070
rect 13537 5067 13603 5070
rect 16481 5130 16547 5133
rect 21725 5130 21791 5133
rect 16481 5128 21791 5130
rect 16481 5072 16486 5128
rect 16542 5072 21730 5128
rect 21786 5072 21791 5128
rect 16481 5070 21791 5072
rect 16481 5067 16547 5070
rect 21725 5067 21791 5070
rect 22001 5130 22067 5133
rect 22200 5130 23000 5160
rect 22001 5128 23000 5130
rect 22001 5072 22006 5128
rect 22062 5072 23000 5128
rect 22001 5070 23000 5072
rect 22001 5067 22067 5070
rect 22200 5040 23000 5070
rect 5092 4992 5184 4994
rect 5134 4936 5184 4992
rect 5092 4934 5184 4936
rect 6269 4992 7114 4994
rect 6269 4936 6274 4992
rect 6330 4936 7114 4992
rect 6269 4934 7114 4936
rect 5092 4932 5139 4934
rect 5073 4931 5139 4932
rect 6269 4931 6335 4934
rect 9438 4932 9444 4996
rect 9508 4994 9514 4996
rect 9581 4994 9647 4997
rect 9508 4992 9647 4994
rect 9508 4936 9586 4992
rect 9642 4936 9647 4992
rect 9508 4934 9647 4936
rect 9508 4932 9514 4934
rect 9581 4931 9647 4934
rect 9857 4994 9923 4997
rect 13813 4994 13879 4997
rect 9857 4992 13879 4994
rect 9857 4936 9862 4992
rect 9918 4936 13818 4992
rect 13874 4936 13879 4992
rect 9857 4934 13879 4936
rect 9857 4931 9923 4934
rect 13813 4931 13879 4934
rect 3545 4928 3861 4929
rect 3545 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3861 4928
rect 3545 4863 3861 4864
rect 8743 4928 9059 4929
rect 8743 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9059 4928
rect 8743 4863 9059 4864
rect 13941 4928 14257 4929
rect 13941 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14257 4928
rect 13941 4863 14257 4864
rect 19139 4928 19455 4929
rect 19139 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19455 4928
rect 19139 4863 19455 4864
rect 4981 4858 5047 4861
rect 5206 4858 5212 4860
rect 4981 4856 5212 4858
rect 4981 4800 4986 4856
rect 5042 4800 5212 4856
rect 4981 4798 5212 4800
rect 4981 4795 5047 4798
rect 5206 4796 5212 4798
rect 5276 4858 5282 4860
rect 5942 4858 5948 4860
rect 5276 4798 5948 4858
rect 5276 4796 5282 4798
rect 5942 4796 5948 4798
rect 6012 4858 6018 4860
rect 6269 4858 6335 4861
rect 6012 4856 6335 4858
rect 6012 4800 6274 4856
rect 6330 4800 6335 4856
rect 6012 4798 6335 4800
rect 6012 4796 6018 4798
rect 6269 4795 6335 4798
rect 12198 4796 12204 4860
rect 12268 4858 12274 4860
rect 12985 4858 13051 4861
rect 12268 4856 13051 4858
rect 12268 4800 12990 4856
rect 13046 4800 13051 4856
rect 12268 4798 13051 4800
rect 12268 4796 12274 4798
rect 12985 4795 13051 4798
rect 15326 4796 15332 4860
rect 15396 4858 15402 4860
rect 15396 4798 16314 4858
rect 15396 4796 15402 4798
rect 0 4722 800 4752
rect 1025 4722 1091 4725
rect 0 4720 1091 4722
rect 0 4664 1030 4720
rect 1086 4664 1091 4720
rect 0 4662 1091 4664
rect 0 4632 800 4662
rect 1025 4659 1091 4662
rect 2262 4660 2268 4724
rect 2332 4722 2338 4724
rect 2497 4722 2563 4725
rect 12433 4722 12499 4725
rect 2332 4720 12499 4722
rect 2332 4664 2502 4720
rect 2558 4664 12438 4720
rect 12494 4664 12499 4720
rect 2332 4662 12499 4664
rect 2332 4660 2338 4662
rect 2497 4659 2563 4662
rect 12433 4659 12499 4662
rect 12709 4722 12775 4725
rect 13721 4722 13787 4725
rect 14457 4724 14523 4725
rect 12709 4720 13787 4722
rect 12709 4664 12714 4720
rect 12770 4664 13726 4720
rect 13782 4664 13787 4720
rect 12709 4662 13787 4664
rect 12709 4659 12775 4662
rect 13721 4659 13787 4662
rect 14406 4660 14412 4724
rect 14476 4722 14523 4724
rect 16113 4722 16179 4725
rect 14476 4720 16179 4722
rect 14518 4664 16118 4720
rect 16174 4664 16179 4720
rect 14476 4662 16179 4664
rect 16254 4722 16314 4798
rect 20989 4722 21055 4725
rect 16254 4720 21055 4722
rect 16254 4664 20994 4720
rect 21050 4664 21055 4720
rect 16254 4662 21055 4664
rect 14476 4660 14523 4662
rect 14457 4659 14523 4660
rect 16113 4659 16179 4662
rect 20989 4659 21055 4662
rect 22001 4722 22067 4725
rect 22200 4722 23000 4752
rect 22001 4720 23000 4722
rect 22001 4664 22006 4720
rect 22062 4664 23000 4720
rect 22001 4662 23000 4664
rect 22001 4659 22067 4662
rect 22200 4632 23000 4662
rect 3877 4586 3943 4589
rect 5625 4586 5691 4589
rect 3877 4584 5691 4586
rect 3877 4528 3882 4584
rect 3938 4528 5630 4584
rect 5686 4528 5691 4584
rect 3877 4526 5691 4528
rect 3877 4523 3943 4526
rect 5625 4523 5691 4526
rect 5809 4586 5875 4589
rect 13118 4586 13124 4588
rect 5809 4584 13124 4586
rect 5809 4528 5814 4584
rect 5870 4528 13124 4584
rect 5809 4526 13124 4528
rect 5809 4523 5875 4526
rect 13118 4524 13124 4526
rect 13188 4586 13194 4588
rect 16757 4586 16823 4589
rect 13188 4584 16823 4586
rect 13188 4528 16762 4584
rect 16818 4528 16823 4584
rect 13188 4526 16823 4528
rect 13188 4524 13194 4526
rect 16757 4523 16823 4526
rect 17217 4586 17283 4589
rect 17902 4586 17908 4588
rect 17217 4584 17908 4586
rect 17217 4528 17222 4584
rect 17278 4528 17908 4584
rect 17217 4526 17908 4528
rect 17217 4523 17283 4526
rect 17902 4524 17908 4526
rect 17972 4524 17978 4588
rect 2865 4450 2931 4453
rect 4286 4450 4292 4452
rect 2865 4448 4292 4450
rect 2865 4392 2870 4448
rect 2926 4392 4292 4448
rect 2865 4390 4292 4392
rect 2865 4387 2931 4390
rect 4286 4388 4292 4390
rect 4356 4388 4362 4452
rect 5073 4450 5139 4453
rect 5901 4452 5967 4453
rect 5390 4450 5396 4452
rect 5073 4448 5396 4450
rect 5073 4392 5078 4448
rect 5134 4392 5396 4448
rect 5073 4390 5396 4392
rect 5073 4387 5139 4390
rect 5390 4388 5396 4390
rect 5460 4388 5466 4452
rect 5901 4448 5948 4452
rect 6012 4450 6018 4452
rect 7557 4450 7623 4453
rect 9029 4450 9095 4453
rect 5901 4392 5906 4448
rect 5901 4388 5948 4392
rect 6012 4390 6058 4450
rect 7557 4448 9095 4450
rect 7557 4392 7562 4448
rect 7618 4392 9034 4448
rect 9090 4392 9095 4448
rect 7557 4390 9095 4392
rect 6012 4388 6018 4390
rect 5901 4387 5967 4388
rect 7557 4387 7623 4390
rect 9029 4387 9095 4390
rect 9254 4388 9260 4452
rect 9324 4450 9330 4452
rect 9949 4450 10015 4453
rect 9324 4448 10015 4450
rect 9324 4392 9954 4448
rect 10010 4392 10015 4448
rect 9324 4390 10015 4392
rect 9324 4388 9330 4390
rect 9949 4387 10015 4390
rect 11973 4450 12039 4453
rect 13629 4450 13695 4453
rect 11973 4448 13695 4450
rect 11973 4392 11978 4448
rect 12034 4392 13634 4448
rect 13690 4392 13695 4448
rect 11973 4390 13695 4392
rect 11973 4387 12039 4390
rect 13629 4387 13695 4390
rect 14549 4450 14615 4453
rect 16297 4450 16363 4453
rect 14549 4448 16363 4450
rect 14549 4392 14554 4448
rect 14610 4392 16302 4448
rect 16358 4392 16363 4448
rect 14549 4390 16363 4392
rect 14549 4387 14615 4390
rect 16297 4387 16363 4390
rect 17769 4450 17835 4453
rect 18638 4450 18644 4452
rect 17769 4448 18644 4450
rect 17769 4392 17774 4448
rect 17830 4392 18644 4448
rect 17769 4390 18644 4392
rect 17769 4387 17835 4390
rect 18638 4388 18644 4390
rect 18708 4388 18714 4452
rect 6144 4384 6460 4385
rect 0 4314 800 4344
rect 6144 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6460 4384
rect 6144 4319 6460 4320
rect 11342 4384 11658 4385
rect 11342 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11658 4384
rect 11342 4319 11658 4320
rect 16540 4384 16856 4385
rect 16540 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16856 4384
rect 16540 4319 16856 4320
rect 21738 4384 22054 4385
rect 21738 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22054 4384
rect 21738 4319 22054 4320
rect 974 4314 980 4316
rect 0 4254 980 4314
rect 0 4224 800 4254
rect 974 4252 980 4254
rect 1044 4314 1050 4316
rect 1393 4314 1459 4317
rect 1761 4316 1827 4317
rect 1710 4314 1716 4316
rect 1044 4312 1459 4314
rect 1044 4256 1398 4312
rect 1454 4256 1459 4312
rect 1044 4254 1459 4256
rect 1634 4254 1716 4314
rect 1780 4314 1827 4316
rect 8477 4316 8543 4317
rect 8477 4314 8524 4316
rect 1780 4312 6010 4314
rect 1822 4256 6010 4312
rect 1044 4252 1050 4254
rect 1393 4251 1459 4254
rect 1710 4252 1716 4254
rect 1780 4254 6010 4256
rect 8396 4312 8524 4314
rect 8588 4314 8594 4316
rect 9029 4314 9095 4317
rect 8588 4312 9095 4314
rect 8396 4256 8482 4312
rect 8588 4256 9034 4312
rect 9090 4256 9095 4312
rect 8396 4254 8524 4256
rect 1780 4252 1827 4254
rect 1761 4251 1827 4252
rect 5950 4178 6010 4254
rect 8477 4252 8524 4254
rect 8588 4254 9095 4256
rect 8588 4252 8594 4254
rect 8477 4251 8543 4252
rect 9029 4251 9095 4254
rect 9438 4252 9444 4316
rect 9508 4314 9514 4316
rect 9581 4314 9647 4317
rect 9508 4312 9647 4314
rect 9508 4256 9586 4312
rect 9642 4256 9647 4312
rect 9508 4254 9647 4256
rect 9508 4252 9514 4254
rect 9581 4251 9647 4254
rect 11973 4314 12039 4317
rect 15009 4314 15075 4317
rect 22200 4314 23000 4344
rect 11973 4312 15075 4314
rect 11973 4256 11978 4312
rect 12034 4256 15014 4312
rect 15070 4256 15075 4312
rect 11973 4254 15075 4256
rect 11973 4251 12039 4254
rect 15009 4251 15075 4254
rect 22142 4224 23000 4314
rect 11881 4178 11947 4181
rect 5950 4176 11947 4178
rect 5950 4120 11886 4176
rect 11942 4120 11947 4176
rect 5950 4118 11947 4120
rect 11881 4115 11947 4118
rect 13537 4178 13603 4181
rect 15285 4178 15351 4181
rect 13537 4176 15351 4178
rect 13537 4120 13542 4176
rect 13598 4120 15290 4176
rect 15346 4120 15351 4176
rect 13537 4118 15351 4120
rect 13537 4115 13603 4118
rect 15285 4115 15351 4118
rect 16021 4178 16087 4181
rect 19149 4178 19215 4181
rect 16021 4176 19215 4178
rect 16021 4120 16026 4176
rect 16082 4120 19154 4176
rect 19210 4120 19215 4176
rect 16021 4118 19215 4120
rect 16021 4115 16087 4118
rect 19149 4115 19215 4118
rect 20805 4178 20871 4181
rect 22142 4178 22202 4224
rect 20805 4176 22202 4178
rect 20805 4120 20810 4176
rect 20866 4120 22202 4176
rect 20805 4118 22202 4120
rect 20805 4115 20871 4118
rect 5758 4042 5764 4044
rect 3420 3982 5764 4042
rect 0 3906 800 3936
rect 3420 3906 3480 3982
rect 5758 3980 5764 3982
rect 5828 3980 5834 4044
rect 6361 4042 6427 4045
rect 8334 4042 8340 4044
rect 6361 4040 8340 4042
rect 6361 3984 6366 4040
rect 6422 3984 8340 4040
rect 6361 3982 8340 3984
rect 6361 3979 6427 3982
rect 8334 3980 8340 3982
rect 8404 3980 8410 4044
rect 9029 4042 9095 4045
rect 15193 4042 15259 4045
rect 20989 4042 21055 4045
rect 9029 4040 14428 4042
rect 9029 3984 9034 4040
rect 9090 3984 14428 4040
rect 9029 3982 14428 3984
rect 9029 3979 9095 3982
rect 0 3846 3480 3906
rect 5993 3906 6059 3909
rect 6678 3906 6684 3908
rect 5993 3904 6684 3906
rect 5993 3848 5998 3904
rect 6054 3848 6684 3904
rect 5993 3846 6684 3848
rect 0 3816 800 3846
rect 5993 3843 6059 3846
rect 6678 3844 6684 3846
rect 6748 3844 6754 3908
rect 7097 3906 7163 3909
rect 7230 3906 7236 3908
rect 7097 3904 7236 3906
rect 7097 3848 7102 3904
rect 7158 3848 7236 3904
rect 7097 3846 7236 3848
rect 7097 3843 7163 3846
rect 7230 3844 7236 3846
rect 7300 3844 7306 3908
rect 14368 3906 14428 3982
rect 15193 4040 21055 4042
rect 15193 3984 15198 4040
rect 15254 3984 20994 4040
rect 21050 3984 21055 4040
rect 15193 3982 21055 3984
rect 15193 3979 15259 3982
rect 20989 3979 21055 3982
rect 15653 3906 15719 3909
rect 14368 3904 15719 3906
rect 14368 3848 15658 3904
rect 15714 3848 15719 3904
rect 14368 3846 15719 3848
rect 15653 3843 15719 3846
rect 19926 3844 19932 3908
rect 19996 3906 20002 3908
rect 20805 3906 20871 3909
rect 19996 3904 20871 3906
rect 19996 3848 20810 3904
rect 20866 3848 20871 3904
rect 19996 3846 20871 3848
rect 19996 3844 20002 3846
rect 20805 3843 20871 3846
rect 21265 3906 21331 3909
rect 22200 3906 23000 3936
rect 21265 3904 23000 3906
rect 21265 3848 21270 3904
rect 21326 3848 23000 3904
rect 21265 3846 23000 3848
rect 21265 3843 21331 3846
rect 3545 3840 3861 3841
rect 3545 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3861 3840
rect 3545 3775 3861 3776
rect 8743 3840 9059 3841
rect 8743 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9059 3840
rect 8743 3775 9059 3776
rect 13941 3840 14257 3841
rect 13941 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14257 3840
rect 13941 3775 14257 3776
rect 19139 3840 19455 3841
rect 19139 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19455 3840
rect 22200 3816 23000 3846
rect 19139 3775 19455 3776
rect 4705 3770 4771 3773
rect 6545 3770 6611 3773
rect 4705 3768 6611 3770
rect 4705 3712 4710 3768
rect 4766 3712 6550 3768
rect 6606 3712 6611 3768
rect 4705 3710 6611 3712
rect 4705 3707 4771 3710
rect 6545 3707 6611 3710
rect 10317 3770 10383 3773
rect 12525 3770 12591 3773
rect 10317 3768 12591 3770
rect 10317 3712 10322 3768
rect 10378 3712 12530 3768
rect 12586 3712 12591 3768
rect 10317 3710 12591 3712
rect 10317 3707 10383 3710
rect 12525 3707 12591 3710
rect 15009 3770 15075 3773
rect 17166 3770 17172 3772
rect 15009 3768 17172 3770
rect 15009 3712 15014 3768
rect 15070 3712 17172 3768
rect 15009 3710 17172 3712
rect 15009 3707 15075 3710
rect 17166 3708 17172 3710
rect 17236 3770 17242 3772
rect 17677 3770 17743 3773
rect 17236 3768 17743 3770
rect 17236 3712 17682 3768
rect 17738 3712 17743 3768
rect 17236 3710 17743 3712
rect 17236 3708 17242 3710
rect 17677 3707 17743 3710
rect 19742 3708 19748 3772
rect 19812 3770 19818 3772
rect 20345 3770 20411 3773
rect 19812 3768 20411 3770
rect 19812 3712 20350 3768
rect 20406 3712 20411 3768
rect 19812 3710 20411 3712
rect 19812 3708 19818 3710
rect 20345 3707 20411 3710
rect 1945 3634 2011 3637
rect 3417 3634 3483 3637
rect 1945 3632 3483 3634
rect 1945 3576 1950 3632
rect 2006 3576 3422 3632
rect 3478 3576 3483 3632
rect 1945 3574 3483 3576
rect 1945 3571 2011 3574
rect 3417 3571 3483 3574
rect 3785 3634 3851 3637
rect 4245 3634 4311 3637
rect 4797 3634 4863 3637
rect 3785 3632 4170 3634
rect 3785 3576 3790 3632
rect 3846 3576 4170 3632
rect 3785 3574 4170 3576
rect 3785 3571 3851 3574
rect 0 3498 800 3528
rect 3918 3498 3924 3500
rect 0 3438 3924 3498
rect 0 3408 800 3438
rect 3918 3436 3924 3438
rect 3988 3436 3994 3500
rect 4110 3498 4170 3574
rect 4245 3632 4863 3634
rect 4245 3576 4250 3632
rect 4306 3576 4802 3632
rect 4858 3576 4863 3632
rect 4245 3574 4863 3576
rect 4245 3571 4311 3574
rect 4797 3571 4863 3574
rect 6862 3572 6868 3636
rect 6932 3634 6938 3636
rect 9489 3634 9555 3637
rect 6932 3632 9555 3634
rect 6932 3576 9494 3632
rect 9550 3576 9555 3632
rect 6932 3574 9555 3576
rect 6932 3572 6938 3574
rect 9489 3571 9555 3574
rect 9857 3634 9923 3637
rect 12934 3634 12940 3636
rect 9857 3632 12940 3634
rect 9857 3576 9862 3632
rect 9918 3576 12940 3632
rect 9857 3574 12940 3576
rect 9857 3571 9923 3574
rect 12934 3572 12940 3574
rect 13004 3572 13010 3636
rect 13813 3634 13879 3637
rect 14733 3634 14799 3637
rect 13813 3632 14799 3634
rect 13813 3576 13818 3632
rect 13874 3576 14738 3632
rect 14794 3576 14799 3632
rect 13813 3574 14799 3576
rect 13813 3571 13879 3574
rect 14733 3571 14799 3574
rect 17309 3634 17375 3637
rect 17309 3632 21098 3634
rect 17309 3576 17314 3632
rect 17370 3576 21098 3632
rect 17309 3574 21098 3576
rect 17309 3571 17375 3574
rect 4110 3438 6608 3498
rect 933 3362 999 3365
rect 5349 3362 5415 3365
rect 6548 3362 6608 3438
rect 6678 3436 6684 3500
rect 6748 3498 6754 3500
rect 20805 3498 20871 3501
rect 6748 3496 20871 3498
rect 6748 3440 20810 3496
rect 20866 3440 20871 3496
rect 6748 3438 20871 3440
rect 21038 3498 21098 3574
rect 22200 3498 23000 3528
rect 21038 3438 23000 3498
rect 6748 3436 6754 3438
rect 20805 3435 20871 3438
rect 22200 3408 23000 3438
rect 6913 3362 6979 3365
rect 8109 3362 8175 3365
rect 9857 3362 9923 3365
rect 933 3360 5964 3362
rect 933 3304 938 3360
rect 994 3304 5354 3360
rect 5410 3304 5964 3360
rect 933 3302 5964 3304
rect 6548 3360 8175 3362
rect 6548 3304 6918 3360
rect 6974 3304 8114 3360
rect 8170 3304 8175 3360
rect 6548 3302 8175 3304
rect 933 3299 999 3302
rect 5349 3299 5415 3302
rect 3366 3226 3372 3228
rect 3190 3166 3372 3226
rect 0 3090 800 3120
rect 3190 3090 3250 3166
rect 3366 3164 3372 3166
rect 3436 3164 3442 3228
rect 3969 3226 4035 3229
rect 4654 3226 4660 3228
rect 3969 3224 4660 3226
rect 3969 3168 3974 3224
rect 4030 3168 4660 3224
rect 3969 3166 4660 3168
rect 3969 3163 4035 3166
rect 4654 3164 4660 3166
rect 4724 3164 4730 3228
rect 0 3030 3250 3090
rect 3417 3090 3483 3093
rect 3417 3088 4722 3090
rect 3417 3032 3422 3088
rect 3478 3032 4722 3088
rect 3417 3030 4722 3032
rect 0 3000 800 3030
rect 3417 3027 3483 3030
rect 2681 2954 2747 2957
rect 4429 2954 4495 2957
rect 2681 2952 4495 2954
rect 2681 2896 2686 2952
rect 2742 2896 4434 2952
rect 4490 2896 4495 2952
rect 2681 2894 4495 2896
rect 4662 2954 4722 3030
rect 5390 3028 5396 3092
rect 5460 3090 5466 3092
rect 5533 3090 5599 3093
rect 5460 3088 5599 3090
rect 5460 3032 5538 3088
rect 5594 3032 5599 3088
rect 5460 3030 5599 3032
rect 5904 3090 5964 3302
rect 6913 3299 6979 3302
rect 8109 3299 8175 3302
rect 9308 3360 9923 3362
rect 9308 3304 9862 3360
rect 9918 3304 9923 3360
rect 9308 3302 9923 3304
rect 6144 3296 6460 3297
rect 6144 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6460 3296
rect 6144 3231 6460 3232
rect 6821 3226 6887 3229
rect 6821 3224 7298 3226
rect 6821 3168 6826 3224
rect 6882 3168 7298 3224
rect 6821 3166 7298 3168
rect 6821 3163 6887 3166
rect 7005 3090 7071 3093
rect 5904 3088 7071 3090
rect 5904 3032 7010 3088
rect 7066 3032 7071 3088
rect 5904 3030 7071 3032
rect 7238 3090 7298 3166
rect 7414 3164 7420 3228
rect 7484 3226 7490 3228
rect 9308 3226 9368 3302
rect 9857 3299 9923 3302
rect 12341 3362 12407 3365
rect 15837 3362 15903 3365
rect 12341 3360 15903 3362
rect 12341 3304 12346 3360
rect 12402 3304 15842 3360
rect 15898 3304 15903 3360
rect 12341 3302 15903 3304
rect 12341 3299 12407 3302
rect 15837 3299 15903 3302
rect 17309 3364 17375 3365
rect 17309 3360 17356 3364
rect 17420 3362 17426 3364
rect 18597 3362 18663 3365
rect 21265 3362 21331 3365
rect 17309 3304 17314 3360
rect 17309 3300 17356 3304
rect 17420 3302 17466 3362
rect 18597 3360 21331 3362
rect 18597 3304 18602 3360
rect 18658 3304 21270 3360
rect 21326 3304 21331 3360
rect 18597 3302 21331 3304
rect 17420 3300 17426 3302
rect 17309 3299 17375 3300
rect 18597 3299 18663 3302
rect 21265 3299 21331 3302
rect 11342 3296 11658 3297
rect 11342 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11658 3296
rect 11342 3231 11658 3232
rect 16540 3296 16856 3297
rect 16540 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16856 3296
rect 16540 3231 16856 3232
rect 21738 3296 22054 3297
rect 21738 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22054 3296
rect 21738 3231 22054 3232
rect 7484 3166 9368 3226
rect 9489 3226 9555 3229
rect 11053 3226 11119 3229
rect 9489 3224 11119 3226
rect 9489 3168 9494 3224
rect 9550 3168 11058 3224
rect 11114 3168 11119 3224
rect 9489 3166 11119 3168
rect 7484 3164 7490 3166
rect 9489 3163 9555 3166
rect 11053 3163 11119 3166
rect 12433 3226 12499 3229
rect 14733 3226 14799 3229
rect 12433 3224 14799 3226
rect 12433 3168 12438 3224
rect 12494 3168 14738 3224
rect 14794 3168 14799 3224
rect 12433 3166 14799 3168
rect 12433 3163 12499 3166
rect 14733 3163 14799 3166
rect 17953 3226 18019 3229
rect 20713 3226 20779 3229
rect 17953 3224 20779 3226
rect 17953 3168 17958 3224
rect 18014 3168 20718 3224
rect 20774 3168 20779 3224
rect 17953 3166 20779 3168
rect 17953 3163 18019 3166
rect 20713 3163 20779 3166
rect 12709 3090 12775 3093
rect 7238 3088 12775 3090
rect 7238 3032 12714 3088
rect 12770 3032 12775 3088
rect 7238 3030 12775 3032
rect 5460 3028 5466 3030
rect 5533 3027 5599 3030
rect 7005 3027 7071 3030
rect 12709 3027 12775 3030
rect 13261 3090 13327 3093
rect 14825 3090 14891 3093
rect 13261 3088 14891 3090
rect 13261 3032 13266 3088
rect 13322 3032 14830 3088
rect 14886 3032 14891 3088
rect 13261 3030 14891 3032
rect 13261 3027 13327 3030
rect 14825 3027 14891 3030
rect 15878 3028 15884 3092
rect 15948 3090 15954 3092
rect 16757 3090 16823 3093
rect 16941 3092 17007 3093
rect 16941 3090 16988 3092
rect 15948 3088 16823 3090
rect 15948 3032 16762 3088
rect 16818 3032 16823 3088
rect 15948 3030 16823 3032
rect 16896 3088 16988 3090
rect 16896 3032 16946 3088
rect 16896 3030 16988 3032
rect 15948 3028 15954 3030
rect 16757 3027 16823 3030
rect 16941 3028 16988 3030
rect 17052 3028 17058 3092
rect 21541 3090 21607 3093
rect 22200 3090 23000 3120
rect 21541 3088 23000 3090
rect 21541 3032 21546 3088
rect 21602 3032 23000 3088
rect 21541 3030 23000 3032
rect 16941 3027 17007 3028
rect 21541 3027 21607 3030
rect 22200 3000 23000 3030
rect 7741 2954 7807 2957
rect 4662 2952 7807 2954
rect 4662 2896 7746 2952
rect 7802 2896 7807 2952
rect 4662 2894 7807 2896
rect 2681 2891 2747 2894
rect 4429 2891 4495 2894
rect 7741 2891 7807 2894
rect 7966 2892 7972 2956
rect 8036 2954 8042 2956
rect 12525 2954 12591 2957
rect 17769 2954 17835 2957
rect 20253 2954 20319 2957
rect 8036 2952 17835 2954
rect 8036 2896 12530 2952
rect 12586 2896 17774 2952
rect 17830 2896 17835 2952
rect 8036 2894 17835 2896
rect 8036 2892 8042 2894
rect 12525 2891 12591 2894
rect 17769 2891 17835 2894
rect 17910 2952 20319 2954
rect 17910 2896 20258 2952
rect 20314 2896 20319 2952
rect 17910 2894 20319 2896
rect 2998 2756 3004 2820
rect 3068 2818 3074 2820
rect 3366 2818 3372 2820
rect 3068 2758 3372 2818
rect 3068 2756 3074 2758
rect 3366 2756 3372 2758
rect 3436 2756 3442 2820
rect 3969 2818 4035 2821
rect 4613 2818 4679 2821
rect 3969 2816 4679 2818
rect 3969 2760 3974 2816
rect 4030 2760 4618 2816
rect 4674 2760 4679 2816
rect 3969 2758 4679 2760
rect 3969 2755 4035 2758
rect 4613 2755 4679 2758
rect 5022 2756 5028 2820
rect 5092 2818 5098 2820
rect 6545 2818 6611 2821
rect 6821 2820 6887 2821
rect 7465 2820 7531 2821
rect 6821 2818 6868 2820
rect 5092 2816 6611 2818
rect 5092 2760 6550 2816
rect 6606 2760 6611 2816
rect 5092 2758 6611 2760
rect 6776 2816 6868 2818
rect 6776 2760 6826 2816
rect 6776 2758 6868 2760
rect 5092 2756 5098 2758
rect 6545 2755 6611 2758
rect 6821 2756 6868 2758
rect 6932 2756 6938 2820
rect 7414 2756 7420 2820
rect 7484 2818 7531 2820
rect 10317 2818 10383 2821
rect 12341 2818 12407 2821
rect 7484 2816 7576 2818
rect 7526 2760 7576 2816
rect 7484 2758 7576 2760
rect 10317 2816 12407 2818
rect 10317 2760 10322 2816
rect 10378 2760 12346 2816
rect 12402 2760 12407 2816
rect 10317 2758 12407 2760
rect 7484 2756 7531 2758
rect 6821 2755 6887 2756
rect 7465 2755 7531 2756
rect 10317 2755 10383 2758
rect 12341 2755 12407 2758
rect 16113 2818 16179 2821
rect 17910 2818 17970 2894
rect 20253 2891 20319 2894
rect 16113 2816 17970 2818
rect 16113 2760 16118 2816
rect 16174 2760 17970 2816
rect 16113 2758 17970 2760
rect 16113 2755 16179 2758
rect 3545 2752 3861 2753
rect 0 2682 800 2712
rect 3545 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3861 2752
rect 3545 2687 3861 2688
rect 8743 2752 9059 2753
rect 8743 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9059 2752
rect 8743 2687 9059 2688
rect 13941 2752 14257 2753
rect 13941 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14257 2752
rect 13941 2687 14257 2688
rect 19139 2752 19455 2753
rect 19139 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19455 2752
rect 19139 2687 19455 2688
rect 2773 2682 2839 2685
rect 0 2680 2839 2682
rect 0 2624 2778 2680
rect 2834 2624 2839 2680
rect 0 2622 2839 2624
rect 0 2592 800 2622
rect 2773 2619 2839 2622
rect 4153 2682 4219 2685
rect 4470 2682 4476 2684
rect 4153 2680 4476 2682
rect 4153 2624 4158 2680
rect 4214 2624 4476 2680
rect 4153 2622 4476 2624
rect 4153 2619 4219 2622
rect 4470 2620 4476 2622
rect 4540 2620 4546 2684
rect 5441 2682 5507 2685
rect 7046 2682 7052 2684
rect 5441 2680 7052 2682
rect 5441 2624 5446 2680
rect 5502 2624 7052 2680
rect 5441 2622 7052 2624
rect 5441 2619 5507 2622
rect 7046 2620 7052 2622
rect 7116 2682 7122 2684
rect 7649 2682 7715 2685
rect 7116 2680 7715 2682
rect 7116 2624 7654 2680
rect 7710 2624 7715 2680
rect 7116 2622 7715 2624
rect 7116 2620 7122 2622
rect 7649 2619 7715 2622
rect 9305 2682 9371 2685
rect 20529 2684 20595 2685
rect 12566 2682 12572 2684
rect 9305 2680 12572 2682
rect 9305 2624 9310 2680
rect 9366 2624 12572 2680
rect 9305 2622 12572 2624
rect 9305 2619 9371 2622
rect 12566 2620 12572 2622
rect 12636 2620 12642 2684
rect 20478 2682 20484 2684
rect 20438 2622 20484 2682
rect 20548 2680 20595 2684
rect 22200 2682 23000 2712
rect 20590 2624 20595 2680
rect 20478 2620 20484 2622
rect 20548 2620 20595 2624
rect 20529 2619 20595 2620
rect 20670 2622 23000 2682
rect 1342 2484 1348 2548
rect 1412 2546 1418 2548
rect 2221 2546 2287 2549
rect 2681 2546 2747 2549
rect 1412 2544 2747 2546
rect 1412 2488 2226 2544
rect 2282 2488 2686 2544
rect 2742 2488 2747 2544
rect 1412 2486 2747 2488
rect 1412 2484 1418 2486
rect 2221 2483 2287 2486
rect 2681 2483 2747 2486
rect 3366 2484 3372 2548
rect 3436 2546 3442 2548
rect 3601 2546 3667 2549
rect 6678 2546 6684 2548
rect 3436 2544 6684 2546
rect 3436 2488 3606 2544
rect 3662 2488 6684 2544
rect 3436 2486 6684 2488
rect 3436 2484 3442 2486
rect 3601 2483 3667 2486
rect 6678 2484 6684 2486
rect 6748 2484 6754 2548
rect 9397 2546 9463 2549
rect 12198 2546 12204 2548
rect 6870 2544 12204 2546
rect 6870 2488 9402 2544
rect 9458 2488 12204 2544
rect 6870 2486 12204 2488
rect 1761 2410 1827 2413
rect 4981 2410 5047 2413
rect 1761 2408 5047 2410
rect 1761 2352 1766 2408
rect 1822 2352 4986 2408
rect 5042 2352 5047 2408
rect 1761 2350 5047 2352
rect 1761 2347 1827 2350
rect 4981 2347 5047 2350
rect 5390 2348 5396 2412
rect 5460 2410 5466 2412
rect 5533 2410 5599 2413
rect 5460 2408 5599 2410
rect 5460 2352 5538 2408
rect 5594 2352 5599 2408
rect 5460 2350 5599 2352
rect 5460 2348 5466 2350
rect 5533 2347 5599 2350
rect 5901 2410 5967 2413
rect 6870 2410 6930 2486
rect 9397 2483 9463 2486
rect 12198 2484 12204 2486
rect 12268 2484 12274 2548
rect 12341 2546 12407 2549
rect 16246 2546 16252 2548
rect 12341 2544 16252 2546
rect 12341 2488 12346 2544
rect 12402 2488 16252 2544
rect 12341 2486 16252 2488
rect 12341 2483 12407 2486
rect 16246 2484 16252 2486
rect 16316 2484 16322 2548
rect 18689 2546 18755 2549
rect 20670 2546 20730 2622
rect 22200 2592 23000 2622
rect 18689 2544 20730 2546
rect 18689 2488 18694 2544
rect 18750 2488 20730 2544
rect 18689 2486 20730 2488
rect 18689 2483 18755 2486
rect 5901 2408 6930 2410
rect 5901 2352 5906 2408
rect 5962 2352 6930 2408
rect 5901 2350 6930 2352
rect 7649 2410 7715 2413
rect 10133 2410 10199 2413
rect 7649 2408 10199 2410
rect 7649 2352 7654 2408
rect 7710 2352 10138 2408
rect 10194 2352 10199 2408
rect 7649 2350 10199 2352
rect 5901 2347 5967 2350
rect 7649 2347 7715 2350
rect 10133 2347 10199 2350
rect 17401 2410 17467 2413
rect 17401 2408 22202 2410
rect 17401 2352 17406 2408
rect 17462 2352 22202 2408
rect 17401 2350 22202 2352
rect 17401 2347 17467 2350
rect 22142 2304 22202 2350
rect 0 2274 800 2304
rect 3785 2274 3851 2277
rect 5901 2276 5967 2277
rect 5901 2274 5948 2276
rect 0 2272 3851 2274
rect 0 2216 3790 2272
rect 3846 2216 3851 2272
rect 0 2214 3851 2216
rect 5856 2272 5948 2274
rect 5856 2216 5906 2272
rect 5856 2214 5948 2216
rect 0 2184 800 2214
rect 3785 2211 3851 2214
rect 5901 2212 5948 2214
rect 6012 2212 6018 2276
rect 22142 2214 23000 2304
rect 5901 2211 5967 2212
rect 6144 2208 6460 2209
rect 6144 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6460 2208
rect 6144 2143 6460 2144
rect 11342 2208 11658 2209
rect 11342 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11658 2208
rect 11342 2143 11658 2144
rect 16540 2208 16856 2209
rect 16540 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16856 2208
rect 16540 2143 16856 2144
rect 21738 2208 22054 2209
rect 21738 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22054 2208
rect 22200 2184 23000 2214
rect 21738 2143 22054 2144
rect 7782 2076 7788 2140
rect 7852 2138 7858 2140
rect 8109 2138 8175 2141
rect 7852 2136 8175 2138
rect 7852 2080 8114 2136
rect 8170 2080 8175 2136
rect 7852 2078 8175 2080
rect 7852 2076 7858 2078
rect 8109 2075 8175 2078
rect 3325 2002 3391 2005
rect 10961 2002 11027 2005
rect 13302 2002 13308 2004
rect 3325 2000 11027 2002
rect 3325 1944 3330 2000
rect 3386 1944 10966 2000
rect 11022 1944 11027 2000
rect 3325 1942 11027 1944
rect 3325 1939 3391 1942
rect 10961 1939 11027 1942
rect 12390 1942 13308 2002
rect 0 1866 800 1896
rect 5533 1868 5599 1869
rect 4654 1866 4660 1868
rect 0 1806 4660 1866
rect 0 1776 800 1806
rect 4654 1804 4660 1806
rect 4724 1804 4730 1868
rect 5533 1866 5580 1868
rect 5488 1864 5580 1866
rect 5488 1808 5538 1864
rect 5488 1806 5580 1808
rect 5533 1804 5580 1806
rect 5644 1804 5650 1868
rect 6729 1866 6795 1869
rect 12390 1866 12450 1942
rect 13302 1940 13308 1942
rect 13372 1940 13378 2004
rect 6729 1864 12450 1866
rect 6729 1808 6734 1864
rect 6790 1808 12450 1864
rect 6729 1806 12450 1808
rect 19241 1866 19307 1869
rect 22200 1866 23000 1896
rect 19241 1864 23000 1866
rect 19241 1808 19246 1864
rect 19302 1808 23000 1864
rect 19241 1806 23000 1808
rect 5533 1803 5599 1804
rect 6729 1803 6795 1806
rect 19241 1803 19307 1806
rect 22200 1776 23000 1806
rect 4838 1668 4844 1732
rect 4908 1730 4914 1732
rect 12065 1730 12131 1733
rect 4908 1728 12131 1730
rect 4908 1672 12070 1728
rect 12126 1672 12131 1728
rect 4908 1670 12131 1672
rect 4908 1668 4914 1670
rect 12065 1667 12131 1670
rect 2957 1594 3023 1597
rect 2730 1592 3023 1594
rect 2730 1536 2962 1592
rect 3018 1536 3023 1592
rect 2730 1534 3023 1536
rect 0 1458 800 1488
rect 2730 1458 2790 1534
rect 2957 1531 3023 1534
rect 3182 1532 3188 1596
rect 3252 1594 3258 1596
rect 9489 1594 9555 1597
rect 3252 1592 9555 1594
rect 3252 1536 9494 1592
rect 9550 1536 9555 1592
rect 3252 1534 9555 1536
rect 3252 1532 3258 1534
rect 9489 1531 9555 1534
rect 0 1398 2790 1458
rect 4981 1458 5047 1461
rect 9305 1458 9371 1461
rect 4981 1456 9371 1458
rect 4981 1400 4986 1456
rect 5042 1400 9310 1456
rect 9366 1400 9371 1456
rect 4981 1398 9371 1400
rect 0 1368 800 1398
rect 4981 1395 5047 1398
rect 9305 1395 9371 1398
rect 19149 1458 19215 1461
rect 22200 1458 23000 1488
rect 19149 1456 23000 1458
rect 19149 1400 19154 1456
rect 19210 1400 23000 1456
rect 19149 1398 23000 1400
rect 19149 1395 19215 1398
rect 22200 1368 23000 1398
rect 1577 1322 1643 1325
rect 12985 1322 13051 1325
rect 1577 1320 13051 1322
rect 1577 1264 1582 1320
rect 1638 1264 12990 1320
rect 13046 1264 13051 1320
rect 1577 1262 13051 1264
rect 1577 1259 1643 1262
rect 12985 1259 13051 1262
rect 3141 1186 3207 1189
rect 3417 1186 3483 1189
rect 3141 1184 3483 1186
rect 3141 1128 3146 1184
rect 3202 1128 3422 1184
rect 3478 1128 3483 1184
rect 3141 1126 3483 1128
rect 3141 1123 3207 1126
rect 3417 1123 3483 1126
rect 3877 1186 3943 1189
rect 11094 1186 11100 1188
rect 3877 1184 11100 1186
rect 3877 1128 3882 1184
rect 3938 1128 11100 1184
rect 3877 1126 11100 1128
rect 3877 1123 3943 1126
rect 11094 1124 11100 1126
rect 11164 1124 11170 1188
rect 11237 1186 11303 1189
rect 14590 1186 14596 1188
rect 11237 1184 14596 1186
rect 11237 1128 11242 1184
rect 11298 1128 14596 1184
rect 11237 1126 14596 1128
rect 11237 1123 11303 1126
rect 14590 1124 14596 1126
rect 14660 1124 14666 1188
rect 0 1050 800 1080
rect 2773 1050 2839 1053
rect 13486 1050 13492 1052
rect 0 1048 13492 1050
rect 0 992 2778 1048
rect 2834 992 13492 1048
rect 0 990 13492 992
rect 0 960 800 990
rect 2773 987 2839 990
rect 13486 988 13492 990
rect 13556 988 13562 1052
rect 16062 988 16068 1052
rect 16132 1050 16138 1052
rect 20713 1050 20779 1053
rect 22200 1050 23000 1080
rect 16132 990 19626 1050
rect 16132 988 16138 990
rect 3417 914 3483 917
rect 11237 914 11303 917
rect 19425 914 19491 917
rect 3417 912 11303 914
rect 3417 856 3422 912
rect 3478 856 11242 912
rect 11298 856 11303 912
rect 3417 854 11303 856
rect 3417 851 3483 854
rect 11237 851 11303 854
rect 16530 912 19491 914
rect 16530 856 19430 912
rect 19486 856 19491 912
rect 16530 854 19491 856
rect 5206 716 5212 780
rect 5276 778 5282 780
rect 16530 778 16590 854
rect 19425 851 19491 854
rect 5276 718 16590 778
rect 5276 716 5282 718
rect 0 642 800 672
rect 1025 642 1091 645
rect 0 640 1091 642
rect 0 584 1030 640
rect 1086 584 1091 640
rect 0 582 1091 584
rect 19566 642 19626 990
rect 20713 1048 23000 1050
rect 20713 992 20718 1048
rect 20774 992 23000 1048
rect 20713 990 23000 992
rect 20713 987 20779 990
rect 22200 960 23000 990
rect 22200 642 23000 672
rect 19566 582 23000 642
rect 0 552 800 582
rect 1025 579 1091 582
rect 22200 552 23000 582
rect 4613 98 4679 101
rect 14774 98 14780 100
rect 4613 96 14780 98
rect 4613 40 4618 96
rect 4674 40 14780 96
rect 4613 38 14780 40
rect 4613 35 4679 38
rect 14774 36 14780 38
rect 14844 36 14850 100
<< via3 >>
rect 60 22476 124 22540
rect 14412 22476 14476 22540
rect 12756 21252 12820 21316
rect 1164 21116 1228 21180
rect 4844 20980 4908 21044
rect 8156 20844 8220 20908
rect 11100 20708 11164 20772
rect 6150 20700 6214 20704
rect 6150 20644 6154 20700
rect 6154 20644 6210 20700
rect 6210 20644 6214 20700
rect 6150 20640 6214 20644
rect 6230 20700 6294 20704
rect 6230 20644 6234 20700
rect 6234 20644 6290 20700
rect 6290 20644 6294 20700
rect 6230 20640 6294 20644
rect 6310 20700 6374 20704
rect 6310 20644 6314 20700
rect 6314 20644 6370 20700
rect 6370 20644 6374 20700
rect 6310 20640 6374 20644
rect 6390 20700 6454 20704
rect 6390 20644 6394 20700
rect 6394 20644 6450 20700
rect 6450 20644 6454 20700
rect 6390 20640 6454 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 16546 20700 16610 20704
rect 16546 20644 16550 20700
rect 16550 20644 16606 20700
rect 16606 20644 16610 20700
rect 16546 20640 16610 20644
rect 16626 20700 16690 20704
rect 16626 20644 16630 20700
rect 16630 20644 16686 20700
rect 16686 20644 16690 20700
rect 16626 20640 16690 20644
rect 16706 20700 16770 20704
rect 16706 20644 16710 20700
rect 16710 20644 16766 20700
rect 16766 20644 16770 20700
rect 16706 20640 16770 20644
rect 16786 20700 16850 20704
rect 16786 20644 16790 20700
rect 16790 20644 16846 20700
rect 16846 20644 16850 20700
rect 16786 20640 16850 20644
rect 21744 20700 21808 20704
rect 21744 20644 21748 20700
rect 21748 20644 21804 20700
rect 21804 20644 21808 20700
rect 21744 20640 21808 20644
rect 21824 20700 21888 20704
rect 21824 20644 21828 20700
rect 21828 20644 21884 20700
rect 21884 20644 21888 20700
rect 21824 20640 21888 20644
rect 21904 20700 21968 20704
rect 21904 20644 21908 20700
rect 21908 20644 21964 20700
rect 21964 20644 21968 20700
rect 21904 20640 21968 20644
rect 21984 20700 22048 20704
rect 21984 20644 21988 20700
rect 21988 20644 22044 20700
rect 22044 20644 22048 20700
rect 21984 20640 22048 20644
rect 14596 20300 14660 20364
rect 2452 20164 2516 20228
rect 3551 20156 3615 20160
rect 3551 20100 3555 20156
rect 3555 20100 3611 20156
rect 3611 20100 3615 20156
rect 3551 20096 3615 20100
rect 3631 20156 3695 20160
rect 3631 20100 3635 20156
rect 3635 20100 3691 20156
rect 3691 20100 3695 20156
rect 3631 20096 3695 20100
rect 3711 20156 3775 20160
rect 3711 20100 3715 20156
rect 3715 20100 3771 20156
rect 3771 20100 3775 20156
rect 3711 20096 3775 20100
rect 3791 20156 3855 20160
rect 3791 20100 3795 20156
rect 3795 20100 3851 20156
rect 3851 20100 3855 20156
rect 3791 20096 3855 20100
rect 8749 20156 8813 20160
rect 8749 20100 8753 20156
rect 8753 20100 8809 20156
rect 8809 20100 8813 20156
rect 8749 20096 8813 20100
rect 8829 20156 8893 20160
rect 8829 20100 8833 20156
rect 8833 20100 8889 20156
rect 8889 20100 8893 20156
rect 8829 20096 8893 20100
rect 8909 20156 8973 20160
rect 8909 20100 8913 20156
rect 8913 20100 8969 20156
rect 8969 20100 8973 20156
rect 8909 20096 8973 20100
rect 8989 20156 9053 20160
rect 8989 20100 8993 20156
rect 8993 20100 9049 20156
rect 9049 20100 9053 20156
rect 8989 20096 9053 20100
rect 13947 20156 14011 20160
rect 13947 20100 13951 20156
rect 13951 20100 14007 20156
rect 14007 20100 14011 20156
rect 13947 20096 14011 20100
rect 14027 20156 14091 20160
rect 14027 20100 14031 20156
rect 14031 20100 14087 20156
rect 14087 20100 14091 20156
rect 14027 20096 14091 20100
rect 14107 20156 14171 20160
rect 14107 20100 14111 20156
rect 14111 20100 14167 20156
rect 14167 20100 14171 20156
rect 14107 20096 14171 20100
rect 14187 20156 14251 20160
rect 14187 20100 14191 20156
rect 14191 20100 14247 20156
rect 14247 20100 14251 20156
rect 14187 20096 14251 20100
rect 19145 20156 19209 20160
rect 19145 20100 19149 20156
rect 19149 20100 19205 20156
rect 19205 20100 19209 20156
rect 19145 20096 19209 20100
rect 19225 20156 19289 20160
rect 19225 20100 19229 20156
rect 19229 20100 19285 20156
rect 19285 20100 19289 20156
rect 19225 20096 19289 20100
rect 19305 20156 19369 20160
rect 19305 20100 19309 20156
rect 19309 20100 19365 20156
rect 19365 20100 19369 20156
rect 19305 20096 19369 20100
rect 19385 20156 19449 20160
rect 19385 20100 19389 20156
rect 19389 20100 19445 20156
rect 19445 20100 19449 20156
rect 19385 20096 19449 20100
rect 8340 20028 8404 20092
rect 6150 19612 6214 19616
rect 6150 19556 6154 19612
rect 6154 19556 6210 19612
rect 6210 19556 6214 19612
rect 6150 19552 6214 19556
rect 6230 19612 6294 19616
rect 6230 19556 6234 19612
rect 6234 19556 6290 19612
rect 6290 19556 6294 19612
rect 6230 19552 6294 19556
rect 6310 19612 6374 19616
rect 6310 19556 6314 19612
rect 6314 19556 6370 19612
rect 6370 19556 6374 19612
rect 6310 19552 6374 19556
rect 6390 19612 6454 19616
rect 6390 19556 6394 19612
rect 6394 19556 6450 19612
rect 6450 19556 6454 19612
rect 6390 19552 6454 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 16546 19612 16610 19616
rect 16546 19556 16550 19612
rect 16550 19556 16606 19612
rect 16606 19556 16610 19612
rect 16546 19552 16610 19556
rect 16626 19612 16690 19616
rect 16626 19556 16630 19612
rect 16630 19556 16686 19612
rect 16686 19556 16690 19612
rect 16626 19552 16690 19556
rect 16706 19612 16770 19616
rect 16706 19556 16710 19612
rect 16710 19556 16766 19612
rect 16766 19556 16770 19612
rect 16706 19552 16770 19556
rect 16786 19612 16850 19616
rect 16786 19556 16790 19612
rect 16790 19556 16846 19612
rect 16846 19556 16850 19612
rect 16786 19552 16850 19556
rect 21744 19612 21808 19616
rect 21744 19556 21748 19612
rect 21748 19556 21804 19612
rect 21804 19556 21808 19612
rect 21744 19552 21808 19556
rect 21824 19612 21888 19616
rect 21824 19556 21828 19612
rect 21828 19556 21884 19612
rect 21884 19556 21888 19612
rect 21824 19552 21888 19556
rect 21904 19612 21968 19616
rect 21904 19556 21908 19612
rect 21908 19556 21964 19612
rect 21964 19556 21968 19612
rect 21904 19552 21968 19556
rect 21984 19612 22048 19616
rect 21984 19556 21988 19612
rect 21988 19556 22044 19612
rect 22044 19556 22048 19612
rect 21984 19552 22048 19556
rect 4476 19544 4540 19548
rect 4476 19488 4526 19544
rect 4526 19488 4540 19544
rect 4476 19484 4540 19488
rect 8524 19484 8588 19548
rect 7420 19348 7484 19412
rect 7788 19348 7852 19412
rect 19564 19272 19628 19276
rect 19564 19216 19614 19272
rect 19614 19216 19628 19272
rect 19564 19212 19628 19216
rect 3551 19068 3615 19072
rect 3551 19012 3555 19068
rect 3555 19012 3611 19068
rect 3611 19012 3615 19068
rect 3551 19008 3615 19012
rect 3631 19068 3695 19072
rect 3631 19012 3635 19068
rect 3635 19012 3691 19068
rect 3691 19012 3695 19068
rect 3631 19008 3695 19012
rect 3711 19068 3775 19072
rect 3711 19012 3715 19068
rect 3715 19012 3771 19068
rect 3771 19012 3775 19068
rect 3711 19008 3775 19012
rect 3791 19068 3855 19072
rect 3791 19012 3795 19068
rect 3795 19012 3851 19068
rect 3851 19012 3855 19068
rect 3791 19008 3855 19012
rect 17908 19076 17972 19140
rect 8749 19068 8813 19072
rect 8749 19012 8753 19068
rect 8753 19012 8809 19068
rect 8809 19012 8813 19068
rect 8749 19008 8813 19012
rect 8829 19068 8893 19072
rect 8829 19012 8833 19068
rect 8833 19012 8889 19068
rect 8889 19012 8893 19068
rect 8829 19008 8893 19012
rect 8909 19068 8973 19072
rect 8909 19012 8913 19068
rect 8913 19012 8969 19068
rect 8969 19012 8973 19068
rect 8909 19008 8973 19012
rect 8989 19068 9053 19072
rect 8989 19012 8993 19068
rect 8993 19012 9049 19068
rect 9049 19012 9053 19068
rect 8989 19008 9053 19012
rect 13947 19068 14011 19072
rect 13947 19012 13951 19068
rect 13951 19012 14007 19068
rect 14007 19012 14011 19068
rect 13947 19008 14011 19012
rect 14027 19068 14091 19072
rect 14027 19012 14031 19068
rect 14031 19012 14087 19068
rect 14087 19012 14091 19068
rect 14027 19008 14091 19012
rect 14107 19068 14171 19072
rect 14107 19012 14111 19068
rect 14111 19012 14167 19068
rect 14167 19012 14171 19068
rect 14107 19008 14171 19012
rect 14187 19068 14251 19072
rect 14187 19012 14191 19068
rect 14191 19012 14247 19068
rect 14247 19012 14251 19068
rect 14187 19008 14251 19012
rect 19145 19068 19209 19072
rect 19145 19012 19149 19068
rect 19149 19012 19205 19068
rect 19205 19012 19209 19068
rect 19145 19008 19209 19012
rect 19225 19068 19289 19072
rect 19225 19012 19229 19068
rect 19229 19012 19285 19068
rect 19285 19012 19289 19068
rect 19225 19008 19289 19012
rect 19305 19068 19369 19072
rect 19305 19012 19309 19068
rect 19309 19012 19365 19068
rect 19365 19012 19369 19068
rect 19305 19008 19369 19012
rect 19385 19068 19449 19072
rect 19385 19012 19389 19068
rect 19389 19012 19445 19068
rect 19445 19012 19449 19068
rect 19385 19008 19449 19012
rect 19932 18940 19996 19004
rect 5764 18804 5828 18868
rect 10732 18804 10796 18868
rect 5580 18456 5644 18460
rect 5580 18400 5594 18456
rect 5594 18400 5644 18456
rect 5580 18396 5644 18400
rect 5764 18320 5828 18324
rect 5764 18264 5814 18320
rect 5814 18264 5828 18320
rect 5764 18260 5828 18264
rect 10548 18592 10612 18596
rect 10548 18536 10598 18592
rect 10598 18536 10612 18592
rect 10548 18532 10612 18536
rect 6150 18524 6214 18528
rect 6150 18468 6154 18524
rect 6154 18468 6210 18524
rect 6210 18468 6214 18524
rect 6150 18464 6214 18468
rect 6230 18524 6294 18528
rect 6230 18468 6234 18524
rect 6234 18468 6290 18524
rect 6290 18468 6294 18524
rect 6230 18464 6294 18468
rect 6310 18524 6374 18528
rect 6310 18468 6314 18524
rect 6314 18468 6370 18524
rect 6370 18468 6374 18524
rect 6310 18464 6374 18468
rect 6390 18524 6454 18528
rect 6390 18468 6394 18524
rect 6394 18468 6450 18524
rect 6450 18468 6454 18524
rect 6390 18464 6454 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 15332 18668 15396 18732
rect 16546 18524 16610 18528
rect 16546 18468 16550 18524
rect 16550 18468 16606 18524
rect 16606 18468 16610 18524
rect 16546 18464 16610 18468
rect 16626 18524 16690 18528
rect 16626 18468 16630 18524
rect 16630 18468 16686 18524
rect 16686 18468 16690 18524
rect 16626 18464 16690 18468
rect 16706 18524 16770 18528
rect 16706 18468 16710 18524
rect 16710 18468 16766 18524
rect 16766 18468 16770 18524
rect 16706 18464 16770 18468
rect 16786 18524 16850 18528
rect 16786 18468 16790 18524
rect 16790 18468 16846 18524
rect 16846 18468 16850 18524
rect 16786 18464 16850 18468
rect 21744 18524 21808 18528
rect 21744 18468 21748 18524
rect 21748 18468 21804 18524
rect 21804 18468 21808 18524
rect 21744 18464 21808 18468
rect 21824 18524 21888 18528
rect 21824 18468 21828 18524
rect 21828 18468 21884 18524
rect 21884 18468 21888 18524
rect 21824 18464 21888 18468
rect 21904 18524 21968 18528
rect 21904 18468 21908 18524
rect 21908 18468 21964 18524
rect 21964 18468 21968 18524
rect 21904 18464 21968 18468
rect 21984 18524 22048 18528
rect 21984 18468 21988 18524
rect 21988 18468 22044 18524
rect 22044 18468 22048 18524
rect 21984 18464 22048 18468
rect 19564 18456 19628 18460
rect 19564 18400 19614 18456
rect 19614 18400 19628 18456
rect 19564 18396 19628 18400
rect 19932 18396 19996 18460
rect 4108 17988 4172 18052
rect 14964 18124 15028 18188
rect 16252 17988 16316 18052
rect 3551 17980 3615 17984
rect 3551 17924 3555 17980
rect 3555 17924 3611 17980
rect 3611 17924 3615 17980
rect 3551 17920 3615 17924
rect 3631 17980 3695 17984
rect 3631 17924 3635 17980
rect 3635 17924 3691 17980
rect 3691 17924 3695 17980
rect 3631 17920 3695 17924
rect 3711 17980 3775 17984
rect 3711 17924 3715 17980
rect 3715 17924 3771 17980
rect 3771 17924 3775 17980
rect 3711 17920 3775 17924
rect 3791 17980 3855 17984
rect 3791 17924 3795 17980
rect 3795 17924 3851 17980
rect 3851 17924 3855 17980
rect 3791 17920 3855 17924
rect 8749 17980 8813 17984
rect 8749 17924 8753 17980
rect 8753 17924 8809 17980
rect 8809 17924 8813 17980
rect 8749 17920 8813 17924
rect 8829 17980 8893 17984
rect 8829 17924 8833 17980
rect 8833 17924 8889 17980
rect 8889 17924 8893 17980
rect 8829 17920 8893 17924
rect 8909 17980 8973 17984
rect 8909 17924 8913 17980
rect 8913 17924 8969 17980
rect 8969 17924 8973 17980
rect 8909 17920 8973 17924
rect 8989 17980 9053 17984
rect 8989 17924 8993 17980
rect 8993 17924 9049 17980
rect 9049 17924 9053 17980
rect 8989 17920 9053 17924
rect 13947 17980 14011 17984
rect 13947 17924 13951 17980
rect 13951 17924 14007 17980
rect 14007 17924 14011 17980
rect 13947 17920 14011 17924
rect 14027 17980 14091 17984
rect 14027 17924 14031 17980
rect 14031 17924 14087 17980
rect 14087 17924 14091 17980
rect 14027 17920 14091 17924
rect 14107 17980 14171 17984
rect 14107 17924 14111 17980
rect 14111 17924 14167 17980
rect 14167 17924 14171 17980
rect 14107 17920 14171 17924
rect 14187 17980 14251 17984
rect 14187 17924 14191 17980
rect 14191 17924 14247 17980
rect 14247 17924 14251 17980
rect 14187 17920 14251 17924
rect 19145 17980 19209 17984
rect 19145 17924 19149 17980
rect 19149 17924 19205 17980
rect 19205 17924 19209 17980
rect 19145 17920 19209 17924
rect 19225 17980 19289 17984
rect 19225 17924 19229 17980
rect 19229 17924 19285 17980
rect 19285 17924 19289 17980
rect 19225 17920 19289 17924
rect 19305 17980 19369 17984
rect 19305 17924 19309 17980
rect 19309 17924 19365 17980
rect 19365 17924 19369 17980
rect 19305 17920 19369 17924
rect 19385 17980 19449 17984
rect 19385 17924 19389 17980
rect 19389 17924 19445 17980
rect 19445 17924 19449 17980
rect 19385 17920 19449 17924
rect 7604 17852 7668 17916
rect 9996 17716 10060 17780
rect 20300 17716 20364 17780
rect 6684 17444 6748 17508
rect 6150 17436 6214 17440
rect 6150 17380 6154 17436
rect 6154 17380 6210 17436
rect 6210 17380 6214 17436
rect 6150 17376 6214 17380
rect 6230 17436 6294 17440
rect 6230 17380 6234 17436
rect 6234 17380 6290 17436
rect 6290 17380 6294 17436
rect 6230 17376 6294 17380
rect 6310 17436 6374 17440
rect 6310 17380 6314 17436
rect 6314 17380 6370 17436
rect 6370 17380 6374 17436
rect 6310 17376 6374 17380
rect 6390 17436 6454 17440
rect 6390 17380 6394 17436
rect 6394 17380 6450 17436
rect 6450 17380 6454 17436
rect 6390 17376 6454 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 16546 17436 16610 17440
rect 16546 17380 16550 17436
rect 16550 17380 16606 17436
rect 16606 17380 16610 17436
rect 16546 17376 16610 17380
rect 16626 17436 16690 17440
rect 16626 17380 16630 17436
rect 16630 17380 16686 17436
rect 16686 17380 16690 17436
rect 16626 17376 16690 17380
rect 16706 17436 16770 17440
rect 16706 17380 16710 17436
rect 16710 17380 16766 17436
rect 16766 17380 16770 17436
rect 16706 17376 16770 17380
rect 16786 17436 16850 17440
rect 16786 17380 16790 17436
rect 16790 17380 16846 17436
rect 16846 17380 16850 17436
rect 16786 17376 16850 17380
rect 21744 17436 21808 17440
rect 21744 17380 21748 17436
rect 21748 17380 21804 17436
rect 21804 17380 21808 17436
rect 21744 17376 21808 17380
rect 21824 17436 21888 17440
rect 21824 17380 21828 17436
rect 21828 17380 21884 17436
rect 21884 17380 21888 17436
rect 21824 17376 21888 17380
rect 21904 17436 21968 17440
rect 21904 17380 21908 17436
rect 21908 17380 21964 17436
rect 21964 17380 21968 17436
rect 21904 17376 21968 17380
rect 21984 17436 22048 17440
rect 21984 17380 21988 17436
rect 21988 17380 22044 17436
rect 22044 17380 22048 17436
rect 21984 17376 22048 17380
rect 3924 17308 3988 17372
rect 3372 17172 3436 17236
rect 15332 17036 15396 17100
rect 13676 16960 13740 16964
rect 13676 16904 13726 16960
rect 13726 16904 13740 16960
rect 3551 16892 3615 16896
rect 3551 16836 3555 16892
rect 3555 16836 3611 16892
rect 3611 16836 3615 16892
rect 3551 16832 3615 16836
rect 3631 16892 3695 16896
rect 3631 16836 3635 16892
rect 3635 16836 3691 16892
rect 3691 16836 3695 16892
rect 3631 16832 3695 16836
rect 3711 16892 3775 16896
rect 3711 16836 3715 16892
rect 3715 16836 3771 16892
rect 3771 16836 3775 16892
rect 3711 16832 3775 16836
rect 3791 16892 3855 16896
rect 3791 16836 3795 16892
rect 3795 16836 3851 16892
rect 3851 16836 3855 16892
rect 3791 16832 3855 16836
rect 8749 16892 8813 16896
rect 8749 16836 8753 16892
rect 8753 16836 8809 16892
rect 8809 16836 8813 16892
rect 8749 16832 8813 16836
rect 8829 16892 8893 16896
rect 8829 16836 8833 16892
rect 8833 16836 8889 16892
rect 8889 16836 8893 16892
rect 8829 16832 8893 16836
rect 8909 16892 8973 16896
rect 8909 16836 8913 16892
rect 8913 16836 8969 16892
rect 8969 16836 8973 16892
rect 8909 16832 8973 16836
rect 8989 16892 9053 16896
rect 8989 16836 8993 16892
rect 8993 16836 9049 16892
rect 9049 16836 9053 16892
rect 8989 16832 9053 16836
rect 7972 16688 8036 16692
rect 7972 16632 7986 16688
rect 7986 16632 8036 16688
rect 7972 16628 8036 16632
rect 8524 16628 8588 16692
rect 13676 16900 13740 16904
rect 13947 16892 14011 16896
rect 13947 16836 13951 16892
rect 13951 16836 14007 16892
rect 14007 16836 14011 16892
rect 13947 16832 14011 16836
rect 14027 16892 14091 16896
rect 14027 16836 14031 16892
rect 14031 16836 14087 16892
rect 14087 16836 14091 16892
rect 14027 16832 14091 16836
rect 14107 16892 14171 16896
rect 14107 16836 14111 16892
rect 14111 16836 14167 16892
rect 14167 16836 14171 16892
rect 14107 16832 14171 16836
rect 14187 16892 14251 16896
rect 14187 16836 14191 16892
rect 14191 16836 14247 16892
rect 14247 16836 14251 16892
rect 14187 16832 14251 16836
rect 19145 16892 19209 16896
rect 19145 16836 19149 16892
rect 19149 16836 19205 16892
rect 19205 16836 19209 16892
rect 19145 16832 19209 16836
rect 19225 16892 19289 16896
rect 19225 16836 19229 16892
rect 19229 16836 19285 16892
rect 19285 16836 19289 16892
rect 19225 16832 19289 16836
rect 19305 16892 19369 16896
rect 19305 16836 19309 16892
rect 19309 16836 19365 16892
rect 19365 16836 19369 16892
rect 19305 16832 19369 16836
rect 19385 16892 19449 16896
rect 19385 16836 19389 16892
rect 19389 16836 19445 16892
rect 19445 16836 19449 16892
rect 19385 16832 19449 16836
rect 10916 16628 10980 16692
rect 6150 16348 6214 16352
rect 6150 16292 6154 16348
rect 6154 16292 6210 16348
rect 6210 16292 6214 16348
rect 6150 16288 6214 16292
rect 6230 16348 6294 16352
rect 6230 16292 6234 16348
rect 6234 16292 6290 16348
rect 6290 16292 6294 16348
rect 6230 16288 6294 16292
rect 6310 16348 6374 16352
rect 6310 16292 6314 16348
rect 6314 16292 6370 16348
rect 6370 16292 6374 16348
rect 6310 16288 6374 16292
rect 6390 16348 6454 16352
rect 6390 16292 6394 16348
rect 6394 16292 6450 16348
rect 6450 16292 6454 16348
rect 6390 16288 6454 16292
rect 8156 16492 8220 16556
rect 8524 16356 8588 16420
rect 15700 16628 15764 16692
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 9812 16220 9876 16284
rect 16546 16348 16610 16352
rect 16546 16292 16550 16348
rect 16550 16292 16606 16348
rect 16606 16292 16610 16348
rect 16546 16288 16610 16292
rect 16626 16348 16690 16352
rect 16626 16292 16630 16348
rect 16630 16292 16686 16348
rect 16686 16292 16690 16348
rect 16626 16288 16690 16292
rect 16706 16348 16770 16352
rect 16706 16292 16710 16348
rect 16710 16292 16766 16348
rect 16766 16292 16770 16348
rect 16706 16288 16770 16292
rect 16786 16348 16850 16352
rect 16786 16292 16790 16348
rect 16790 16292 16846 16348
rect 16846 16292 16850 16348
rect 16786 16288 16850 16292
rect 21744 16348 21808 16352
rect 21744 16292 21748 16348
rect 21748 16292 21804 16348
rect 21804 16292 21808 16348
rect 21744 16288 21808 16292
rect 21824 16348 21888 16352
rect 21824 16292 21828 16348
rect 21828 16292 21884 16348
rect 21884 16292 21888 16348
rect 21824 16288 21888 16292
rect 21904 16348 21968 16352
rect 21904 16292 21908 16348
rect 21908 16292 21964 16348
rect 21964 16292 21968 16348
rect 21904 16288 21968 16292
rect 21984 16348 22048 16352
rect 21984 16292 21988 16348
rect 21988 16292 22044 16348
rect 22044 16292 22048 16348
rect 21984 16288 22048 16292
rect 10180 16084 10244 16148
rect 16252 15948 16316 16012
rect 3551 15804 3615 15808
rect 3551 15748 3555 15804
rect 3555 15748 3611 15804
rect 3611 15748 3615 15804
rect 3551 15744 3615 15748
rect 3631 15804 3695 15808
rect 3631 15748 3635 15804
rect 3635 15748 3691 15804
rect 3691 15748 3695 15804
rect 3631 15744 3695 15748
rect 3711 15804 3775 15808
rect 3711 15748 3715 15804
rect 3715 15748 3771 15804
rect 3771 15748 3775 15804
rect 3711 15744 3775 15748
rect 3791 15804 3855 15808
rect 3791 15748 3795 15804
rect 3795 15748 3851 15804
rect 3851 15748 3855 15804
rect 3791 15744 3855 15748
rect 8749 15804 8813 15808
rect 8749 15748 8753 15804
rect 8753 15748 8809 15804
rect 8809 15748 8813 15804
rect 8749 15744 8813 15748
rect 8829 15804 8893 15808
rect 8829 15748 8833 15804
rect 8833 15748 8889 15804
rect 8889 15748 8893 15804
rect 8829 15744 8893 15748
rect 8909 15804 8973 15808
rect 8909 15748 8913 15804
rect 8913 15748 8969 15804
rect 8969 15748 8973 15804
rect 8909 15744 8973 15748
rect 8989 15804 9053 15808
rect 8989 15748 8993 15804
rect 8993 15748 9049 15804
rect 9049 15748 9053 15804
rect 8989 15744 9053 15748
rect 13947 15804 14011 15808
rect 13947 15748 13951 15804
rect 13951 15748 14007 15804
rect 14007 15748 14011 15804
rect 13947 15744 14011 15748
rect 14027 15804 14091 15808
rect 14027 15748 14031 15804
rect 14031 15748 14087 15804
rect 14087 15748 14091 15804
rect 14027 15744 14091 15748
rect 14107 15804 14171 15808
rect 14107 15748 14111 15804
rect 14111 15748 14167 15804
rect 14167 15748 14171 15804
rect 14107 15744 14171 15748
rect 14187 15804 14251 15808
rect 14187 15748 14191 15804
rect 14191 15748 14247 15804
rect 14247 15748 14251 15804
rect 14187 15744 14251 15748
rect 10732 15540 10796 15604
rect 8156 15404 8220 15468
rect 19145 15804 19209 15808
rect 19145 15748 19149 15804
rect 19149 15748 19205 15804
rect 19205 15748 19209 15804
rect 19145 15744 19209 15748
rect 19225 15804 19289 15808
rect 19225 15748 19229 15804
rect 19229 15748 19285 15804
rect 19285 15748 19289 15804
rect 19225 15744 19289 15748
rect 19305 15804 19369 15808
rect 19305 15748 19309 15804
rect 19309 15748 19365 15804
rect 19365 15748 19369 15804
rect 19305 15744 19369 15748
rect 19385 15804 19449 15808
rect 19385 15748 19389 15804
rect 19389 15748 19445 15804
rect 19445 15748 19449 15804
rect 19385 15744 19449 15748
rect 5948 15328 6012 15332
rect 5948 15272 5962 15328
rect 5962 15272 6012 15328
rect 5948 15268 6012 15272
rect 6150 15260 6214 15264
rect 6150 15204 6154 15260
rect 6154 15204 6210 15260
rect 6210 15204 6214 15260
rect 6150 15200 6214 15204
rect 6230 15260 6294 15264
rect 6230 15204 6234 15260
rect 6234 15204 6290 15260
rect 6290 15204 6294 15260
rect 6230 15200 6294 15204
rect 6310 15260 6374 15264
rect 6310 15204 6314 15260
rect 6314 15204 6370 15260
rect 6370 15204 6374 15260
rect 6310 15200 6374 15204
rect 6390 15260 6454 15264
rect 6390 15204 6394 15260
rect 6394 15204 6450 15260
rect 6450 15204 6454 15260
rect 6390 15200 6454 15204
rect 9444 15268 9508 15332
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 10548 15132 10612 15196
rect 19932 15268 19996 15332
rect 16546 15260 16610 15264
rect 16546 15204 16550 15260
rect 16550 15204 16606 15260
rect 16606 15204 16610 15260
rect 16546 15200 16610 15204
rect 16626 15260 16690 15264
rect 16626 15204 16630 15260
rect 16630 15204 16686 15260
rect 16686 15204 16690 15260
rect 16626 15200 16690 15204
rect 16706 15260 16770 15264
rect 16706 15204 16710 15260
rect 16710 15204 16766 15260
rect 16766 15204 16770 15260
rect 16706 15200 16770 15204
rect 16786 15260 16850 15264
rect 16786 15204 16790 15260
rect 16790 15204 16846 15260
rect 16846 15204 16850 15260
rect 16786 15200 16850 15204
rect 21744 15260 21808 15264
rect 21744 15204 21748 15260
rect 21748 15204 21804 15260
rect 21804 15204 21808 15260
rect 21744 15200 21808 15204
rect 21824 15260 21888 15264
rect 21824 15204 21828 15260
rect 21828 15204 21884 15260
rect 21884 15204 21888 15260
rect 21824 15200 21888 15204
rect 21904 15260 21968 15264
rect 21904 15204 21908 15260
rect 21908 15204 21964 15260
rect 21964 15204 21968 15260
rect 21904 15200 21968 15204
rect 21984 15260 22048 15264
rect 21984 15204 21988 15260
rect 21988 15204 22044 15260
rect 22044 15204 22048 15260
rect 21984 15200 22048 15204
rect 12572 15132 12636 15196
rect 15516 14996 15580 15060
rect 3924 14860 3988 14924
rect 10916 14860 10980 14924
rect 13124 14920 13188 14924
rect 13124 14864 13174 14920
rect 13174 14864 13188 14920
rect 13124 14860 13188 14864
rect 10548 14784 10612 14788
rect 10548 14728 10598 14784
rect 10598 14728 10612 14784
rect 10548 14724 10612 14728
rect 20116 14784 20180 14788
rect 20116 14728 20130 14784
rect 20130 14728 20180 14784
rect 20116 14724 20180 14728
rect 3551 14716 3615 14720
rect 3551 14660 3555 14716
rect 3555 14660 3611 14716
rect 3611 14660 3615 14716
rect 3551 14656 3615 14660
rect 3631 14716 3695 14720
rect 3631 14660 3635 14716
rect 3635 14660 3691 14716
rect 3691 14660 3695 14716
rect 3631 14656 3695 14660
rect 3711 14716 3775 14720
rect 3711 14660 3715 14716
rect 3715 14660 3771 14716
rect 3771 14660 3775 14716
rect 3711 14656 3775 14660
rect 3791 14716 3855 14720
rect 3791 14660 3795 14716
rect 3795 14660 3851 14716
rect 3851 14660 3855 14716
rect 3791 14656 3855 14660
rect 8749 14716 8813 14720
rect 8749 14660 8753 14716
rect 8753 14660 8809 14716
rect 8809 14660 8813 14716
rect 8749 14656 8813 14660
rect 8829 14716 8893 14720
rect 8829 14660 8833 14716
rect 8833 14660 8889 14716
rect 8889 14660 8893 14716
rect 8829 14656 8893 14660
rect 8909 14716 8973 14720
rect 8909 14660 8913 14716
rect 8913 14660 8969 14716
rect 8969 14660 8973 14716
rect 8909 14656 8973 14660
rect 8989 14716 9053 14720
rect 8989 14660 8993 14716
rect 8993 14660 9049 14716
rect 9049 14660 9053 14716
rect 8989 14656 9053 14660
rect 13947 14716 14011 14720
rect 13947 14660 13951 14716
rect 13951 14660 14007 14716
rect 14007 14660 14011 14716
rect 13947 14656 14011 14660
rect 14027 14716 14091 14720
rect 14027 14660 14031 14716
rect 14031 14660 14087 14716
rect 14087 14660 14091 14716
rect 14027 14656 14091 14660
rect 14107 14716 14171 14720
rect 14107 14660 14111 14716
rect 14111 14660 14167 14716
rect 14167 14660 14171 14716
rect 14107 14656 14171 14660
rect 14187 14716 14251 14720
rect 14187 14660 14191 14716
rect 14191 14660 14247 14716
rect 14247 14660 14251 14716
rect 14187 14656 14251 14660
rect 19145 14716 19209 14720
rect 19145 14660 19149 14716
rect 19149 14660 19205 14716
rect 19205 14660 19209 14716
rect 19145 14656 19209 14660
rect 19225 14716 19289 14720
rect 19225 14660 19229 14716
rect 19229 14660 19285 14716
rect 19285 14660 19289 14716
rect 19225 14656 19289 14660
rect 19305 14716 19369 14720
rect 19305 14660 19309 14716
rect 19309 14660 19365 14716
rect 19365 14660 19369 14716
rect 19305 14656 19369 14660
rect 19385 14716 19449 14720
rect 19385 14660 19389 14716
rect 19389 14660 19445 14716
rect 19445 14660 19449 14716
rect 19385 14656 19449 14660
rect 11100 14588 11164 14652
rect 11836 14588 11900 14652
rect 12020 14588 12084 14652
rect 1164 14316 1228 14380
rect 14412 14452 14476 14516
rect 8340 14180 8404 14244
rect 9260 14180 9324 14244
rect 11836 14180 11900 14244
rect 6150 14172 6214 14176
rect 6150 14116 6154 14172
rect 6154 14116 6210 14172
rect 6210 14116 6214 14172
rect 6150 14112 6214 14116
rect 6230 14172 6294 14176
rect 6230 14116 6234 14172
rect 6234 14116 6290 14172
rect 6290 14116 6294 14172
rect 6230 14112 6294 14116
rect 6310 14172 6374 14176
rect 6310 14116 6314 14172
rect 6314 14116 6370 14172
rect 6370 14116 6374 14172
rect 6310 14112 6374 14116
rect 6390 14172 6454 14176
rect 6390 14116 6394 14172
rect 6394 14116 6450 14172
rect 6450 14116 6454 14172
rect 6390 14112 6454 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 16546 14172 16610 14176
rect 16546 14116 16550 14172
rect 16550 14116 16606 14172
rect 16606 14116 16610 14172
rect 16546 14112 16610 14116
rect 16626 14172 16690 14176
rect 16626 14116 16630 14172
rect 16630 14116 16686 14172
rect 16686 14116 16690 14172
rect 16626 14112 16690 14116
rect 16706 14172 16770 14176
rect 16706 14116 16710 14172
rect 16710 14116 16766 14172
rect 16766 14116 16770 14172
rect 16706 14112 16770 14116
rect 16786 14172 16850 14176
rect 16786 14116 16790 14172
rect 16790 14116 16846 14172
rect 16846 14116 16850 14172
rect 16786 14112 16850 14116
rect 21744 14172 21808 14176
rect 21744 14116 21748 14172
rect 21748 14116 21804 14172
rect 21804 14116 21808 14172
rect 21744 14112 21808 14116
rect 21824 14172 21888 14176
rect 21824 14116 21828 14172
rect 21828 14116 21884 14172
rect 21884 14116 21888 14172
rect 21824 14112 21888 14116
rect 21904 14172 21968 14176
rect 21904 14116 21908 14172
rect 21908 14116 21964 14172
rect 21964 14116 21968 14172
rect 21904 14112 21968 14116
rect 21984 14172 22048 14176
rect 21984 14116 21988 14172
rect 21988 14116 22044 14172
rect 22044 14116 22048 14172
rect 21984 14112 22048 14116
rect 5580 14104 5644 14108
rect 5580 14048 5630 14104
rect 5630 14048 5644 14104
rect 5580 14044 5644 14048
rect 10364 14044 10428 14108
rect 2268 13772 2332 13836
rect 5028 13772 5092 13836
rect 11100 13772 11164 13836
rect 2636 13636 2700 13700
rect 4476 13636 4540 13700
rect 11836 13772 11900 13836
rect 13492 13832 13556 13836
rect 13492 13776 13506 13832
rect 13506 13776 13556 13832
rect 13492 13772 13556 13776
rect 12940 13636 13004 13700
rect 3551 13628 3615 13632
rect 3551 13572 3555 13628
rect 3555 13572 3611 13628
rect 3611 13572 3615 13628
rect 3551 13568 3615 13572
rect 3631 13628 3695 13632
rect 3631 13572 3635 13628
rect 3635 13572 3691 13628
rect 3691 13572 3695 13628
rect 3631 13568 3695 13572
rect 3711 13628 3775 13632
rect 3711 13572 3715 13628
rect 3715 13572 3771 13628
rect 3771 13572 3775 13628
rect 3711 13568 3775 13572
rect 3791 13628 3855 13632
rect 3791 13572 3795 13628
rect 3795 13572 3851 13628
rect 3851 13572 3855 13628
rect 3791 13568 3855 13572
rect 8749 13628 8813 13632
rect 8749 13572 8753 13628
rect 8753 13572 8809 13628
rect 8809 13572 8813 13628
rect 8749 13568 8813 13572
rect 8829 13628 8893 13632
rect 8829 13572 8833 13628
rect 8833 13572 8889 13628
rect 8889 13572 8893 13628
rect 8829 13568 8893 13572
rect 8909 13628 8973 13632
rect 8909 13572 8913 13628
rect 8913 13572 8969 13628
rect 8969 13572 8973 13628
rect 8909 13568 8973 13572
rect 8989 13628 9053 13632
rect 8989 13572 8993 13628
rect 8993 13572 9049 13628
rect 9049 13572 9053 13628
rect 8989 13568 9053 13572
rect 13947 13628 14011 13632
rect 13947 13572 13951 13628
rect 13951 13572 14007 13628
rect 14007 13572 14011 13628
rect 13947 13568 14011 13572
rect 14027 13628 14091 13632
rect 14027 13572 14031 13628
rect 14031 13572 14087 13628
rect 14087 13572 14091 13628
rect 14027 13568 14091 13572
rect 14107 13628 14171 13632
rect 14107 13572 14111 13628
rect 14111 13572 14167 13628
rect 14167 13572 14171 13628
rect 14107 13568 14171 13572
rect 14187 13628 14251 13632
rect 14187 13572 14191 13628
rect 14191 13572 14247 13628
rect 14247 13572 14251 13628
rect 14187 13568 14251 13572
rect 19145 13628 19209 13632
rect 19145 13572 19149 13628
rect 19149 13572 19205 13628
rect 19205 13572 19209 13628
rect 19145 13568 19209 13572
rect 19225 13628 19289 13632
rect 19225 13572 19229 13628
rect 19229 13572 19285 13628
rect 19285 13572 19289 13628
rect 19225 13568 19289 13572
rect 19305 13628 19369 13632
rect 19305 13572 19309 13628
rect 19309 13572 19365 13628
rect 19365 13572 19369 13628
rect 19305 13568 19369 13572
rect 19385 13628 19449 13632
rect 19385 13572 19389 13628
rect 19389 13572 19445 13628
rect 19445 13572 19449 13628
rect 19385 13568 19449 13572
rect 5580 13500 5644 13564
rect 10732 13560 10796 13564
rect 10732 13504 10782 13560
rect 10782 13504 10796 13560
rect 10732 13500 10796 13504
rect 12756 13500 12820 13564
rect 21588 13364 21652 13428
rect 1716 12956 1780 13020
rect 10916 13092 10980 13156
rect 14596 13092 14660 13156
rect 20484 13092 20548 13156
rect 6150 13084 6214 13088
rect 6150 13028 6154 13084
rect 6154 13028 6210 13084
rect 6210 13028 6214 13084
rect 6150 13024 6214 13028
rect 6230 13084 6294 13088
rect 6230 13028 6234 13084
rect 6234 13028 6290 13084
rect 6290 13028 6294 13084
rect 6230 13024 6294 13028
rect 6310 13084 6374 13088
rect 6310 13028 6314 13084
rect 6314 13028 6370 13084
rect 6370 13028 6374 13084
rect 6310 13024 6374 13028
rect 6390 13084 6454 13088
rect 6390 13028 6394 13084
rect 6394 13028 6450 13084
rect 6450 13028 6454 13084
rect 6390 13024 6454 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 16546 13084 16610 13088
rect 16546 13028 16550 13084
rect 16550 13028 16606 13084
rect 16606 13028 16610 13084
rect 16546 13024 16610 13028
rect 16626 13084 16690 13088
rect 16626 13028 16630 13084
rect 16630 13028 16686 13084
rect 16686 13028 16690 13084
rect 16626 13024 16690 13028
rect 16706 13084 16770 13088
rect 16706 13028 16710 13084
rect 16710 13028 16766 13084
rect 16766 13028 16770 13084
rect 16706 13024 16770 13028
rect 16786 13084 16850 13088
rect 16786 13028 16790 13084
rect 16790 13028 16846 13084
rect 16846 13028 16850 13084
rect 16786 13024 16850 13028
rect 21744 13084 21808 13088
rect 21744 13028 21748 13084
rect 21748 13028 21804 13084
rect 21804 13028 21808 13084
rect 21744 13024 21808 13028
rect 21824 13084 21888 13088
rect 21824 13028 21828 13084
rect 21828 13028 21884 13084
rect 21884 13028 21888 13084
rect 21824 13024 21888 13028
rect 21904 13084 21968 13088
rect 21904 13028 21908 13084
rect 21908 13028 21964 13084
rect 21964 13028 21968 13084
rect 21904 13024 21968 13028
rect 21984 13084 22048 13088
rect 21984 13028 21988 13084
rect 21988 13028 22044 13084
rect 22044 13028 22048 13084
rect 21984 13024 22048 13028
rect 8340 12956 8404 13020
rect 13308 12880 13372 12884
rect 13308 12824 13358 12880
rect 13358 12824 13372 12880
rect 13308 12820 13372 12824
rect 14780 12820 14844 12884
rect 21220 12684 21284 12748
rect 9444 12548 9508 12612
rect 3551 12540 3615 12544
rect 3551 12484 3555 12540
rect 3555 12484 3611 12540
rect 3611 12484 3615 12540
rect 3551 12480 3615 12484
rect 3631 12540 3695 12544
rect 3631 12484 3635 12540
rect 3635 12484 3691 12540
rect 3691 12484 3695 12540
rect 3631 12480 3695 12484
rect 3711 12540 3775 12544
rect 3711 12484 3715 12540
rect 3715 12484 3771 12540
rect 3771 12484 3775 12540
rect 3711 12480 3775 12484
rect 3791 12540 3855 12544
rect 3791 12484 3795 12540
rect 3795 12484 3851 12540
rect 3851 12484 3855 12540
rect 3791 12480 3855 12484
rect 8749 12540 8813 12544
rect 8749 12484 8753 12540
rect 8753 12484 8809 12540
rect 8809 12484 8813 12540
rect 8749 12480 8813 12484
rect 8829 12540 8893 12544
rect 8829 12484 8833 12540
rect 8833 12484 8889 12540
rect 8889 12484 8893 12540
rect 8829 12480 8893 12484
rect 8909 12540 8973 12544
rect 8909 12484 8913 12540
rect 8913 12484 8969 12540
rect 8969 12484 8973 12540
rect 8909 12480 8973 12484
rect 8989 12540 9053 12544
rect 8989 12484 8993 12540
rect 8993 12484 9049 12540
rect 9049 12484 9053 12540
rect 8989 12480 9053 12484
rect 9444 12412 9508 12476
rect 10364 12412 10428 12476
rect 13947 12540 14011 12544
rect 13947 12484 13951 12540
rect 13951 12484 14007 12540
rect 14007 12484 14011 12540
rect 13947 12480 14011 12484
rect 14027 12540 14091 12544
rect 14027 12484 14031 12540
rect 14031 12484 14087 12540
rect 14087 12484 14091 12540
rect 14027 12480 14091 12484
rect 14107 12540 14171 12544
rect 14107 12484 14111 12540
rect 14111 12484 14167 12540
rect 14167 12484 14171 12540
rect 14107 12480 14171 12484
rect 14187 12540 14251 12544
rect 14187 12484 14191 12540
rect 14191 12484 14247 12540
rect 14247 12484 14251 12540
rect 14187 12480 14251 12484
rect 19145 12540 19209 12544
rect 19145 12484 19149 12540
rect 19149 12484 19205 12540
rect 19205 12484 19209 12540
rect 19145 12480 19209 12484
rect 19225 12540 19289 12544
rect 19225 12484 19229 12540
rect 19229 12484 19285 12540
rect 19285 12484 19289 12540
rect 19225 12480 19289 12484
rect 19305 12540 19369 12544
rect 19305 12484 19309 12540
rect 19309 12484 19365 12540
rect 19365 12484 19369 12540
rect 19305 12480 19369 12484
rect 19385 12540 19449 12544
rect 19385 12484 19389 12540
rect 19389 12484 19445 12540
rect 19445 12484 19449 12540
rect 19385 12480 19449 12484
rect 4108 12276 4172 12340
rect 8524 12276 8588 12340
rect 12572 12276 12636 12340
rect 17724 12276 17788 12340
rect 21220 12276 21284 12340
rect 21588 12276 21652 12340
rect 7420 12064 7484 12068
rect 7420 12008 7434 12064
rect 7434 12008 7484 12064
rect 7420 12004 7484 12008
rect 10548 12004 10612 12068
rect 6150 11996 6214 12000
rect 6150 11940 6154 11996
rect 6154 11940 6210 11996
rect 6210 11940 6214 11996
rect 6150 11936 6214 11940
rect 6230 11996 6294 12000
rect 6230 11940 6234 11996
rect 6234 11940 6290 11996
rect 6290 11940 6294 11996
rect 6230 11936 6294 11940
rect 6310 11996 6374 12000
rect 6310 11940 6314 11996
rect 6314 11940 6370 11996
rect 6370 11940 6374 11996
rect 6310 11936 6374 11940
rect 6390 11996 6454 12000
rect 6390 11940 6394 11996
rect 6394 11940 6450 11996
rect 6450 11940 6454 11996
rect 6390 11936 6454 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 5764 11792 5828 11796
rect 11836 11868 11900 11932
rect 5764 11736 5778 11792
rect 5778 11736 5828 11792
rect 5764 11732 5828 11736
rect 16546 11996 16610 12000
rect 16546 11940 16550 11996
rect 16550 11940 16606 11996
rect 16606 11940 16610 11996
rect 16546 11936 16610 11940
rect 16626 11996 16690 12000
rect 16626 11940 16630 11996
rect 16630 11940 16686 11996
rect 16686 11940 16690 11996
rect 16626 11936 16690 11940
rect 16706 11996 16770 12000
rect 16706 11940 16710 11996
rect 16710 11940 16766 11996
rect 16766 11940 16770 11996
rect 16706 11936 16770 11940
rect 16786 11996 16850 12000
rect 16786 11940 16790 11996
rect 16790 11940 16846 11996
rect 16846 11940 16850 11996
rect 16786 11936 16850 11940
rect 21744 11996 21808 12000
rect 21744 11940 21748 11996
rect 21748 11940 21804 11996
rect 21804 11940 21808 11996
rect 21744 11936 21808 11940
rect 21824 11996 21888 12000
rect 21824 11940 21828 11996
rect 21828 11940 21884 11996
rect 21884 11940 21888 11996
rect 21824 11936 21888 11940
rect 21904 11996 21968 12000
rect 21904 11940 21908 11996
rect 21908 11940 21964 11996
rect 21964 11940 21968 11996
rect 21904 11936 21968 11940
rect 21984 11996 22048 12000
rect 21984 11940 21988 11996
rect 21988 11940 22044 11996
rect 22044 11940 22048 11996
rect 21984 11936 22048 11940
rect 17172 11868 17236 11932
rect 4844 11520 4908 11524
rect 4844 11464 4858 11520
rect 4858 11464 4908 11520
rect 4844 11460 4908 11464
rect 7604 11460 7668 11524
rect 9812 11460 9876 11524
rect 10732 11460 10796 11524
rect 15148 11520 15212 11524
rect 15148 11464 15198 11520
rect 15198 11464 15212 11520
rect 15148 11460 15212 11464
rect 15516 11460 15580 11524
rect 3551 11452 3615 11456
rect 3551 11396 3555 11452
rect 3555 11396 3611 11452
rect 3611 11396 3615 11452
rect 3551 11392 3615 11396
rect 3631 11452 3695 11456
rect 3631 11396 3635 11452
rect 3635 11396 3691 11452
rect 3691 11396 3695 11452
rect 3631 11392 3695 11396
rect 3711 11452 3775 11456
rect 3711 11396 3715 11452
rect 3715 11396 3771 11452
rect 3771 11396 3775 11452
rect 3711 11392 3775 11396
rect 3791 11452 3855 11456
rect 3791 11396 3795 11452
rect 3795 11396 3851 11452
rect 3851 11396 3855 11452
rect 3791 11392 3855 11396
rect 8749 11452 8813 11456
rect 8749 11396 8753 11452
rect 8753 11396 8809 11452
rect 8809 11396 8813 11452
rect 8749 11392 8813 11396
rect 8829 11452 8893 11456
rect 8829 11396 8833 11452
rect 8833 11396 8889 11452
rect 8889 11396 8893 11452
rect 8829 11392 8893 11396
rect 8909 11452 8973 11456
rect 8909 11396 8913 11452
rect 8913 11396 8969 11452
rect 8969 11396 8973 11452
rect 8909 11392 8973 11396
rect 8989 11452 9053 11456
rect 8989 11396 8993 11452
rect 8993 11396 9049 11452
rect 9049 11396 9053 11452
rect 8989 11392 9053 11396
rect 13947 11452 14011 11456
rect 13947 11396 13951 11452
rect 13951 11396 14007 11452
rect 14007 11396 14011 11452
rect 13947 11392 14011 11396
rect 14027 11452 14091 11456
rect 14027 11396 14031 11452
rect 14031 11396 14087 11452
rect 14087 11396 14091 11452
rect 14027 11392 14091 11396
rect 14107 11452 14171 11456
rect 14107 11396 14111 11452
rect 14111 11396 14167 11452
rect 14167 11396 14171 11452
rect 14107 11392 14171 11396
rect 14187 11452 14251 11456
rect 14187 11396 14191 11452
rect 14191 11396 14247 11452
rect 14247 11396 14251 11452
rect 14187 11392 14251 11396
rect 19145 11452 19209 11456
rect 19145 11396 19149 11452
rect 19149 11396 19205 11452
rect 19205 11396 19209 11452
rect 19145 11392 19209 11396
rect 19225 11452 19289 11456
rect 19225 11396 19229 11452
rect 19229 11396 19285 11452
rect 19285 11396 19289 11452
rect 19225 11392 19289 11396
rect 19305 11452 19369 11456
rect 19305 11396 19309 11452
rect 19309 11396 19365 11452
rect 19365 11396 19369 11452
rect 19305 11392 19369 11396
rect 19385 11452 19449 11456
rect 19385 11396 19389 11452
rect 19389 11396 19445 11452
rect 19445 11396 19449 11452
rect 19385 11392 19449 11396
rect 5396 11052 5460 11116
rect 9444 11052 9508 11116
rect 6150 10908 6214 10912
rect 6150 10852 6154 10908
rect 6154 10852 6210 10908
rect 6210 10852 6214 10908
rect 6150 10848 6214 10852
rect 6230 10908 6294 10912
rect 6230 10852 6234 10908
rect 6234 10852 6290 10908
rect 6290 10852 6294 10908
rect 6230 10848 6294 10852
rect 6310 10908 6374 10912
rect 6310 10852 6314 10908
rect 6314 10852 6370 10908
rect 6370 10852 6374 10908
rect 6310 10848 6374 10852
rect 6390 10908 6454 10912
rect 6390 10852 6394 10908
rect 6394 10852 6450 10908
rect 6450 10852 6454 10908
rect 6390 10848 6454 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 16546 10908 16610 10912
rect 16546 10852 16550 10908
rect 16550 10852 16606 10908
rect 16606 10852 16610 10908
rect 16546 10848 16610 10852
rect 16626 10908 16690 10912
rect 16626 10852 16630 10908
rect 16630 10852 16686 10908
rect 16686 10852 16690 10908
rect 16626 10848 16690 10852
rect 16706 10908 16770 10912
rect 16706 10852 16710 10908
rect 16710 10852 16766 10908
rect 16766 10852 16770 10908
rect 16706 10848 16770 10852
rect 16786 10908 16850 10912
rect 16786 10852 16790 10908
rect 16790 10852 16846 10908
rect 16846 10852 16850 10908
rect 16786 10848 16850 10852
rect 21744 10908 21808 10912
rect 21744 10852 21748 10908
rect 21748 10852 21804 10908
rect 21804 10852 21808 10908
rect 21744 10848 21808 10852
rect 21824 10908 21888 10912
rect 21824 10852 21828 10908
rect 21828 10852 21884 10908
rect 21884 10852 21888 10908
rect 21824 10848 21888 10852
rect 21904 10908 21968 10912
rect 21904 10852 21908 10908
rect 21908 10852 21964 10908
rect 21964 10852 21968 10908
rect 21904 10848 21968 10852
rect 21984 10908 22048 10912
rect 21984 10852 21988 10908
rect 21988 10852 22044 10908
rect 22044 10852 22048 10908
rect 21984 10848 22048 10852
rect 9444 10780 9508 10844
rect 10180 10780 10244 10844
rect 13124 10780 13188 10844
rect 9996 10644 10060 10708
rect 9628 10372 9692 10436
rect 3551 10364 3615 10368
rect 3551 10308 3555 10364
rect 3555 10308 3611 10364
rect 3611 10308 3615 10364
rect 3551 10304 3615 10308
rect 3631 10364 3695 10368
rect 3631 10308 3635 10364
rect 3635 10308 3691 10364
rect 3691 10308 3695 10364
rect 3631 10304 3695 10308
rect 3711 10364 3775 10368
rect 3711 10308 3715 10364
rect 3715 10308 3771 10364
rect 3771 10308 3775 10364
rect 3711 10304 3775 10308
rect 3791 10364 3855 10368
rect 3791 10308 3795 10364
rect 3795 10308 3851 10364
rect 3851 10308 3855 10364
rect 3791 10304 3855 10308
rect 8749 10364 8813 10368
rect 8749 10308 8753 10364
rect 8753 10308 8809 10364
rect 8809 10308 8813 10364
rect 8749 10304 8813 10308
rect 8829 10364 8893 10368
rect 8829 10308 8833 10364
rect 8833 10308 8889 10364
rect 8889 10308 8893 10364
rect 8829 10304 8893 10308
rect 8909 10364 8973 10368
rect 8909 10308 8913 10364
rect 8913 10308 8969 10364
rect 8969 10308 8973 10364
rect 8909 10304 8973 10308
rect 8989 10364 9053 10368
rect 8989 10308 8993 10364
rect 8993 10308 9049 10364
rect 9049 10308 9053 10364
rect 8989 10304 9053 10308
rect 13947 10364 14011 10368
rect 13947 10308 13951 10364
rect 13951 10308 14007 10364
rect 14007 10308 14011 10364
rect 13947 10304 14011 10308
rect 14027 10364 14091 10368
rect 14027 10308 14031 10364
rect 14031 10308 14087 10364
rect 14087 10308 14091 10364
rect 14027 10304 14091 10308
rect 14107 10364 14171 10368
rect 14107 10308 14111 10364
rect 14111 10308 14167 10364
rect 14167 10308 14171 10364
rect 14107 10304 14171 10308
rect 14187 10364 14251 10368
rect 14187 10308 14191 10364
rect 14191 10308 14247 10364
rect 14247 10308 14251 10364
rect 14187 10304 14251 10308
rect 19145 10364 19209 10368
rect 19145 10308 19149 10364
rect 19149 10308 19205 10364
rect 19205 10308 19209 10364
rect 19145 10304 19209 10308
rect 19225 10364 19289 10368
rect 19225 10308 19229 10364
rect 19229 10308 19285 10364
rect 19285 10308 19289 10364
rect 19225 10304 19289 10308
rect 19305 10364 19369 10368
rect 19305 10308 19309 10364
rect 19309 10308 19365 10364
rect 19365 10308 19369 10364
rect 19305 10304 19369 10308
rect 19385 10364 19449 10368
rect 19385 10308 19389 10364
rect 19389 10308 19445 10364
rect 19445 10308 19449 10364
rect 19385 10304 19449 10308
rect 4660 10236 4724 10300
rect 13124 10236 13188 10300
rect 11100 10100 11164 10164
rect 11836 10100 11900 10164
rect 12940 10100 13004 10164
rect 19748 9964 19812 10028
rect 20116 9964 20180 10028
rect 13676 9888 13740 9892
rect 13676 9832 13690 9888
rect 13690 9832 13740 9888
rect 13676 9828 13740 9832
rect 15332 9828 15396 9892
rect 16252 9828 16316 9892
rect 17908 9828 17972 9892
rect 6150 9820 6214 9824
rect 6150 9764 6154 9820
rect 6154 9764 6210 9820
rect 6210 9764 6214 9820
rect 6150 9760 6214 9764
rect 6230 9820 6294 9824
rect 6230 9764 6234 9820
rect 6234 9764 6290 9820
rect 6290 9764 6294 9820
rect 6230 9760 6294 9764
rect 6310 9820 6374 9824
rect 6310 9764 6314 9820
rect 6314 9764 6370 9820
rect 6370 9764 6374 9820
rect 6310 9760 6374 9764
rect 6390 9820 6454 9824
rect 6390 9764 6394 9820
rect 6394 9764 6450 9820
rect 6450 9764 6454 9820
rect 6390 9760 6454 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 16546 9820 16610 9824
rect 16546 9764 16550 9820
rect 16550 9764 16606 9820
rect 16606 9764 16610 9820
rect 16546 9760 16610 9764
rect 16626 9820 16690 9824
rect 16626 9764 16630 9820
rect 16630 9764 16686 9820
rect 16686 9764 16690 9820
rect 16626 9760 16690 9764
rect 16706 9820 16770 9824
rect 16706 9764 16710 9820
rect 16710 9764 16766 9820
rect 16766 9764 16770 9820
rect 16706 9760 16770 9764
rect 16786 9820 16850 9824
rect 16786 9764 16790 9820
rect 16790 9764 16846 9820
rect 16846 9764 16850 9820
rect 16786 9760 16850 9764
rect 21744 9820 21808 9824
rect 21744 9764 21748 9820
rect 21748 9764 21804 9820
rect 21804 9764 21808 9820
rect 21744 9760 21808 9764
rect 21824 9820 21888 9824
rect 21824 9764 21828 9820
rect 21828 9764 21884 9820
rect 21884 9764 21888 9820
rect 21824 9760 21888 9764
rect 21904 9820 21968 9824
rect 21904 9764 21908 9820
rect 21908 9764 21964 9820
rect 21964 9764 21968 9820
rect 21904 9760 21968 9764
rect 21984 9820 22048 9824
rect 21984 9764 21988 9820
rect 21988 9764 22044 9820
rect 22044 9764 22048 9820
rect 21984 9760 22048 9764
rect 8156 9752 8220 9756
rect 8156 9696 8206 9752
rect 8206 9696 8220 9752
rect 8156 9692 8220 9696
rect 8340 9692 8404 9756
rect 9260 9692 9324 9756
rect 12204 9692 12268 9756
rect 17540 9752 17604 9756
rect 17540 9696 17554 9752
rect 17554 9696 17604 9752
rect 9628 9556 9692 9620
rect 3924 9420 3988 9484
rect 4292 9480 4356 9484
rect 4292 9424 4306 9480
rect 4306 9424 4356 9480
rect 4292 9420 4356 9424
rect 7788 9420 7852 9484
rect 17540 9692 17604 9696
rect 16988 9556 17052 9620
rect 18276 9556 18340 9620
rect 3551 9276 3615 9280
rect 3551 9220 3555 9276
rect 3555 9220 3611 9276
rect 3611 9220 3615 9276
rect 3551 9216 3615 9220
rect 3631 9276 3695 9280
rect 3631 9220 3635 9276
rect 3635 9220 3691 9276
rect 3691 9220 3695 9276
rect 3631 9216 3695 9220
rect 3711 9276 3775 9280
rect 3711 9220 3715 9276
rect 3715 9220 3771 9276
rect 3771 9220 3775 9276
rect 3711 9216 3775 9220
rect 3791 9276 3855 9280
rect 3791 9220 3795 9276
rect 3795 9220 3851 9276
rect 3851 9220 3855 9276
rect 3791 9216 3855 9220
rect 7972 9284 8036 9348
rect 14412 9284 14476 9348
rect 8749 9276 8813 9280
rect 8749 9220 8753 9276
rect 8753 9220 8809 9276
rect 8809 9220 8813 9276
rect 8749 9216 8813 9220
rect 8829 9276 8893 9280
rect 8829 9220 8833 9276
rect 8833 9220 8889 9276
rect 8889 9220 8893 9276
rect 8829 9216 8893 9220
rect 8909 9276 8973 9280
rect 8909 9220 8913 9276
rect 8913 9220 8969 9276
rect 8969 9220 8973 9276
rect 8909 9216 8973 9220
rect 8989 9276 9053 9280
rect 8989 9220 8993 9276
rect 8993 9220 9049 9276
rect 9049 9220 9053 9276
rect 8989 9216 9053 9220
rect 13947 9276 14011 9280
rect 13947 9220 13951 9276
rect 13951 9220 14007 9276
rect 14007 9220 14011 9276
rect 13947 9216 14011 9220
rect 14027 9276 14091 9280
rect 14027 9220 14031 9276
rect 14031 9220 14087 9276
rect 14087 9220 14091 9276
rect 14027 9216 14091 9220
rect 14107 9276 14171 9280
rect 14107 9220 14111 9276
rect 14111 9220 14167 9276
rect 14167 9220 14171 9276
rect 14107 9216 14171 9220
rect 14187 9276 14251 9280
rect 14187 9220 14191 9276
rect 14191 9220 14247 9276
rect 14247 9220 14251 9276
rect 14187 9216 14251 9220
rect 7788 9208 7852 9212
rect 7788 9152 7838 9208
rect 7838 9152 7852 9208
rect 7788 9148 7852 9152
rect 8156 9208 8220 9212
rect 8156 9152 8170 9208
rect 8170 9152 8220 9208
rect 8156 9148 8220 9152
rect 11100 9148 11164 9212
rect 15700 9148 15764 9212
rect 17908 9148 17972 9212
rect 18644 9344 18708 9348
rect 18644 9288 18694 9344
rect 18694 9288 18708 9344
rect 18644 9284 18708 9288
rect 20668 9284 20732 9348
rect 19145 9276 19209 9280
rect 19145 9220 19149 9276
rect 19149 9220 19205 9276
rect 19205 9220 19209 9276
rect 19145 9216 19209 9220
rect 19225 9276 19289 9280
rect 19225 9220 19229 9276
rect 19229 9220 19285 9276
rect 19285 9220 19289 9276
rect 19225 9216 19289 9220
rect 19305 9276 19369 9280
rect 19305 9220 19309 9276
rect 19309 9220 19365 9276
rect 19365 9220 19369 9276
rect 19305 9216 19369 9220
rect 19385 9276 19449 9280
rect 19385 9220 19389 9276
rect 19389 9220 19445 9276
rect 19445 9220 19449 9276
rect 19385 9216 19449 9220
rect 4292 9012 4356 9076
rect 12388 9012 12452 9076
rect 4292 8876 4356 8940
rect 6684 8936 6748 8940
rect 6684 8880 6698 8936
rect 6698 8880 6748 8936
rect 5580 8740 5644 8804
rect 6684 8876 6748 8880
rect 6868 8740 6932 8804
rect 7604 8740 7668 8804
rect 7972 8740 8036 8804
rect 10916 8740 10980 8804
rect 12572 8740 12636 8804
rect 20300 8740 20364 8804
rect 6150 8732 6214 8736
rect 6150 8676 6154 8732
rect 6154 8676 6210 8732
rect 6210 8676 6214 8732
rect 6150 8672 6214 8676
rect 6230 8732 6294 8736
rect 6230 8676 6234 8732
rect 6234 8676 6290 8732
rect 6290 8676 6294 8732
rect 6230 8672 6294 8676
rect 6310 8732 6374 8736
rect 6310 8676 6314 8732
rect 6314 8676 6370 8732
rect 6370 8676 6374 8732
rect 6310 8672 6374 8676
rect 6390 8732 6454 8736
rect 6390 8676 6394 8732
rect 6394 8676 6450 8732
rect 6450 8676 6454 8732
rect 6390 8672 6454 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 16546 8732 16610 8736
rect 16546 8676 16550 8732
rect 16550 8676 16606 8732
rect 16606 8676 16610 8732
rect 16546 8672 16610 8676
rect 16626 8732 16690 8736
rect 16626 8676 16630 8732
rect 16630 8676 16686 8732
rect 16686 8676 16690 8732
rect 16626 8672 16690 8676
rect 16706 8732 16770 8736
rect 16706 8676 16710 8732
rect 16710 8676 16766 8732
rect 16766 8676 16770 8732
rect 16706 8672 16770 8676
rect 16786 8732 16850 8736
rect 16786 8676 16790 8732
rect 16790 8676 16846 8732
rect 16846 8676 16850 8732
rect 16786 8672 16850 8676
rect 21744 8732 21808 8736
rect 21744 8676 21748 8732
rect 21748 8676 21804 8732
rect 21804 8676 21808 8732
rect 21744 8672 21808 8676
rect 21824 8732 21888 8736
rect 21824 8676 21828 8732
rect 21828 8676 21884 8732
rect 21884 8676 21888 8732
rect 21824 8672 21888 8676
rect 21904 8732 21968 8736
rect 21904 8676 21908 8732
rect 21908 8676 21964 8732
rect 21964 8676 21968 8732
rect 21904 8672 21968 8676
rect 21984 8732 22048 8736
rect 21984 8676 21988 8732
rect 21988 8676 22044 8732
rect 22044 8676 22048 8732
rect 21984 8672 22048 8676
rect 6868 8528 6932 8532
rect 6868 8472 6918 8528
rect 6918 8472 6932 8528
rect 6868 8468 6932 8472
rect 7604 8528 7668 8532
rect 7604 8472 7618 8528
rect 7618 8472 7668 8528
rect 7604 8468 7668 8472
rect 14412 8604 14476 8668
rect 15332 8604 15396 8668
rect 13124 8468 13188 8532
rect 3924 8332 3988 8396
rect 2636 8196 2700 8260
rect 10916 8332 10980 8396
rect 19564 8332 19628 8396
rect 7420 8196 7484 8260
rect 3551 8188 3615 8192
rect 3551 8132 3555 8188
rect 3555 8132 3611 8188
rect 3611 8132 3615 8188
rect 3551 8128 3615 8132
rect 3631 8188 3695 8192
rect 3631 8132 3635 8188
rect 3635 8132 3691 8188
rect 3691 8132 3695 8188
rect 3631 8128 3695 8132
rect 3711 8188 3775 8192
rect 3711 8132 3715 8188
rect 3715 8132 3771 8188
rect 3771 8132 3775 8188
rect 3711 8128 3775 8132
rect 3791 8188 3855 8192
rect 3791 8132 3795 8188
rect 3795 8132 3851 8188
rect 3851 8132 3855 8188
rect 3791 8128 3855 8132
rect 8749 8188 8813 8192
rect 8749 8132 8753 8188
rect 8753 8132 8809 8188
rect 8809 8132 8813 8188
rect 8749 8128 8813 8132
rect 8829 8188 8893 8192
rect 8829 8132 8833 8188
rect 8833 8132 8889 8188
rect 8889 8132 8893 8188
rect 8829 8128 8893 8132
rect 8909 8188 8973 8192
rect 8909 8132 8913 8188
rect 8913 8132 8969 8188
rect 8969 8132 8973 8188
rect 8909 8128 8973 8132
rect 8989 8188 9053 8192
rect 8989 8132 8993 8188
rect 8993 8132 9049 8188
rect 9049 8132 9053 8188
rect 8989 8128 9053 8132
rect 10732 8060 10796 8124
rect 4108 7924 4172 7988
rect 10916 7924 10980 7988
rect 9628 7652 9692 7716
rect 9996 7712 10060 7716
rect 9996 7656 10010 7712
rect 10010 7656 10060 7712
rect 9996 7652 10060 7656
rect 15148 8196 15212 8260
rect 17356 8196 17420 8260
rect 18276 8196 18340 8260
rect 13947 8188 14011 8192
rect 13947 8132 13951 8188
rect 13951 8132 14007 8188
rect 14007 8132 14011 8188
rect 13947 8128 14011 8132
rect 14027 8188 14091 8192
rect 14027 8132 14031 8188
rect 14031 8132 14087 8188
rect 14087 8132 14091 8188
rect 14027 8128 14091 8132
rect 14107 8188 14171 8192
rect 14107 8132 14111 8188
rect 14111 8132 14167 8188
rect 14167 8132 14171 8188
rect 14107 8128 14171 8132
rect 14187 8188 14251 8192
rect 14187 8132 14191 8188
rect 14191 8132 14247 8188
rect 14247 8132 14251 8188
rect 14187 8128 14251 8132
rect 19145 8188 19209 8192
rect 19145 8132 19149 8188
rect 19149 8132 19205 8188
rect 19205 8132 19209 8188
rect 19145 8128 19209 8132
rect 19225 8188 19289 8192
rect 19225 8132 19229 8188
rect 19229 8132 19285 8188
rect 19285 8132 19289 8188
rect 19225 8128 19289 8132
rect 19305 8188 19369 8192
rect 19305 8132 19309 8188
rect 19309 8132 19365 8188
rect 19365 8132 19369 8188
rect 19305 8128 19369 8132
rect 19385 8188 19449 8192
rect 19385 8132 19389 8188
rect 19389 8132 19445 8188
rect 19445 8132 19449 8188
rect 19385 8128 19449 8132
rect 17540 7924 17604 7988
rect 14412 7788 14476 7852
rect 20116 7652 20180 7716
rect 6150 7644 6214 7648
rect 6150 7588 6154 7644
rect 6154 7588 6210 7644
rect 6210 7588 6214 7644
rect 6150 7584 6214 7588
rect 6230 7644 6294 7648
rect 6230 7588 6234 7644
rect 6234 7588 6290 7644
rect 6290 7588 6294 7644
rect 6230 7584 6294 7588
rect 6310 7644 6374 7648
rect 6310 7588 6314 7644
rect 6314 7588 6370 7644
rect 6370 7588 6374 7644
rect 6310 7584 6374 7588
rect 6390 7644 6454 7648
rect 6390 7588 6394 7644
rect 6394 7588 6450 7644
rect 6450 7588 6454 7644
rect 6390 7584 6454 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 16546 7644 16610 7648
rect 16546 7588 16550 7644
rect 16550 7588 16606 7644
rect 16606 7588 16610 7644
rect 16546 7584 16610 7588
rect 16626 7644 16690 7648
rect 16626 7588 16630 7644
rect 16630 7588 16686 7644
rect 16686 7588 16690 7644
rect 16626 7584 16690 7588
rect 16706 7644 16770 7648
rect 16706 7588 16710 7644
rect 16710 7588 16766 7644
rect 16766 7588 16770 7644
rect 16706 7584 16770 7588
rect 16786 7644 16850 7648
rect 16786 7588 16790 7644
rect 16790 7588 16846 7644
rect 16846 7588 16850 7644
rect 16786 7584 16850 7588
rect 21744 7644 21808 7648
rect 21744 7588 21748 7644
rect 21748 7588 21804 7644
rect 21804 7588 21808 7644
rect 21744 7584 21808 7588
rect 21824 7644 21888 7648
rect 21824 7588 21828 7644
rect 21828 7588 21884 7644
rect 21884 7588 21888 7644
rect 21824 7584 21888 7588
rect 21904 7644 21968 7648
rect 21904 7588 21908 7644
rect 21908 7588 21964 7644
rect 21964 7588 21968 7644
rect 21904 7584 21968 7588
rect 21984 7644 22048 7648
rect 21984 7588 21988 7644
rect 21988 7588 22044 7644
rect 22044 7588 22048 7644
rect 21984 7584 22048 7588
rect 3551 7100 3615 7104
rect 3551 7044 3555 7100
rect 3555 7044 3611 7100
rect 3611 7044 3615 7100
rect 3551 7040 3615 7044
rect 3631 7100 3695 7104
rect 3631 7044 3635 7100
rect 3635 7044 3691 7100
rect 3691 7044 3695 7100
rect 3631 7040 3695 7044
rect 3711 7100 3775 7104
rect 3711 7044 3715 7100
rect 3715 7044 3771 7100
rect 3771 7044 3775 7100
rect 3711 7040 3775 7044
rect 3791 7100 3855 7104
rect 3791 7044 3795 7100
rect 3795 7044 3851 7100
rect 3851 7044 3855 7100
rect 3791 7040 3855 7044
rect 4476 7032 4540 7036
rect 4476 6976 4490 7032
rect 4490 6976 4540 7032
rect 4476 6972 4540 6976
rect 16068 7108 16132 7172
rect 8749 7100 8813 7104
rect 8749 7044 8753 7100
rect 8753 7044 8809 7100
rect 8809 7044 8813 7100
rect 8749 7040 8813 7044
rect 8829 7100 8893 7104
rect 8829 7044 8833 7100
rect 8833 7044 8889 7100
rect 8889 7044 8893 7100
rect 8829 7040 8893 7044
rect 8909 7100 8973 7104
rect 8909 7044 8913 7100
rect 8913 7044 8969 7100
rect 8969 7044 8973 7100
rect 8909 7040 8973 7044
rect 8989 7100 9053 7104
rect 8989 7044 8993 7100
rect 8993 7044 9049 7100
rect 9049 7044 9053 7100
rect 8989 7040 9053 7044
rect 13947 7100 14011 7104
rect 13947 7044 13951 7100
rect 13951 7044 14007 7100
rect 14007 7044 14011 7100
rect 13947 7040 14011 7044
rect 14027 7100 14091 7104
rect 14027 7044 14031 7100
rect 14031 7044 14087 7100
rect 14087 7044 14091 7100
rect 14027 7040 14091 7044
rect 14107 7100 14171 7104
rect 14107 7044 14111 7100
rect 14111 7044 14167 7100
rect 14167 7044 14171 7100
rect 14107 7040 14171 7044
rect 14187 7100 14251 7104
rect 14187 7044 14191 7100
rect 14191 7044 14247 7100
rect 14247 7044 14251 7100
rect 14187 7040 14251 7044
rect 8156 6972 8220 7036
rect 12020 7032 12084 7036
rect 12020 6976 12034 7032
rect 12034 6976 12084 7032
rect 12020 6972 12084 6976
rect 19145 7100 19209 7104
rect 19145 7044 19149 7100
rect 19149 7044 19205 7100
rect 19205 7044 19209 7100
rect 19145 7040 19209 7044
rect 19225 7100 19289 7104
rect 19225 7044 19229 7100
rect 19229 7044 19285 7100
rect 19285 7044 19289 7100
rect 19225 7040 19289 7044
rect 19305 7100 19369 7104
rect 19305 7044 19309 7100
rect 19309 7044 19365 7100
rect 19365 7044 19369 7100
rect 19305 7040 19369 7044
rect 19385 7100 19449 7104
rect 19385 7044 19389 7100
rect 19389 7044 19445 7100
rect 19445 7044 19449 7100
rect 19385 7040 19449 7044
rect 4108 6836 4172 6900
rect 5580 6836 5644 6900
rect 7788 6836 7852 6900
rect 8156 6836 8220 6900
rect 8524 6836 8588 6900
rect 14964 6836 15028 6900
rect 17724 6836 17788 6900
rect 3372 6564 3436 6628
rect 7604 6564 7668 6628
rect 6150 6556 6214 6560
rect 6150 6500 6154 6556
rect 6154 6500 6210 6556
rect 6210 6500 6214 6556
rect 6150 6496 6214 6500
rect 6230 6556 6294 6560
rect 6230 6500 6234 6556
rect 6234 6500 6290 6556
rect 6290 6500 6294 6556
rect 6230 6496 6294 6500
rect 6310 6556 6374 6560
rect 6310 6500 6314 6556
rect 6314 6500 6370 6556
rect 6370 6500 6374 6556
rect 6310 6496 6374 6500
rect 6390 6556 6454 6560
rect 6390 6500 6394 6556
rect 6394 6500 6450 6556
rect 6450 6500 6454 6556
rect 6390 6496 6454 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 5764 6428 5828 6492
rect 15884 6564 15948 6628
rect 16546 6556 16610 6560
rect 16546 6500 16550 6556
rect 16550 6500 16606 6556
rect 16606 6500 16610 6556
rect 16546 6496 16610 6500
rect 16626 6556 16690 6560
rect 16626 6500 16630 6556
rect 16630 6500 16686 6556
rect 16686 6500 16690 6556
rect 16626 6496 16690 6500
rect 16706 6556 16770 6560
rect 16706 6500 16710 6556
rect 16710 6500 16766 6556
rect 16766 6500 16770 6556
rect 16706 6496 16770 6500
rect 16786 6556 16850 6560
rect 16786 6500 16790 6556
rect 16790 6500 16846 6556
rect 16846 6500 16850 6556
rect 16786 6496 16850 6500
rect 21744 6556 21808 6560
rect 21744 6500 21748 6556
rect 21748 6500 21804 6556
rect 21804 6500 21808 6556
rect 21744 6496 21808 6500
rect 21824 6556 21888 6560
rect 21824 6500 21828 6556
rect 21828 6500 21884 6556
rect 21884 6500 21888 6556
rect 21824 6496 21888 6500
rect 21904 6556 21968 6560
rect 21904 6500 21908 6556
rect 21908 6500 21964 6556
rect 21964 6500 21968 6556
rect 21904 6496 21968 6500
rect 21984 6556 22048 6560
rect 21984 6500 21988 6556
rect 21988 6500 22044 6556
rect 22044 6500 22048 6556
rect 21984 6496 22048 6500
rect 20668 6428 20732 6492
rect 4292 6156 4356 6220
rect 5764 6156 5828 6220
rect 8524 6292 8588 6356
rect 9260 6292 9324 6356
rect 12756 6292 12820 6356
rect 13676 6292 13740 6356
rect 19564 6156 19628 6220
rect 20668 6216 20732 6220
rect 20668 6160 20718 6216
rect 20718 6160 20732 6216
rect 20668 6156 20732 6160
rect 3551 6012 3615 6016
rect 3551 5956 3555 6012
rect 3555 5956 3611 6012
rect 3611 5956 3615 6012
rect 3551 5952 3615 5956
rect 3631 6012 3695 6016
rect 3631 5956 3635 6012
rect 3635 5956 3691 6012
rect 3691 5956 3695 6012
rect 3631 5952 3695 5956
rect 3711 6012 3775 6016
rect 3711 5956 3715 6012
rect 3715 5956 3771 6012
rect 3771 5956 3775 6012
rect 3711 5952 3775 5956
rect 3791 6012 3855 6016
rect 3791 5956 3795 6012
rect 3795 5956 3851 6012
rect 3851 5956 3855 6012
rect 3791 5952 3855 5956
rect 8749 6012 8813 6016
rect 8749 5956 8753 6012
rect 8753 5956 8809 6012
rect 8809 5956 8813 6012
rect 8749 5952 8813 5956
rect 8829 6012 8893 6016
rect 8829 5956 8833 6012
rect 8833 5956 8889 6012
rect 8889 5956 8893 6012
rect 8829 5952 8893 5956
rect 8909 6012 8973 6016
rect 8909 5956 8913 6012
rect 8913 5956 8969 6012
rect 8969 5956 8973 6012
rect 8909 5952 8973 5956
rect 8989 6012 9053 6016
rect 8989 5956 8993 6012
rect 8993 5956 9049 6012
rect 9049 5956 9053 6012
rect 8989 5952 9053 5956
rect 1164 5884 1228 5948
rect 6684 5884 6748 5948
rect 9996 6020 10060 6084
rect 12572 6020 12636 6084
rect 13947 6012 14011 6016
rect 13947 5956 13951 6012
rect 13951 5956 14007 6012
rect 14007 5956 14011 6012
rect 13947 5952 14011 5956
rect 14027 6012 14091 6016
rect 14027 5956 14031 6012
rect 14031 5956 14087 6012
rect 14087 5956 14091 6012
rect 14027 5952 14091 5956
rect 14107 6012 14171 6016
rect 14107 5956 14111 6012
rect 14111 5956 14167 6012
rect 14167 5956 14171 6012
rect 14107 5952 14171 5956
rect 14187 6012 14251 6016
rect 14187 5956 14191 6012
rect 14191 5956 14247 6012
rect 14247 5956 14251 6012
rect 14187 5952 14251 5956
rect 19145 6012 19209 6016
rect 19145 5956 19149 6012
rect 19149 5956 19205 6012
rect 19205 5956 19209 6012
rect 19145 5952 19209 5956
rect 19225 6012 19289 6016
rect 19225 5956 19229 6012
rect 19229 5956 19285 6012
rect 19285 5956 19289 6012
rect 19225 5952 19289 5956
rect 19305 6012 19369 6016
rect 19305 5956 19309 6012
rect 19309 5956 19365 6012
rect 19365 5956 19369 6012
rect 19305 5952 19369 5956
rect 19385 6012 19449 6016
rect 19385 5956 19389 6012
rect 19389 5956 19445 6012
rect 19445 5956 19449 6012
rect 19385 5952 19449 5956
rect 5580 5612 5644 5676
rect 6868 5612 6932 5676
rect 12756 5748 12820 5812
rect 12940 5748 13004 5812
rect 20116 5808 20180 5812
rect 20116 5752 20166 5808
rect 20166 5752 20180 5808
rect 20116 5748 20180 5752
rect 3004 5476 3068 5540
rect 6150 5468 6214 5472
rect 6150 5412 6154 5468
rect 6154 5412 6210 5468
rect 6210 5412 6214 5468
rect 6150 5408 6214 5412
rect 6230 5468 6294 5472
rect 6230 5412 6234 5468
rect 6234 5412 6290 5468
rect 6290 5412 6294 5468
rect 6230 5408 6294 5412
rect 6310 5468 6374 5472
rect 6310 5412 6314 5468
rect 6314 5412 6370 5468
rect 6370 5412 6374 5468
rect 6310 5408 6374 5412
rect 6390 5468 6454 5472
rect 6390 5412 6394 5468
rect 6394 5412 6450 5468
rect 6450 5412 6454 5468
rect 6390 5408 6454 5412
rect 7236 5536 7300 5540
rect 7236 5480 7286 5536
rect 7286 5480 7300 5536
rect 7236 5476 7300 5480
rect 2820 5340 2884 5404
rect 7052 5400 7116 5404
rect 7052 5344 7066 5400
rect 7066 5344 7116 5400
rect 7052 5340 7116 5344
rect 9628 5476 9692 5540
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 16546 5468 16610 5472
rect 16546 5412 16550 5468
rect 16550 5412 16606 5468
rect 16606 5412 16610 5468
rect 16546 5408 16610 5412
rect 16626 5468 16690 5472
rect 16626 5412 16630 5468
rect 16630 5412 16686 5468
rect 16686 5412 16690 5468
rect 16626 5408 16690 5412
rect 16706 5468 16770 5472
rect 16706 5412 16710 5468
rect 16710 5412 16766 5468
rect 16766 5412 16770 5468
rect 16706 5408 16770 5412
rect 16786 5468 16850 5472
rect 16786 5412 16790 5468
rect 16790 5412 16846 5468
rect 16846 5412 16850 5468
rect 16786 5408 16850 5412
rect 21744 5468 21808 5472
rect 21744 5412 21748 5468
rect 21748 5412 21804 5468
rect 21804 5412 21808 5468
rect 21744 5408 21808 5412
rect 21824 5468 21888 5472
rect 21824 5412 21828 5468
rect 21828 5412 21884 5468
rect 21884 5412 21888 5468
rect 21824 5408 21888 5412
rect 21904 5468 21968 5472
rect 21904 5412 21908 5468
rect 21908 5412 21964 5468
rect 21964 5412 21968 5468
rect 21904 5408 21968 5412
rect 21984 5468 22048 5472
rect 21984 5412 21988 5468
rect 21988 5412 22044 5468
rect 22044 5412 22048 5468
rect 21984 5408 22048 5412
rect 10916 5340 10980 5404
rect 3188 5204 3252 5268
rect 8156 5204 8220 5268
rect 5028 4992 5092 4996
rect 5028 4936 5078 4992
rect 5078 4936 5092 4992
rect 5028 4932 5092 4936
rect 9444 4932 9508 4996
rect 3551 4924 3615 4928
rect 3551 4868 3555 4924
rect 3555 4868 3611 4924
rect 3611 4868 3615 4924
rect 3551 4864 3615 4868
rect 3631 4924 3695 4928
rect 3631 4868 3635 4924
rect 3635 4868 3691 4924
rect 3691 4868 3695 4924
rect 3631 4864 3695 4868
rect 3711 4924 3775 4928
rect 3711 4868 3715 4924
rect 3715 4868 3771 4924
rect 3771 4868 3775 4924
rect 3711 4864 3775 4868
rect 3791 4924 3855 4928
rect 3791 4868 3795 4924
rect 3795 4868 3851 4924
rect 3851 4868 3855 4924
rect 3791 4864 3855 4868
rect 8749 4924 8813 4928
rect 8749 4868 8753 4924
rect 8753 4868 8809 4924
rect 8809 4868 8813 4924
rect 8749 4864 8813 4868
rect 8829 4924 8893 4928
rect 8829 4868 8833 4924
rect 8833 4868 8889 4924
rect 8889 4868 8893 4924
rect 8829 4864 8893 4868
rect 8909 4924 8973 4928
rect 8909 4868 8913 4924
rect 8913 4868 8969 4924
rect 8969 4868 8973 4924
rect 8909 4864 8973 4868
rect 8989 4924 9053 4928
rect 8989 4868 8993 4924
rect 8993 4868 9049 4924
rect 9049 4868 9053 4924
rect 8989 4864 9053 4868
rect 13947 4924 14011 4928
rect 13947 4868 13951 4924
rect 13951 4868 14007 4924
rect 14007 4868 14011 4924
rect 13947 4864 14011 4868
rect 14027 4924 14091 4928
rect 14027 4868 14031 4924
rect 14031 4868 14087 4924
rect 14087 4868 14091 4924
rect 14027 4864 14091 4868
rect 14107 4924 14171 4928
rect 14107 4868 14111 4924
rect 14111 4868 14167 4924
rect 14167 4868 14171 4924
rect 14107 4864 14171 4868
rect 14187 4924 14251 4928
rect 14187 4868 14191 4924
rect 14191 4868 14247 4924
rect 14247 4868 14251 4924
rect 14187 4864 14251 4868
rect 19145 4924 19209 4928
rect 19145 4868 19149 4924
rect 19149 4868 19205 4924
rect 19205 4868 19209 4924
rect 19145 4864 19209 4868
rect 19225 4924 19289 4928
rect 19225 4868 19229 4924
rect 19229 4868 19285 4924
rect 19285 4868 19289 4924
rect 19225 4864 19289 4868
rect 19305 4924 19369 4928
rect 19305 4868 19309 4924
rect 19309 4868 19365 4924
rect 19365 4868 19369 4924
rect 19305 4864 19369 4868
rect 19385 4924 19449 4928
rect 19385 4868 19389 4924
rect 19389 4868 19445 4924
rect 19445 4868 19449 4924
rect 19385 4864 19449 4868
rect 5212 4796 5276 4860
rect 5948 4796 6012 4860
rect 12204 4796 12268 4860
rect 15332 4796 15396 4860
rect 2268 4660 2332 4724
rect 14412 4720 14476 4724
rect 14412 4664 14462 4720
rect 14462 4664 14476 4720
rect 14412 4660 14476 4664
rect 13124 4524 13188 4588
rect 17908 4524 17972 4588
rect 4292 4388 4356 4452
rect 5396 4388 5460 4452
rect 5948 4448 6012 4452
rect 5948 4392 5962 4448
rect 5962 4392 6012 4448
rect 5948 4388 6012 4392
rect 9260 4388 9324 4452
rect 18644 4388 18708 4452
rect 6150 4380 6214 4384
rect 6150 4324 6154 4380
rect 6154 4324 6210 4380
rect 6210 4324 6214 4380
rect 6150 4320 6214 4324
rect 6230 4380 6294 4384
rect 6230 4324 6234 4380
rect 6234 4324 6290 4380
rect 6290 4324 6294 4380
rect 6230 4320 6294 4324
rect 6310 4380 6374 4384
rect 6310 4324 6314 4380
rect 6314 4324 6370 4380
rect 6370 4324 6374 4380
rect 6310 4320 6374 4324
rect 6390 4380 6454 4384
rect 6390 4324 6394 4380
rect 6394 4324 6450 4380
rect 6450 4324 6454 4380
rect 6390 4320 6454 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 16546 4380 16610 4384
rect 16546 4324 16550 4380
rect 16550 4324 16606 4380
rect 16606 4324 16610 4380
rect 16546 4320 16610 4324
rect 16626 4380 16690 4384
rect 16626 4324 16630 4380
rect 16630 4324 16686 4380
rect 16686 4324 16690 4380
rect 16626 4320 16690 4324
rect 16706 4380 16770 4384
rect 16706 4324 16710 4380
rect 16710 4324 16766 4380
rect 16766 4324 16770 4380
rect 16706 4320 16770 4324
rect 16786 4380 16850 4384
rect 16786 4324 16790 4380
rect 16790 4324 16846 4380
rect 16846 4324 16850 4380
rect 16786 4320 16850 4324
rect 21744 4380 21808 4384
rect 21744 4324 21748 4380
rect 21748 4324 21804 4380
rect 21804 4324 21808 4380
rect 21744 4320 21808 4324
rect 21824 4380 21888 4384
rect 21824 4324 21828 4380
rect 21828 4324 21884 4380
rect 21884 4324 21888 4380
rect 21824 4320 21888 4324
rect 21904 4380 21968 4384
rect 21904 4324 21908 4380
rect 21908 4324 21964 4380
rect 21964 4324 21968 4380
rect 21904 4320 21968 4324
rect 21984 4380 22048 4384
rect 21984 4324 21988 4380
rect 21988 4324 22044 4380
rect 22044 4324 22048 4380
rect 21984 4320 22048 4324
rect 980 4252 1044 4316
rect 1716 4312 1780 4316
rect 1716 4256 1766 4312
rect 1766 4256 1780 4312
rect 1716 4252 1780 4256
rect 8524 4312 8588 4316
rect 8524 4256 8538 4312
rect 8538 4256 8588 4312
rect 8524 4252 8588 4256
rect 9444 4252 9508 4316
rect 5764 3980 5828 4044
rect 8340 3980 8404 4044
rect 6684 3844 6748 3908
rect 7236 3844 7300 3908
rect 19932 3844 19996 3908
rect 3551 3836 3615 3840
rect 3551 3780 3555 3836
rect 3555 3780 3611 3836
rect 3611 3780 3615 3836
rect 3551 3776 3615 3780
rect 3631 3836 3695 3840
rect 3631 3780 3635 3836
rect 3635 3780 3691 3836
rect 3691 3780 3695 3836
rect 3631 3776 3695 3780
rect 3711 3836 3775 3840
rect 3711 3780 3715 3836
rect 3715 3780 3771 3836
rect 3771 3780 3775 3836
rect 3711 3776 3775 3780
rect 3791 3836 3855 3840
rect 3791 3780 3795 3836
rect 3795 3780 3851 3836
rect 3851 3780 3855 3836
rect 3791 3776 3855 3780
rect 8749 3836 8813 3840
rect 8749 3780 8753 3836
rect 8753 3780 8809 3836
rect 8809 3780 8813 3836
rect 8749 3776 8813 3780
rect 8829 3836 8893 3840
rect 8829 3780 8833 3836
rect 8833 3780 8889 3836
rect 8889 3780 8893 3836
rect 8829 3776 8893 3780
rect 8909 3836 8973 3840
rect 8909 3780 8913 3836
rect 8913 3780 8969 3836
rect 8969 3780 8973 3836
rect 8909 3776 8973 3780
rect 8989 3836 9053 3840
rect 8989 3780 8993 3836
rect 8993 3780 9049 3836
rect 9049 3780 9053 3836
rect 8989 3776 9053 3780
rect 13947 3836 14011 3840
rect 13947 3780 13951 3836
rect 13951 3780 14007 3836
rect 14007 3780 14011 3836
rect 13947 3776 14011 3780
rect 14027 3836 14091 3840
rect 14027 3780 14031 3836
rect 14031 3780 14087 3836
rect 14087 3780 14091 3836
rect 14027 3776 14091 3780
rect 14107 3836 14171 3840
rect 14107 3780 14111 3836
rect 14111 3780 14167 3836
rect 14167 3780 14171 3836
rect 14107 3776 14171 3780
rect 14187 3836 14251 3840
rect 14187 3780 14191 3836
rect 14191 3780 14247 3836
rect 14247 3780 14251 3836
rect 14187 3776 14251 3780
rect 19145 3836 19209 3840
rect 19145 3780 19149 3836
rect 19149 3780 19205 3836
rect 19205 3780 19209 3836
rect 19145 3776 19209 3780
rect 19225 3836 19289 3840
rect 19225 3780 19229 3836
rect 19229 3780 19285 3836
rect 19285 3780 19289 3836
rect 19225 3776 19289 3780
rect 19305 3836 19369 3840
rect 19305 3780 19309 3836
rect 19309 3780 19365 3836
rect 19365 3780 19369 3836
rect 19305 3776 19369 3780
rect 19385 3836 19449 3840
rect 19385 3780 19389 3836
rect 19389 3780 19445 3836
rect 19445 3780 19449 3836
rect 19385 3776 19449 3780
rect 17172 3708 17236 3772
rect 19748 3708 19812 3772
rect 3924 3436 3988 3500
rect 6868 3572 6932 3636
rect 12940 3572 13004 3636
rect 6684 3436 6748 3500
rect 3372 3164 3436 3228
rect 4660 3164 4724 3228
rect 5396 3028 5460 3092
rect 6150 3292 6214 3296
rect 6150 3236 6154 3292
rect 6154 3236 6210 3292
rect 6210 3236 6214 3292
rect 6150 3232 6214 3236
rect 6230 3292 6294 3296
rect 6230 3236 6234 3292
rect 6234 3236 6290 3292
rect 6290 3236 6294 3292
rect 6230 3232 6294 3236
rect 6310 3292 6374 3296
rect 6310 3236 6314 3292
rect 6314 3236 6370 3292
rect 6370 3236 6374 3292
rect 6310 3232 6374 3236
rect 6390 3292 6454 3296
rect 6390 3236 6394 3292
rect 6394 3236 6450 3292
rect 6450 3236 6454 3292
rect 6390 3232 6454 3236
rect 7420 3164 7484 3228
rect 17356 3360 17420 3364
rect 17356 3304 17370 3360
rect 17370 3304 17420 3360
rect 17356 3300 17420 3304
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 16546 3292 16610 3296
rect 16546 3236 16550 3292
rect 16550 3236 16606 3292
rect 16606 3236 16610 3292
rect 16546 3232 16610 3236
rect 16626 3292 16690 3296
rect 16626 3236 16630 3292
rect 16630 3236 16686 3292
rect 16686 3236 16690 3292
rect 16626 3232 16690 3236
rect 16706 3292 16770 3296
rect 16706 3236 16710 3292
rect 16710 3236 16766 3292
rect 16766 3236 16770 3292
rect 16706 3232 16770 3236
rect 16786 3292 16850 3296
rect 16786 3236 16790 3292
rect 16790 3236 16846 3292
rect 16846 3236 16850 3292
rect 16786 3232 16850 3236
rect 21744 3292 21808 3296
rect 21744 3236 21748 3292
rect 21748 3236 21804 3292
rect 21804 3236 21808 3292
rect 21744 3232 21808 3236
rect 21824 3292 21888 3296
rect 21824 3236 21828 3292
rect 21828 3236 21884 3292
rect 21884 3236 21888 3292
rect 21824 3232 21888 3236
rect 21904 3292 21968 3296
rect 21904 3236 21908 3292
rect 21908 3236 21964 3292
rect 21964 3236 21968 3292
rect 21904 3232 21968 3236
rect 21984 3292 22048 3296
rect 21984 3236 21988 3292
rect 21988 3236 22044 3292
rect 22044 3236 22048 3292
rect 21984 3232 22048 3236
rect 15884 3028 15948 3092
rect 16988 3088 17052 3092
rect 16988 3032 17002 3088
rect 17002 3032 17052 3088
rect 16988 3028 17052 3032
rect 7972 2892 8036 2956
rect 3004 2756 3068 2820
rect 3372 2756 3436 2820
rect 5028 2756 5092 2820
rect 6868 2816 6932 2820
rect 6868 2760 6882 2816
rect 6882 2760 6932 2816
rect 6868 2756 6932 2760
rect 7420 2816 7484 2820
rect 7420 2760 7470 2816
rect 7470 2760 7484 2816
rect 7420 2756 7484 2760
rect 3551 2748 3615 2752
rect 3551 2692 3555 2748
rect 3555 2692 3611 2748
rect 3611 2692 3615 2748
rect 3551 2688 3615 2692
rect 3631 2748 3695 2752
rect 3631 2692 3635 2748
rect 3635 2692 3691 2748
rect 3691 2692 3695 2748
rect 3631 2688 3695 2692
rect 3711 2748 3775 2752
rect 3711 2692 3715 2748
rect 3715 2692 3771 2748
rect 3771 2692 3775 2748
rect 3711 2688 3775 2692
rect 3791 2748 3855 2752
rect 3791 2692 3795 2748
rect 3795 2692 3851 2748
rect 3851 2692 3855 2748
rect 3791 2688 3855 2692
rect 8749 2748 8813 2752
rect 8749 2692 8753 2748
rect 8753 2692 8809 2748
rect 8809 2692 8813 2748
rect 8749 2688 8813 2692
rect 8829 2748 8893 2752
rect 8829 2692 8833 2748
rect 8833 2692 8889 2748
rect 8889 2692 8893 2748
rect 8829 2688 8893 2692
rect 8909 2748 8973 2752
rect 8909 2692 8913 2748
rect 8913 2692 8969 2748
rect 8969 2692 8973 2748
rect 8909 2688 8973 2692
rect 8989 2748 9053 2752
rect 8989 2692 8993 2748
rect 8993 2692 9049 2748
rect 9049 2692 9053 2748
rect 8989 2688 9053 2692
rect 13947 2748 14011 2752
rect 13947 2692 13951 2748
rect 13951 2692 14007 2748
rect 14007 2692 14011 2748
rect 13947 2688 14011 2692
rect 14027 2748 14091 2752
rect 14027 2692 14031 2748
rect 14031 2692 14087 2748
rect 14087 2692 14091 2748
rect 14027 2688 14091 2692
rect 14107 2748 14171 2752
rect 14107 2692 14111 2748
rect 14111 2692 14167 2748
rect 14167 2692 14171 2748
rect 14107 2688 14171 2692
rect 14187 2748 14251 2752
rect 14187 2692 14191 2748
rect 14191 2692 14247 2748
rect 14247 2692 14251 2748
rect 14187 2688 14251 2692
rect 19145 2748 19209 2752
rect 19145 2692 19149 2748
rect 19149 2692 19205 2748
rect 19205 2692 19209 2748
rect 19145 2688 19209 2692
rect 19225 2748 19289 2752
rect 19225 2692 19229 2748
rect 19229 2692 19285 2748
rect 19285 2692 19289 2748
rect 19225 2688 19289 2692
rect 19305 2748 19369 2752
rect 19305 2692 19309 2748
rect 19309 2692 19365 2748
rect 19365 2692 19369 2748
rect 19305 2688 19369 2692
rect 19385 2748 19449 2752
rect 19385 2692 19389 2748
rect 19389 2692 19445 2748
rect 19445 2692 19449 2748
rect 19385 2688 19449 2692
rect 4476 2620 4540 2684
rect 7052 2620 7116 2684
rect 12572 2620 12636 2684
rect 20484 2680 20548 2684
rect 20484 2624 20534 2680
rect 20534 2624 20548 2680
rect 20484 2620 20548 2624
rect 1348 2484 1412 2548
rect 3372 2484 3436 2548
rect 6684 2484 6748 2548
rect 5396 2348 5460 2412
rect 12204 2484 12268 2548
rect 16252 2484 16316 2548
rect 5948 2272 6012 2276
rect 5948 2216 5962 2272
rect 5962 2216 6012 2272
rect 5948 2212 6012 2216
rect 6150 2204 6214 2208
rect 6150 2148 6154 2204
rect 6154 2148 6210 2204
rect 6210 2148 6214 2204
rect 6150 2144 6214 2148
rect 6230 2204 6294 2208
rect 6230 2148 6234 2204
rect 6234 2148 6290 2204
rect 6290 2148 6294 2204
rect 6230 2144 6294 2148
rect 6310 2204 6374 2208
rect 6310 2148 6314 2204
rect 6314 2148 6370 2204
rect 6370 2148 6374 2204
rect 6310 2144 6374 2148
rect 6390 2204 6454 2208
rect 6390 2148 6394 2204
rect 6394 2148 6450 2204
rect 6450 2148 6454 2204
rect 6390 2144 6454 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 16546 2204 16610 2208
rect 16546 2148 16550 2204
rect 16550 2148 16606 2204
rect 16606 2148 16610 2204
rect 16546 2144 16610 2148
rect 16626 2204 16690 2208
rect 16626 2148 16630 2204
rect 16630 2148 16686 2204
rect 16686 2148 16690 2204
rect 16626 2144 16690 2148
rect 16706 2204 16770 2208
rect 16706 2148 16710 2204
rect 16710 2148 16766 2204
rect 16766 2148 16770 2204
rect 16706 2144 16770 2148
rect 16786 2204 16850 2208
rect 16786 2148 16790 2204
rect 16790 2148 16846 2204
rect 16846 2148 16850 2204
rect 16786 2144 16850 2148
rect 21744 2204 21808 2208
rect 21744 2148 21748 2204
rect 21748 2148 21804 2204
rect 21804 2148 21808 2204
rect 21744 2144 21808 2148
rect 21824 2204 21888 2208
rect 21824 2148 21828 2204
rect 21828 2148 21884 2204
rect 21884 2148 21888 2204
rect 21824 2144 21888 2148
rect 21904 2204 21968 2208
rect 21904 2148 21908 2204
rect 21908 2148 21964 2204
rect 21964 2148 21968 2204
rect 21904 2144 21968 2148
rect 21984 2204 22048 2208
rect 21984 2148 21988 2204
rect 21988 2148 22044 2204
rect 22044 2148 22048 2204
rect 21984 2144 22048 2148
rect 7788 2076 7852 2140
rect 4660 1804 4724 1868
rect 5580 1864 5644 1868
rect 5580 1808 5594 1864
rect 5594 1808 5644 1864
rect 5580 1804 5644 1808
rect 13308 1940 13372 2004
rect 4844 1668 4908 1732
rect 3188 1532 3252 1596
rect 11100 1124 11164 1188
rect 14596 1124 14660 1188
rect 13492 988 13556 1052
rect 16068 988 16132 1052
rect 5212 716 5276 780
rect 14780 36 14844 100
<< metal4 >>
rect 59 22540 125 22541
rect 59 22476 60 22540
rect 124 22476 125 22540
rect 59 22475 125 22476
rect 14411 22540 14477 22541
rect 14411 22476 14412 22540
rect 14476 22476 14477 22540
rect 14411 22475 14477 22476
rect 62 16590 122 22475
rect 12755 21316 12821 21317
rect 12755 21252 12756 21316
rect 12820 21252 12821 21316
rect 12755 21251 12821 21252
rect 1163 21180 1229 21181
rect 1163 21116 1164 21180
rect 1228 21116 1229 21180
rect 1163 21115 1229 21116
rect 1166 16590 1226 21115
rect 4843 21044 4909 21045
rect 4843 20980 4844 21044
rect 4908 20980 4909 21044
rect 4843 20979 4909 20980
rect 2451 20228 2517 20229
rect 2451 20164 2452 20228
rect 2516 20164 2517 20228
rect 2451 20163 2517 20164
rect 62 16530 1042 16590
rect 1166 16530 1410 16590
rect 982 4317 1042 16530
rect 1163 14380 1229 14381
rect 1163 14316 1164 14380
rect 1228 14316 1229 14380
rect 1163 14315 1229 14316
rect 1166 5949 1226 14315
rect 1163 5948 1229 5949
rect 1163 5884 1164 5948
rect 1228 5884 1229 5948
rect 1163 5883 1229 5884
rect 979 4316 1045 4317
rect 979 4252 980 4316
rect 1044 4252 1045 4316
rect 979 4251 1045 4252
rect 1350 2549 1410 16530
rect 2267 13836 2333 13837
rect 2267 13772 2268 13836
rect 2332 13772 2333 13836
rect 2267 13771 2333 13772
rect 1715 13020 1781 13021
rect 1715 12956 1716 13020
rect 1780 12956 1781 13020
rect 1715 12955 1781 12956
rect 1718 4317 1778 12955
rect 2270 4725 2330 13771
rect 2454 7850 2514 20163
rect 3543 20160 3863 20720
rect 3543 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3863 20160
rect 3543 19072 3863 20096
rect 4475 19548 4541 19549
rect 4475 19484 4476 19548
rect 4540 19484 4541 19548
rect 4475 19483 4541 19484
rect 3543 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3863 19072
rect 3543 17984 3863 19008
rect 4107 18052 4173 18053
rect 4107 17988 4108 18052
rect 4172 17988 4173 18052
rect 4107 17987 4173 17988
rect 3543 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3863 17984
rect 3371 17236 3437 17237
rect 3371 17172 3372 17236
rect 3436 17172 3437 17236
rect 3371 17171 3437 17172
rect 2635 13700 2701 13701
rect 2635 13636 2636 13700
rect 2700 13636 2701 13700
rect 2635 13635 2701 13636
rect 2638 8261 2698 13635
rect 3374 12450 3434 17171
rect 3006 12390 3434 12450
rect 3543 16896 3863 17920
rect 3923 17372 3989 17373
rect 3923 17308 3924 17372
rect 3988 17308 3989 17372
rect 3923 17307 3989 17308
rect 3543 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3863 16896
rect 3543 15808 3863 16832
rect 3543 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3863 15808
rect 3543 14720 3863 15744
rect 3926 14925 3986 17307
rect 3923 14924 3989 14925
rect 3923 14860 3924 14924
rect 3988 14860 3989 14924
rect 3923 14859 3989 14860
rect 3543 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3863 14720
rect 3543 13632 3863 14656
rect 3543 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3863 13632
rect 3543 12544 3863 13568
rect 3543 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3863 12544
rect 2635 8260 2701 8261
rect 2635 8196 2636 8260
rect 2700 8196 2701 8260
rect 2635 8195 2701 8196
rect 2454 7790 2882 7850
rect 2822 5405 2882 7790
rect 3006 5541 3066 12390
rect 3543 11456 3863 12480
rect 3543 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3863 11456
rect 3543 10368 3863 11392
rect 3543 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3863 10368
rect 3543 9280 3863 10304
rect 3926 9485 3986 14859
rect 4110 12341 4170 17987
rect 4478 13701 4538 19483
rect 4475 13700 4541 13701
rect 4475 13636 4476 13700
rect 4540 13636 4541 13700
rect 4475 13635 4541 13636
rect 4107 12340 4173 12341
rect 4107 12276 4108 12340
rect 4172 12276 4173 12340
rect 4107 12275 4173 12276
rect 3923 9484 3989 9485
rect 3923 9420 3924 9484
rect 3988 9420 3989 9484
rect 3923 9419 3989 9420
rect 3543 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3863 9280
rect 3543 8192 3863 9216
rect 3923 8396 3989 8397
rect 3923 8332 3924 8396
rect 3988 8332 3989 8396
rect 3923 8331 3989 8332
rect 3543 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3863 8192
rect 3543 7104 3863 8128
rect 3543 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3863 7104
rect 3371 6628 3437 6629
rect 3371 6564 3372 6628
rect 3436 6564 3437 6628
rect 3371 6563 3437 6564
rect 3003 5540 3069 5541
rect 3003 5476 3004 5540
rect 3068 5476 3069 5540
rect 3003 5475 3069 5476
rect 2819 5404 2885 5405
rect 2819 5340 2820 5404
rect 2884 5340 2885 5404
rect 2819 5339 2885 5340
rect 2267 4724 2333 4725
rect 2267 4660 2268 4724
rect 2332 4660 2333 4724
rect 2267 4659 2333 4660
rect 1715 4316 1781 4317
rect 1715 4252 1716 4316
rect 1780 4252 1781 4316
rect 1715 4251 1781 4252
rect 3006 2821 3066 5475
rect 3187 5268 3253 5269
rect 3187 5204 3188 5268
rect 3252 5204 3253 5268
rect 3187 5203 3253 5204
rect 3003 2820 3069 2821
rect 3003 2756 3004 2820
rect 3068 2756 3069 2820
rect 3003 2755 3069 2756
rect 1347 2548 1413 2549
rect 1347 2484 1348 2548
rect 1412 2484 1413 2548
rect 1347 2483 1413 2484
rect 3190 1597 3250 5203
rect 3374 3229 3434 6563
rect 3543 6016 3863 7040
rect 3543 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3863 6016
rect 3543 4928 3863 5952
rect 3543 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3863 4928
rect 3543 3840 3863 4864
rect 3543 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3863 3840
rect 3371 3228 3437 3229
rect 3371 3164 3372 3228
rect 3436 3164 3437 3228
rect 3371 3163 3437 3164
rect 3371 2820 3437 2821
rect 3371 2756 3372 2820
rect 3436 2756 3437 2820
rect 3371 2755 3437 2756
rect 3374 2549 3434 2755
rect 3543 2752 3863 3776
rect 3926 3501 3986 8331
rect 4110 7989 4170 12275
rect 4291 9484 4357 9485
rect 4291 9420 4292 9484
rect 4356 9420 4357 9484
rect 4291 9419 4357 9420
rect 4294 9077 4354 9419
rect 4291 9076 4357 9077
rect 4291 9012 4292 9076
rect 4356 9012 4357 9076
rect 4291 9011 4357 9012
rect 4291 8940 4357 8941
rect 4291 8876 4292 8940
rect 4356 8876 4357 8940
rect 4291 8875 4357 8876
rect 4107 7988 4173 7989
rect 4107 7924 4108 7988
rect 4172 7924 4173 7988
rect 4107 7923 4173 7924
rect 4294 6930 4354 8875
rect 4478 7037 4538 13635
rect 4846 11525 4906 20979
rect 8155 20908 8221 20909
rect 8155 20844 8156 20908
rect 8220 20844 8221 20908
rect 8155 20843 8221 20844
rect 6142 20704 6462 20720
rect 6142 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6462 20704
rect 6142 19616 6462 20640
rect 6142 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6462 19616
rect 5763 18868 5829 18869
rect 5763 18804 5764 18868
rect 5828 18804 5829 18868
rect 5763 18803 5829 18804
rect 5579 18460 5645 18461
rect 5579 18396 5580 18460
rect 5644 18396 5645 18460
rect 5579 18395 5645 18396
rect 5582 14109 5642 18395
rect 5766 18325 5826 18803
rect 6142 18528 6462 19552
rect 7419 19412 7485 19413
rect 7419 19348 7420 19412
rect 7484 19348 7485 19412
rect 7419 19347 7485 19348
rect 7787 19412 7853 19413
rect 7787 19348 7788 19412
rect 7852 19348 7853 19412
rect 7787 19347 7853 19348
rect 6142 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6462 18528
rect 5763 18324 5829 18325
rect 5763 18260 5764 18324
rect 5828 18260 5829 18324
rect 5763 18259 5829 18260
rect 6142 17440 6462 18464
rect 6683 17508 6749 17509
rect 6683 17444 6684 17508
rect 6748 17444 6749 17508
rect 6683 17443 6749 17444
rect 6142 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6462 17440
rect 6142 16352 6462 17376
rect 6142 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6462 16352
rect 5947 15332 6013 15333
rect 5947 15268 5948 15332
rect 6012 15268 6013 15332
rect 5947 15267 6013 15268
rect 5579 14108 5645 14109
rect 5579 14044 5580 14108
rect 5644 14044 5645 14108
rect 5579 14043 5645 14044
rect 5027 13836 5093 13837
rect 5027 13772 5028 13836
rect 5092 13772 5093 13836
rect 5027 13771 5093 13772
rect 4843 11524 4909 11525
rect 4843 11460 4844 11524
rect 4908 11460 4909 11524
rect 4843 11459 4909 11460
rect 4659 10300 4725 10301
rect 4659 10236 4660 10300
rect 4724 10236 4725 10300
rect 4659 10235 4725 10236
rect 4475 7036 4541 7037
rect 4475 6972 4476 7036
rect 4540 6972 4541 7036
rect 4475 6971 4541 6972
rect 4110 6901 4354 6930
rect 4107 6900 4354 6901
rect 4107 6836 4108 6900
rect 4172 6870 4354 6900
rect 4172 6836 4173 6870
rect 4107 6835 4173 6836
rect 4291 6220 4357 6221
rect 4291 6156 4292 6220
rect 4356 6156 4357 6220
rect 4291 6155 4357 6156
rect 4294 4453 4354 6155
rect 4291 4452 4357 4453
rect 4291 4388 4292 4452
rect 4356 4388 4357 4452
rect 4291 4387 4357 4388
rect 3923 3500 3989 3501
rect 3923 3436 3924 3500
rect 3988 3436 3989 3500
rect 4662 3498 4722 10235
rect 3923 3435 3989 3436
rect 4478 3438 4722 3498
rect 3543 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3863 2752
rect 3371 2548 3437 2549
rect 3371 2484 3372 2548
rect 3436 2484 3437 2548
rect 3371 2483 3437 2484
rect 3543 2128 3863 2688
rect 4478 2685 4538 3438
rect 4659 3228 4725 3229
rect 4659 3164 4660 3228
rect 4724 3164 4725 3228
rect 4659 3163 4725 3164
rect 4475 2684 4541 2685
rect 4475 2620 4476 2684
rect 4540 2620 4541 2684
rect 4475 2619 4541 2620
rect 4662 1869 4722 3163
rect 4659 1868 4725 1869
rect 4659 1804 4660 1868
rect 4724 1804 4725 1868
rect 4659 1803 4725 1804
rect 4846 1733 4906 11459
rect 5030 4997 5090 13771
rect 5579 13564 5645 13565
rect 5579 13500 5580 13564
rect 5644 13500 5645 13564
rect 5579 13499 5645 13500
rect 5395 11116 5461 11117
rect 5395 11052 5396 11116
rect 5460 11052 5461 11116
rect 5395 11051 5461 11052
rect 5027 4996 5093 4997
rect 5027 4932 5028 4996
rect 5092 4932 5093 4996
rect 5027 4931 5093 4932
rect 5030 2821 5090 4931
rect 5211 4860 5277 4861
rect 5211 4796 5212 4860
rect 5276 4796 5277 4860
rect 5211 4795 5277 4796
rect 5027 2820 5093 2821
rect 5027 2756 5028 2820
rect 5092 2756 5093 2820
rect 5027 2755 5093 2756
rect 4843 1732 4909 1733
rect 4843 1668 4844 1732
rect 4908 1668 4909 1732
rect 4843 1667 4909 1668
rect 3187 1596 3253 1597
rect 3187 1532 3188 1596
rect 3252 1532 3253 1596
rect 3187 1531 3253 1532
rect 5214 781 5274 4795
rect 5398 4453 5458 11051
rect 5582 8805 5642 13499
rect 5763 11796 5829 11797
rect 5763 11732 5764 11796
rect 5828 11732 5829 11796
rect 5763 11731 5829 11732
rect 5579 8804 5645 8805
rect 5579 8740 5580 8804
rect 5644 8740 5645 8804
rect 5579 8739 5645 8740
rect 5579 6900 5645 6901
rect 5579 6836 5580 6900
rect 5644 6836 5645 6900
rect 5579 6835 5645 6836
rect 5582 5946 5642 6835
rect 5766 6493 5826 11731
rect 5763 6492 5829 6493
rect 5763 6428 5764 6492
rect 5828 6428 5829 6492
rect 5763 6427 5829 6428
rect 5766 6221 5826 6427
rect 5763 6220 5829 6221
rect 5763 6156 5764 6220
rect 5828 6156 5829 6220
rect 5763 6155 5829 6156
rect 5582 5886 5826 5946
rect 5579 5676 5645 5677
rect 5579 5612 5580 5676
rect 5644 5612 5645 5676
rect 5579 5611 5645 5612
rect 5395 4452 5461 4453
rect 5395 4388 5396 4452
rect 5460 4388 5461 4452
rect 5395 4387 5461 4388
rect 5395 3092 5461 3093
rect 5395 3028 5396 3092
rect 5460 3028 5461 3092
rect 5395 3027 5461 3028
rect 5398 2413 5458 3027
rect 5395 2412 5461 2413
rect 5395 2348 5396 2412
rect 5460 2348 5461 2412
rect 5395 2347 5461 2348
rect 5582 1869 5642 5611
rect 5766 4045 5826 5886
rect 5950 4861 6010 15267
rect 6142 15264 6462 16288
rect 6142 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6462 15264
rect 6142 14176 6462 15200
rect 6142 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6462 14176
rect 6142 13088 6462 14112
rect 6142 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6462 13088
rect 6142 12000 6462 13024
rect 6686 12450 6746 17443
rect 6686 12390 6930 12450
rect 6142 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6462 12000
rect 6142 10912 6462 11936
rect 6142 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6462 10912
rect 6142 9824 6462 10848
rect 6142 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6462 9824
rect 6142 8736 6462 9760
rect 6683 8940 6749 8941
rect 6683 8876 6684 8940
rect 6748 8876 6749 8940
rect 6683 8875 6749 8876
rect 6142 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6462 8736
rect 6142 7648 6462 8672
rect 6142 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6462 7648
rect 6142 6560 6462 7584
rect 6142 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6462 6560
rect 6142 5472 6462 6496
rect 6686 5949 6746 8875
rect 6870 8805 6930 12390
rect 7422 12069 7482 19347
rect 7603 17916 7669 17917
rect 7603 17852 7604 17916
rect 7668 17852 7669 17916
rect 7603 17851 7669 17852
rect 7419 12068 7485 12069
rect 7419 12004 7420 12068
rect 7484 12004 7485 12068
rect 7419 12003 7485 12004
rect 7606 11525 7666 17851
rect 7603 11524 7669 11525
rect 7603 11460 7604 11524
rect 7668 11460 7669 11524
rect 7603 11459 7669 11460
rect 7790 9485 7850 19347
rect 7971 16692 8037 16693
rect 7971 16628 7972 16692
rect 8036 16628 8037 16692
rect 7971 16627 8037 16628
rect 7787 9484 7853 9485
rect 7787 9420 7788 9484
rect 7852 9420 7853 9484
rect 7787 9419 7853 9420
rect 7790 9213 7850 9419
rect 7974 9349 8034 16627
rect 8158 16557 8218 20843
rect 11099 20772 11165 20773
rect 8741 20160 9061 20720
rect 11099 20708 11100 20772
rect 11164 20708 11165 20772
rect 11099 20707 11165 20708
rect 8741 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9061 20160
rect 8339 20092 8405 20093
rect 8339 20028 8340 20092
rect 8404 20028 8405 20092
rect 8339 20027 8405 20028
rect 8155 16556 8221 16557
rect 8155 16492 8156 16556
rect 8220 16492 8221 16556
rect 8155 16491 8221 16492
rect 8155 15468 8221 15469
rect 8155 15404 8156 15468
rect 8220 15404 8221 15468
rect 8155 15403 8221 15404
rect 8158 9757 8218 15403
rect 8342 14245 8402 20027
rect 8523 19548 8589 19549
rect 8523 19484 8524 19548
rect 8588 19484 8589 19548
rect 8523 19483 8589 19484
rect 8526 16693 8586 19483
rect 8741 19072 9061 20096
rect 8741 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9061 19072
rect 8741 17984 9061 19008
rect 10731 18868 10797 18869
rect 10731 18804 10732 18868
rect 10796 18804 10797 18868
rect 10731 18803 10797 18804
rect 10547 18596 10613 18597
rect 10547 18532 10548 18596
rect 10612 18532 10613 18596
rect 10547 18531 10613 18532
rect 8741 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9061 17984
rect 8741 16896 9061 17920
rect 9995 17780 10061 17781
rect 9995 17716 9996 17780
rect 10060 17716 10061 17780
rect 9995 17715 10061 17716
rect 8741 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9061 16896
rect 8523 16692 8589 16693
rect 8523 16628 8524 16692
rect 8588 16628 8589 16692
rect 8523 16627 8589 16628
rect 8523 16420 8589 16421
rect 8523 16356 8524 16420
rect 8588 16356 8589 16420
rect 8523 16355 8589 16356
rect 8339 14244 8405 14245
rect 8339 14180 8340 14244
rect 8404 14180 8405 14244
rect 8339 14179 8405 14180
rect 8339 13020 8405 13021
rect 8339 12956 8340 13020
rect 8404 12956 8405 13020
rect 8339 12955 8405 12956
rect 8342 9890 8402 12955
rect 8526 12341 8586 16355
rect 8741 15808 9061 16832
rect 9811 16284 9877 16285
rect 9811 16220 9812 16284
rect 9876 16220 9877 16284
rect 9811 16219 9877 16220
rect 8741 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9061 15808
rect 8741 14720 9061 15744
rect 9443 15332 9509 15333
rect 9443 15268 9444 15332
rect 9508 15268 9509 15332
rect 9443 15267 9509 15268
rect 8741 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9061 14720
rect 8741 13632 9061 14656
rect 9259 14244 9325 14245
rect 9259 14180 9260 14244
rect 9324 14180 9325 14244
rect 9259 14179 9325 14180
rect 8741 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9061 13632
rect 8741 12544 9061 13568
rect 8741 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9061 12544
rect 8523 12340 8589 12341
rect 8523 12276 8524 12340
rect 8588 12276 8589 12340
rect 8523 12275 8589 12276
rect 8741 11456 9061 12480
rect 8741 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9061 11456
rect 8741 10368 9061 11392
rect 8741 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9061 10368
rect 8342 9830 8586 9890
rect 8155 9756 8221 9757
rect 8155 9692 8156 9756
rect 8220 9692 8221 9756
rect 8155 9691 8221 9692
rect 8339 9756 8405 9757
rect 8339 9692 8340 9756
rect 8404 9692 8405 9756
rect 8339 9691 8405 9692
rect 7971 9348 8037 9349
rect 7971 9284 7972 9348
rect 8036 9284 8037 9348
rect 7971 9283 8037 9284
rect 7787 9212 7853 9213
rect 7787 9148 7788 9212
rect 7852 9148 7853 9212
rect 7787 9147 7853 9148
rect 7974 8805 8034 9283
rect 8155 9212 8221 9213
rect 8155 9148 8156 9212
rect 8220 9148 8221 9212
rect 8155 9147 8221 9148
rect 6867 8804 6933 8805
rect 6867 8740 6868 8804
rect 6932 8740 6933 8804
rect 6867 8739 6933 8740
rect 7603 8804 7669 8805
rect 7603 8740 7604 8804
rect 7668 8802 7669 8804
rect 7971 8804 8037 8805
rect 7668 8742 7850 8802
rect 7668 8740 7669 8742
rect 7603 8739 7669 8740
rect 6867 8532 6933 8533
rect 6867 8468 6868 8532
rect 6932 8468 6933 8532
rect 6867 8467 6933 8468
rect 7603 8532 7669 8533
rect 7603 8468 7604 8532
rect 7668 8468 7669 8532
rect 7603 8467 7669 8468
rect 6683 5948 6749 5949
rect 6683 5884 6684 5948
rect 6748 5884 6749 5948
rect 6683 5883 6749 5884
rect 6870 5810 6930 8467
rect 7419 8260 7485 8261
rect 7419 8196 7420 8260
rect 7484 8196 7485 8260
rect 7419 8195 7485 8196
rect 6142 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6462 5472
rect 5947 4860 6013 4861
rect 5947 4796 5948 4860
rect 6012 4796 6013 4860
rect 5947 4795 6013 4796
rect 5947 4452 6013 4453
rect 5947 4388 5948 4452
rect 6012 4388 6013 4452
rect 5947 4387 6013 4388
rect 5763 4044 5829 4045
rect 5763 3980 5764 4044
rect 5828 3980 5829 4044
rect 5763 3979 5829 3980
rect 5950 2277 6010 4387
rect 6142 4384 6462 5408
rect 6142 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6462 4384
rect 6142 3296 6462 4320
rect 6686 5750 6930 5810
rect 6686 3909 6746 5750
rect 6867 5676 6933 5677
rect 6867 5612 6868 5676
rect 6932 5612 6933 5676
rect 6867 5611 6933 5612
rect 6683 3908 6749 3909
rect 6683 3844 6684 3908
rect 6748 3844 6749 3908
rect 6683 3843 6749 3844
rect 6870 3637 6930 5611
rect 7235 5540 7301 5541
rect 7235 5476 7236 5540
rect 7300 5476 7301 5540
rect 7235 5475 7301 5476
rect 7051 5404 7117 5405
rect 7051 5340 7052 5404
rect 7116 5340 7117 5404
rect 7051 5339 7117 5340
rect 6867 3636 6933 3637
rect 6867 3572 6868 3636
rect 6932 3572 6933 3636
rect 6867 3571 6933 3572
rect 6683 3500 6749 3501
rect 6683 3436 6684 3500
rect 6748 3436 6749 3500
rect 6683 3435 6749 3436
rect 6142 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6462 3296
rect 5947 2276 6013 2277
rect 5947 2212 5948 2276
rect 6012 2212 6013 2276
rect 5947 2211 6013 2212
rect 6142 2208 6462 3232
rect 6686 2549 6746 3435
rect 6870 2821 6930 3571
rect 6867 2820 6933 2821
rect 6867 2756 6868 2820
rect 6932 2756 6933 2820
rect 6867 2755 6933 2756
rect 7054 2685 7114 5339
rect 7238 3909 7298 5475
rect 7235 3908 7301 3909
rect 7235 3844 7236 3908
rect 7300 3844 7301 3908
rect 7235 3843 7301 3844
rect 7422 3229 7482 8195
rect 7606 6629 7666 8467
rect 7790 8258 7850 8742
rect 7971 8740 7972 8804
rect 8036 8740 8037 8804
rect 7971 8739 8037 8740
rect 7790 8198 8034 8258
rect 7787 6900 7853 6901
rect 7787 6836 7788 6900
rect 7852 6836 7853 6900
rect 7787 6835 7853 6836
rect 7603 6628 7669 6629
rect 7603 6564 7604 6628
rect 7668 6564 7669 6628
rect 7603 6563 7669 6564
rect 7419 3228 7485 3229
rect 7419 3164 7420 3228
rect 7484 3164 7485 3228
rect 7419 3163 7485 3164
rect 7422 2821 7482 3163
rect 7419 2820 7485 2821
rect 7419 2756 7420 2820
rect 7484 2756 7485 2820
rect 7419 2755 7485 2756
rect 7051 2684 7117 2685
rect 7051 2620 7052 2684
rect 7116 2620 7117 2684
rect 7051 2619 7117 2620
rect 6683 2548 6749 2549
rect 6683 2484 6684 2548
rect 6748 2484 6749 2548
rect 6683 2483 6749 2484
rect 6142 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6462 2208
rect 6142 2128 6462 2144
rect 7790 2141 7850 6835
rect 7974 2957 8034 8198
rect 8158 7037 8218 9147
rect 8155 7036 8221 7037
rect 8155 6972 8156 7036
rect 8220 6972 8221 7036
rect 8155 6971 8221 6972
rect 8155 6900 8221 6901
rect 8155 6836 8156 6900
rect 8220 6836 8221 6900
rect 8155 6835 8221 6836
rect 8158 5269 8218 6835
rect 8155 5268 8221 5269
rect 8155 5204 8156 5268
rect 8220 5204 8221 5268
rect 8155 5203 8221 5204
rect 8342 4045 8402 9691
rect 8526 6901 8586 9830
rect 8741 9280 9061 10304
rect 9262 9757 9322 14179
rect 9446 12613 9506 15267
rect 9443 12612 9509 12613
rect 9443 12548 9444 12612
rect 9508 12548 9509 12612
rect 9443 12547 9509 12548
rect 9443 12476 9509 12477
rect 9443 12412 9444 12476
rect 9508 12412 9509 12476
rect 9443 12411 9509 12412
rect 9446 11117 9506 12411
rect 9814 11525 9874 16219
rect 9811 11524 9877 11525
rect 9811 11460 9812 11524
rect 9876 11460 9877 11524
rect 9811 11459 9877 11460
rect 9443 11116 9509 11117
rect 9443 11052 9444 11116
rect 9508 11052 9509 11116
rect 9443 11051 9509 11052
rect 9443 10844 9509 10845
rect 9443 10780 9444 10844
rect 9508 10780 9509 10844
rect 9443 10779 9509 10780
rect 9259 9756 9325 9757
rect 9259 9692 9260 9756
rect 9324 9692 9325 9756
rect 9259 9691 9325 9692
rect 8741 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9061 9280
rect 8741 8192 9061 9216
rect 8741 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9061 8192
rect 8741 7104 9061 8128
rect 8741 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9061 7104
rect 8523 6900 8589 6901
rect 8523 6836 8524 6900
rect 8588 6836 8589 6900
rect 8523 6835 8589 6836
rect 8523 6356 8589 6357
rect 8523 6292 8524 6356
rect 8588 6292 8589 6356
rect 8523 6291 8589 6292
rect 8526 4317 8586 6291
rect 8741 6016 9061 7040
rect 9259 6356 9325 6357
rect 9259 6292 9260 6356
rect 9324 6354 9325 6356
rect 9446 6354 9506 10779
rect 9998 10709 10058 17715
rect 10179 16148 10245 16149
rect 10179 16084 10180 16148
rect 10244 16084 10245 16148
rect 10179 16083 10245 16084
rect 10182 10845 10242 16083
rect 10550 15197 10610 18531
rect 10734 15605 10794 18803
rect 10915 16692 10981 16693
rect 10915 16628 10916 16692
rect 10980 16628 10981 16692
rect 10915 16627 10981 16628
rect 10731 15604 10797 15605
rect 10731 15540 10732 15604
rect 10796 15540 10797 15604
rect 10731 15539 10797 15540
rect 10547 15196 10613 15197
rect 10547 15132 10548 15196
rect 10612 15132 10613 15196
rect 10547 15131 10613 15132
rect 10547 14788 10613 14789
rect 10547 14724 10548 14788
rect 10612 14724 10613 14788
rect 10547 14723 10613 14724
rect 10363 14108 10429 14109
rect 10363 14044 10364 14108
rect 10428 14044 10429 14108
rect 10363 14043 10429 14044
rect 10366 12477 10426 14043
rect 10363 12476 10429 12477
rect 10363 12412 10364 12476
rect 10428 12412 10429 12476
rect 10363 12411 10429 12412
rect 10550 12069 10610 14723
rect 10734 13565 10794 15539
rect 10918 14925 10978 16627
rect 10915 14924 10981 14925
rect 10915 14860 10916 14924
rect 10980 14860 10981 14924
rect 10915 14859 10981 14860
rect 11102 14653 11162 20707
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11099 14652 11165 14653
rect 11099 14588 11100 14652
rect 11164 14588 11165 14652
rect 11099 14587 11165 14588
rect 11340 14176 11660 15200
rect 12571 15196 12637 15197
rect 12571 15132 12572 15196
rect 12636 15132 12637 15196
rect 12571 15131 12637 15132
rect 11835 14652 11901 14653
rect 11835 14588 11836 14652
rect 11900 14588 11901 14652
rect 11835 14587 11901 14588
rect 12019 14652 12085 14653
rect 12019 14588 12020 14652
rect 12084 14588 12085 14652
rect 12019 14587 12085 14588
rect 11838 14245 11898 14587
rect 11835 14244 11901 14245
rect 11835 14180 11836 14244
rect 11900 14180 11901 14244
rect 11835 14179 11901 14180
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11099 13836 11165 13837
rect 11099 13772 11100 13836
rect 11164 13772 11165 13836
rect 11099 13771 11165 13772
rect 10731 13564 10797 13565
rect 10731 13500 10732 13564
rect 10796 13500 10797 13564
rect 10731 13499 10797 13500
rect 10915 13156 10981 13157
rect 10915 13092 10916 13156
rect 10980 13092 10981 13156
rect 10915 13091 10981 13092
rect 10547 12068 10613 12069
rect 10547 12004 10548 12068
rect 10612 12004 10613 12068
rect 10547 12003 10613 12004
rect 10731 11524 10797 11525
rect 10731 11460 10732 11524
rect 10796 11460 10797 11524
rect 10731 11459 10797 11460
rect 10179 10844 10245 10845
rect 10179 10780 10180 10844
rect 10244 10780 10245 10844
rect 10179 10779 10245 10780
rect 9995 10708 10061 10709
rect 9995 10644 9996 10708
rect 10060 10644 10061 10708
rect 9995 10643 10061 10644
rect 9627 10436 9693 10437
rect 9627 10372 9628 10436
rect 9692 10372 9693 10436
rect 9627 10371 9693 10372
rect 9630 9621 9690 10371
rect 9627 9620 9693 9621
rect 9627 9556 9628 9620
rect 9692 9556 9693 9620
rect 9627 9555 9693 9556
rect 10734 8125 10794 11459
rect 10918 9890 10978 13091
rect 11102 10165 11162 13771
rect 11340 13088 11660 14112
rect 11838 13837 11898 14179
rect 11835 13836 11901 13837
rect 11835 13772 11836 13836
rect 11900 13772 11901 13836
rect 11835 13771 11901 13772
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11835 11932 11901 11933
rect 11835 11868 11836 11932
rect 11900 11868 11901 11932
rect 11835 11867 11901 11868
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11099 10164 11165 10165
rect 11099 10100 11100 10164
rect 11164 10100 11165 10164
rect 11099 10099 11165 10100
rect 10918 9830 11162 9890
rect 11102 9213 11162 9830
rect 11340 9824 11660 10848
rect 11838 10165 11898 11867
rect 11835 10164 11901 10165
rect 11835 10100 11836 10164
rect 11900 10100 11901 10164
rect 11835 10099 11901 10100
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11099 9212 11165 9213
rect 11099 9148 11100 9212
rect 11164 9148 11165 9212
rect 11099 9147 11165 9148
rect 10915 8804 10981 8805
rect 10915 8740 10916 8804
rect 10980 8740 10981 8804
rect 10915 8739 10981 8740
rect 10918 8397 10978 8739
rect 10915 8396 10981 8397
rect 10915 8332 10916 8396
rect 10980 8332 10981 8396
rect 10915 8331 10981 8332
rect 10731 8124 10797 8125
rect 10731 8060 10732 8124
rect 10796 8060 10797 8124
rect 10731 8059 10797 8060
rect 10915 7988 10981 7989
rect 10915 7924 10916 7988
rect 10980 7924 10981 7988
rect 10915 7923 10981 7924
rect 9627 7716 9693 7717
rect 9627 7652 9628 7716
rect 9692 7652 9693 7716
rect 9627 7651 9693 7652
rect 9995 7716 10061 7717
rect 9995 7652 9996 7716
rect 10060 7652 10061 7716
rect 9995 7651 10061 7652
rect 9324 6294 9506 6354
rect 9324 6292 9325 6294
rect 9259 6291 9325 6292
rect 8741 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9061 6016
rect 8741 4928 9061 5952
rect 8741 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9061 4928
rect 8523 4316 8589 4317
rect 8523 4252 8524 4316
rect 8588 4252 8589 4316
rect 8523 4251 8589 4252
rect 8339 4044 8405 4045
rect 8339 3980 8340 4044
rect 8404 3980 8405 4044
rect 8339 3979 8405 3980
rect 8741 3840 9061 4864
rect 9262 4453 9322 6291
rect 9630 5541 9690 7651
rect 9998 6085 10058 7651
rect 9995 6084 10061 6085
rect 9995 6020 9996 6084
rect 10060 6020 10061 6084
rect 9995 6019 10061 6020
rect 9627 5540 9693 5541
rect 9627 5476 9628 5540
rect 9692 5476 9693 5540
rect 9627 5475 9693 5476
rect 10918 5405 10978 7923
rect 10915 5404 10981 5405
rect 10915 5340 10916 5404
rect 10980 5340 10981 5404
rect 10915 5339 10981 5340
rect 9443 4996 9509 4997
rect 9443 4932 9444 4996
rect 9508 4932 9509 4996
rect 9443 4931 9509 4932
rect 9259 4452 9325 4453
rect 9259 4388 9260 4452
rect 9324 4388 9325 4452
rect 9259 4387 9325 4388
rect 9446 4317 9506 4931
rect 9443 4316 9509 4317
rect 9443 4252 9444 4316
rect 9508 4252 9509 4316
rect 9443 4251 9509 4252
rect 8741 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9061 3840
rect 7971 2956 8037 2957
rect 7971 2892 7972 2956
rect 8036 2892 8037 2956
rect 7971 2891 8037 2892
rect 8741 2752 9061 3776
rect 8741 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9061 2752
rect 7787 2140 7853 2141
rect 7787 2076 7788 2140
rect 7852 2076 7853 2140
rect 8741 2128 9061 2688
rect 7787 2075 7853 2076
rect 5579 1868 5645 1869
rect 5579 1804 5580 1868
rect 5644 1804 5645 1868
rect 5579 1803 5645 1804
rect 11102 1189 11162 9147
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 12022 7037 12082 14587
rect 12574 12341 12634 15131
rect 12758 13565 12818 21251
rect 13939 20160 14259 20720
rect 13939 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14259 20160
rect 13939 19072 14259 20096
rect 13939 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14259 19072
rect 13939 17984 14259 19008
rect 13939 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14259 17984
rect 13675 16964 13741 16965
rect 13675 16900 13676 16964
rect 13740 16900 13741 16964
rect 13675 16899 13741 16900
rect 13123 14924 13189 14925
rect 13123 14860 13124 14924
rect 13188 14860 13189 14924
rect 13123 14859 13189 14860
rect 12939 13700 13005 13701
rect 12939 13636 12940 13700
rect 13004 13636 13005 13700
rect 12939 13635 13005 13636
rect 12755 13564 12821 13565
rect 12755 13500 12756 13564
rect 12820 13500 12821 13564
rect 12755 13499 12821 13500
rect 12571 12340 12637 12341
rect 12571 12276 12572 12340
rect 12636 12276 12637 12340
rect 12571 12275 12637 12276
rect 12942 10165 13002 13635
rect 13126 10845 13186 14859
rect 13491 13836 13557 13837
rect 13491 13772 13492 13836
rect 13556 13772 13557 13836
rect 13491 13771 13557 13772
rect 13307 12884 13373 12885
rect 13307 12820 13308 12884
rect 13372 12820 13373 12884
rect 13307 12819 13373 12820
rect 13123 10844 13189 10845
rect 13123 10780 13124 10844
rect 13188 10780 13189 10844
rect 13123 10779 13189 10780
rect 13126 10301 13186 10779
rect 13123 10300 13189 10301
rect 13123 10236 13124 10300
rect 13188 10236 13189 10300
rect 13123 10235 13189 10236
rect 12939 10164 13005 10165
rect 12939 10100 12940 10164
rect 13004 10100 13005 10164
rect 12939 10099 13005 10100
rect 12203 9756 12269 9757
rect 12203 9692 12204 9756
rect 12268 9692 12269 9756
rect 12203 9691 12269 9692
rect 12019 7036 12085 7037
rect 12019 6972 12020 7036
rect 12084 6972 12085 7036
rect 12019 6971 12085 6972
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 12206 4861 12266 9691
rect 12390 9150 12634 9210
rect 12390 9077 12450 9150
rect 12387 9076 12453 9077
rect 12387 9012 12388 9076
rect 12452 9012 12453 9076
rect 12387 9011 12453 9012
rect 12574 8805 12634 9150
rect 12571 8804 12637 8805
rect 12571 8740 12572 8804
rect 12636 8740 12637 8804
rect 12571 8739 12637 8740
rect 13123 8532 13189 8533
rect 13123 8468 13124 8532
rect 13188 8468 13189 8532
rect 13123 8467 13189 8468
rect 12755 6356 12821 6357
rect 12755 6292 12756 6356
rect 12820 6292 12821 6356
rect 12755 6291 12821 6292
rect 12571 6084 12637 6085
rect 12571 6020 12572 6084
rect 12636 6020 12637 6084
rect 12571 6019 12637 6020
rect 12203 4860 12269 4861
rect 12203 4796 12204 4860
rect 12268 4796 12269 4860
rect 12203 4795 12269 4796
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 2208 11660 3232
rect 12206 2549 12266 4795
rect 12574 2685 12634 6019
rect 12758 5813 12818 6291
rect 12755 5812 12821 5813
rect 12755 5748 12756 5812
rect 12820 5748 12821 5812
rect 12755 5747 12821 5748
rect 12939 5812 13005 5813
rect 12939 5748 12940 5812
rect 13004 5748 13005 5812
rect 12939 5747 13005 5748
rect 12942 3637 13002 5747
rect 13126 4589 13186 8467
rect 13123 4588 13189 4589
rect 13123 4524 13124 4588
rect 13188 4524 13189 4588
rect 13123 4523 13189 4524
rect 12939 3636 13005 3637
rect 12939 3572 12940 3636
rect 13004 3572 13005 3636
rect 12939 3571 13005 3572
rect 12571 2684 12637 2685
rect 12571 2620 12572 2684
rect 12636 2620 12637 2684
rect 12571 2619 12637 2620
rect 12203 2548 12269 2549
rect 12203 2484 12204 2548
rect 12268 2484 12269 2548
rect 12203 2483 12269 2484
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 13310 2005 13370 12819
rect 13307 2004 13373 2005
rect 13307 1940 13308 2004
rect 13372 1940 13373 2004
rect 13307 1939 13373 1940
rect 11099 1188 11165 1189
rect 11099 1124 11100 1188
rect 11164 1124 11165 1188
rect 11099 1123 11165 1124
rect 13494 1053 13554 13771
rect 13678 9893 13738 16899
rect 13939 16896 14259 17920
rect 13939 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14259 16896
rect 13939 15808 14259 16832
rect 13939 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14259 15808
rect 13939 14720 14259 15744
rect 13939 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14259 14720
rect 13939 13632 14259 14656
rect 14414 14517 14474 22475
rect 16538 20704 16858 20720
rect 16538 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16858 20704
rect 14595 20364 14661 20365
rect 14595 20300 14596 20364
rect 14660 20300 14661 20364
rect 14595 20299 14661 20300
rect 14411 14516 14477 14517
rect 14411 14452 14412 14516
rect 14476 14452 14477 14516
rect 14411 14451 14477 14452
rect 14598 13970 14658 20299
rect 16538 19616 16858 20640
rect 16538 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16858 19616
rect 15331 18732 15397 18733
rect 15331 18668 15332 18732
rect 15396 18668 15397 18732
rect 15331 18667 15397 18668
rect 14963 18188 15029 18189
rect 14963 18124 14964 18188
rect 15028 18124 15029 18188
rect 14963 18123 15029 18124
rect 13939 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14259 13632
rect 13939 12544 14259 13568
rect 13939 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14259 12544
rect 13939 11456 14259 12480
rect 13939 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14259 11456
rect 13939 10368 14259 11392
rect 13939 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14259 10368
rect 13675 9892 13741 9893
rect 13675 9828 13676 9892
rect 13740 9828 13741 9892
rect 13675 9827 13741 9828
rect 13678 6357 13738 9827
rect 13939 9280 14259 10304
rect 14414 13910 14658 13970
rect 14414 9349 14474 13910
rect 14595 13156 14661 13157
rect 14595 13092 14596 13156
rect 14660 13092 14661 13156
rect 14595 13091 14661 13092
rect 14411 9348 14477 9349
rect 14411 9284 14412 9348
rect 14476 9284 14477 9348
rect 14411 9283 14477 9284
rect 13939 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14259 9280
rect 13939 8192 14259 9216
rect 14414 8669 14474 9283
rect 14411 8668 14477 8669
rect 14411 8604 14412 8668
rect 14476 8604 14477 8668
rect 14411 8603 14477 8604
rect 13939 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14259 8192
rect 13939 7104 14259 8128
rect 14411 7852 14477 7853
rect 14411 7788 14412 7852
rect 14476 7788 14477 7852
rect 14411 7787 14477 7788
rect 13939 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14259 7104
rect 13675 6356 13741 6357
rect 13675 6292 13676 6356
rect 13740 6292 13741 6356
rect 13675 6291 13741 6292
rect 13939 6016 14259 7040
rect 13939 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14259 6016
rect 13939 4928 14259 5952
rect 13939 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14259 4928
rect 13939 3840 14259 4864
rect 14414 4725 14474 7787
rect 14411 4724 14477 4725
rect 14411 4660 14412 4724
rect 14476 4660 14477 4724
rect 14411 4659 14477 4660
rect 13939 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14259 3840
rect 13939 2752 14259 3776
rect 13939 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14259 2752
rect 13939 2128 14259 2688
rect 14598 1189 14658 13091
rect 14779 12884 14845 12885
rect 14779 12820 14780 12884
rect 14844 12820 14845 12884
rect 14779 12819 14845 12820
rect 14595 1188 14661 1189
rect 14595 1124 14596 1188
rect 14660 1124 14661 1188
rect 14595 1123 14661 1124
rect 13491 1052 13557 1053
rect 13491 988 13492 1052
rect 13556 988 13557 1052
rect 13491 987 13557 988
rect 5211 780 5277 781
rect 5211 716 5212 780
rect 5276 716 5277 780
rect 5211 715 5277 716
rect 14782 101 14842 12819
rect 14966 6901 15026 18123
rect 15334 17101 15394 18667
rect 16538 18528 16858 19552
rect 19137 20160 19457 20720
rect 19137 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19457 20160
rect 17907 19140 17973 19141
rect 17907 19076 17908 19140
rect 17972 19076 17973 19140
rect 17907 19075 17973 19076
rect 16538 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16858 18528
rect 16251 18052 16317 18053
rect 16251 17988 16252 18052
rect 16316 17988 16317 18052
rect 16251 17987 16317 17988
rect 15331 17100 15397 17101
rect 15331 17036 15332 17100
rect 15396 17036 15397 17100
rect 15331 17035 15397 17036
rect 15147 11524 15213 11525
rect 15147 11460 15148 11524
rect 15212 11460 15213 11524
rect 15147 11459 15213 11460
rect 15150 8261 15210 11459
rect 15334 9893 15394 17035
rect 15699 16692 15765 16693
rect 15699 16628 15700 16692
rect 15764 16628 15765 16692
rect 15699 16627 15765 16628
rect 15515 15060 15581 15061
rect 15515 14996 15516 15060
rect 15580 14996 15581 15060
rect 15515 14995 15581 14996
rect 15518 11525 15578 14995
rect 15515 11524 15581 11525
rect 15515 11460 15516 11524
rect 15580 11460 15581 11524
rect 15515 11459 15581 11460
rect 15331 9892 15397 9893
rect 15331 9828 15332 9892
rect 15396 9828 15397 9892
rect 15331 9827 15397 9828
rect 15702 9213 15762 16627
rect 16254 16013 16314 17987
rect 16538 17440 16858 18464
rect 16538 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16858 17440
rect 16538 16352 16858 17376
rect 16538 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16858 16352
rect 16251 16012 16317 16013
rect 16251 15948 16252 16012
rect 16316 15948 16317 16012
rect 16251 15947 16317 15948
rect 16254 9893 16314 15947
rect 16538 15264 16858 16288
rect 16538 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16858 15264
rect 16538 14176 16858 15200
rect 16538 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16858 14176
rect 16538 13088 16858 14112
rect 16538 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16858 13088
rect 16538 12000 16858 13024
rect 17723 12340 17789 12341
rect 17723 12276 17724 12340
rect 17788 12276 17789 12340
rect 17723 12275 17789 12276
rect 16538 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16858 12000
rect 16538 10912 16858 11936
rect 17171 11932 17237 11933
rect 17171 11868 17172 11932
rect 17236 11868 17237 11932
rect 17171 11867 17237 11868
rect 16538 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16858 10912
rect 16251 9892 16317 9893
rect 16251 9828 16252 9892
rect 16316 9828 16317 9892
rect 16251 9827 16317 9828
rect 15699 9212 15765 9213
rect 15699 9148 15700 9212
rect 15764 9148 15765 9212
rect 15699 9147 15765 9148
rect 15331 8668 15397 8669
rect 15331 8604 15332 8668
rect 15396 8604 15397 8668
rect 15331 8603 15397 8604
rect 15147 8260 15213 8261
rect 15147 8196 15148 8260
rect 15212 8196 15213 8260
rect 15147 8195 15213 8196
rect 14963 6900 15029 6901
rect 14963 6836 14964 6900
rect 15028 6836 15029 6900
rect 14963 6835 15029 6836
rect 15334 4861 15394 8603
rect 16067 7172 16133 7173
rect 16067 7108 16068 7172
rect 16132 7108 16133 7172
rect 16067 7107 16133 7108
rect 15883 6628 15949 6629
rect 15883 6564 15884 6628
rect 15948 6564 15949 6628
rect 15883 6563 15949 6564
rect 15331 4860 15397 4861
rect 15331 4796 15332 4860
rect 15396 4796 15397 4860
rect 15331 4795 15397 4796
rect 15886 3093 15946 6563
rect 15883 3092 15949 3093
rect 15883 3028 15884 3092
rect 15948 3028 15949 3092
rect 15883 3027 15949 3028
rect 16070 1053 16130 7107
rect 16254 2549 16314 9827
rect 16538 9824 16858 10848
rect 16538 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16858 9824
rect 16538 8736 16858 9760
rect 16987 9620 17053 9621
rect 16987 9556 16988 9620
rect 17052 9556 17053 9620
rect 16987 9555 17053 9556
rect 16538 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16858 8736
rect 16538 7648 16858 8672
rect 16538 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16858 7648
rect 16538 6560 16858 7584
rect 16538 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16858 6560
rect 16538 5472 16858 6496
rect 16538 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16858 5472
rect 16538 4384 16858 5408
rect 16538 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16858 4384
rect 16538 3296 16858 4320
rect 16538 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16858 3296
rect 16251 2548 16317 2549
rect 16251 2484 16252 2548
rect 16316 2484 16317 2548
rect 16251 2483 16317 2484
rect 16538 2208 16858 3232
rect 16990 3093 17050 9555
rect 17174 3773 17234 11867
rect 17539 9756 17605 9757
rect 17539 9692 17540 9756
rect 17604 9692 17605 9756
rect 17539 9691 17605 9692
rect 17355 8260 17421 8261
rect 17355 8196 17356 8260
rect 17420 8196 17421 8260
rect 17355 8195 17421 8196
rect 17171 3772 17237 3773
rect 17171 3708 17172 3772
rect 17236 3708 17237 3772
rect 17171 3707 17237 3708
rect 17358 3365 17418 8195
rect 17542 7989 17602 9691
rect 17539 7988 17605 7989
rect 17539 7924 17540 7988
rect 17604 7924 17605 7988
rect 17539 7923 17605 7924
rect 17726 6901 17786 12275
rect 17910 9893 17970 19075
rect 19137 19072 19457 20096
rect 21736 20704 22056 20720
rect 21736 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22056 20704
rect 21736 19616 22056 20640
rect 21736 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22056 19616
rect 19563 19276 19629 19277
rect 19563 19212 19564 19276
rect 19628 19212 19629 19276
rect 19563 19211 19629 19212
rect 19137 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19457 19072
rect 19137 17984 19457 19008
rect 19566 18461 19626 19211
rect 19931 19004 19997 19005
rect 19931 18940 19932 19004
rect 19996 18940 19997 19004
rect 19931 18939 19997 18940
rect 19934 18461 19994 18939
rect 21736 18528 22056 19552
rect 21736 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22056 18528
rect 19563 18460 19629 18461
rect 19563 18396 19564 18460
rect 19628 18396 19629 18460
rect 19563 18395 19629 18396
rect 19931 18460 19997 18461
rect 19931 18396 19932 18460
rect 19996 18396 19997 18460
rect 19931 18395 19997 18396
rect 19137 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19457 17984
rect 19137 16896 19457 17920
rect 20299 17780 20365 17781
rect 20299 17716 20300 17780
rect 20364 17716 20365 17780
rect 20299 17715 20365 17716
rect 19137 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19457 16896
rect 19137 15808 19457 16832
rect 19137 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19457 15808
rect 19137 14720 19457 15744
rect 19931 15332 19997 15333
rect 19931 15268 19932 15332
rect 19996 15268 19997 15332
rect 19931 15267 19997 15268
rect 19137 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19457 14720
rect 19137 13632 19457 14656
rect 19137 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19457 13632
rect 19137 12544 19457 13568
rect 19137 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19457 12544
rect 19137 11456 19457 12480
rect 19137 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19457 11456
rect 19137 10368 19457 11392
rect 19137 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19457 10368
rect 17907 9892 17973 9893
rect 17907 9828 17908 9892
rect 17972 9828 17973 9892
rect 17907 9827 17973 9828
rect 18275 9620 18341 9621
rect 18275 9556 18276 9620
rect 18340 9556 18341 9620
rect 18275 9555 18341 9556
rect 17907 9212 17973 9213
rect 17907 9148 17908 9212
rect 17972 9148 17973 9212
rect 17907 9147 17973 9148
rect 17723 6900 17789 6901
rect 17723 6836 17724 6900
rect 17788 6836 17789 6900
rect 17723 6835 17789 6836
rect 17910 4589 17970 9147
rect 18278 8261 18338 9555
rect 18643 9348 18709 9349
rect 18643 9284 18644 9348
rect 18708 9284 18709 9348
rect 18643 9283 18709 9284
rect 18275 8260 18341 8261
rect 18275 8196 18276 8260
rect 18340 8196 18341 8260
rect 18275 8195 18341 8196
rect 17907 4588 17973 4589
rect 17907 4524 17908 4588
rect 17972 4524 17973 4588
rect 17907 4523 17973 4524
rect 18646 4453 18706 9283
rect 19137 9280 19457 10304
rect 19747 10028 19813 10029
rect 19747 9964 19748 10028
rect 19812 9964 19813 10028
rect 19747 9963 19813 9964
rect 19137 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19457 9280
rect 19137 8192 19457 9216
rect 19563 8396 19629 8397
rect 19563 8332 19564 8396
rect 19628 8332 19629 8396
rect 19563 8331 19629 8332
rect 19137 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19457 8192
rect 19137 7104 19457 8128
rect 19137 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19457 7104
rect 19137 6016 19457 7040
rect 19566 6221 19626 8331
rect 19563 6220 19629 6221
rect 19563 6156 19564 6220
rect 19628 6156 19629 6220
rect 19563 6155 19629 6156
rect 19137 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19457 6016
rect 19137 4928 19457 5952
rect 19137 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19457 4928
rect 18643 4452 18709 4453
rect 18643 4388 18644 4452
rect 18708 4388 18709 4452
rect 18643 4387 18709 4388
rect 19137 3840 19457 4864
rect 19137 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19457 3840
rect 17355 3364 17421 3365
rect 17355 3300 17356 3364
rect 17420 3300 17421 3364
rect 17355 3299 17421 3300
rect 16987 3092 17053 3093
rect 16987 3028 16988 3092
rect 17052 3028 17053 3092
rect 16987 3027 17053 3028
rect 16538 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16858 2208
rect 16538 2128 16858 2144
rect 19137 2752 19457 3776
rect 19750 3773 19810 9963
rect 19934 3909 19994 15267
rect 20115 14788 20181 14789
rect 20115 14724 20116 14788
rect 20180 14724 20181 14788
rect 20115 14723 20181 14724
rect 20118 10029 20178 14723
rect 20115 10028 20181 10029
rect 20115 9964 20116 10028
rect 20180 9964 20181 10028
rect 20115 9963 20181 9964
rect 20302 8805 20362 17715
rect 21736 17440 22056 18464
rect 21736 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22056 17440
rect 21736 16352 22056 17376
rect 21736 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22056 16352
rect 21736 15264 22056 16288
rect 21736 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22056 15264
rect 21736 14176 22056 15200
rect 21736 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22056 14176
rect 21587 13428 21653 13429
rect 21587 13364 21588 13428
rect 21652 13364 21653 13428
rect 21587 13363 21653 13364
rect 20483 13156 20549 13157
rect 20483 13092 20484 13156
rect 20548 13092 20549 13156
rect 20483 13091 20549 13092
rect 20299 8804 20365 8805
rect 20299 8740 20300 8804
rect 20364 8740 20365 8804
rect 20299 8739 20365 8740
rect 20115 7716 20181 7717
rect 20115 7652 20116 7716
rect 20180 7652 20181 7716
rect 20115 7651 20181 7652
rect 20118 5813 20178 7651
rect 20115 5812 20181 5813
rect 20115 5748 20116 5812
rect 20180 5748 20181 5812
rect 20115 5747 20181 5748
rect 19931 3908 19997 3909
rect 19931 3844 19932 3908
rect 19996 3844 19997 3908
rect 19931 3843 19997 3844
rect 19747 3772 19813 3773
rect 19747 3708 19748 3772
rect 19812 3708 19813 3772
rect 19747 3707 19813 3708
rect 19137 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19457 2752
rect 19137 2128 19457 2688
rect 20486 2685 20546 13091
rect 21219 12748 21285 12749
rect 21219 12684 21220 12748
rect 21284 12684 21285 12748
rect 21219 12683 21285 12684
rect 21222 12341 21282 12683
rect 21590 12341 21650 13363
rect 21736 13088 22056 14112
rect 21736 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22056 13088
rect 21219 12340 21285 12341
rect 21219 12276 21220 12340
rect 21284 12276 21285 12340
rect 21219 12275 21285 12276
rect 21587 12340 21653 12341
rect 21587 12276 21588 12340
rect 21652 12276 21653 12340
rect 21587 12275 21653 12276
rect 21736 12000 22056 13024
rect 21736 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22056 12000
rect 21736 10912 22056 11936
rect 21736 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22056 10912
rect 21736 9824 22056 10848
rect 21736 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22056 9824
rect 20667 9348 20733 9349
rect 20667 9284 20668 9348
rect 20732 9284 20733 9348
rect 20667 9283 20733 9284
rect 20670 6493 20730 9283
rect 21736 8736 22056 9760
rect 21736 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22056 8736
rect 21736 7648 22056 8672
rect 21736 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22056 7648
rect 21736 6560 22056 7584
rect 21736 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22056 6560
rect 20667 6492 20733 6493
rect 20667 6428 20668 6492
rect 20732 6428 20733 6492
rect 20667 6427 20733 6428
rect 20670 6221 20730 6427
rect 20667 6220 20733 6221
rect 20667 6156 20668 6220
rect 20732 6156 20733 6220
rect 20667 6155 20733 6156
rect 21736 5472 22056 6496
rect 21736 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22056 5472
rect 21736 4384 22056 5408
rect 21736 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22056 4384
rect 21736 3296 22056 4320
rect 21736 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22056 3296
rect 20483 2684 20549 2685
rect 20483 2620 20484 2684
rect 20548 2620 20549 2684
rect 20483 2619 20549 2620
rect 21736 2208 22056 3232
rect 21736 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22056 2208
rect 21736 2128 22056 2144
rect 16067 1052 16133 1053
rect 16067 988 16068 1052
rect 16132 988 16133 1052
rect 16067 987 16133 988
rect 14779 100 14845 101
rect 14779 36 14780 100
rect 14844 36 14845 100
rect 14779 35 14845 36
use sky130_fd_sc_hd__diode_2  ANTENNA__059__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__061__A
timestamp 1649977179
transform 1 0 4232 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__062__A
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__A
timestamp 1649977179
transform 1 0 5888 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__065__A
timestamp 1649977179
transform 1 0 8280 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A
timestamp 1649977179
transform 1 0 11868 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A
timestamp 1649977179
transform 1 0 2116 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__A
timestamp 1649977179
transform 1 0 13156 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1649977179
transform 1 0 11684 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1649977179
transform 1 0 15180 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1649977179
transform -1 0 6532 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1649977179
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1649977179
transform -1 0 2852 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A
timestamp 1649977179
transform 1 0 19964 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1649977179
transform -1 0 21252 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1649977179
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1649977179
transform -1 0 21252 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A
timestamp 1649977179
transform 1 0 19412 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1649977179
transform 1 0 19780 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1649977179
transform 1 0 19596 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1649977179
transform -1 0 20332 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1649977179
transform 1 0 20608 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1649977179
transform 1 0 21068 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1649977179
transform 1 0 20424 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1649977179
transform 1 0 19688 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1649977179
transform 1 0 19504 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1649977179
transform 1 0 14352 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1649977179
transform 1 0 14168 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1649977179
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1649977179
transform 1 0 15916 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1649977179
transform 1 0 14904 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1649977179
transform 1 0 18768 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1649977179
transform 1 0 14720 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1649977179
transform 1 0 19964 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1649977179
transform 1 0 18400 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1649977179
transform -1 0 10764 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1649977179
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__A
timestamp 1649977179
transform 1 0 11776 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A
timestamp 1649977179
transform -1 0 13984 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A
timestamp 1649977179
transform -1 0 16376 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__A
timestamp 1649977179
transform 1 0 16376 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__127__A
timestamp 1649977179
transform -1 0 16008 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__A
timestamp 1649977179
transform -1 0 17572 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__130__A
timestamp 1649977179
transform -1 0 16192 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__131__A
timestamp 1649977179
transform 1 0 17572 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__133__A
timestamp 1649977179
transform 1 0 17204 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__134__A
timestamp 1649977179
transform -1 0 17388 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__A
timestamp 1649977179
transform 1 0 18032 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 15272 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 5152 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform 1 0 6992 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 14168 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 2852 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 10580 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 13892 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 13340 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 14444 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 14260 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 10764 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 4600 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 12236 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 4784 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 10764 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 7820 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 12420 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 8004 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 6256 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 5336 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 13984 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 12788 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 14168 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 13708 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 10488 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 11684 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 11868 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 10948 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 14628 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 15456 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 17388 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 16560 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 20332 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 15088 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 17572 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 18124 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 21620 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 17940 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 17756 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 19228 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 18400 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 19412 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1649977179
transform -1 0 14444 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1649977179
transform -1 0 17204 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1649977179
transform -1 0 19964 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1649977179
transform -1 0 14352 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1649977179
transform -1 0 14444 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1649977179
transform -1 0 13616 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1649977179
transform -1 0 12052 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1649977179
transform -1 0 11868 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1649977179
transform -1 0 9936 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1649977179
transform -1 0 10856 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1649977179
transform -1 0 14260 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1649977179
transform -1 0 9936 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1649977179
transform -1 0 11776 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1649977179
transform -1 0 16560 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1649977179
transform -1 0 10672 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1649977179
transform -1 0 11132 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1649977179
transform -1 0 10580 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1649977179
transform -1 0 13708 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1649977179
transform -1 0 11132 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1649977179
transform -1 0 10672 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1649977179
transform -1 0 13524 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1649977179
transform -1 0 10304 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1649977179
transform -1 0 13156 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1649977179
transform -1 0 12972 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1649977179
transform -1 0 10396 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1649977179
transform -1 0 4232 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1649977179
transform -1 0 13984 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1649977179
transform -1 0 8004 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1649977179
transform -1 0 2300 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1649977179
transform -1 0 13984 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1649977179
transform -1 0 9016 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1649977179
transform -1 0 13432 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1649977179
transform -1 0 3956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1649977179
transform -1 0 9476 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1649977179
transform -1 0 14168 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1649977179
transform -1 0 9108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1649977179
transform -1 0 8832 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1649977179
transform -1 0 12420 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1649977179
transform -1 0 13156 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1649977179
transform -1 0 15732 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1649977179
transform -1 0 14352 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1649977179
transform -1 0 12236 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 1649977179
transform -1 0 2852 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input89_A
timestamp 1649977179
transform -1 0 15548 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input90_A
timestamp 1649977179
transform -1 0 2576 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input91_A
timestamp 1649977179
transform -1 0 19044 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input92_A
timestamp 1649977179
transform 1 0 19228 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input93_A
timestamp 1649977179
transform -1 0 18860 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input94_A
timestamp 1649977179
transform -1 0 1932 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input95_A
timestamp 1649977179
transform -1 0 13616 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input96_A
timestamp 1649977179
transform -1 0 3956 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input97_A
timestamp 1649977179
transform -1 0 6808 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input98_A
timestamp 1649977179
transform -1 0 8740 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input99_A
timestamp 1649977179
transform -1 0 10120 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input100_A
timestamp 1649977179
transform -1 0 10304 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input101_A
timestamp 1649977179
transform -1 0 10488 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input102_A
timestamp 1649977179
transform -1 0 18032 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input103_A
timestamp 1649977179
transform -1 0 19412 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input104_A
timestamp 1649977179
transform -1 0 20332 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input105_A
timestamp 1649977179
transform -1 0 16284 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input106_A
timestamp 1649977179
transform -1 0 18216 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input107_A
timestamp 1649977179
transform -1 0 14904 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input108_A
timestamp 1649977179
transform -1 0 13984 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input109_A
timestamp 1649977179
transform -1 0 17020 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input110_A
timestamp 1649977179
transform 1 0 18768 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input111_A
timestamp 1649977179
transform 1 0 21436 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input112_A
timestamp 1649977179
transform -1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input113_A
timestamp 1649977179
transform -1 0 4232 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input114_A
timestamp 1649977179
transform 1 0 4324 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input115_A
timestamp 1649977179
transform -1 0 8464 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input116_A
timestamp 1649977179
transform 1 0 1748 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input117_A
timestamp 1649977179
transform -1 0 6256 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input118_A
timestamp 1649977179
transform -1 0 3588 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input119_A
timestamp 1649977179
transform -1 0 4232 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input120_A
timestamp 1649977179
transform -1 0 6716 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 21252 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 16652 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 13616 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 13616 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 12420 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_4__A0
timestamp 1649977179
transform 1 0 12880 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 12052 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 12144 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 7360 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 11408 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 12328 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 10488 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_4__A0
timestamp 1649977179
transform 1 0 11776 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 11960 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 10948 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 10304 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 10120 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 9936 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 10764 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_6__A0
timestamp 1649977179
transform 1 0 11040 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_6__A1
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_7__A1
timestamp 1649977179
transform 1 0 7820 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 12696 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 13248 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 13984 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 13800 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 13432 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 10396 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 12512 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8188 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8004 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 10856 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 10672 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 10396 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 6992 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 10120 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 12512 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 13524 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 13800 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 10856 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 12236 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 13708 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 11040 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 16100 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 14904 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 15824 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 10672 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 10304 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 10764 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 9936 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 10856 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__A1
timestamp 1649977179
transform -1 0 5888 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 3220 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 7452 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 10120 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 2852 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 8188 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 10948 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A0
timestamp 1649977179
transform -1 0 1564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 11132 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 7728 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 10028 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 6808 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 7084 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 7268 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 8924 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 8280 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 6440 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 6256 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6716 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 9752 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 6716 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 6164 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 10028 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 11316 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 11500 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 8740 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 10396 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 4784 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6072 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 1564 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 10212 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 15456 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 14536 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_3__A0
timestamp 1649977179
transform 1 0 14444 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_4__A1
timestamp 1649977179
transform 1 0 16008 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 16836 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 15088 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 13432 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 13524 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 16652 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__A0
timestamp 1649977179
transform 1 0 18584 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_4__A0
timestamp 1649977179
transform 1 0 14536 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 14168 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_5__A1
timestamp 1649977179
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_6__A0
timestamp 1649977179
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_6__A1
timestamp 1649977179
transform 1 0 18400 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_7__A1
timestamp 1649977179
transform 1 0 14260 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 17388 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 14352 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 16100 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 16468 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 16652 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 14168 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 16100 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 14444 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 16284 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 16284 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 18032 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 17204 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 17020 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 18124 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 17664 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 19412 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 18860 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 19504 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 14812 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 14812 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 14352 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 17020 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 6348 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 4508 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_3__A0
timestamp 1649977179
transform 1 0 6440 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_4__A1
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 2576 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 9016 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 8096 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 7912 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A0
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 6716 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_4__A0
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_4__A1
timestamp 1649977179
transform 1 0 7636 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 8464 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__A0
timestamp 1649977179
transform -1 0 8464 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_4__A0
timestamp 1649977179
transform 1 0 8832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_4__A1
timestamp 1649977179
transform -1 0 10028 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_5__A0
timestamp 1649977179
transform 1 0 7544 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_5__A1
timestamp 1649977179
transform 1 0 8464 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_6__A0
timestamp 1649977179
transform 1 0 7820 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_6__A1
timestamp 1649977179
transform 1 0 8096 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 11132 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 12052 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 11868 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 9292 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 13616 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 12052 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 13248 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 11684 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 10488 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 11500 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 18032 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 17480 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 16836 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 14352 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 14536 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 16192 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 13616 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 11868 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 11684 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 12052 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output217_A
timestamp 1649977179
transform 1 0 16376 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_2_E_FTB01_A
timestamp 1649977179
transform 1 0 19320 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_2_N_FTB01_A
timestamp 1649977179
transform -1 0 20424 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_2_S_FTB01_A
timestamp 1649977179
transform -1 0 17848 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_2_W_FTB01_A
timestamp 1649977179
transform -1 0 19964 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3220 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1649977179
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_39
timestamp 1649977179
transform 1 0 4692 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_126
timestamp 1649977179
transform 1 0 12696 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_156
timestamp 1649977179
transform 1 0 15456 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1649977179
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_74
timestamp 1649977179
transform 1 0 7912 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_174
timestamp 1649977179
transform 1 0 17112 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_80
timestamp 1649977179
transform 1 0 8464 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_212
timestamp 1649977179
transform 1 0 20608 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_32
timestamp 1649977179
transform 1 0 4048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_79
timestamp 1649977179
transform 1 0 8372 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_121
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_66
timestamp 1649977179
transform 1 0 7176 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_134
timestamp 1649977179
transform 1 0 13432 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1649977179
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_125
timestamp 1649977179
transform 1 0 12604 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_169
timestamp 1649977179
transform 1 0 16652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_218
timestamp 1649977179
transform 1 0 21160 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_7
timestamp 1649977179
transform 1 0 1748 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_45
timestamp 1649977179
transform 1 0 5244 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1649977179
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_66
timestamp 1649977179
transform 1 0 7176 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_124
timestamp 1649977179
transform 1 0 12512 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_164
timestamp 1649977179
transform 1 0 16192 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_172
timestamp 1649977179
transform 1 0 16928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_94
timestamp 1649977179
transform 1 0 9752 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_122
timestamp 1649977179
transform 1 0 12328 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_7
timestamp 1649977179
transform 1 0 1748 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_69
timestamp 1649977179
transform 1 0 7452 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_106
timestamp 1649977179
transform 1 0 10856 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_125
timestamp 1649977179
transform 1 0 12604 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_71
timestamp 1649977179
transform 1 0 7636 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1649977179
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_200
timestamp 1649977179
transform 1 0 19504 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_210
timestamp 1649977179
transform 1 0 20424 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_142
timestamp 1649977179
transform 1 0 14168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_44
timestamp 1649977179
transform 1 0 5152 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_74
timestamp 1649977179
transform 1 0 7912 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_133
timestamp 1649977179
transform 1 0 13340 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_157
timestamp 1649977179
transform 1 0 15548 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_222
timestamp 1649977179
transform 1 0 21528 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_7
timestamp 1649977179
transform 1 0 1748 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_34
timestamp 1649977179
transform 1 0 4232 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_165
timestamp 1649977179
transform 1 0 16284 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_35
timestamp 1649977179
transform 1 0 4324 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_118
timestamp 1649977179
transform 1 0 11960 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_137
timestamp 1649977179
transform 1 0 13708 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_157
timestamp 1649977179
transform 1 0 15548 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_39
timestamp 1649977179
transform 1 0 4692 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_43
timestamp 1649977179
transform 1 0 5060 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1649977179
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_59
timestamp 1649977179
transform 1 0 6532 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_81
timestamp 1649977179
transform 1 0 8556 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_105
timestamp 1649977179
transform 1 0 10764 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1649977179
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_179
timestamp 1649977179
transform 1 0 17572 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_222
timestamp 1649977179
transform 1 0 21528 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_22
timestamp 1649977179
transform 1 0 3128 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_46
timestamp 1649977179
transform 1 0 5336 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_149
timestamp 1649977179
transform 1 0 14812 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_165
timestamp 1649977179
transform 1 0 16284 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_77
timestamp 1649977179
transform 1 0 8188 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_107
timestamp 1649977179
transform 1 0 10948 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_137
timestamp 1649977179
transform 1 0 13708 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_172
timestamp 1649977179
transform 1 0 16928 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_177
timestamp 1649977179
transform 1 0 17388 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_192
timestamp 1649977179
transform 1 0 18768 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_201
timestamp 1649977179
transform 1 0 19596 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_7
timestamp 1649977179
transform 1 0 1748 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_17
timestamp 1649977179
transform 1 0 2668 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_82
timestamp 1649977179
transform 1 0 8648 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_142
timestamp 1649977179
transform 1 0 14168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_203
timestamp 1649977179
transform 1 0 19780 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_34
timestamp 1649977179
transform 1 0 4232 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_121
timestamp 1649977179
transform 1 0 12236 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_176
timestamp 1649977179
transform 1 0 17296 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1649977179
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_211
timestamp 1649977179
transform 1 0 20516 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_34
timestamp 1649977179
transform 1 0 4232 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_117
timestamp 1649977179
transform 1 0 11868 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_153 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15180 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1649977179
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_18
timestamp 1649977179
transform 1 0 2760 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_32
timestamp 1649977179
transform 1 0 4048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_65
timestamp 1649977179
transform 1 0 7084 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_157 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15548 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_186
timestamp 1649977179
transform 1 0 18216 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1649977179
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_218
timestamp 1649977179
transform 1 0 21160 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_14
timestamp 1649977179
transform 1 0 2392 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_40
timestamp 1649977179
transform 1 0 4784 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_88
timestamp 1649977179
transform 1 0 9200 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1649977179
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_164
timestamp 1649977179
transform 1 0 16192 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_172
timestamp 1649977179
transform 1 0 16928 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_214
timestamp 1649977179
transform 1 0 20792 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_7
timestamp 1649977179
transform 1 0 1748 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_60
timestamp 1649977179
transform 1 0 6624 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_121
timestamp 1649977179
transform 1 0 12236 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_134 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13432 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_148
timestamp 1649977179
transform 1 0 14720 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_199
timestamp 1649977179
transform 1 0 19412 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_7
timestamp 1649977179
transform 1 0 1748 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_92
timestamp 1649977179
transform 1 0 9568 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_157
timestamp 1649977179
transform 1 0 15548 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_163
timestamp 1649977179
transform 1 0 16100 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_179 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_191
timestamp 1649977179
transform 1 0 18676 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_11
timestamp 1649977179
transform 1 0 2116 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_88
timestamp 1649977179
transform 1 0 9200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1649977179
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_186 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18216 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1649977179
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1649977179
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_133
timestamp 1649977179
transform 1 0 13340 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_180
timestamp 1649977179
transform 1 0 17664 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_192
timestamp 1649977179
transform 1 0 18768 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_200
timestamp 1649977179
transform 1 0 19504 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_60
timestamp 1649977179
transform 1 0 6624 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_94
timestamp 1649977179
transform 1 0 9752 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_118
timestamp 1649977179
transform 1 0 11960 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_134
timestamp 1649977179
transform 1 0 13432 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_151
timestamp 1649977179
transform 1 0 14996 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_173
timestamp 1649977179
transform 1 0 17020 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_185
timestamp 1649977179
transform 1 0 18124 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_193
timestamp 1649977179
transform 1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_11
timestamp 1649977179
transform 1 0 2116 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_46
timestamp 1649977179
transform 1 0 5336 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_66
timestamp 1649977179
transform 1 0 7176 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_71
timestamp 1649977179
transform 1 0 7636 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_90
timestamp 1649977179
transform 1 0 9384 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_104
timestamp 1649977179
transform 1 0 10672 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1649977179
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_159
timestamp 1649977179
transform 1 0 15732 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1649977179
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_181
timestamp 1649977179
transform 1 0 17756 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_189
timestamp 1649977179
transform 1 0 18492 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_7
timestamp 1649977179
transform 1 0 1748 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_168
timestamp 1649977179
transform 1 0 16560 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_174
timestamp 1649977179
transform 1 0 17112 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_177
timestamp 1649977179
transform 1 0 17388 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_218
timestamp 1649977179
transform 1 0 21160 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_141
timestamp 1649977179
transform 1 0 14076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1649977179
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_208
timestamp 1649977179
transform 1 0 20240 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_110
timestamp 1649977179
transform 1 0 11224 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_186
timestamp 1649977179
transform 1 0 18216 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_191
timestamp 1649977179
transform 1 0 18676 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_212
timestamp 1649977179
transform 1 0 20608 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_11
timestamp 1649977179
transform 1 0 2116 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_97
timestamp 1649977179
transform 1 0 10028 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_139
timestamp 1649977179
transform 1 0 13892 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 21896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 21896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 21896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 21896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 21896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 21896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 21896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 21896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 21896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 21896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 21896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 21896 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 21896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 21896 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 21896 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 21896 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 21896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 21896 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 21896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 21896 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 21896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 21896 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 21896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 21896 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 21896 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 21896 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 21896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 21896 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 21896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 21896 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 21896 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 21896 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 3680 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 8832 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 13984 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  Test_en_N_FTB01 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18768 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _056_
timestamp 1649977179
transform 1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _057_
timestamp 1649977179
transform 1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _058_
timestamp 1649977179
transform 1 0 3128 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _059_
timestamp 1649977179
transform 1 0 3220 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _060_
timestamp 1649977179
transform 1 0 2116 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _061_
timestamp 1649977179
transform 1 0 2208 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _062_
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _063_
timestamp 1649977179
transform 1 0 2116 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _064_
timestamp 1649977179
transform 1 0 2392 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _065_
timestamp 1649977179
transform 1 0 4048 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _066_
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _067_
timestamp 1649977179
transform 1 0 1840 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _068_
timestamp 1649977179
transform 1 0 2116 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _069_
timestamp 1649977179
transform 1 0 2116 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _070_
timestamp 1649977179
transform 1 0 2484 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp 1649977179
transform 1 0 2116 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp 1649977179
transform 1 0 1840 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp 1649977179
transform 1 0 4048 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp 1649977179
transform -1 0 19504 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1649977179
transform -1 0 17940 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1649977179
transform -1 0 18584 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp 1649977179
transform -1 0 20424 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1649977179
transform -1 0 19688 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp 1649977179
transform -1 0 20884 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp 1649977179
transform -1 0 21068 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp 1649977179
transform -1 0 20792 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1649977179
transform -1 0 21068 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1649977179
transform -1 0 20792 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp 1649977179
transform -1 0 20240 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1649977179
transform -1 0 20516 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp 1649977179
transform -1 0 20884 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp 1649977179
transform -1 0 20608 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp 1649977179
transform -1 0 21068 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp 1649977179
transform 1 0 20976 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1649977179
transform -1 0 20240 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1649977179
transform -1 0 20884 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp 1649977179
transform -1 0 20608 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 1649977179
transform -1 0 20240 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp 1649977179
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 1649977179
transform -1 0 12144 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 1649977179
transform -1 0 12604 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp 1649977179
transform 1 0 15916 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp 1649977179
transform -1 0 15180 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp 1649977179
transform 1 0 16192 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp 1649977179
transform -1 0 11776 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _104_
timestamp 1649977179
transform -1 0 10948 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp 1649977179
transform 1 0 17204 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1649977179
transform 1 0 19596 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _107_
timestamp 1649977179
transform 1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1649977179
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1649977179
transform 1 0 19872 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _110_
timestamp 1649977179
transform -1 0 18124 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 1649977179
transform -1 0 11408 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp 1649977179
transform -1 0 17848 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 1649977179
transform 1 0 20148 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1649977179
transform 1 0 20424 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1649977179
transform 1 0 20332 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp 1649977179
transform 1 0 10120 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1649977179
transform -1 0 11316 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1649977179
transform -1 0 11040 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 1649977179
transform -1 0 11316 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _120_
timestamp 1649977179
transform -1 0 11040 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp 1649977179
transform 1 0 13800 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _122_
timestamp 1649977179
transform -1 0 11408 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1649977179
transform 1 0 15456 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp 1649977179
transform 1 0 15180 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1649977179
transform 1 0 15640 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _126_
timestamp 1649977179
transform 1 0 16284 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _127_
timestamp 1649977179
transform -1 0 15548 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _128_
timestamp 1649977179
transform 1 0 16560 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _129_
timestamp 1649977179
transform 1 0 16836 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1649977179
transform -1 0 15824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _131_
timestamp 1649977179
transform 1 0 17112 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _132_
timestamp 1649977179
transform -1 0 16468 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1649977179
transform -1 0 17664 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _134_
timestamp 1649977179
transform -1 0 17204 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _135_
timestamp 1649977179
transform -1 0 18032 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_1_E_FTB01
timestamp 1649977179
transform -1 0 19136 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_1_W_FTB01
timestamp 1649977179
transform 1 0 17664 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_2_E_FTB01
timestamp 1649977179
transform -1 0 19872 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_2_N_FTB01
timestamp 1649977179
transform -1 0 20700 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_2_S_FTB01
timestamp 1649977179
transform -1 0 20148 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_2_W_FTB01
timestamp 1649977179
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_3_E_FTB01
timestamp 1649977179
transform 1 0 19872 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_3_N_FTB01
timestamp 1649977179
transform -1 0 19136 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_3_S_FTB01
timestamp 1649977179
transform -1 0 20424 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_3_W_FTB01
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform -1 0 17296 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1649977179
transform -1 0 5152 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform -1 0 7452 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 3220 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform -1 0 6808 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform -1 0 5244 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform -1 0 1932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1649977179
transform -1 0 4692 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1649977179
transform -1 0 1840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1649977179
transform -1 0 2116 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1649977179
transform 1 0 6256 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input12 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3220 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform -1 0 4048 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input14 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input15
timestamp 1649977179
transform 1 0 3864 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform -1 0 2944 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1649977179
transform 1 0 1748 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp 1649977179
transform -1 0 2300 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1649977179
transform -1 0 1656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1649977179
transform 1 0 2300 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1649977179
transform -1 0 2300 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1649977179
transform 1 0 2668 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1649977179
transform 1 0 2300 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input28
timestamp 1649977179
transform -1 0 2300 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1649977179
transform 1 0 3128 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1649977179
transform 1 0 18032 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1649977179
transform -1 0 21620 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp 1649977179
transform 1 0 20700 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1649977179
transform -1 0 19136 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1649977179
transform -1 0 18952 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1649977179
transform -1 0 20700 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input37
timestamp 1649977179
transform 1 0 20700 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1649977179
transform -1 0 20056 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1649977179
transform -1 0 20700 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1649977179
transform -1 0 21252 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input41
timestamp 1649977179
transform 1 0 20700 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input42
timestamp 1649977179
transform 1 0 20700 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1649977179
transform -1 0 21620 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input44
timestamp 1649977179
transform 1 0 20700 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1649977179
transform -1 0 20700 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1649977179
transform -1 0 19136 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1649977179
transform -1 0 21620 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input48
timestamp 1649977179
transform 1 0 20700 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1649977179
transform -1 0 21620 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1649977179
transform -1 0 20424 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input51
timestamp 1649977179
transform -1 0 7268 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input52
timestamp 1649977179
transform -1 0 6256 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1649977179
transform -1 0 9200 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input54
timestamp 1649977179
transform -1 0 9752 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1649977179
transform -1 0 7912 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input56
timestamp 1649977179
transform 1 0 12328 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1649977179
transform 1 0 11316 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input58
timestamp 1649977179
transform -1 0 12604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input59
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input60
timestamp 1649977179
transform 1 0 11868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1649977179
transform -1 0 11868 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1649977179
transform -1 0 5980 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1649977179
transform 1 0 6072 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1649977179
transform -1 0 5244 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input65
timestamp 1649977179
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input66
timestamp 1649977179
transform 1 0 5244 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1649977179
transform 1 0 3864 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1649977179
transform -1 0 3680 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1649977179
transform -1 0 6992 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input70
timestamp 1649977179
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input71
timestamp 1649977179
transform -1 0 4692 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input72
timestamp 1649977179
transform -1 0 7636 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1649977179
transform -1 0 6532 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input74
timestamp 1649977179
transform -1 0 6900 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input75
timestamp 1649977179
transform -1 0 6808 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input76
timestamp 1649977179
transform -1 0 8832 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input77
timestamp 1649977179
transform 1 0 9108 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input78
timestamp 1649977179
transform 1 0 9476 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input79
timestamp 1649977179
transform 1 0 7544 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input80
timestamp 1649977179
transform 1 0 11684 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input81
timestamp 1649977179
transform 1 0 10488 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1649977179
transform -1 0 4876 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input83
timestamp 1649977179
transform 1 0 2208 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1649977179
transform -1 0 4232 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input85
timestamp 1649977179
transform 1 0 2576 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input86
timestamp 1649977179
transform -1 0 7268 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input87
timestamp 1649977179
transform 1 0 2944 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 1649977179
transform -1 0 6256 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input89
timestamp 1649977179
transform 1 0 3312 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input90
timestamp 1649977179
transform 1 0 6532 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1649977179
transform 1 0 19044 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input92
timestamp 1649977179
transform -1 0 19596 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1649977179
transform -1 0 19872 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1649977179
transform -1 0 4324 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input95
timestamp 1649977179
transform -1 0 2300 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 1649977179
transform 1 0 3404 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input97
timestamp 1649977179
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input98
timestamp 1649977179
transform -1 0 8832 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input99
timestamp 1649977179
transform 1 0 6532 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input100
timestamp 1649977179
transform 1 0 6256 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input101
timestamp 1649977179
transform 1 0 5980 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input102
timestamp 1649977179
transform 1 0 19412 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input103
timestamp 1649977179
transform 1 0 18492 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input104
timestamp 1649977179
transform 1 0 19044 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input105
timestamp 1649977179
transform -1 0 16560 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input106
timestamp 1649977179
transform 1 0 20700 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input107
timestamp 1649977179
transform -1 0 14352 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input108
timestamp 1649977179
transform -1 0 13984 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input109
timestamp 1649977179
transform 1 0 17204 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input110
timestamp 1649977179
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input111
timestamp 1649977179
transform -1 0 17296 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input112
timestamp 1649977179
transform -1 0 17020 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input113
timestamp 1649977179
transform -1 0 4048 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input114
timestamp 1649977179
transform -1 0 5612 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input115
timestamp 1649977179
transform -1 0 8004 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input116
timestamp 1649977179
transform -1 0 3680 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input117
timestamp 1649977179
transform 1 0 7452 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input118
timestamp 1649977179
transform -1 0 3404 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input119
timestamp 1649977179
transform -1 0 3128 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input120
timestamp 1649977179
transform -1 0 6072 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 18032 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 14996 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 12512 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 14260 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12052 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10120 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 10672 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 11316 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 8280 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 9016 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 7912 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 6992 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  mem_bottom_track_9.delay_buf dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9752 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9936 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11500 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 12972 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 12512 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  mem_bottom_track_17.delay_buf
timestamp 1649977179
transform -1 0 9200 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 8372 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 9292 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 10488 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  mem_bottom_track_25.delay_buf
timestamp 1649977179
transform -1 0 9936 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9936 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11040 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 13892 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  mem_bottom_track_33.delay_buf_2
timestamp 1649977179
transform 1 0 13340 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 14444 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 16652 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 4784 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 1932 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 2760 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 4232 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 2852 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 3220 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4784 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 3680 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 1932 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform 1 0 1748 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  mem_left_track_9.delay_buf
timestamp 1649977179
transform -1 0 3128 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 3220 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 7820 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 4232 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 6256 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  mem_left_track_17.delay_buf
timestamp 1649977179
transform -1 0 5888 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 8648 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 5612 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 5612 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  mem_left_track_25.delay_buf
timestamp 1649977179
transform -1 0 7544 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8004 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9016 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 2760 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 3220 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  mem_left_track_33.delay_buf_2
timestamp 1649977179
transform 1 0 1840 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 1656 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 3312 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 3312 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 17112 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 16928 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 18124 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19596 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18768 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 17296 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 18308 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20148 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 16836 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 17664 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  mem_right_track_8.delay_buf
timestamp 1649977179
transform 1 0 20056 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20332 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 14260 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 15456 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  mem_right_track_16.delay_buf
timestamp 1649977179
transform 1 0 15732 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18124 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14444 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 14720 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 15732 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  mem_right_track_24.delay_buf
timestamp 1649977179
transform -1 0 17572 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 17020 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 18492 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 19780 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 19780 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  mem_right_track_32.delay_buf_2
timestamp 1649977179
transform 1 0 20424 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21620 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 15640 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 18124 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4232 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 3128 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 2208 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 3128 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 4324 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 5980 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 5060 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 3956 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 4784 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 4968 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 6808 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  mem_top_track_8.delay_buf
timestamp 1649977179
transform 1 0 10396 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 11132 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 6624 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 8096 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 10488 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  mem_top_track_16.delay_buf
timestamp 1649977179
transform 1 0 10488 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 10028 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 13800 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  mem_top_track_24.delay_buf
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14168 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 16560 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 13432 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 15548 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  mem_top_track_32.delay_buf_2
timestamp 1649977179
transform -1 0 14720 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13892 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 10488 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 11960 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15824 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1649977179
transform 1 0 16652 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1649977179
transform 1 0 12696 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_3_
timestamp 1649977179
transform -1 0 13156 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_4_
timestamp 1649977179
transform 1 0 13156 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 14720 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1649977179
transform -1 0 13432 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_2_
timestamp 1649977179
transform -1 0 13892 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_1.mux_l2_in_3__293 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_3_
timestamp 1649977179
transform -1 0 14904 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1649977179
transform -1 0 14720 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_1_
timestamp 1649977179
transform 1 0 14260 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l4_in_0_
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 12880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1649977179
transform 1 0 11408 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1649977179
transform -1 0 11408 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_2_
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_3_
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_4_
timestamp 1649977179
transform -1 0 12236 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 10580 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1649977179
transform -1 0 8832 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_2_
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_3.mux_l2_in_3__296
timestamp 1649977179
transform -1 0 11408 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_3_
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1649977179
transform -1 0 9752 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_1_
timestamp 1649977179
transform 1 0 10396 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l4_in_0_
timestamp 1649977179
transform -1 0 10580 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 10396 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8096 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_2_
timestamp 1649977179
transform -1 0 8096 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_3_
timestamp 1649977179
transform 1 0 8096 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_4_
timestamp 1649977179
transform 1 0 6440 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_5_
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_6_
timestamp 1649977179
transform 1 0 7820 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_7_
timestamp 1649977179
transform 1 0 7728 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_5.mux_l2_in_7__298
timestamp 1649977179
transform 1 0 8280 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1649977179
transform -1 0 8096 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_1_
timestamp 1649977179
transform -1 0 8740 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_2_
timestamp 1649977179
transform -1 0 6440 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_3_
timestamp 1649977179
transform -1 0 8004 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_0_
timestamp 1649977179
transform -1 0 8832 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_1_
timestamp 1649977179
transform -1 0 8372 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l5_in_0_
timestamp 1649977179
transform 1 0 8924 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 7544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1649977179
transform -1 0 13708 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_1_
timestamp 1649977179
transform 1 0 12972 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_2_
timestamp 1649977179
transform -1 0 13248 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 12972 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1649977179
transform 1 0 13708 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_2_
timestamp 1649977179
transform -1 0 11408 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_9.mux_l2_in_3__299
timestamp 1649977179
transform 1 0 13248 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_3_
timestamp 1649977179
transform -1 0 13340 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1649977179
transform 1 0 11776 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_1_
timestamp 1649977179
transform 1 0 12512 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l4_in_0_
timestamp 1649977179
transform -1 0 11500 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 12420 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9200 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1649977179
transform 1 0 9844 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_2_
timestamp 1649977179
transform 1 0 8004 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7544 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1649977179
transform -1 0 7544 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_2_
timestamp 1649977179
transform -1 0 8832 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_17.mux_l2_in_3__294
timestamp 1649977179
transform 1 0 10488 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_3_
timestamp 1649977179
transform -1 0 10120 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1649977179
transform -1 0 8004 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_1_
timestamp 1649977179
transform 1 0 10120 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l4_in_0_
timestamp 1649977179
transform 1 0 9108 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 6624 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1649977179
transform -1 0 13524 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1649977179
transform -1 0 13800 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_2_
timestamp 1649977179
transform -1 0 12052 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1649977179
transform 1 0 13156 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1649977179
transform -1 0 12420 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_2_
timestamp 1649977179
transform 1 0 12328 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_25.mux_l2_in_3__295
timestamp 1649977179
transform 1 0 12328 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_3_
timestamp 1649977179
transform -1 0 12328 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1649977179
transform 1 0 12880 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_1_
timestamp 1649977179
transform -1 0 12880 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l4_in_0_
timestamp 1649977179
transform -1 0 13248 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 17204 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1649977179
transform -1 0 15916 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1649977179
transform -1 0 16100 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_2_
timestamp 1649977179
transform -1 0 13432 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_3_
timestamp 1649977179
transform 1 0 15640 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_33.mux_l1_in_3__297
timestamp 1649977179
transform -1 0 14812 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_1_
timestamp 1649977179
transform 1 0 15548 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l3_in_0_
timestamp 1649977179
transform -1 0 15824 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 17756 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1649977179
transform 1 0 3680 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1649977179
transform 1 0 5428 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1649977179
transform 1 0 4600 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_3_
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_4_
timestamp 1649977179
transform -1 0 10580 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 2852 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1649977179
transform 1 0 2944 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1649977179
transform 1 0 10580 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1649977179
transform 1 0 9752 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_1.mux_l2_in_3__300
timestamp 1649977179
transform -1 0 4048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1649977179
transform -1 0 2944 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1649977179
transform -1 0 7176 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1649977179
transform 1 0 10580 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1649977179
transform 1 0 6164 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_2_
timestamp 1649977179
transform 1 0 5428 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_3_
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_4_
timestamp 1649977179
transform 1 0 2852 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5336 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1649977179
transform 1 0 5244 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_2_
timestamp 1649977179
transform 1 0 2024 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_3_
timestamp 1649977179
transform 1 0 5428 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_3.mux_l2_in_3__303
timestamp 1649977179
transform -1 0 2024 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4140 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_1_
timestamp 1649977179
transform -1 0 2760 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l4_in_0_
timestamp 1649977179
transform -1 0 3680 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 4600 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1649977179
transform -1 0 7636 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6900 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1649977179
transform 1 0 5244 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1649977179
transform 1 0 6072 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1649977179
transform 1 0 5244 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_4_
timestamp 1649977179
transform 1 0 2392 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_5_
timestamp 1649977179
transform 1 0 1472 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_6_
timestamp 1649977179
transform 1 0 2300 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_5.mux_l2_in_7__277
timestamp 1649977179
transform 1 0 4600 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_7_
timestamp 1649977179
transform 1 0 1840 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4324 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1649977179
transform 1 0 5152 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_2_
timestamp 1649977179
transform -1 0 2208 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_3_
timestamp 1649977179
transform -1 0 2392 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_1_
timestamp 1649977179
transform -1 0 2668 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l5_in_0_
timestamp 1649977179
transform -1 0 3128 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3404 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7268 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1649977179
transform 1 0 8096 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_2_
timestamp 1649977179
transform 1 0 7452 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6440 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1649977179
transform 1 0 6624 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1649977179
transform -1 0 6256 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_9.mux_l2_in_3__278
timestamp 1649977179
transform 1 0 4784 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1649977179
transform -1 0 5244 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1649977179
transform -1 0 6256 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1649977179
transform -1 0 6532 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1649977179
transform 1 0 6256 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 1656 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7728 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1649977179
transform 1 0 7820 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7176 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1649977179
transform 1 0 6900 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_2_
timestamp 1649977179
transform 1 0 5336 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_17.mux_l2_in_3__301
timestamp 1649977179
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_3_
timestamp 1649977179
transform -1 0 5336 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_1_
timestamp 1649977179
transform -1 0 5980 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l4_in_0_
timestamp 1649977179
transform 1 0 5244 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2116 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9568 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1649977179
transform 1 0 10488 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1649977179
transform -1 0 9568 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9476 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_2_
timestamp 1649977179
transform 1 0 3956 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_3_
timestamp 1649977179
transform 1 0 3404 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_25.mux_l2_in_3__302
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4232 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_1_
timestamp 1649977179
transform 1 0 3220 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l4_in_0_
timestamp 1649977179
transform 1 0 2576 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2208 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5244 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1649977179
transform 1 0 4416 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_2_
timestamp 1649977179
transform -1 0 3680 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_3_
timestamp 1649977179
transform 1 0 4600 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_33.mux_l1_in_3__276
timestamp 1649977179
transform -1 0 4048 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1649977179
transform -1 0 4416 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2392 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 14996 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1649977179
transform -1 0 18308 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_3_
timestamp 1649977179
transform 1 0 18952 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_4_
timestamp 1649977179
transform -1 0 16376 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 18308 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1649977179
transform 1 0 18124 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1649977179
transform -1 0 18032 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_0.mux_l2_in_3__279
timestamp 1649977179
transform 1 0 20056 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1649977179
transform 1 0 19228 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1649977179
transform -1 0 18860 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1649977179
transform -1 0 19228 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1649977179
transform -1 0 20056 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 20056 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1649977179
transform -1 0 14444 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1649977179
transform 1 0 17480 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_2_
timestamp 1649977179
transform -1 0 18308 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_3_
timestamp 1649977179
transform 1 0 20424 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_4_
timestamp 1649977179
transform -1 0 15180 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1649977179
transform -1 0 17572 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1649977179
transform 1 0 20332 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1649977179
transform -1 0 19136 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_2.mux_l2_in_3__281
timestamp 1649977179
transform 1 0 20056 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1649977179
transform 1 0 19504 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1649977179
transform 1 0 19780 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1649977179
transform -1 0 19780 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1649977179
transform -1 0 20056 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 19780 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1649977179
transform -1 0 11132 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1649977179
transform -1 0 11960 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1649977179
transform 1 0 19780 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1649977179
transform -1 0 21436 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1649977179
transform -1 0 21344 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_4_
timestamp 1649977179
transform -1 0 21252 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_5_
timestamp 1649977179
transform -1 0 12328 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_6_
timestamp 1649977179
transform -1 0 19136 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_4.mux_l2_in_7__284
timestamp 1649977179
transform 1 0 21344 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_7_
timestamp 1649977179
transform -1 0 20424 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1649977179
transform -1 0 19136 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1649977179
transform 1 0 20700 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_2_
timestamp 1649977179
transform 1 0 20700 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_3_
timestamp 1649977179
transform 1 0 20608 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_1_
timestamp 1649977179
transform -1 0 19780 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l5_in_0_
timestamp 1649977179
transform 1 0 19136 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 18584 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1649977179
transform -1 0 14812 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1649977179
transform 1 0 17480 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_2_
timestamp 1649977179
transform 1 0 15272 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1649977179
transform 1 0 16560 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1649977179
transform -1 0 15364 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1649977179
transform 1 0 15640 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_8.mux_l2_in_3__285
timestamp 1649977179
transform -1 0 16468 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1649977179
transform 1 0 15732 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1649977179
transform -1 0 16192 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1649977179
transform -1 0 16284 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 19872 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1649977179
transform -1 0 15180 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1649977179
transform 1 0 16468 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1649977179
transform -1 0 15456 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1649977179
transform 1 0 15456 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1649977179
transform -1 0 15456 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_2_
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_16.mux_l2_in_3__280
timestamp 1649977179
transform -1 0 16928 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_3_
timestamp 1649977179
transform 1 0 17204 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1649977179
transform -1 0 16100 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_1_
timestamp 1649977179
transform -1 0 16928 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l4_in_0_
timestamp 1649977179
transform -1 0 17756 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 20516 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1649977179
transform -1 0 18216 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1649977179
transform 1 0 18952 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1649977179
transform -1 0 18768 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1649977179
transform 1 0 18124 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1649977179
transform 1 0 18216 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_2_
timestamp 1649977179
transform -1 0 20056 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_24.mux_l2_in_3__282
timestamp 1649977179
transform -1 0 20240 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_3_
timestamp 1649977179
transform -1 0 20792 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1649977179
transform -1 0 18308 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_1_
timestamp 1649977179
transform 1 0 20056 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l4_in_0_
timestamp 1649977179
transform 1 0 19688 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 19964 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1649977179
transform -1 0 15824 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1649977179
transform 1 0 18308 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_2_
timestamp 1649977179
transform -1 0 15640 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_3_
timestamp 1649977179
transform 1 0 17940 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_32.mux_l1_in_3__283
timestamp 1649977179
transform -1 0 18400 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1649977179
transform 1 0 17572 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1649977179
transform 1 0 17112 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1649977179
transform -1 0 17572 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 19044 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 3128 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 2852 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 4324 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_3_
timestamp 1649977179
transform 1 0 4508 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_4_
timestamp 1649977179
transform 1 0 5152 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 3588 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1649977179
transform -1 0 3680 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1649977179
transform 1 0 3956 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_0.mux_l2_in_3__286
timestamp 1649977179
transform 1 0 3772 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1649977179
transform 1 0 2944 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1649977179
transform -1 0 2944 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1649977179
transform -1 0 3680 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 8832 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1649977179
transform -1 0 6256 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_2_
timestamp 1649977179
transform 1 0 6900 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_3_
timestamp 1649977179
transform 1 0 6624 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_4_
timestamp 1649977179
transform 1 0 6532 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5428 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1649977179
transform 1 0 5704 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_2_
timestamp 1649977179
transform 1 0 5428 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_2.mux_l2_in_3__288
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_3_
timestamp 1649977179
transform 1 0 5612 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4876 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_1_
timestamp 1649977179
transform 1 0 4600 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l4_in_0_
timestamp 1649977179
transform -1 0 5428 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 10120 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1649977179
transform -1 0 3956 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1649977179
transform 1 0 5428 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_2_
timestamp 1649977179
transform 1 0 9752 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_3_
timestamp 1649977179
transform 1 0 7728 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_4_
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_5_
timestamp 1649977179
transform -1 0 9384 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_6_
timestamp 1649977179
transform 1 0 8004 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_4.mux_l2_in_7__291
timestamp 1649977179
transform -1 0 8004 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_7_
timestamp 1649977179
transform 1 0 8004 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1649977179
transform -1 0 3680 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_1_
timestamp 1649977179
transform 1 0 6900 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_2_
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_3_
timestamp 1649977179
transform -1 0 8556 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_0_
timestamp 1649977179
transform -1 0 7728 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_1_
timestamp 1649977179
transform -1 0 8556 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l5_in_0_
timestamp 1649977179
transform -1 0 9384 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 10672 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1649977179
transform -1 0 4784 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1649977179
transform 1 0 10304 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_2_
timestamp 1649977179
transform 1 0 10764 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1649977179
transform -1 0 9936 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1649977179
transform -1 0 10488 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_2_
timestamp 1649977179
transform -1 0 10304 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_8.mux_l2_in_3__292
timestamp 1649977179
transform 1 0 11592 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_3_
timestamp 1649977179
transform 1 0 9936 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1649977179
transform 1 0 10488 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_1_
timestamp 1649977179
transform 1 0 9476 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l4_in_0_
timestamp 1649977179
transform -1 0 8832 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 9660 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1649977179
transform -1 0 7544 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1649977179
transform 1 0 12328 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_2_
timestamp 1649977179
transform -1 0 13064 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1649977179
transform 1 0 11868 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1649977179
transform 1 0 12696 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_2_
timestamp 1649977179
transform -1 0 12328 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_3_
timestamp 1649977179
transform -1 0 12972 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_16.mux_l2_in_3__287
timestamp 1649977179
transform 1 0 13524 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1649977179
transform -1 0 12144 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_1_
timestamp 1649977179
transform -1 0 13800 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l4_in_0_
timestamp 1649977179
transform 1 0 12972 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 12328 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1649977179
transform -1 0 14996 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1649977179
transform 1 0 15548 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_2_
timestamp 1649977179
transform 1 0 17204 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1649977179
transform -1 0 15180 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_2_
timestamp 1649977179
transform -1 0 15548 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_24.mux_l2_in_3__289
timestamp 1649977179
transform -1 0 16836 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_3_
timestamp 1649977179
transform 1 0 16376 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1649977179
transform 1 0 15732 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_1_
timestamp 1649977179
transform 1 0 14904 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l4_in_0_
timestamp 1649977179
transform -1 0 14996 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 15272 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1649977179
transform -1 0 11316 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_1_
timestamp 1649977179
transform -1 0 13616 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_2_
timestamp 1649977179
transform 1 0 12236 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_32.mux_l1_in_3__290
timestamp 1649977179
transform -1 0 13432 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_3_
timestamp 1649977179
transform 1 0 13064 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1649977179
transform 1 0 13892 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1649977179
transform -1 0 12788 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1649977179
transform -1 0 13156 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 16192 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1649977179
transform -1 0 18676 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1649977179
transform 1 0 4232 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1649977179
transform -1 0 1748 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1649977179
transform -1 0 2116 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1649977179
transform -1 0 1748 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1649977179
transform -1 0 2116 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1649977179
transform -1 0 1748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1649977179
transform -1 0 2116 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1649977179
transform -1 0 1748 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1649977179
transform -1 0 1748 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1649977179
transform -1 0 1748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1649977179
transform -1 0 2116 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1649977179
transform -1 0 2116 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 1649977179
transform -1 0 1748 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 1649977179
transform -1 0 1748 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 1649977179
transform -1 0 1748 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1649977179
transform -1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1649977179
transform -1 0 1748 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1649977179
transform -1 0 2116 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1649977179
transform -1 0 1748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 1649977179
transform -1 0 1748 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp 1649977179
transform 1 0 21252 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 1649977179
transform 1 0 21252 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 1649977179
transform 1 0 20884 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 1649977179
transform 1 0 21252 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp 1649977179
transform 1 0 21252 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp 1649977179
transform 1 0 21252 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp 1649977179
transform 1 0 20884 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp 1649977179
transform 1 0 21252 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output151
timestamp 1649977179
transform 1 0 21252 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output152
timestamp 1649977179
transform 1 0 21252 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output153
timestamp 1649977179
transform 1 0 20884 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output154
timestamp 1649977179
transform 1 0 21252 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output155
timestamp 1649977179
transform 1 0 20884 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output156
timestamp 1649977179
transform 1 0 21252 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output157
timestamp 1649977179
transform 1 0 21252 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output158
timestamp 1649977179
transform 1 0 21252 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output159
timestamp 1649977179
transform 1 0 21252 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output160
timestamp 1649977179
transform 1 0 20884 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output161
timestamp 1649977179
transform 1 0 21252 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output162
timestamp 1649977179
transform 1 0 21252 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output163
timestamp 1649977179
transform -1 0 12972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output164
timestamp 1649977179
transform -1 0 17388 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output165
timestamp 1649977179
transform -1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output166
timestamp 1649977179
transform -1 0 18124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output167
timestamp 1649977179
transform -1 0 18492 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output168
timestamp 1649977179
transform 1 0 18492 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output169
timestamp 1649977179
transform 1 0 17756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output170
timestamp 1649977179
transform 1 0 20056 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output171
timestamp 1649977179
transform -1 0 19596 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output172
timestamp 1649977179
transform -1 0 20148 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output173
timestamp 1649977179
transform -1 0 20516 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output174
timestamp 1649977179
transform 1 0 12972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output175
timestamp 1649977179
transform 1 0 13340 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output176
timestamp 1649977179
transform -1 0 15272 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output177
timestamp 1649977179
transform 1 0 15272 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output178
timestamp 1649977179
transform -1 0 15456 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output179
timestamp 1649977179
transform 1 0 15640 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output180
timestamp 1649977179
transform -1 0 16376 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output181
timestamp 1649977179
transform 1 0 15548 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output182
timestamp 1649977179
transform -1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output183
timestamp 1649977179
transform 1 0 10120 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output184
timestamp 1649977179
transform -1 0 15180 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output185
timestamp 1649977179
transform -1 0 15548 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output186
timestamp 1649977179
transform -1 0 15916 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output187
timestamp 1649977179
transform -1 0 16284 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output188
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output189
timestamp 1649977179
transform -1 0 17388 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output190
timestamp 1649977179
transform 1 0 17388 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output191
timestamp 1649977179
transform 1 0 17756 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output192
timestamp 1649977179
transform 1 0 18124 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output193
timestamp 1649977179
transform 1 0 18492 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output194
timestamp 1649977179
transform 1 0 11316 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output195
timestamp 1649977179
transform 1 0 11684 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output196
timestamp 1649977179
transform 1 0 12052 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output197
timestamp 1649977179
transform 1 0 12420 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output198
timestamp 1649977179
transform -1 0 13156 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output199
timestamp 1649977179
transform 1 0 13156 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output200
timestamp 1649977179
transform -1 0 13892 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output201
timestamp 1649977179
transform -1 0 14444 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output202
timestamp 1649977179
transform -1 0 14812 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output203
timestamp 1649977179
transform 1 0 20148 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output204
timestamp 1649977179
transform -1 0 1748 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output205
timestamp 1649977179
transform 1 0 19780 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output206
timestamp 1649977179
transform 1 0 21252 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output207
timestamp 1649977179
transform 1 0 20516 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output208
timestamp 1649977179
transform -1 0 2116 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output209
timestamp 1649977179
transform -1 0 19780 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output210
timestamp 1649977179
transform 1 0 20516 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output211
timestamp 1649977179
transform 1 0 20884 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output212
timestamp 1649977179
transform -1 0 2484 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output213
timestamp 1649977179
transform 1 0 20332 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output214
timestamp 1649977179
transform -1 0 2116 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output215
timestamp 1649977179
transform -1 0 18584 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output216
timestamp 1649977179
transform -1 0 18308 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output217
timestamp 1649977179
transform -1 0 15272 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output218
timestamp 1649977179
transform 1 0 7360 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output219
timestamp 1649977179
transform -1 0 19136 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output220
timestamp 1649977179
transform 1 0 20240 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output221
timestamp 1649977179
transform 1 0 21252 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output222
timestamp 1649977179
transform -1 0 2852 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  prog_clk_0_FTB00
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_1_E_FTB01
timestamp 1649977179
transform -1 0 19964 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_1_W_FTB01
timestamp 1649977179
transform 1 0 18216 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_E_FTB01 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20700 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_N_FTB01
timestamp 1649977179
transform 1 0 20700 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_S_FTB01
timestamp 1649977179
transform 1 0 20608 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_W_FTB01
timestamp 1649977179
transform -1 0 20608 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_3_E_FTB01
timestamp 1649977179
transform 1 0 19320 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_3_N_FTB01
timestamp 1649977179
transform -1 0 18860 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_3_S_FTB01
timestamp 1649977179
transform -1 0 20976 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_3_W_FTB01
timestamp 1649977179
transform 1 0 17940 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater223
timestamp 1649977179
transform -1 0 8832 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater224
timestamp 1649977179
transform -1 0 4968 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater225
timestamp 1649977179
transform 1 0 6256 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater226
timestamp 1649977179
transform -1 0 5244 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater227
timestamp 1649977179
transform -1 0 20424 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater228
timestamp 1649977179
transform -1 0 20700 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater229
timestamp 1649977179
transform -1 0 20700 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater230
timestamp 1649977179
transform -1 0 16928 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater231
timestamp 1649977179
transform -1 0 3864 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  repeater232
timestamp 1649977179
transform 1 0 6440 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater233
timestamp 1649977179
transform 1 0 4508 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater234
timestamp 1649977179
transform 1 0 6440 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  repeater235
timestamp 1649977179
transform 1 0 7268 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater236
timestamp 1649977179
transform 1 0 9016 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  repeater237
timestamp 1649977179
transform -1 0 12604 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater238
timestamp 1649977179
transform -1 0 16468 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater239
timestamp 1649977179
transform -1 0 2484 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater240
timestamp 1649977179
transform 1 0 2576 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater241
timestamp 1649977179
transform 1 0 5060 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater242
timestamp 1649977179
transform 1 0 4232 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater243
timestamp 1649977179
transform 1 0 7268 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater244
timestamp 1649977179
transform 1 0 14904 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater245
timestamp 1649977179
transform 1 0 3956 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater246
timestamp 1649977179
transform 1 0 7544 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater247
timestamp 1649977179
transform -1 0 8280 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater248
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater249
timestamp 1649977179
transform 1 0 11500 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater250
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater251
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater252
timestamp 1649977179
transform 1 0 5152 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater253
timestamp 1649977179
transform -1 0 8556 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater254
timestamp 1649977179
transform 1 0 9752 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater255
timestamp 1649977179
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater256
timestamp 1649977179
transform 1 0 13156 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater257
timestamp 1649977179
transform -1 0 13800 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater258
timestamp 1649977179
transform 1 0 15732 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater259
timestamp 1649977179
transform 1 0 16008 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater260
timestamp 1649977179
transform 1 0 10764 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater261
timestamp 1649977179
transform -1 0 14168 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater262
timestamp 1649977179
transform 1 0 15456 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater263
timestamp 1649977179
transform 1 0 17756 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater264
timestamp 1649977179
transform -1 0 18584 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater265
timestamp 1649977179
transform 1 0 18584 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater266
timestamp 1649977179
transform 1 0 7544 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater267
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater268
timestamp 1649977179
transform 1 0 15916 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater269
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater270
timestamp 1649977179
transform -1 0 18676 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater271
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater272
timestamp 1649977179
transform -1 0 19136 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater273
timestamp 1649977179
transform -1 0 19596 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater274
timestamp 1649977179
transform -1 0 21160 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater275
timestamp 1649977179
transform 1 0 19872 0 -1 19584
box -38 -48 406 592
<< labels >>
flabel metal2 s 18234 22200 18290 23000 0 FreeSans 224 90 0 0 Test_en_N_out
port 0 nsew signal tristate
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 Test_en_S_in
port 1 nsew signal input
flabel metal4 s 6142 2128 6462 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 11340 2128 11660 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 16538 2128 16858 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 21736 2128 22056 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 3543 2128 3863 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal4 s 8741 2128 9061 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal4 s 13939 2128 14259 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal4 s 19137 2128 19457 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal2 s 1490 0 1546 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_42_
port 4 nsew signal input
flabel metal2 s 1858 0 1914 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_43_
port 5 nsew signal input
flabel metal2 s 2226 0 2282 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_44_
port 6 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_45_
port 7 nsew signal input
flabel metal2 s 2962 0 3018 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_46_
port 8 nsew signal input
flabel metal2 s 3330 0 3386 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_47_
port 9 nsew signal input
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_48_
port 10 nsew signal input
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_49_
port 11 nsew signal input
flabel metal2 s 4434 0 4490 800 0 FreeSans 224 90 0 0 ccff_head
port 12 nsew signal input
flabel metal2 s 4802 0 4858 800 0 FreeSans 224 90 0 0 ccff_tail
port 13 nsew signal tristate
flabel metal3 s 0 3816 800 3936 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 14 nsew signal input
flabel metal3 s 0 7896 800 8016 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 15 nsew signal input
flabel metal3 s 0 8304 800 8424 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 16 nsew signal input
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 17 nsew signal input
flabel metal3 s 0 9120 800 9240 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 18 nsew signal input
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 19 nsew signal input
flabel metal3 s 0 9936 800 10056 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 20 nsew signal input
flabel metal3 s 0 10344 800 10464 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 21 nsew signal input
flabel metal3 s 0 10752 800 10872 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 22 nsew signal input
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 23 nsew signal input
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 chanx_left_in[19]
port 24 nsew signal input
flabel metal3 s 0 4224 800 4344 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 25 nsew signal input
flabel metal3 s 0 4632 800 4752 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 26 nsew signal input
flabel metal3 s 0 5040 800 5160 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 27 nsew signal input
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 28 nsew signal input
flabel metal3 s 0 5856 800 5976 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 29 nsew signal input
flabel metal3 s 0 6264 800 6384 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 30 nsew signal input
flabel metal3 s 0 6672 800 6792 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 31 nsew signal input
flabel metal3 s 0 7080 800 7200 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 32 nsew signal input
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 33 nsew signal input
flabel metal3 s 0 11976 800 12096 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 34 nsew signal tristate
flabel metal3 s 0 16056 800 16176 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 35 nsew signal tristate
flabel metal3 s 0 16464 800 16584 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 36 nsew signal tristate
flabel metal3 s 0 16872 800 16992 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 37 nsew signal tristate
flabel metal3 s 0 17280 800 17400 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 38 nsew signal tristate
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 39 nsew signal tristate
flabel metal3 s 0 18096 800 18216 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 40 nsew signal tristate
flabel metal3 s 0 18504 800 18624 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 41 nsew signal tristate
flabel metal3 s 0 18912 800 19032 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 42 nsew signal tristate
flabel metal3 s 0 19320 800 19440 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 43 nsew signal tristate
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 chanx_left_out[19]
port 44 nsew signal tristate
flabel metal3 s 0 12384 800 12504 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 45 nsew signal tristate
flabel metal3 s 0 12792 800 12912 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 46 nsew signal tristate
flabel metal3 s 0 13200 800 13320 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 47 nsew signal tristate
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 48 nsew signal tristate
flabel metal3 s 0 14016 800 14136 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 49 nsew signal tristate
flabel metal3 s 0 14424 800 14544 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 50 nsew signal tristate
flabel metal3 s 0 14832 800 14952 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 51 nsew signal tristate
flabel metal3 s 0 15240 800 15360 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 52 nsew signal tristate
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 53 nsew signal tristate
flabel metal3 s 22200 3816 23000 3936 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 54 nsew signal input
flabel metal3 s 22200 7896 23000 8016 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 55 nsew signal input
flabel metal3 s 22200 8304 23000 8424 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 56 nsew signal input
flabel metal3 s 22200 8712 23000 8832 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 57 nsew signal input
flabel metal3 s 22200 9120 23000 9240 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 58 nsew signal input
flabel metal3 s 22200 9528 23000 9648 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 59 nsew signal input
flabel metal3 s 22200 9936 23000 10056 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 60 nsew signal input
flabel metal3 s 22200 10344 23000 10464 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 61 nsew signal input
flabel metal3 s 22200 10752 23000 10872 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 62 nsew signal input
flabel metal3 s 22200 11160 23000 11280 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 63 nsew signal input
flabel metal3 s 22200 11568 23000 11688 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 64 nsew signal input
flabel metal3 s 22200 4224 23000 4344 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 65 nsew signal input
flabel metal3 s 22200 4632 23000 4752 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 66 nsew signal input
flabel metal3 s 22200 5040 23000 5160 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 67 nsew signal input
flabel metal3 s 22200 5448 23000 5568 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 68 nsew signal input
flabel metal3 s 22200 5856 23000 5976 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 69 nsew signal input
flabel metal3 s 22200 6264 23000 6384 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 70 nsew signal input
flabel metal3 s 22200 6672 23000 6792 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 71 nsew signal input
flabel metal3 s 22200 7080 23000 7200 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 72 nsew signal input
flabel metal3 s 22200 7488 23000 7608 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 73 nsew signal input
flabel metal3 s 22200 11976 23000 12096 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 74 nsew signal tristate
flabel metal3 s 22200 16056 23000 16176 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 75 nsew signal tristate
flabel metal3 s 22200 16464 23000 16584 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 76 nsew signal tristate
flabel metal3 s 22200 16872 23000 16992 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 77 nsew signal tristate
flabel metal3 s 22200 17280 23000 17400 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 78 nsew signal tristate
flabel metal3 s 22200 17688 23000 17808 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 79 nsew signal tristate
flabel metal3 s 22200 18096 23000 18216 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 80 nsew signal tristate
flabel metal3 s 22200 18504 23000 18624 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 81 nsew signal tristate
flabel metal3 s 22200 18912 23000 19032 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 82 nsew signal tristate
flabel metal3 s 22200 19320 23000 19440 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 83 nsew signal tristate
flabel metal3 s 22200 19728 23000 19848 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 84 nsew signal tristate
flabel metal3 s 22200 12384 23000 12504 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 85 nsew signal tristate
flabel metal3 s 22200 12792 23000 12912 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 86 nsew signal tristate
flabel metal3 s 22200 13200 23000 13320 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 87 nsew signal tristate
flabel metal3 s 22200 13608 23000 13728 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 88 nsew signal tristate
flabel metal3 s 22200 14016 23000 14136 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 89 nsew signal tristate
flabel metal3 s 22200 14424 23000 14544 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 90 nsew signal tristate
flabel metal3 s 22200 14832 23000 14952 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 91 nsew signal tristate
flabel metal3 s 22200 15240 23000 15360 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 92 nsew signal tristate
flabel metal3 s 22200 15648 23000 15768 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 93 nsew signal tristate
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 94 nsew signal input
flabel metal2 s 8850 0 8906 800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 95 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 96 nsew signal input
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 97 nsew signal input
flabel metal2 s 9954 0 10010 800 0 FreeSans 224 90 0 0 chany_bottom_in[13]
port 98 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 99 nsew signal input
flabel metal2 s 10690 0 10746 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 100 nsew signal input
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 chany_bottom_in[16]
port 101 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 102 nsew signal input
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 103 nsew signal input
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 chany_bottom_in[19]
port 104 nsew signal input
flabel metal2 s 5538 0 5594 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 105 nsew signal input
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 106 nsew signal input
flabel metal2 s 6274 0 6330 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 107 nsew signal input
flabel metal2 s 6642 0 6698 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 108 nsew signal input
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 109 nsew signal input
flabel metal2 s 7378 0 7434 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 110 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 111 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 112 nsew signal input
flabel metal2 s 8482 0 8538 800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 113 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 114 nsew signal tristate
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 chany_bottom_out[10]
port 115 nsew signal tristate
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 chany_bottom_out[11]
port 116 nsew signal tristate
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 chany_bottom_out[12]
port 117 nsew signal tristate
flabel metal2 s 17314 0 17370 800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 118 nsew signal tristate
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 chany_bottom_out[14]
port 119 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 120 nsew signal tristate
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 chany_bottom_out[16]
port 121 nsew signal tristate
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 122 nsew signal tristate
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 123 nsew signal tristate
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 chany_bottom_out[19]
port 124 nsew signal tristate
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 125 nsew signal tristate
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 126 nsew signal tristate
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 127 nsew signal tristate
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 128 nsew signal tristate
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 129 nsew signal tristate
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 130 nsew signal tristate
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 131 nsew signal tristate
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 chany_bottom_out[8]
port 132 nsew signal tristate
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 133 nsew signal tristate
flabel metal2 s 3514 22200 3570 23000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 134 nsew signal input
flabel metal2 s 7194 22200 7250 23000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 135 nsew signal input
flabel metal2 s 7562 22200 7618 23000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 136 nsew signal input
flabel metal2 s 7930 22200 7986 23000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 137 nsew signal input
flabel metal2 s 8298 22200 8354 23000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 138 nsew signal input
flabel metal2 s 8666 22200 8722 23000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 139 nsew signal input
flabel metal2 s 9034 22200 9090 23000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 140 nsew signal input
flabel metal2 s 9402 22200 9458 23000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 141 nsew signal input
flabel metal2 s 9770 22200 9826 23000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 142 nsew signal input
flabel metal2 s 10138 22200 10194 23000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 143 nsew signal input
flabel metal2 s 10506 22200 10562 23000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 144 nsew signal input
flabel metal2 s 3882 22200 3938 23000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 145 nsew signal input
flabel metal2 s 4250 22200 4306 23000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 146 nsew signal input
flabel metal2 s 4618 22200 4674 23000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 147 nsew signal input
flabel metal2 s 4986 22200 5042 23000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 148 nsew signal input
flabel metal2 s 5354 22200 5410 23000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 149 nsew signal input
flabel metal2 s 5722 22200 5778 23000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 150 nsew signal input
flabel metal2 s 6090 22200 6146 23000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 151 nsew signal input
flabel metal2 s 6458 22200 6514 23000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 152 nsew signal input
flabel metal2 s 6826 22200 6882 23000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 153 nsew signal input
flabel metal2 s 10874 22200 10930 23000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 154 nsew signal tristate
flabel metal2 s 14554 22200 14610 23000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 155 nsew signal tristate
flabel metal2 s 14922 22200 14978 23000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 156 nsew signal tristate
flabel metal2 s 15290 22200 15346 23000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 157 nsew signal tristate
flabel metal2 s 15658 22200 15714 23000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 158 nsew signal tristate
flabel metal2 s 16026 22200 16082 23000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 159 nsew signal tristate
flabel metal2 s 16394 22200 16450 23000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 160 nsew signal tristate
flabel metal2 s 16762 22200 16818 23000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 161 nsew signal tristate
flabel metal2 s 17130 22200 17186 23000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 162 nsew signal tristate
flabel metal2 s 17498 22200 17554 23000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 163 nsew signal tristate
flabel metal2 s 17866 22200 17922 23000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 164 nsew signal tristate
flabel metal2 s 11242 22200 11298 23000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 165 nsew signal tristate
flabel metal2 s 11610 22200 11666 23000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 166 nsew signal tristate
flabel metal2 s 11978 22200 12034 23000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 167 nsew signal tristate
flabel metal2 s 12346 22200 12402 23000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 168 nsew signal tristate
flabel metal2 s 12714 22200 12770 23000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 169 nsew signal tristate
flabel metal2 s 13082 22200 13138 23000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 170 nsew signal tristate
flabel metal2 s 13450 22200 13506 23000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 171 nsew signal tristate
flabel metal2 s 13818 22200 13874 23000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 172 nsew signal tristate
flabel metal2 s 14186 22200 14242 23000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 173 nsew signal tristate
flabel metal3 s 22200 20136 23000 20256 0 FreeSans 480 0 0 0 clk_1_E_out
port 174 nsew signal tristate
flabel metal2 s 18602 22200 18658 23000 0 FreeSans 224 90 0 0 clk_1_N_in
port 175 nsew signal input
flabel metal3 s 0 20136 800 20256 0 FreeSans 480 0 0 0 clk_1_W_out
port 176 nsew signal tristate
flabel metal3 s 22200 20544 23000 20664 0 FreeSans 480 0 0 0 clk_2_E_out
port 177 nsew signal tristate
flabel metal2 s 18970 22200 19026 23000 0 FreeSans 224 90 0 0 clk_2_N_in
port 178 nsew signal input
flabel metal2 s 21178 22200 21234 23000 0 FreeSans 224 90 0 0 clk_2_N_out
port 179 nsew signal tristate
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 clk_2_S_out
port 180 nsew signal tristate
flabel metal3 s 0 20544 800 20664 0 FreeSans 480 0 0 0 clk_2_W_out
port 181 nsew signal tristate
flabel metal3 s 22200 20952 23000 21072 0 FreeSans 480 0 0 0 clk_3_E_out
port 182 nsew signal tristate
flabel metal2 s 19338 22200 19394 23000 0 FreeSans 224 90 0 0 clk_3_N_in
port 183 nsew signal input
flabel metal2 s 21546 22200 21602 23000 0 FreeSans 224 90 0 0 clk_3_N_out
port 184 nsew signal tristate
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 clk_3_S_out
port 185 nsew signal tristate
flabel metal3 s 0 20952 800 21072 0 FreeSans 480 0 0 0 clk_3_W_out
port 186 nsew signal tristate
flabel metal3 s 0 552 800 672 0 FreeSans 480 0 0 0 left_bottom_grid_pin_34_
port 187 nsew signal input
flabel metal3 s 0 960 800 1080 0 FreeSans 480 0 0 0 left_bottom_grid_pin_35_
port 188 nsew signal input
flabel metal3 s 0 1368 800 1488 0 FreeSans 480 0 0 0 left_bottom_grid_pin_36_
port 189 nsew signal input
flabel metal3 s 0 1776 800 1896 0 FreeSans 480 0 0 0 left_bottom_grid_pin_37_
port 190 nsew signal input
flabel metal3 s 0 2184 800 2304 0 FreeSans 480 0 0 0 left_bottom_grid_pin_38_
port 191 nsew signal input
flabel metal3 s 0 2592 800 2712 0 FreeSans 480 0 0 0 left_bottom_grid_pin_39_
port 192 nsew signal input
flabel metal3 s 0 3000 800 3120 0 FreeSans 480 0 0 0 left_bottom_grid_pin_40_
port 193 nsew signal input
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 left_bottom_grid_pin_41_
port 194 nsew signal input
flabel metal2 s 19706 22200 19762 23000 0 FreeSans 224 90 0 0 prog_clk_0_N_in
port 195 nsew signal input
flabel metal3 s 22200 21360 23000 21480 0 FreeSans 480 0 0 0 prog_clk_1_E_out
port 196 nsew signal tristate
flabel metal2 s 20074 22200 20130 23000 0 FreeSans 224 90 0 0 prog_clk_1_N_in
port 197 nsew signal input
flabel metal3 s 0 21360 800 21480 0 FreeSans 480 0 0 0 prog_clk_1_W_out
port 198 nsew signal tristate
flabel metal3 s 22200 21768 23000 21888 0 FreeSans 480 0 0 0 prog_clk_2_E_out
port 199 nsew signal tristate
flabel metal2 s 20442 22200 20498 23000 0 FreeSans 224 90 0 0 prog_clk_2_N_in
port 200 nsew signal input
flabel metal2 s 21914 22200 21970 23000 0 FreeSans 224 90 0 0 prog_clk_2_N_out
port 201 nsew signal tristate
flabel metal2 s 20994 0 21050 800 0 FreeSans 224 90 0 0 prog_clk_2_S_out
port 202 nsew signal tristate
flabel metal3 s 0 21768 800 21888 0 FreeSans 480 0 0 0 prog_clk_2_W_out
port 203 nsew signal tristate
flabel metal3 s 22200 22176 23000 22296 0 FreeSans 480 0 0 0 prog_clk_3_E_out
port 204 nsew signal tristate
flabel metal2 s 20810 22200 20866 23000 0 FreeSans 224 90 0 0 prog_clk_3_N_in
port 205 nsew signal input
flabel metal2 s 22282 22200 22338 23000 0 FreeSans 224 90 0 0 prog_clk_3_N_out
port 206 nsew signal tristate
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 prog_clk_3_S_out
port 207 nsew signal tristate
flabel metal3 s 0 22176 800 22296 0 FreeSans 480 0 0 0 prog_clk_3_W_out
port 208 nsew signal tristate
flabel metal3 s 22200 552 23000 672 0 FreeSans 480 0 0 0 right_bottom_grid_pin_34_
port 209 nsew signal input
flabel metal3 s 22200 960 23000 1080 0 FreeSans 480 0 0 0 right_bottom_grid_pin_35_
port 210 nsew signal input
flabel metal3 s 22200 1368 23000 1488 0 FreeSans 480 0 0 0 right_bottom_grid_pin_36_
port 211 nsew signal input
flabel metal3 s 22200 1776 23000 1896 0 FreeSans 480 0 0 0 right_bottom_grid_pin_37_
port 212 nsew signal input
flabel metal3 s 22200 2184 23000 2304 0 FreeSans 480 0 0 0 right_bottom_grid_pin_38_
port 213 nsew signal input
flabel metal3 s 22200 2592 23000 2712 0 FreeSans 480 0 0 0 right_bottom_grid_pin_39_
port 214 nsew signal input
flabel metal3 s 22200 3000 23000 3120 0 FreeSans 480 0 0 0 right_bottom_grid_pin_40_
port 215 nsew signal input
flabel metal3 s 22200 3408 23000 3528 0 FreeSans 480 0 0 0 right_bottom_grid_pin_41_
port 216 nsew signal input
flabel metal2 s 570 22200 626 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_42_
port 217 nsew signal input
flabel metal2 s 938 22200 994 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_43_
port 218 nsew signal input
flabel metal2 s 1306 22200 1362 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_44_
port 219 nsew signal input
flabel metal2 s 1674 22200 1730 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_45_
port 220 nsew signal input
flabel metal2 s 2042 22200 2098 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_46_
port 221 nsew signal input
flabel metal2 s 2410 22200 2466 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_47_
port 222 nsew signal input
flabel metal2 s 2778 22200 2834 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_48_
port 223 nsew signal input
flabel metal2 s 3146 22200 3202 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_49_
port 224 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
