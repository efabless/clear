* NGSPICE file created from left_tile.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_1 abstract view
.subckt sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

.subckt left_tile VGND VPWR ccff_head ccff_head_0 ccff_tail ccff_tail_0 chanx_right_in[0]
+ chanx_right_in[10] chanx_right_in[11] chanx_right_in[12] chanx_right_in[13] chanx_right_in[14]
+ chanx_right_in[15] chanx_right_in[16] chanx_right_in[17] chanx_right_in[18] chanx_right_in[19]
+ chanx_right_in[1] chanx_right_in[20] chanx_right_in[21] chanx_right_in[22] chanx_right_in[23]
+ chanx_right_in[24] chanx_right_in[25] chanx_right_in[26] chanx_right_in[27] chanx_right_in[28]
+ chanx_right_in[29] chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5]
+ chanx_right_in[6] chanx_right_in[7] chanx_right_in[8] chanx_right_in[9] chanx_right_out[0]
+ chanx_right_out[10] chanx_right_out[11] chanx_right_out[12] chanx_right_out[13]
+ chanx_right_out[14] chanx_right_out[15] chanx_right_out[16] chanx_right_out[17]
+ chanx_right_out[18] chanx_right_out[19] chanx_right_out[1] chanx_right_out[20] chanx_right_out[21]
+ chanx_right_out[22] chanx_right_out[23] chanx_right_out[24] chanx_right_out[25]
+ chanx_right_out[26] chanx_right_out[27] chanx_right_out[28] chanx_right_out[29]
+ chanx_right_out[2] chanx_right_out[3] chanx_right_out[4] chanx_right_out[5] chanx_right_out[6]
+ chanx_right_out[7] chanx_right_out[8] chanx_right_out[9] chany_bottom_in[0] chany_bottom_in[10]
+ chany_bottom_in[11] chany_bottom_in[12] chany_bottom_in[13] chany_bottom_in[14]
+ chany_bottom_in[15] chany_bottom_in[16] chany_bottom_in[17] chany_bottom_in[18]
+ chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[20] chany_bottom_in[21] chany_bottom_in[22]
+ chany_bottom_in[23] chany_bottom_in[24] chany_bottom_in[25] chany_bottom_in[26]
+ chany_bottom_in[27] chany_bottom_in[28] chany_bottom_in[29] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[20] chany_bottom_out[21] chany_bottom_out[22]
+ chany_bottom_out[23] chany_bottom_out[24] chany_bottom_out[25] chany_bottom_out[26]
+ chany_bottom_out[27] chany_bottom_out[28] chany_bottom_out[29] chany_bottom_out[2]
+ chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6]
+ chany_bottom_out[7] chany_bottom_out[8] chany_bottom_out[9] chany_top_in_0[0] chany_top_in_0[10]
+ chany_top_in_0[11] chany_top_in_0[12] chany_top_in_0[13] chany_top_in_0[14] chany_top_in_0[15]
+ chany_top_in_0[16] chany_top_in_0[17] chany_top_in_0[18] chany_top_in_0[19] chany_top_in_0[1]
+ chany_top_in_0[20] chany_top_in_0[21] chany_top_in_0[22] chany_top_in_0[23] chany_top_in_0[24]
+ chany_top_in_0[25] chany_top_in_0[26] chany_top_in_0[27] chany_top_in_0[28] chany_top_in_0[29]
+ chany_top_in_0[2] chany_top_in_0[3] chany_top_in_0[4] chany_top_in_0[5] chany_top_in_0[6]
+ chany_top_in_0[7] chany_top_in_0[8] chany_top_in_0[9] chany_top_out_0[0] chany_top_out_0[10]
+ chany_top_out_0[11] chany_top_out_0[12] chany_top_out_0[13] chany_top_out_0[14]
+ chany_top_out_0[15] chany_top_out_0[16] chany_top_out_0[17] chany_top_out_0[18]
+ chany_top_out_0[19] chany_top_out_0[1] chany_top_out_0[20] chany_top_out_0[21] chany_top_out_0[22]
+ chany_top_out_0[23] chany_top_out_0[24] chany_top_out_0[25] chany_top_out_0[26]
+ chany_top_out_0[27] chany_top_out_0[28] chany_top_out_0[29] chany_top_out_0[2] chany_top_out_0[3]
+ chany_top_out_0[4] chany_top_out_0[5] chany_top_out_0[6] chany_top_out_0[7] chany_top_out_0[8]
+ chany_top_out_0[9] gfpga_pad_io_soc_dir[0] gfpga_pad_io_soc_dir[1] gfpga_pad_io_soc_dir[2]
+ gfpga_pad_io_soc_dir[3] gfpga_pad_io_soc_in[0] gfpga_pad_io_soc_in[1] gfpga_pad_io_soc_in[2]
+ gfpga_pad_io_soc_in[3] gfpga_pad_io_soc_out[0] gfpga_pad_io_soc_out[1] gfpga_pad_io_soc_out[2]
+ gfpga_pad_io_soc_out[3] isol_n prog_clk prog_reset_bottom_in prog_reset_bottom_out
+ prog_reset_left_in prog_reset_right_out prog_reset_top_in prog_reset_top_out reset_bottom_in
+ reset_bottom_out reset_right_in reset_top_in reset_top_out right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_ right_width_0_height_0_subtile_0__pin_inpad_0_
+ right_width_0_height_0_subtile_1__pin_inpad_0_ right_width_0_height_0_subtile_2__pin_inpad_0_
+ right_width_0_height_0_subtile_3__pin_inpad_0_ test_enable_bottom_in test_enable_bottom_out
+ test_enable_right_in test_enable_top_in test_enable_top_out top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
+ top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_ top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
+ top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
XANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4_ net65 net34 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_0__A1 net116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input92_A chany_top_in_0[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_right_track_16.mux_l2_in_1__A1 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l4_in_0_ cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X cby_0__1_.cby_0__1_.mem_right_ipin_1.ccff_tail
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xcby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_1_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[0\] net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_0__1_.mux_bottom_track_45.mux_l1_in_0__A1 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_14.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_14.out sky130_fd_sc_hd__clkbuf_1
Xsb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_9_0_prog_clk sb_0__1_.mem_right_track_22.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_22.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_0__1_.mux_right_track_34.mux_l1_in_0__A0 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__214__A net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_0__A0 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput220 net220 VGND VGND VPWR VPWR prog_reset_top_out sky130_fd_sc_hd__buf_12
XFILLER_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__209__A net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3__272 VGND VGND VPWR VPWR net272
+ cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3__272/LO sky130_fd_sc_hd__conb_1
Xsb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_5_0_prog_clk sb_0__1_.mem_right_track_54.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_54.ccff_tail sky130_fd_sc_hd__dfrtp_1
X_200_ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__clkbuf_1
Xsb_0__1_.mux_right_track_8.mux_l1_in_0_ net73 net80 sb_0__1_.mem_right_track_8.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
X_131_ sb_0__1_.mux_right_track_12.out VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_0__1_.mux_right_track_26.mux_l1_in_0__A1 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input55_A chany_bottom_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l3_in_1_ cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_bottom_track_11.mux_l1_in_0_ net88 net73 sb_0__1_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_64_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_114_ sb_0__1_.mux_right_track_46.out VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_1
XFILLER_78_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_14.mux_l3_in_0_ sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_1_X sb_0__1_.mem_right_track_14.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_69_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_56.mux_l1_in_0_ net54 net110 sb_0__1_.mem_right_track_56.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_2_ net57 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input18_A chanx_right_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_45.out sky130_fd_sc_hd__clkbuf_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_2__A0 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__217__A net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_8_0_prog_clk sb_0__1_.mem_top_track_10.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_10.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_31_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_right_track_14.mux_l2_in_1_ net235 net39 sb_0__1_.mem_right_track_14.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mux_bottom_track_53.mux_l1_in_0__A1 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3_ net71 net40 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input85_A chany_top_in_0[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_0_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_1.ccff_tail net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xsb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_9_0_prog_clk sb_0__1_.mem_right_track_22.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_22.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_0__1_.mux_right_track_34.mux_l1_in_0__A1 net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_6_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_6_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_0__A1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__140__A net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_top_track_12.mux_l3_in_0_ sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_4_X
+ sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_3_X sb_0__1_.mem_top_track_12.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput221 net221 VGND VGND VPWR VPWR reset_bottom_out sky130_fd_sc_hd__buf_12
Xoutput210 net210 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[0] sky130_fd_sc_hd__buf_12
XFILLER_82_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_top_track_6.mux_l1_in_3_ net270 net59 sb_0__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
X_130_ sb_0__1_.mux_right_track_14.out VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_2
Xsb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_5_0_prog_clk sb_0__1_.mem_right_track_52.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_54.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_65_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input48_A chany_bottom_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_36.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_36.out sky130_fd_sc_hd__clkbuf_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l3_in_0_ cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input102_A reset_right_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_113_ sb_0__1_.mux_right_track_48.out VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_top_track_12.mux_l2_in_1_ net262 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mem_top_track_12.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_1__S sb_0__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_1_ cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2__A0 net76 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_bottom_track_45.mux_l2_in_1__228 VGND VGND VPWR VPWR net228 sb_0__1_.mux_bottom_track_45.mux_l2_in_1__228/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_0__1_.mux_right_track_50.mux_l1_in_0__A0 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_top_track_6.mux_l3_in_0_ sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_5_X
+ sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X sb_0__1_.mem_top_track_10.ccff_head
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_2__A1 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_8_0_prog_clk sb_0__1_.mem_top_track_10.ccff_head
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_10.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xsb_0__1_.mux_top_track_12.mux_l1_in_2_ net56 net42 sb_0__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_40_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput110 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_ VGND VGND VPWR
+ VPWR net110 sky130_fd_sc_hd__buf_2
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input30_A chanx_right_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_right_track_14.mux_l2_in_0_ net105 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_14.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4__A0 net65 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__143__A net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_3.out sky130_fd_sc_hd__clkbuf_1
XFILLER_39_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2_ net78 net47 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_24.mux_l1_in_1__241 VGND VGND VPWR VPWR net241 sb_0__1_.mux_right_track_24.mux_l1_in_1__241/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_22_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_0__A0 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input78_A chany_top_in_0[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_6.mux_l2_in_1__258 VGND VGND VPWR VPWR net258 sb_0__1_.mux_right_track_6.mux_l2_in_1__258/LO
+ sky130_fd_sc_hd__conb_1
Xsb_0__1_.mux_top_track_6.mux_l2_in_1_ sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X sb_0__1_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__138__A net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_9_0_prog_clk sb_0__1_.mem_right_track_20.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_22.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_6_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_ cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_
+ sky130_fd_sc_hd__clkbuf_1
Xoutput200 net200 VGND VGND VPWR VPWR chany_top_out_0[28] sky130_fd_sc_hd__buf_12
Xoutput222 net222 VGND VGND VPWR VPWR reset_top_out sky130_fd_sc_hd__buf_12
XANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput211 net211 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[1] sky130_fd_sc_hd__buf_12
XFILLER_82_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mux_top_track_6.mux_l1_in_2_ net46 net26 sb_0__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_189_ net47 VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__151__A net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_36.mux_l2_in_1__266 VGND VGND VPWR VPWR net266 sb_0__1_.mux_top_track_36.mux_l2_in_1__266/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_47_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_112_ sb_0__1_.mux_right_track_50.out VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_2
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_2_0_prog_clk sb_0__1_.mem_right_track_28.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_28.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_input60_A chany_bottom_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_top_track_12.mux_l2_in_0_ sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_top_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_46_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__146__A net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_0_ cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_75_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_top_track_0.mux_l1_in_3__260 VGND VGND VPWR VPWR net260 sb_0__1_.mux_top_track_0.mux_l1_in_3__260/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2__A1 net45 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_right_track_50.mux_l1_in_0__A1 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_top_track_12.mux_l1_in_1_ net14 net6 sb_0__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_31_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput111 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_ VGND VGND VPWR
+ VPWR net111 sky130_fd_sc_hd__clkbuf_2
Xinput100 prog_reset_top_in VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_3__A1 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input23_A chanx_right_in[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_6_0_prog_clk sb_0__1_.mem_bottom_track_11.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_11.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4__A1 net34 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1_ net81 net50 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_62_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_0__A1 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mux_right_track_28.mux_l1_in_1__A1 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_6.mux_l2_in_0_ sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_21_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__154__A net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mux_right_track_36.mux_l2_in_0__A0 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_14.mux_l1_in_0_ net69 net70 sb_0__1_.mem_right_track_14.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_7_0_prog_clk sb_0__1_.mem_bottom_track_5.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_5.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3__A1 net88 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input90_A chany_top_in_0[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_26.mux_l2_in_0_ sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_26.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_32_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput201 net201 VGND VGND VPWR VPWR chany_top_out_0[29] sky130_fd_sc_hd__buf_12
Xoutput223 net223 VGND VGND VPWR VPWR test_enable_bottom_out sky130_fd_sc_hd__buf_12
Xoutput212 net212 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[2] sky130_fd_sc_hd__buf_12
XFILLER_59_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_4_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_top_track_6.mux_l1_in_1_ net8 net20 sb_0__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_23_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_188_ net46 VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_2
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_bottom_track_3.mux_l3_in_0_ sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X sb_0__1_.mem_bottom_track_3.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_70_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_right_track_26.mux_l1_in_1_ net242 net60 sb_0__1_.mem_right_track_26.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
X_111_ sb_0__1_.mux_right_track_52.out VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_1
XFILLER_78_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_3_0_prog_clk sb_0__1_.mem_right_track_26.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_28.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_input53_A chany_bottom_in[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_bottom_track_3.mux_l2_in_1_ net226 right_width_0_height_0_subtile_1__pin_inpad_0_
+ sb_0__1_.mem_bottom_track_3.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_4_0_prog_clk sb_0__1_.mem_right_track_40.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_40.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mux_top_track_12.mux_l1_in_0_ net18 net115 sb_0__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_31_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput112 test_enable_bottom_in VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__buf_2
Xinput101 reset_bottom_in VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__buf_2
XANTENNA_input16_A chanx_right_in[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_6_0_prog_clk sb_0__1_.mem_bottom_track_11.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_11.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_4_9_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_0_ sb_0__1_.mux_bottom_track_3.out
+ net53 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_top_track_36.mux_l3_in_0_ sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X sb_0__1_.mem_top_track_36.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_89_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input8_A chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net94 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR right_width_0_height_0_subtile_2__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__170__A net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mux_right_track_0.mux_l1_in_0__A0 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_3__A1 right_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_7_0_prog_clk sb_0__1_.mem_bottom_track_5.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_5.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_37_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input118_A top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input83_A chany_top_in_0[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_36.mux_l2_in_1_ net266 net38 sb_0__1_.mem_top_track_36.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_32_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput224 net224 VGND VGND VPWR VPWR test_enable_top_out sky130_fd_sc_hd__buf_12
Xoutput202 net202 VGND VGND VPWR VPWR chany_top_out_0[2] sky130_fd_sc_hd__buf_12
Xoutput213 net213 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[3] sky130_fd_sc_hd__buf_12
XFILLER_82_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_top_track_6.mux_l1_in_0_ net117 net115 sb_0__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_23_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ net119 net97 VGND VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_1
X_187_ sb_0__1_.mux_top_track_20.out VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__clkbuf_1
XFILLER_80_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_4.mux_l3_in_0_ sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X sb_0__1_.mem_right_track_4.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_55_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_5_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_5_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_70_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_110_ sb_0__1_.mux_right_track_54.out VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_1
Xsb_0__1_.mux_right_track_26.mux_l1_in_0_ net111 net90 sb_0__1_.mem_right_track_26.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_93_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input46_A chany_bottom_in[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_right_track_38.mux_l2_in_0_ net248 sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_38.ccff_tail VGND VGND VPWR VPWR sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_52_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input100_A prog_reset_top_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_right_track_40.mux_l2_in_0_ net250 sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_40.ccff_tail VGND VGND VPWR VPWR sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mux_right_track_10.mux_l1_in_1__A0 net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_4.mux_l2_in_1_ net249 net47 sb_0__1_.mem_right_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__173__A net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_bottom_track_3.mux_l2_in_0_ sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_bottom_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XFILLER_72_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_1_0_prog_clk sb_0__1_.mem_right_track_38.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_40.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_25_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput113 test_enable_right_in VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__clkbuf_1
Xinput102 reset_right_in VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_6_0_prog_clk sb_0__1_.mem_bottom_track_11.ccff_head
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_11.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__168__A net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_14_0_prog_clk sb_0__1_.mem_right_track_14.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_14.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mux_bottom_track_3.mux_l1_in_1_ net4 net16 sb_0__1_.mem_bottom_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_36_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__1_.mux_right_track_0.mux_l1_in_0__A1 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_20.out sky130_fd_sc_hd__clkbuf_1
XFILLER_94_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_7_0_prog_clk sb_0__1_.mem_bottom_track_3.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_5.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_85_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input76_A chany_top_in_0[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_5_0_prog_clk sb_0__1_.mem_right_track_46.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_46.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_top_track_36.mux_l2_in_0_ net32 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_top_track_36.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput203 net203 VGND VGND VPWR VPWR chany_top_out_0[3] sky130_fd_sc_hd__buf_12
XANTENNA__181__A net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput214 net214 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[0] sky130_fd_sc_hd__buf_12
XANTENNA_sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_186_ net43 VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__176__A net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input39_A chany_bottom_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_169_ net55 VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__clkbuf_2
XFILLER_69_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.ccff_tail net97 VGND
+ VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_1
XFILLER_20_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_right_track_10.mux_l1_in_1__A1 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_4.mux_l2_in_0_ sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_13_0_prog_clk sb_0__1_.mem_right_track_0.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput103 reset_top_in VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_1
Xinput114 test_enable_top_in VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_1
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_right_track_38.mux_l1_in_0_ net57 net109 sb_0__1_.mem_right_track_38.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_31_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_right_track_36.mux_l2_in_1__247 VGND VGND VPWR VPWR net247 sb_0__1_.mux_right_track_36.mux_l2_in_1__247/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA__184__A net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_40.mux_l1_in_0_ net61 net110 sb_0__1_.mem_right_track_40.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_38_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_14_0_prog_clk sb_0__1_.mem_right_track_14.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_14.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mux_right_track_4.mux_l1_in_1_ net109 net106 sb_0__1_.mem_right_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_67_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_52.mux_l2_in_0_ net255 sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_52.ccff_tail VGND VGND VPWR VPWR sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input21_A chanx_right_in[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_bottom_track_3.mux_l1_in_0_ net92 net78 sb_0__1_.mem_bottom_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mux_right_track_48.mux_l1_in_0__A0 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_13_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__A0 net72 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input69_A chany_top_in_0[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_4_0_prog_clk sb_0__1_.mem_right_track_44.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_46.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_78_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_4_2_0_prog_clk cby_0__1_.cby_0__1_.ccff_tail net98 VGND VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput204 net204 VGND VGND VPWR VPWR chany_top_out_0[4] sky130_fd_sc_hd__buf_12
Xoutput215 net215 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[1] sky130_fd_sc_hd__buf_12
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_13.out sky130_fd_sc_hd__clkbuf_1
XFILLER_82_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_2__A0 net58 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_185_ net42 VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_top_track_36.mux_l1_in_0_ net15 net118 sb_0__1_.mem_top_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_78_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_168_ net44 VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_2
Xsb_0__1_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_36.out sky130_fd_sc_hd__clkbuf_1
Xsb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_12_0_prog_clk sb_0__1_.mem_top_track_52.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_0.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_10.out sky130_fd_sc_hd__clkbuf_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input51_A chany_bottom_in[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_13_0_prog_clk sb_0__1_.mem_right_track_0.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_0.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_34_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_1__A0 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput104 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_ VGND VGND VPWR
+ VPWR net104 sky130_fd_sc_hd__buf_2
Xinput115 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_ VGND VGND VPWR
+ VPWR net115 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input99_A prog_reset_left_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1__A1 net49 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3_ net273 sb_0__1_.mux_bottom_track_53.out
+ cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_4.mux_l1_in_0_ net77 net83 sb_0__1_.mem_right_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_14_0_prog_clk sb_0__1_.mem_right_track_12.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_14.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_0__1_.mux_right_track_48.mux_l1_in_0__A1 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_8_0_prog_clk sb_0__1_.mem_top_track_4.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_4.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_input14_A chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__A1 net41 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_0__A0 net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_13_0_prog_clk sb_0__1_.mem_right_track_6.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_6.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mux_bottom_track_29.mux_l3_in_0_ sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_4_X
+ sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_3_X sb_0__1_.mem_bottom_track_29.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mux_right_track_14.mux_l1_in_0__A0 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input6_A chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput205 net205 VGND VGND VPWR VPWR chany_top_out_0[5] sky130_fd_sc_hd__buf_12
Xsb_0__1_.mux_right_track_8.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_8.out sky130_fd_sc_hd__clkbuf_1
XFILLER_57_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput216 net216 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[2] sky130_fd_sc_hd__buf_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4_ net64 net62 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mux_right_track_10.mux_l3_in_0_ sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X sb_0__1_.mem_right_track_10.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_67_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_52.mux_l1_in_0_ net52 net108 sb_0__1_.mem_right_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_23_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_bottom_track_5.mux_l1_in_2__A0 right_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input116_A top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input81_A chany_top_in_0[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_184_ net41 VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__clkbuf_2
XFILLER_89_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l4_in_0_ cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X cby_0__1_.cby_0__1_.mem_right_ipin_2.ccff_tail
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_64_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_8_0_prog_clk sb_0__1_.mem_top_track_20.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_20.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_49_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_bottom_track_29.mux_l2_in_1_ net279 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mem_bottom_track_29.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_56.mux_l2_in_0__257 VGND VGND VPWR VPWR net257 sb_0__1_.mux_right_track_56.mux_l2_in_0__257/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_93_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_12_0_prog_clk sb_0__1_.mem_top_track_52.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_52.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mux_right_track_10.mux_l2_in_1_ net233 net42 sb_0__1_.mem_right_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_6_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_167_ sb_0__1_.mux_bottom_track_1.out VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__clkbuf_1
XFILLER_69_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l3_in_1_ cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_bottom_track_29.mux_l1_in_2_ right_width_0_height_0_subtile_2__pin_inpad_0_
+ net28 sb_0__1_.mem_bottom_track_29.mem_out\[0\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input44_A chany_bottom_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_12_0_prog_clk sb_0__1_.mem_right_track_0.ccff_head
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_0.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_34_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_1__A1 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_top_track_20.mux_l2_in_1__264 VGND VGND VPWR VPWR net264 sb_0__1_.mux_top_track_20.mux_l2_in_1__264/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_42_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_29.out sky130_fd_sc_hd__clkbuf_1
Xclkbuf_4_4_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_4_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_57_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_40.mux_l2_in_0__250 VGND VGND VPWR VPWR net250 sb_0__1_.mux_right_track_40.mux_l2_in_0__250/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_31_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput105 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_ VGND VGND VPWR
+ VPWR net105 sky130_fd_sc_hd__buf_2
Xinput116 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_ VGND VGND VPWR
+ VPWR net116 sky130_fd_sc_hd__clkbuf_2
XFILLER_48_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_0__1_.mux_right_track_56.mux_l1_in_0__A1 net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_right_track_32.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_32.out sky130_fd_sc_hd__clkbuf_1
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2_ net56 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_9_0_prog_clk sb_0__1_.mem_top_track_4.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_4.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_0__A1 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_26.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_26.out sky130_fd_sc_hd__clkbuf_1
Xsb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_13_0_prog_clk sb_0__1_.mem_right_track_6.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_6.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3_ sb_0__1_.mux_bottom_track_29.out
+ net39 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xoutput206 net206 VGND VGND VPWR VPWR chany_top_out_0[6] sky130_fd_sc_hd__buf_12
Xoutput217 net217 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[3] sky130_fd_sc_hd__buf_12
XFILLER_4_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input109_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input74_A chany_top_in_0[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_183_ sb_0__1_.mux_top_track_28.out VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__clkbuf_1
Xsb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_8_0_prog_clk sb_0__1_.mem_top_track_20.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_20.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_49_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_bottom_track_29.mux_l2_in_0_ sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_bottom_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_38_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_right_track_18.mux_l2_in_1__237 VGND VGND VPWR VPWR net237 sb_0__1_.mux_right_track_18.mux_l2_in_1__237/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_87_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_top_track_2.mux_l3_in_0_ sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
+ sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X sb_0__1_.mem_top_track_2.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_95_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_3__A1 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_10.mux_l2_in_0_ sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_14_0_prog_clk sb_0__1_.mem_top_track_44.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_52.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
X_166_ sb_0__1_.mux_bottom_track_3.out VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__1_.mux_right_track_12.mux_l2_in_1__A1 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_22.mux_l3_in_0_ sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_1_X sb_0__1_.mem_right_track_22.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_68_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l3_in_0_ cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_bottom_track_29.mux_l1_in_1_ net10 net22 sb_0__1_.mem_bottom_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_2_0_prog_clk sb_0__1_.mem_right_track_32.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_32.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_input37_A chany_bottom_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_top_track_2.mux_l2_in_1_ net263 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mem_top_track_2.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mux_right_track_30.mux_l1_in_0__A0 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4__A0 net64 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_218_ net112 VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__clkbuf_2
XFILLER_51_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_149_ sb_0__1_.mux_bottom_track_37.out VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_2
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput117 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_ VGND VGND VPWR
+ VPWR net117 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput106 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_ VGND VGND VPWR
+ VPWR net106 sky130_fd_sc_hd__buf_2
XFILLER_56_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_right_track_10.mux_l1_in_1_ net109 net106 sb_0__1_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mux_right_track_22.mux_l1_in_0__A1 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_22.mux_l2_in_1_ net240 net34 sb_0__1_.mem_right_track_22.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_46_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_1_ cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mux_top_track_2.mux_l1_in_2_ net62 net48 sb_0__1_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_88_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_11_0_prog_clk sb_0__1_.mem_top_track_2.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_4.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_67_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mux_right_track_54.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_54.out sky130_fd_sc_hd__clkbuf_1
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_top_track_4.mux_l2_in_1__267 VGND VGND VPWR VPWR net267 sb_0__1_.mux_top_track_4.mux_l2_in_1__267/LO
+ sky130_fd_sc_hd__conb_1
Xsb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_13_0_prog_clk sb_0__1_.mem_right_track_4.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_6.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_0__A0 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2_ net77 net46 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xoutput207 net207 VGND VGND VPWR VPWR chany_top_out_0[7] sky130_fd_sc_hd__buf_12
Xoutput218 net218 VGND VGND VPWR VPWR prog_reset_bottom_out sky130_fd_sc_hd__buf_12
XFILLER_4_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_20.mux_l3_in_0_ sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_4_X
+ sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_3_X sb_0__1_.mem_top_track_20.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_48_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_right_track_48.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_48.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_182_ net39 VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input67_A chany_top_in_0[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_77 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_8_0_prog_clk sb_0__1_.mem_top_track_12.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_20.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_49_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_right_track_20.mux_l2_in_1__A1 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_165_ sb_0__1_.mux_bottom_track_5.out VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_1
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_top_track_20.mux_l2_in_1_ net264 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mem_top_track_20.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_bottom_track_29.mux_l1_in_0_ net74 net69 sb_0__1_.mem_bottom_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_2_0_prog_clk sb_0__1_.mem_right_track_30.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_32.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_2.mux_l2_in_0_ sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mux_right_track_30.mux_l1_in_0__A1 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4__A1 net62 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_217_ net112 VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_1
X_148_ net65 VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__clkbuf_2
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_0__A0 net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput118 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_ VGND VGND VPWR
+ VPWR net118 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput107 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_ VGND VGND VPWR
+ VPWR net107 sky130_fd_sc_hd__buf_2
XFILLER_56_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_10.mux_l1_in_0_ net72 net79 sb_0__1_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_top_track_20.mux_l1_in_2_ net55 net41 sb_0__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_4_0_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[2\] net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mux_right_track_22.mux_l2_in_0_ net109 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_22.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_0_ cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_0_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_2.mux_l1_in_1_ net28 net10 sb_0__1_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mux_top_track_4.mux_l1_in_2__A0 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input97_A isol_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_right_track_16.mux_l2_in_0__A0 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_1_0_prog_clk sb_0__1_.mem_right_track_38.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_38.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input12_A chanx_right_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1_ sb_0__1_.mux_bottom_track_11.out
+ net49 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xoutput208 net208 VGND VGND VPWR VPWR chany_top_out_0[8] sky130_fd_sc_hd__buf_12
Xoutput219 net219 VGND VGND VPWR VPWR prog_reset_right_out sky130_fd_sc_hd__buf_12
XFILLER_4_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input4_A chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_181_ net38 VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__clkbuf_2
XFILLER_89_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_7_0_prog_clk sb_0__1_.mem_bottom_track_21.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_21.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_63_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input114_A test_enable_top_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_164_ sb_0__1_.mux_bottom_track_7.out VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_2
Xsb_0__1_.mux_top_track_20.mux_l2_in_0_ sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_top_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_41_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_4.out sky130_fd_sc_hd__clkbuf_1
XFILLER_45_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_5_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_11_0_prog_clk sb_0__1_.mem_bottom_track_53.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__dfrtp_2
XFILLER_83_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mux_right_track_4.mux_l2_in_1__A1 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_216_ net112 VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__clkbuf_1
X_147_ net64 VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__clkbuf_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput108 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_ VGND VGND VPWR
+ VPWR net108 sky130_fd_sc_hd__buf_2
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_top_track_20.mux_l1_in_1_ net3 net5 sb_0__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_1_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[1\] net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input42_A chany_bottom_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mux_top_track_52.mux_l2_in_1__269 VGND VGND VPWR VPWR net269 sb_0__1_.mux_top_track_52.mux_l2_in_1__269/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_3__A1 right_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput90 chany_top_in_0[7] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_2
Xsb_0__1_.mux_top_track_2.mux_l1_in_0_ net22 net116 sb_0__1_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mux_top_track_4.mux_l1_in_2__A1 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_4.mux_l2_in_1__249 VGND VGND VPWR VPWR net249 sb_0__1_.mux_right_track_4.mux_l2_in_1__249/LO
+ sky130_fd_sc_hd__conb_1
Xclkbuf_4_3_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_3_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_16_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_38.mux_l2_in_0__248 VGND VGND VPWR VPWR net248 sb_0__1_.mux_right_track_38.mux_l2_in_0__248/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_29_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_1_0_prog_clk sb_0__1_.mem_right_track_36.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_38.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mux_right_track_0.mux_l3_in_0_ sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X sb_0__1_.mem_right_track_0.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_41_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_22.mux_l1_in_0_ net63 net64 sb_0__1_.mem_right_track_22.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0_ sb_0__1_.mux_bottom_track_5.out
+ net52 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xoutput209 net209 VGND VGND VPWR VPWR chany_top_out_0[9] sky130_fd_sc_hd__buf_12
XFILLER_68_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_34.mux_l2_in_0_ sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_34.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_180_ net37 VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__clkbuf_2
XFILLER_22_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_5_0_prog_clk sb_0__1_.mem_right_track_50.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_50.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_64_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_right_track_0.mux_l2_in_1_ net232 net51 sb_0__1_.mem_right_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mux_bottom_track_29.mux_l1_in_2__A0 right_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_7_0_prog_clk sb_0__1_.mem_bottom_track_21.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_21.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_95_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mux_top_track_28.mux_l2_in_1__A1 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input107_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input72_A chany_top_in_0[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_34.mux_l1_in_1_ net246 net55 sb_0__1_.mem_right_track_34.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_40_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_163_ net81 VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__clkbuf_2
XFILLER_77_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_right_track_24.mux_l1_in_1__A1 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_12_0_prog_clk sb_0__1_.mem_bottom_track_45.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_53.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_68_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__212__A net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_215_ net112 VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__clkbuf_2
X_146_ net92 VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__clkbuf_2
XFILLER_76_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput109 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_ VGND VGND VPWR
+ VPWR net109 sky130_fd_sc_hd__buf_2
XANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_1__A0 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__207__A net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_top_track_20.mux_l1_in_0_ net17 net116 sb_0__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_10.out sky130_fd_sc_hd__clkbuf_1
XFILLER_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_1_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[0\] net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input35_A chany_bottom_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_129_ sb_0__1_.mux_right_track_16.out VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_2
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput91 chany_top_in_0[8] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_1
Xinput80 chany_top_in_0[25] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_2.mux_l2_in_1__263 VGND VGND VPWR VPWR net263 sb_0__1_.mux_top_track_2.mux_l2_in_1__263/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_7_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_top_track_36.mux_l2_in_1__A1 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_8_0_prog_clk sb_0__1_.mem_top_track_12.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_12.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_58_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__215__A net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_5_0_prog_clk sb_0__1_.mem_right_track_48.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_50.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_0__1_.mux_right_track_32.mux_l1_in_1__A1 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_right_track_0.mux_l2_in_0_ sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_7_0_prog_clk sb_0__1_.mem_bottom_track_13.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_21.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_48_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_11_0_prog_clk sb_0__1_.mem_top_track_44.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_44.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mux_bottom_track_13.mux_l3_in_0_ sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_4_X
+ sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_3_X sb_0__1_.mem_bottom_track_13.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_86_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_162_ sb_0__1_.mux_bottom_track_11.out VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input65_A chany_top_in_0[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_34.mux_l1_in_0_ net107 net85 sb_0__1_.mem_right_track_34.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_46.mux_l2_in_0_ net252 sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_46.ccff_tail VGND VGND VPWR VPWR sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xinput1 ccff_head VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_51_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_prog_clk prog_clk VGND VGND VPWR VPWR clknet_0_prog_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_86_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_0.mux_l1_in_1_ net110 net107 sb_0__1_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_27_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_214_ net101 VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__clkbuf_2
XFILLER_51_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_145_ sb_0__1_.mux_bottom_track_45.out VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__clkbuf_2
Xsb_0__1_.mux_bottom_track_13.mux_l2_in_1_ net277 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mem_bottom_track_13.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_4_0_prog_clk sb_0__1_.mem_right_track_56.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_1.ccff_head sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XFILLER_72_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_1__A1 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_ cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_21_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_0_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_0.ccff_tail net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xoutput190 net190 VGND VGND VPWR VPWR chany_top_out_0[19] sky130_fd_sc_hd__buf_12
XANTENNA_sb_0__1_.mux_top_track_10.mux_l1_in_2__A0 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input28_A chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3__A0 net71 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_128_ sb_0__1_.mux_right_track_18.out VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_2
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput70 chany_top_in_0[16] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_1
Xinput92 chany_top_in_0[9] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__buf_2
Xinput81 chany_top_in_0[26] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__buf_2
XFILLER_29_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__218__A net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_right_track_28.mux_l1_in_0__A0 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_4_1_0_prog_clk cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.ccff_tail
+ net98 VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__dfrtp_2
Xsb_0__1_.mux_bottom_track_13.mux_l1_in_2_ right_width_0_height_0_subtile_0__pin_inpad_0_
+ net26 sb_0__1_.mem_bottom_track_13.mem_out\[0\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xleft_tile_225 VGND VGND VPWR VPWR left_tile_225/HI chanx_right_out[0] sky130_fd_sc_hd__conb_1
XFILLER_93_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input95_A gfpga_pad_io_soc_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_44.mux_l2_in_0_ sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_top_track_44.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_9_0_prog_clk sb_0__1_.mem_top_track_12.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_12.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_14_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input10_A chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_10_0_prog_clk sb_0__1_.mem_top_track_36.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_44.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_63_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_bottom_track_37.mux_l2_in_1__A1 right_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input2_A ccff_head_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_54.mux_l2_in_0__256 VGND VGND VPWR VPWR net256 sb_0__1_.mux_right_track_54.mux_l2_in_0__256/LO
+ sky130_fd_sc_hd__conb_1
Xsb_0__1_.mux_top_track_10.mux_l1_in_3__261 VGND VGND VPWR VPWR net261 sb_0__1_.mux_top_track_10.mux_l1_in_3__261/LO
+ sky130_fd_sc_hd__conb_1
X_161_ sb_0__1_.mux_bottom_track_13.out VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__clkbuf_2
Xsb_0__1_.mux_top_track_44.mux_l1_in_1_ net268 net37 sb_0__1_.mem_top_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_input58_A chany_bottom_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_3_0_prog_clk sb_0__1_.mem_right_track_24.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_24.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_3__A1 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput2 ccff_head_0 VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_3_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_right_track_18.mux_l2_in_1__A1 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_0.mux_l1_in_0_ net104 net81 sb_0__1_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_42_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input112_A test_enable_bottom_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1__A1 net51 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_213_ net101 VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_1
X_144_ net90 VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_2
Xsb_0__1_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_4.out sky130_fd_sc_hd__clkbuf_1
Xsb_0__1_.mux_bottom_track_13.mux_l2_in_0_ sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_bottom_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_76_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_4_0_prog_clk sb_0__1_.mem_right_track_54.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_56.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_33_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_2__S sb_0__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_0__1_.mux_right_track_36.mux_l1_in_0__A0 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__1_.mux_top_track_52.mux_l2_in_1__A1 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput191 net191 VGND VGND VPWR VPWR chany_top_out_0[1] sky130_fd_sc_hd__buf_12
Xoutput180 net180 VGND VGND VPWR VPWR chany_top_out_0[0] sky130_fd_sc_hd__buf_12
XFILLER_21_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_right_track_46.mux_l1_in_0_ net45 net105 sb_0__1_.mem_right_track_46.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mux_bottom_track_13.mux_l1_in_0__A0 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_127_ sb_0__1_.mux_right_track_20.out VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput71 chany_top_in_0[17] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__buf_2
Xinput82 chany_top_in_0[27] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput93 gfpga_pad_io_soc_in[0] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_1
Xinput60 chany_bottom_in[7] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_2
XFILLER_83_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_bottom_track_13.mux_l1_in_1_ net8 net20 sb_0__1_.mem_bottom_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_52_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_right_track_28.mux_l1_in_0__A1 net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input40_A chany_bottom_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__144__A net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_0__1_.mux_bottom_track_11.mux_l1_in_2__A0 right_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input88_A chany_top_in_0[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_3_0_prog_clk sb_0__1_.mem_bottom_track_1.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_4_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_8_0_prog_clk sb_0__1_.mem_top_track_10.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_12.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3_ net274 net86 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__139__A net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_2_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_2_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_31_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_82 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_16.mux_l2_in_1__236 VGND VGND VPWR VPWR net236 sb_0__1_.mux_right_track_16.mux_l2_in_1__236/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_0__1_.mux_top_track_20.mux_l1_in_0__A1 net116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_13_0_prog_clk sb_0__1_.mem_bottom_track_45.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_45.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_39_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_160_ net78 VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_2
XFILLER_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_top_track_44.mux_l1_in_0_ net31 net13 sb_0__1_.mem_top_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4_ net92 net61 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_3_0_prog_clk sb_0__1_.mem_right_track_22.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_24.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_45_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_22.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_22.out sky130_fd_sc_hd__clkbuf_1
XANTENNA__152__A net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput3 chanx_right_in[0] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input105_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_212_ net101 VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_0__1_.mux_bottom_track_21.mux_l1_in_0__A0 net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l4_in_0_ cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X cby_0__1_.cby_0__1_.ccff_tail
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input70_A chany_top_in_0[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_143_ net89 VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_2
XFILLER_76_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__147__A net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_right_track_36.mux_l1_in_0__A1 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput192 net192 VGND VGND VPWR VPWR chany_top_out_0[20] sky130_fd_sc_hd__buf_12
Xoutput181 net181 VGND VGND VPWR VPWR chany_top_out_0[10] sky130_fd_sc_hd__buf_12
Xclkbuf_4_15_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_15_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
Xsb_0__1_.mux_right_track_16.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_16.out sky130_fd_sc_hd__clkbuf_1
Xoutput170 net170 VGND VGND VPWR VPWR chany_bottom_out[28] sky130_fd_sc_hd__buf_12
XFILLER_62_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_0__1_.mux_bottom_track_13.mux_l1_in_0__A1 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_126_ sb_0__1_.mux_right_track_22.out VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput72 chany_top_in_0[18] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__buf_2
Xinput61 chany_bottom_in[8] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput50 chany_bottom_in[25] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput83 chany_top_in_0[28] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput94 gfpga_pad_io_soc_in[1] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l3_in_1_ cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_bottom_track_13.mux_l1_in_0_ net86 net72 sb_0__1_.mem_bottom_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_20_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input33_A chany_bottom_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_109_ sb_0__1_.mux_right_track_56.out VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_1
XANTENNA__160__A net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_37.mux_l3_in_0_ sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_2_X sb_0__1_.mem_bottom_track_37.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_69_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_53.out sky130_fd_sc_hd__clkbuf_2
XFILLER_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_3_0_prog_clk sb_0__1_.mem_bottom_track_1.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_1.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_43_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_16.mux_l3_in_0_ sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X sb_0__1_.mem_right_track_16.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2_ net55 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__155__A net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_7_0_prog_clk sb_0__1_.mem_bottom_track_13.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_13.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_right_track_52.mux_l1_in_0__A0 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_bottom_track_37.mux_l2_in_1_ net227 right_width_0_height_0_subtile_3__pin_inpad_0_
+ sb_0__1_.mem_bottom_track_37.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_13_0_prog_clk sb_0__1_.mem_bottom_track_45.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_45.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mux_right_track_16.mux_l2_in_1_ net236 net38 sb_0__1_.mem_right_track_16.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_10_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mux_right_track_50.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_50.out sky130_fd_sc_hd__clkbuf_1
XFILLER_49_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3_ net69 net38 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4__A0 net92 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_7_0_prog_clk sb_0__1_.mem_bottom_track_7.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_11.ccff_head sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_0__1_.mux_right_track_44.mux_l1_in_0__A1 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput4 chanx_right_in[10] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_0__1_.mux_bottom_track_3.mux_l1_in_0__A0 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_right_track_10.mux_l1_in_0__A0 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mux_bottom_track_21.mux_l1_in_0__A1 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_211_ net101 VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__clkbuf_1
X_142_ net88 VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input63_A chany_top_in_0[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__163__A net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__273 VGND VGND VPWR VPWR net273
+ cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__273/LO sky130_fd_sc_hd__conb_1
XFILLER_71_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_44.out sky130_fd_sc_hd__clkbuf_1
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput182 net182 VGND VGND VPWR VPWR chany_top_out_0[11] sky130_fd_sc_hd__buf_12
Xoutput193 net193 VGND VGND VPWR VPWR chany_top_out_0[21] sky130_fd_sc_hd__buf_12
Xoutput160 net160 VGND VGND VPWR VPWR chany_bottom_out[19] sky130_fd_sc_hd__buf_12
Xoutput171 net171 VGND VGND VPWR VPWR chany_bottom_out[29] sky130_fd_sc_hd__buf_12
XFILLER_46_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_2__A0 right_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_125_ sb_0__1_.mux_right_track_24.out VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_2
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_bottom_track_37.mux_l2_in_1__227 VGND VGND VPWR VPWR net227 sb_0__1_.mux_bottom_track_37.mux_l2_in_1__227/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_38_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__158__A net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput73 chany_top_in_0[19] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_2
Xinput84 chany_top_in_0[29] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_1
Xinput95 gfpga_pad_io_soc_in[2] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_1
Xinput51 chany_bottom_in[26] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__buf_2
Xinput62 chany_bottom_in[9] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_2
Xinput40 chany_bottom_in[16] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l3_in_0_ cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input26_A chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_14_0_prog_clk sb_0__1_.mem_right_track_10.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_10.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mux_right_track_38.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_38.out sky130_fd_sc_hd__clkbuf_1
XFILLER_7_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_20.mux_l2_in_1__239 VGND VGND VPWR VPWR net239 sb_0__1_.mux_right_track_20.mux_l2_in_1__239/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_4_0_prog_clk sb_0__1_.mem_bottom_track_1.ccff_head
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_1.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_68_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_1_ cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_7_0_prog_clk sb_0__1_.mem_bottom_track_13.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_13.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_22_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_10_0_prog_clk sb_0__1_.mem_top_track_36.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_36.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_57_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input93_A gfpga_pad_io_soc_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_right_track_52.mux_l1_in_0__A1 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net95 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR right_width_0_height_0_subtile_1__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_63_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_bottom_track_37.mux_l2_in_0_ sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_bottom_track_37.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_5_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_12_0_prog_clk sb_0__1_.mem_bottom_track_37.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_45.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_54_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_right_track_16.mux_l2_in_0_ net106 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_16.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_24_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_0_prog_clk_A prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2_ net76 net45 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_6_0_prog_clk sb_0__1_.mem_bottom_track_7.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_7.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xinput5 chanx_right_in[11] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
Xsb_0__1_.mux_top_track_6.mux_l1_in_3__270 VGND VGND VPWR VPWR net270 sb_0__1_.mux_top_track_6.mux_l1_in_3__270/LO
+ sky130_fd_sc_hd__conb_1
Xsb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_5.out sky130_fd_sc_hd__clkbuf_1
XFILLER_51_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_bottom_track_3.mux_l1_in_0__A1 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_210_ net98 VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__clkbuf_1
Xsb_0__1_.mux_top_track_28.mux_l2_in_1__265 VGND VGND VPWR VPWR net265 sb_0__1_.mux_top_track_28.mux_l2_in_1__265/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_141_ sb_0__1_.mux_bottom_track_53.out VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__clkbuf_2
Xsb_0__1_.mux_bottom_track_37.mux_l1_in_1_ net29 net11 sb_0__1_.mem_bottom_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_input56_A chany_bottom_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__A1 net86 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput161 net161 VGND VGND VPWR VPWR chany_bottom_out[1] sky130_fd_sc_hd__buf_12
Xoutput150 net150 VGND VGND VPWR VPWR chany_bottom_out[0] sky130_fd_sc_hd__buf_12
XFILLER_21_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput194 net194 VGND VGND VPWR VPWR chany_top_out_0[22] sky130_fd_sc_hd__buf_12
Xoutput183 net183 VGND VGND VPWR VPWR chany_top_out_0[12] sky130_fd_sc_hd__buf_12
Xoutput172 net172 VGND VGND VPWR VPWR chany_bottom_out[2] sky130_fd_sc_hd__buf_12
XANTENNA_input110_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_0__1_.mux_bottom_track_1.mux_l1_in_2__A1 right_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_124_ sb_0__1_.mux_right_track_26.out VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__174__A net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput74 chany_top_in_0[1] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_2
Xinput63 chany_top_in_0[0] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_1
Xinput85 chany_top_in_0[2] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_2
Xinput96 gfpga_pad_io_soc_in[3] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_1
Xinput30 chanx_right_in[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_ cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_
+ sky130_fd_sc_hd__clkbuf_1
Xinput41 chany_bottom_in[17] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__buf_2
Xinput52 chany_bottom_in[27] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input19_A chanx_right_in[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_0.out sky130_fd_sc_hd__clkbuf_1
Xsb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk sb_0__1_.mem_right_track_10.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_10.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_73_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__169__A net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_0_ cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_1_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_6_0_prog_clk sb_0__1_.mem_bottom_track_11.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_13.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_10_0_prog_clk sb_0__1_.mem_top_track_36.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_36.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input86_A chany_top_in_0[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__182__A net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_11_0_prog_clk sb_0__1_.mem_right_track_16.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_16.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_5_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1_ sb_0__1_.mux_bottom_track_7.out
+ net51 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_1_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_1_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
Xsb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_7_0_prog_clk sb_0__1_.mem_bottom_track_5.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_7.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__177__A net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput6 chanx_right_in[12] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_5_0_prog_clk sb_0__1_.mem_right_track_48.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_48.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_bottom_track_37.mux_l1_in_0_ net23 net68 sb_0__1_.mem_bottom_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
X_140_ net86 VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__clkbuf_2
XFILLER_2_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input49_A chany_bottom_in[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_0__A0 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
Xsb_0__1_.mux_right_track_16.mux_l1_in_0_ net66 net68 sb_0__1_.mem_right_track_16.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_44_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput195 net195 VGND VGND VPWR VPWR chany_top_out_0[23] sky130_fd_sc_hd__buf_12
Xoutput184 net184 VGND VGND VPWR VPWR chany_top_out_0[13] sky130_fd_sc_hd__buf_12
Xoutput140 net140 VGND VGND VPWR VPWR chanx_right_out[28] sky130_fd_sc_hd__buf_12
Xoutput162 net162 VGND VGND VPWR VPWR chany_bottom_out[20] sky130_fd_sc_hd__buf_12
Xoutput173 net173 VGND VGND VPWR VPWR chany_bottom_out[3] sky130_fd_sc_hd__buf_12
Xoutput151 net151 VGND VGND VPWR VPWR chany_bottom_out[10] sky130_fd_sc_hd__buf_12
Xsb_0__1_.mux_right_track_28.mux_l2_in_0_ sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_28.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_input103_A reset_top_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0__A1 net52 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_123_ sb_0__1_.mux_right_track_28.out VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_6_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput20 chanx_right_in[25] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_1
Xinput31 chanx_right_in[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_1
Xsb_0__1_.mux_right_track_30.mux_l2_in_0_ sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_30.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_21_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput64 chany_top_in_0[10] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__buf_2
Xinput75 chany_top_in_0[20] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_1
Xinput86 chany_top_in_0[3] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__buf_2
XANTENNA__190__A net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput97 isol_n VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_2
Xinput42 chany_bottom_in[18] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_2
Xinput53 chany_bottom_in[28] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_2.mux_l2_in_1__238 VGND VGND VPWR VPWR net238 sb_0__1_.mux_right_track_2.mux_l2_in_1__238/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_32_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_11_0_prog_clk sb_0__1_.mem_top_track_0.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_15_0_prog_clk sb_0__1_.mem_right_track_10.ccff_head
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_10.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_43_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2__A1 net48 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mux_bottom_track_5.mux_l3_in_0_ sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X
+ sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X sb_0__1_.mem_bottom_track_5.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_93_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__185__A net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_14_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_14_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
Xsb_0__1_.mux_right_track_28.mux_l1_in_1_ net243 net59 sb_0__1_.mem_right_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_69_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_15_0_prog_clk sb_0__1_.mem_right_track_2.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input31_A chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_30.mux_l1_in_1_ net244 net58 sb_0__1_.mem_right_track_30.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_84_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_10_0_prog_clk sb_0__1_.mem_top_track_28.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_36.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_57_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_bottom_track_5.mux_l2_in_1_ net229 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mem_bottom_track_5.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input79_A chany_top_in_0[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_14_0_prog_clk sb_0__1_.mem_right_track_16.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_16.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_74_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_0_ sb_0__1_.mux_bottom_track_1.out
+ net54 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_2__A0 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput7 chanx_right_in[13] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__193__A net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mux_right_track_12.mux_l2_in_0__A0 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_5_0_prog_clk sb_0__1_.mem_right_track_46.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_48.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_74_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_bottom_track_5.mux_l1_in_2_ right_width_0_height_0_subtile_2__pin_inpad_0_
+ net3 sb_0__1_.mem_bottom_track_5.mem_out\[0\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XFILLER_76_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_48.mux_l2_in_0__253 VGND VGND VPWR VPWR net253 sb_0__1_.mux_right_track_48.mux_l2_in_0__253/LO
+ sky130_fd_sc_hd__conb_1
X_199_ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__clkbuf_1
XANTENNA__188__A net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput196 net196 VGND VGND VPWR VPWR chany_top_out_0[24] sky130_fd_sc_hd__buf_12
Xoutput185 net185 VGND VGND VPWR VPWR chany_top_out_0[14] sky130_fd_sc_hd__buf_12
Xoutput141 net141 VGND VGND VPWR VPWR chanx_right_out[29] sky130_fd_sc_hd__buf_12
Xoutput163 net163 VGND VGND VPWR VPWR chany_bottom_out[21] sky130_fd_sc_hd__buf_12
Xoutput152 net152 VGND VGND VPWR VPWR chany_bottom_out[11] sky130_fd_sc_hd__buf_12
Xoutput174 net174 VGND VGND VPWR VPWR chany_bottom_out[4] sky130_fd_sc_hd__buf_12
Xoutput130 net130 VGND VGND VPWR VPWR chanx_right_out[19] sky130_fd_sc_hd__buf_12
XFILLER_55_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input61_A chany_bottom_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_122_ sb_0__1_.mux_right_track_30.out VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_2
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput21 chanx_right_in[26] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput10 chanx_right_in[16] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_1
Xinput32 chanx_right_in[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput43 chany_bottom_in[19] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__buf_2
Xinput54 chany_bottom_in[29] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput76 chany_top_in_0[21] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_2
Xinput65 chany_top_in_0[11] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_2
Xinput87 chany_top_in_0[4] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_1
Xinput98 prog_reset_bottom_in VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_16
XANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_0.mux_l2_in_1__232 VGND VGND VPWR VPWR net232 sb_0__1_.mux_right_track_0.mux_l2_in_1__232/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_43_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_10_0_prog_clk sb_0__1_.mem_top_track_0.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_0.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mux_right_track_6.mux_l3_in_0_ sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X
+ sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X sb_0__1_.mem_right_track_6.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_right_track_28.mux_l1_in_0_ net104 net89 sb_0__1_.mem_right_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_34_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk sb_0__1_.mem_right_track_2.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_2.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_84_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_30.mux_l1_in_0_ net105 net88 sb_0__1_.mem_right_track_30.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_84_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input24_A chanx_right_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_right_track_0.mux_l2_in_1__A1 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_bottom_track_21.mux_l2_in_1__278 VGND VGND VPWR VPWR net278 sb_0__1_.mux_bottom_track_21.mux_l2_in_1__278/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_90_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_top_track_2.mux_l1_in_0__A1 net116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_6.mux_l2_in_1_ net258 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mem_right_track_6.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_54_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_9_0_prog_clk sb_0__1_.mem_bottom_track_37.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_37.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mux_bottom_track_5.mux_l2_in_0_ sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_bottom_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_79_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mux_right_track_20.mux_l2_in_0__A0 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_14_0_prog_clk sb_0__1_.mem_right_track_14.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_16.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_10_0_prog_clk sb_0__1_.mem_top_track_6.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_10.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_39_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_52.mux_l2_in_0__255 VGND VGND VPWR VPWR net255 sb_0__1_.mux_right_track_52.mux_l2_in_0__255/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_49_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input91_A chany_top_in_0[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_15_0_prog_clk sb_0__1_.mem_right_track_8.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_10.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_60_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput8 chanx_right_in[14] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
XFILLER_91_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_6.mux_l1_in_2_ net46 net110 sb_0__1_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_bottom_track_5.mux_l1_in_1_ net5 net17 sb_0__1_.mem_bottom_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_19_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_198_ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__clkbuf_2
XFILLER_56_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput197 net197 VGND VGND VPWR VPWR chany_top_out_0[25] sky130_fd_sc_hd__buf_12
Xoutput186 net186 VGND VGND VPWR VPWR chany_top_out_0[15] sky130_fd_sc_hd__buf_12
Xoutput120 net120 VGND VGND VPWR VPWR ccff_tail_0 sky130_fd_sc_hd__buf_12
Xoutput131 net131 VGND VGND VPWR VPWR chanx_right_out[1] sky130_fd_sc_hd__buf_12
Xoutput164 net164 VGND VGND VPWR VPWR chany_bottom_out[22] sky130_fd_sc_hd__buf_12
Xoutput175 net175 VGND VGND VPWR VPWR chany_bottom_out[5] sky130_fd_sc_hd__buf_12
Xoutput153 net153 VGND VGND VPWR VPWR chany_bottom_out[12] sky130_fd_sc_hd__buf_12
Xoutput142 net142 VGND VGND VPWR VPWR chanx_right_out[2] sky130_fd_sc_hd__buf_12
XFILLER_70_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_121_ sb_0__1_.mux_right_track_32.out VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input54_A chany_bottom_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_76 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput77 chany_top_in_0[22] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__buf_2
Xinput66 chany_top_in_0[12] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_1
Xinput88 chany_top_in_0[5] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__buf_2
Xinput22 chanx_right_in[27] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput11 chanx_right_in[17] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_1
Xinput33 chany_bottom_in[0] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_1
Xinput44 chany_bottom_in[1] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_2
Xinput55 chany_bottom_in[2] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__buf_2
Xinput99 prog_reset_left_in VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_top_track_52.mux_l3_in_0_ sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_1_X sb_0__1_.mem_right_track_0.ccff_head
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2__A0 net56 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_10_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_10_0_prog_clk net1
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_0.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_7_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_13_0_prog_clk sb_0__1_.mem_right_track_0.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_2.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_27_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input17_A chanx_right_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_0.out sky130_fd_sc_hd__clkbuf_1
XFILLER_17_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_top_track_52.mux_l2_in_1_ net269 net35 sb_0__1_.mem_top_track_52.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_89_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input9_A chanx_right_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_6.mux_l2_in_0_ sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_57_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_12_0_prog_clk sb_0__1_.mem_bottom_track_37.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_37.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_95_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_right_track_4.mux_l1_in_1__A0 net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_14.mux_l2_in_1__235 VGND VGND VPWR VPWR net235 sb_0__1_.mux_right_track_14.mux_l2_in_1__235/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_48_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_8_0_prog_clk sb_0__1_.mem_top_track_6.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_6.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_94_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_bottom_track_21.mux_l3_in_0_ sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_4_X
+ sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_3_X sb_0__1_.mem_bottom_track_21.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_40_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input84_A chany_top_in_0[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk sb_0__1_.mem_right_track_8.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_8.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput9 chanx_right_in[15] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_right_track_54.mux_l2_in_0_ net256 sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_54.ccff_tail VGND VGND VPWR VPWR sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_right_track_6.mux_l1_in_1_ net107 net104 sb_0__1_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_right_track_34.mux_l1_in_1__246 VGND VGND VPWR VPWR net246 sb_0__1_.mux_right_track_34.mux_l1_in_1__246/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_82_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_bottom_track_5.mux_l1_in_0_ net90 net77 sb_0__1_.mem_bottom_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_15_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_5 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_21.out sky130_fd_sc_hd__clkbuf_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3__A1 net39 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_197_ sb_0__1_.mux_top_track_0.out VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__clkbuf_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_bottom_track_21.mux_l2_in_1_ net278 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mem_bottom_track_21.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_64_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__271 VGND VGND VPWR VPWR net271
+ cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__271/LO sky130_fd_sc_hd__conb_1
XFILLER_2_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput143 net143 VGND VGND VPWR VPWR chanx_right_out[3] sky130_fd_sc_hd__buf_12
Xoutput121 net121 VGND VGND VPWR VPWR chanx_right_out[10] sky130_fd_sc_hd__buf_12
Xoutput132 net132 VGND VGND VPWR VPWR chanx_right_out[20] sky130_fd_sc_hd__buf_12
Xclkbuf_4_0_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_0_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
Xoutput198 net198 VGND VGND VPWR VPWR chany_top_out_0[26] sky130_fd_sc_hd__buf_12
Xoutput187 net187 VGND VGND VPWR VPWR chany_top_out_0[16] sky130_fd_sc_hd__buf_12
Xoutput165 net165 VGND VGND VPWR VPWR chany_bottom_out[23] sky130_fd_sc_hd__buf_12
Xoutput154 net154 VGND VGND VPWR VPWR chany_bottom_out[13] sky130_fd_sc_hd__buf_12
Xoutput176 net176 VGND VGND VPWR VPWR chany_bottom_out[6] sky130_fd_sc_hd__buf_12
XFILLER_55_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_120_ sb_0__1_.mux_right_track_34.out VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_2
XFILLER_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input47_A chany_bottom_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput67 chany_top_in_0[13] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_2
Xinput89 chany_top_in_0[6] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_2
Xinput78 chany_top_in_0[23] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__buf_2
Xinput23 chanx_right_in[28] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_1
Xinput12 chanx_right_in[18] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
Xinput34 chany_bottom_in[10] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__buf_2
Xinput56 chany_bottom_in[3] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__buf_2
Xinput45 chany_bottom_in[20] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dlymetal6s2s_1
Xsb_0__1_.mux_top_track_12.mux_l2_in_1__262 VGND VGND VPWR VPWR net262 sb_0__1_.mux_top_track_12.mux_l2_in_1__262/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_0__1_.mux_bottom_track_7.mux_l1_in_2__A0 right_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_44.out sky130_fd_sc_hd__clkbuf_1
XFILLER_57_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_21.mux_l1_in_2_ right_width_0_height_0_subtile_1__pin_inpad_0_
+ net27 sb_0__1_.mem_bottom_track_21.mem_out\[0\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input101_A reset_bottom_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_3_0_prog_clk sb_0__1_.mem_right_track_34.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_34.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_top_track_28.mux_l1_in_1__A0 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_8_0_prog_clk sb_0__1_.mem_top_track_28.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_28.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_16_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mux_top_track_52.mux_l2_in_0_ net30 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_top_track_52.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_12.out sky130_fd_sc_hd__clkbuf_1
XFILLER_70_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_12_0_prog_clk sb_0__1_.mem_bottom_track_29.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_37.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_13_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_13_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_13_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_sb_0__1_.mux_right_track_4.mux_l1_in_1__A1 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_10_0_prog_clk sb_0__1_.mem_top_track_4.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_6.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_94_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_13_0_prog_clk sb_0__1_.mem_right_track_6.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_8.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_65_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input77_A chany_top_in_0[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_right_track_24.mux_l1_in_0__A0 net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_4_2_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[2\] net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mux_right_track_6.mux_l1_in_0_ net76 net82 sb_0__1_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_196_ sb_0__1_.mux_top_track_2.out VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__clkbuf_1
XFILLER_41_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_21.mux_l2_in_0_ sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_bottom_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_64_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mux_right_track_16.mux_l1_in_0__A1 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput166 net166 VGND VGND VPWR VPWR chany_bottom_out[24] sky130_fd_sc_hd__buf_12
Xoutput155 net155 VGND VGND VPWR VPWR chany_bottom_out[14] sky130_fd_sc_hd__buf_12
Xoutput177 net177 VGND VGND VPWR VPWR chany_bottom_out[7] sky130_fd_sc_hd__buf_12
Xoutput144 net144 VGND VGND VPWR VPWR chanx_right_out[4] sky130_fd_sc_hd__buf_12
Xoutput122 net122 VGND VGND VPWR VPWR chanx_right_out[11] sky130_fd_sc_hd__buf_12
Xoutput133 net133 VGND VGND VPWR VPWR chanx_right_out[21] sky130_fd_sc_hd__buf_12
Xoutput188 net188 VGND VGND VPWR VPWR chany_top_out_0[17] sky130_fd_sc_hd__buf_12
Xoutput199 net199 VGND VGND VPWR VPWR chany_top_out_0[27] sky130_fd_sc_hd__buf_12
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_12.mux_l3_in_0_ sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X sb_0__1_.mem_right_track_12.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_61_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_54.mux_l1_in_0_ net53 net109 sb_0__1_.mem_right_track_54.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xinput13 chanx_right_in[19] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput79 chany_top_in_0[24] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_1
Xinput68 chany_top_in_0[14] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_2
X_179_ sb_0__1_.mux_top_track_36.out VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_1
Xinput24 chanx_right_in[29] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_1
Xinput46 chany_bottom_in[21] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_2
Xinput57 chany_bottom_in[4] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput35 chany_bottom_in[11] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_2
XFILLER_37_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_bottom_track_21.mux_l1_in_1_ net9 net21 sb_0__1_.mem_bottom_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_43_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_2_0_prog_clk sb_0__1_.mem_right_track_32.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_34.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_8_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_10.mux_l1_in_3_ net261 net58 sb_0__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_25_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_bottom_track_53.mux_l1_in_1__230 VGND VGND VPWR VPWR net230 sb_0__1_.mux_bottom_track_53.mux_l1_in_1__230/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_right_track_12.mux_l2_in_1_ net234 net41 sb_0__1_.mem_right_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_37.out sky130_fd_sc_hd__clkbuf_1
XFILLER_90_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_8_0_prog_clk sb_0__1_.mem_top_track_28.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_28.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_0__1_.mux_right_track_14.mux_l2_in_1__A1 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_40.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_40.out sky130_fd_sc_hd__clkbuf_1
XFILLER_74_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_4_2_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[2\] net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_0__1_.mux_right_track_32.mux_l1_in_0__A0 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input22_A chanx_right_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mux_top_track_52.mux_l1_in_0_ net12 net24 sb_0__1_.mem_top_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_top_track_10.mux_l3_in_0_ sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_5_X
+ sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X sb_0__1_.mem_top_track_10.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_14_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_34.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_34.out sky130_fd_sc_hd__clkbuf_1
XFILLER_68_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_right_track_24.mux_l1_in_0__A1 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_0_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[1\] net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_4_2_0_prog_clk cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.ccff_tail
+ net98 VGND VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_195_ sb_0__1_.mux_top_track_4.out VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__clkbuf_1
XFILLER_41_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__D sb_0__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput189 net189 VGND VGND VPWR VPWR chany_top_out_0[18] sky130_fd_sc_hd__buf_12
Xsb_0__1_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_28.out sky130_fd_sc_hd__clkbuf_1
Xoutput167 net167 VGND VGND VPWR VPWR chany_bottom_out[25] sky130_fd_sc_hd__buf_12
Xoutput156 net156 VGND VGND VPWR VPWR chany_bottom_out[15] sky130_fd_sc_hd__buf_12
Xoutput178 net178 VGND VGND VPWR VPWR chany_bottom_out[8] sky130_fd_sc_hd__buf_12
Xoutput145 net145 VGND VGND VPWR VPWR chanx_right_out[5] sky130_fd_sc_hd__buf_12
Xoutput123 net123 VGND VGND VPWR VPWR chanx_right_out[12] sky130_fd_sc_hd__buf_12
Xoutput134 net134 VGND VGND VPWR VPWR chanx_right_out[22] sky130_fd_sc_hd__buf_12
Xsb_0__1_.mux_top_track_10.mux_l2_in_1_ sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X sb_0__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_55_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mux_right_track_8.mux_l1_in_0__A0 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput25 chanx_right_in[2] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_1
Xinput14 chanx_right_in[1] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_1
Xinput36 chany_bottom_in[12] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput69 chany_top_in_0[15] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_2
X_178_ net35 VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_2
Xinput47 chany_bottom_in[22] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_2
Xinput58 chany_bottom_in[5] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_2
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.ccff_tail net97 VGND
+ VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_4.mux_l3_in_0_ sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
+ sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X sb_0__1_.mem_top_track_4.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_2__A0 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_bottom_track_21.mux_l1_in_0_ net85 net71 sb_0__1_.mem_bottom_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mux_right_track_22.mux_l2_in_1__A1 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input52_A chany_bottom_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_1.out sky130_fd_sc_hd__clkbuf_2
XFILLER_8_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_10.mux_l1_in_2_ net43 net25 sb_0__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_right_track_50.mux_l1_in_1__254 VGND VGND VPWR VPWR net254 sb_0__1_.mux_right_track_50.mux_l1_in_1__254/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_bottom_track_45.mux_l3_in_0_ sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X sb_0__1_.mem_bottom_track_45.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_right_track_12.mux_l2_in_0_ net104 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_12.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_68_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__210__A net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_8_0_prog_clk sb_0__1_.mem_top_track_20.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_28.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_16_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_2_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[1\] net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mux_top_track_4.mux_l2_in_1_ net267 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mem_top_track_4.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mux_right_track_32.mux_l1_in_0__A1 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input15_A chanx_right_in[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_45.mux_l2_in_1_ net228 net30 sb_0__1_.mem_bottom_track_45.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_54_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input7_A chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_1_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[0\] net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_29_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_top_track_4.mux_l1_in_2_ net60 net47 sb_0__1_.mem_top_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_9_0_prog_clk sb_0__1_.mem_right_track_20.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_20.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_58_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mux_top_track_6.mux_l1_in_2__A0 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input117_A top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input82_A chany_top_in_0[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mux_right_track_18.mux_l2_in_0__A0 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_194_ sb_0__1_.mux_top_track_6.out VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__clkbuf_2
XFILLER_2_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_56.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_56.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mux_top_track_44.mux_l1_in_1__A1 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_5_0_prog_clk sb_0__1_.mem_right_track_52.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_52.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xoutput135 net135 VGND VGND VPWR VPWR chanx_right_out[23] sky130_fd_sc_hd__buf_12
Xoutput168 net168 VGND VGND VPWR VPWR chany_bottom_out[26] sky130_fd_sc_hd__buf_12
Xoutput157 net157 VGND VGND VPWR VPWR chany_bottom_out[16] sky130_fd_sc_hd__buf_12
Xoutput179 net179 VGND VGND VPWR VPWR chany_bottom_out[9] sky130_fd_sc_hd__buf_12
Xoutput146 net146 VGND VGND VPWR VPWR chanx_right_out[6] sky130_fd_sc_hd__buf_12
Xoutput124 net124 VGND VGND VPWR VPWR chanx_right_out[13] sky130_fd_sc_hd__buf_12
XFILLER_70_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_top_track_10.mux_l2_in_0_ sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__213__A net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_177_ net34 VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__clkbuf_2
Xinput15 chanx_right_in[20] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput26 chanx_right_in[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2__A0 net78 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xinput48 chany_bottom_in[23] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_2
Xinput59 chany_bottom_in[6] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_2
Xinput37 chany_bottom_in[13] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__208__A net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_2__A1 net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input45_A chany_bottom_in[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_top_track_10.mux_l1_in_1_ net7 net19 sb_0__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_right_track_40.mux_l1_in_0__A1 net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.ccff_tail net97 VGND
+ VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_1
XFILLER_16_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_9_0_prog_clk sb_0__1_.mem_bottom_track_29.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_29.ccff_tail sky130_fd_sc_hd__dfrtp_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_2_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[0\] net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xsb_0__1_.mux_top_track_4.mux_l2_in_0_ sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_top_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_bottom_track_45.mux_l2_in_0_ net12 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_bottom_track_45.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_39_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_12.mux_l1_in_0_ net71 net75 sb_0__1_.mem_right_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_62_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_24.mux_l2_in_0_ sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_24.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_81_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__216__A net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_2_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_0_0_prog_clk
+ net2 net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xsb_0__1_.mux_right_track_36.mux_l3_in_0_ sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X sb_0__1_.mem_right_track_36.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_top_track_4.mux_l1_in_1_ net27 net9 sb_0__1_.mem_top_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_14_0_prog_clk sb_0__1_.mem_right_track_20.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_20.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_67_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_12_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_12_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_193_ net51 VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__clkbuf_2
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_right_track_46.mux_l2_in_0__252 VGND VGND VPWR VPWR net252 sb_0__1_.mux_right_track_46.mux_l2_in_0__252/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_input75_A chany_top_in_0[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_bottom_track_1.mux_l3_in_0_ sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X
+ sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X sb_0__1_.mem_bottom_track_1.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_17_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_5_0_prog_clk sb_0__1_.mem_right_track_50.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_52.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_70_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput125 net125 VGND VGND VPWR VPWR chanx_right_out[14] sky130_fd_sc_hd__buf_12
Xsb_0__1_.mux_right_track_24.mux_l1_in_1_ net241 net62 sb_0__1_.mem_right_track_24.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xoutput169 net169 VGND VGND VPWR VPWR chany_bottom_out[27] sky130_fd_sc_hd__buf_12
Xoutput158 net158 VGND VGND VPWR VPWR chany_bottom_out[17] sky130_fd_sc_hd__buf_12
Xoutput147 net147 VGND VGND VPWR VPWR chanx_right_out[7] sky130_fd_sc_hd__buf_12
Xoutput136 net136 VGND VGND VPWR VPWR chanx_right_out[24] sky130_fd_sc_hd__buf_12
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_36.mux_l2_in_1_ net247 net33 sb_0__1_.mem_right_track_36.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_36_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_176_ net62 VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__clkbuf_2
Xinput16 chanx_right_in[21] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput27 chanx_right_in[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_1
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2__A1 net47 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xinput49 chany_bottom_in[24] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput38 chany_bottom_in[14] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_2
XANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_1.mux_l2_in_1_ net275 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mem_bottom_track_1.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input38_A chany_bottom_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_top_track_10.mux_l1_in_0_ net118 net116 sb_0__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_159_ net77 VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__clkbuf_2
XFILLER_88_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_7_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_right_track_26.mux_l1_in_1__A1 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_12_0_prog_clk sb_0__1_.mem_bottom_track_29.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_29.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_3_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_6.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_0_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_2.ccff_tail net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_0__S sb_0__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_1.mux_l1_in_2_ right_width_0_height_0_subtile_3__pin_inpad_0_
+ right_width_0_height_0_subtile_0__pin_inpad_0_ sb_0__1_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_21_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input20_A chanx_right_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_14_0_prog_clk sb_0__1_.mem_right_track_18.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_20.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_71_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_top_track_4.mux_l1_in_0_ net21 net117 sb_0__1_.mem_top_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA__142__A net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_192_ sb_0__1_.mux_top_track_10.out VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__clkbuf_2
Xsb_0__1_.mux_bottom_track_45.mux_l1_in_0_ net24 net67 sb_0__1_.mem_bottom_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_41_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input68_A chany_top_in_0[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_2.mux_l3_in_0_ sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
+ sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X sb_0__1_.mem_right_track_2.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_24.mux_l1_in_0_ net110 net92 sb_0__1_.mem_right_track_24.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xoutput137 net137 VGND VGND VPWR VPWR chanx_right_out[25] sky130_fd_sc_hd__buf_12
Xoutput159 net159 VGND VGND VPWR VPWR chany_bottom_out[18] sky130_fd_sc_hd__buf_12
Xoutput148 net148 VGND VGND VPWR VPWR chanx_right_out[8] sky130_fd_sc_hd__buf_12
Xoutput126 net126 VGND VGND VPWR VPWR chanx_right_out[15] sky130_fd_sc_hd__buf_12
XFILLER_55_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_36.mux_l2_in_0_ net44 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_36.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_46_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_right_track_28.mux_l1_in_1__243 VGND VGND VPWR VPWR net243 sb_0__1_.mux_right_track_28.mux_l1_in_1__243/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_36_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_175_ sb_0__1_.mux_top_track_44.out VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__clkbuf_1
Xinput17 chanx_right_in[22] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_1
Xinput28 chanx_right_in[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_1
Xinput39 chany_bottom_in[15] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_2
XFILLER_9_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_top_track_0.mux_l1_in_3__S sb_0__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_bottom_track_11.mux_l1_in_3__276 VGND VGND VPWR VPWR net276 sb_0__1_.mux_bottom_track_11.mux_l1_in_3__276/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_87_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_3_0_prog_clk sb_0__1_.mem_right_track_26.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_26.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_0__1_.mux_right_track_34.mux_l1_in_1__A1 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_2.mux_l2_in_1_ net238 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mem_right_track_2.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_bottom_track_1.mux_l2_in_0_ sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_bottom_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_42_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_158_ net76 VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__clkbuf_2
XANTENNA__150__A net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input50_A chany_bottom_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_7_0_prog_clk sb_0__1_.mem_bottom_track_21.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_29.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_2.mux_l1_in_2_ net48 net111 sb_0__1_.mem_right_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_bottom_track_1.mux_l1_in_1_ net32 net15 sb_0__1_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_79_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_12.mux_l2_in_1__234 VGND VGND VPWR VPWR net234 sb_0__1_.mux_right_track_12.mux_l2_in_1__234/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input98_A prog_reset_bottom_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mux_top_track_12.mux_l1_in_2__A0 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_12.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_input13_A chanx_right_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3__A0 net69 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_32.mux_l1_in_1__245 VGND VGND VPWR VPWR net245 sb_0__1_.mux_right_track_32.mux_l1_in_1__245/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_35_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_6_0_prog_clk sb_0__1_.mem_bottom_track_3.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_3.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_76_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input5_A chanx_right_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_191_ sb_0__1_.mux_top_track_12.out VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XFILLER_1_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput138 net138 VGND VGND VPWR VPWR chanx_right_out[26] sky130_fd_sc_hd__buf_12
Xoutput149 net149 VGND VGND VPWR VPWR chanx_right_out[9] sky130_fd_sc_hd__buf_12
Xoutput127 net127 VGND VGND VPWR VPWR chanx_right_out[16] sky130_fd_sc_hd__buf_12
XFILLER_70_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2__A0 net55 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input115_A top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input80_A chany_top_in_0[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput18 chanx_right_in[23] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_174_ net60 VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__clkbuf_2
Xinput29 chanx_right_in[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_93_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__148__A net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_3_0_prog_clk sb_0__1_.mem_right_track_24.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_26.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_28_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_2.mux_l2_in_0_ sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_51_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_157_ sb_0__1_.mux_bottom_track_21.out VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__clkbuf_2
XFILLER_88_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_36.mux_l1_in_0_ net108 net74 sb_0__1_.mem_right_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_84_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_48.mux_l2_in_0_ net253 sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_48.ccff_tail VGND VGND VPWR VPWR sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input43_A chany_bottom_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_209_ net98 VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_1
XFILLER_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_50.mux_l2_in_0_ sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_50.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_80_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_right_track_2.mux_l1_in_1_ net108 net105 sb_0__1_.mem_right_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xclkbuf_4_9_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_9_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_sb_0__1_.mux_top_track_20.mux_l1_in_2__A0 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_11_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_bottom_track_1.mux_l1_in_0_ net64 net81 sb_0__1_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_21_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__156__A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_11.out sky130_fd_sc_hd__clkbuf_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net93 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR right_width_0_height_0_subtile_3__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XANTENNA_sb_0__1_.mux_top_track_12.mux_l1_in_2__A1 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_ cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_91_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3__A1 net38 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_50.mux_l1_in_1_ net254 net50 sb_0__1_.mem_right_track_50.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_6_0_prog_clk sb_0__1_.mem_bottom_track_3.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_3.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_35_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_190_ net48 VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__clkbuf_2
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_bottom_track_13.mux_l1_in_2__A0 right_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput139 net139 VGND VGND VPWR VPWR chanx_right_out[27] sky130_fd_sc_hd__buf_12
Xoutput128 net128 VGND VGND VPWR VPWR chanx_right_out[17] sky130_fd_sc_hd__buf_12
XFILLER_55_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input108_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput19 chanx_right_in[24] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_1
X_173_ net59 VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input73_A chany_top_in_0[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_11_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_11_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_77_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_28.out sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_156_ net73 VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_2
XFILLER_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__159__A net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_bottom_track_29.mux_l2_in_1__279 VGND VGND VPWR VPWR net279 sb_0__1_.mux_bottom_track_29.mux_l2_in_1__279/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_68_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3_ net271 net89 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input36_A chany_bottom_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_right_track_46.mux_l1_in_0__A0 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_208_ net98 VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__clkbuf_1
X_139_ net85 VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__clkbuf_2
Xsb_0__1_.mux_right_track_2.mux_l1_in_0_ net78 net84 sb_0__1_.mem_right_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_57_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_top_track_20.mux_l1_in_2__A1 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_6.out sky130_fd_sc_hd__clkbuf_1
XANTENNA__172__A net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_0__1_.mux_right_track_38.mux_l1_in_0__A1 net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_14_0_prog_clk sb_0__1_.mem_right_track_12.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_12.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_38_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_48.mux_l1_in_0_ net49 net106 sb_0__1_.mem_right_track_48.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_30_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4_ sb_0__1_.mux_bottom_track_37.out
+ net35 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mux_bottom_track_21.mux_l1_in_2__A0 right_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_50.mux_l1_in_0_ net111 net107 sb_0__1_.mem_right_track_50.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_6_0_prog_clk sb_0__1_.mem_bottom_track_1.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_bottom_track_3.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l4_in_0_ cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X cby_0__1_.cby_0__1_.mem_right_ipin_0.ccff_tail
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_4_0_prog_clk sb_0__1_.mem_right_track_44.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_44.ccff_tail sky130_fd_sc_hd__dfrtp_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_5.mux_l2_in_1__229 VGND VGND VPWR VPWR net229 sb_0__1_.mux_bottom_track_5.mux_l2_in_1__229/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_17_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput129 net129 VGND VGND VPWR VPWR chanx_right_out[18] sky130_fd_sc_hd__buf_12
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net96 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_23_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_172_ net58 VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input66_A chany_top_in_0[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l3_in_1_ cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__180__A net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_right_track_0.mux_l1_in_1__A0 net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_30.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_30.out sky130_fd_sc_hd__clkbuf_1
XFILLER_11_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_155_ net72 VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1__A1 net51 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input29_A chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_2_ net58 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_207_ net98 VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_0__1_.mux_right_track_46.mux_l1_in_0__A1 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_138_ net74 VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_2
Xsb_0__1_.mux_top_track_0.mux_l1_in_3_ net260 net34 sb_0__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_right_track_24.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_24.out sky130_fd_sc_hd__clkbuf_1
XFILLER_2_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_bottom_track_5.mux_l1_in_0__A0 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mux_right_track_12.mux_l1_in_0__A0 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk sb_0__1_.mem_right_track_12.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_12.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3_ net72 net41 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_right_track_18.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_18.out sky130_fd_sc_hd__clkbuf_1
XFILLER_29_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input96_A gfpga_pad_io_soc_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_4_0_prog_clk sb_0__1_.mem_right_track_40.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_44.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mux_top_track_0.mux_l3_in_0_ sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X
+ sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X sb_0__1_.mem_top_track_0.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_49_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input11_A chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput119 net119 VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__buf_12
XANTENNA__178__A net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_18.mux_l3_in_0_ sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_1_X sb_0__1_.mem_right_track_18.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_31_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input3_A chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_171_ sb_0__1_.mux_top_track_52.out VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__clkbuf_2
Xsb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_11_0_prog_clk sb_0__1_.mem_right_track_18.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_18.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_22_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_20.mux_l3_in_0_ sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X sb_0__1_.mem_right_track_20.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_input59_A chany_bottom_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l3_in_0_ cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mux_right_track_0.mux_l1_in_1__A1 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_top_track_0.mux_l2_in_1_ sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X sb_0__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_51_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input113_A test_enable_right_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mux_right_track_54.mux_l1_in_0__A1 net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_154_ net71 VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_2
XFILLER_92_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_18.mux_l2_in_1_ net237 net37 sb_0__1_.mem_right_track_18.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_33_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_20.mux_l2_in_1_ net239 net35 sb_0__1_.mem_right_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_74_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_1_ cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_right_track_52.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_52.out sky130_fd_sc_hd__clkbuf_1
XFILLER_74_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_137_ sb_0__1_.mux_right_track_0.out VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_1
X_206_ net98 VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__dlymetal6s2s_1
Xsb_0__1_.mux_top_track_0.mux_l1_in_2_ net51 net29 sb_0__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_65_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__186__A net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mux_bottom_track_5.mux_l1_in_0__A1 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input41_A chany_bottom_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_5 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_14_0_prog_clk sb_0__1_.mem_right_track_10.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_12.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_10_0_prog_clk sb_0__1_.mem_top_track_2.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_46.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_46.out sky130_fd_sc_hd__clkbuf_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2_ sb_0__1_.mux_bottom_track_13.out
+ net48 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_55_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input89_A chany_top_in_0[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_8_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_8_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
Xsb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_13_0_prog_clk sb_0__1_.mem_right_track_4.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_4.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_90_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_right_track_44.mux_l2_in_0__251 VGND VGND VPWR VPWR net251 sb_0__1_.mux_right_track_44.mux_l2_in_0__251/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_72_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2__A0 net77 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_bottom_track_3.mux_l2_in_1__A1 right_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mux_right_track_10.mux_l2_in_1__A1 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_14_0_prog_clk sb_0__1_.mem_right_track_18.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_18.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
X_170_ net56 VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkbuf_2
XFILLER_54_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__189__A net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_top_track_0.mux_l2_in_0_ sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input106_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_153_ sb_0__1_.mux_bottom_track_29.out VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input71_A chany_top_in_0[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_18.mux_l2_in_0_ net107 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_18.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mux_right_track_20.mux_l1_in_0__A1 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_10_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_10_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
Xsb_0__1_.mux_right_track_20.mux_l2_in_0_ net108 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_20.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__274 VGND VGND VPWR VPWR net274
+ cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__274/LO sky130_fd_sc_hd__conb_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_0_ cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_136_ sb_0__1_.mux_right_track_2.out VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_2
X_205_ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__clkbuf_1
XFILLER_23_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_top_track_0.mux_l1_in_1_ net11 net23 sb_0__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_80_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_7.out sky130_fd_sc_hd__clkbuf_2
XFILLER_56_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mux_right_track_4.mux_l1_in_0__A0 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input34_A chany_bottom_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_119_ sb_0__1_.mux_right_track_36.out VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_11_0_prog_clk sb_0__1_.mem_top_track_2.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_2.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_53_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1_ sb_0__1_.mux_bottom_track_7.out
+ net51 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk sb_0__1_.mem_right_track_4.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_4.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_20_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_2__A0 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2__A1 net46 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_2.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_top_track_28.mux_l3_in_0_ sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_2_X sb_0__1_.mem_top_track_28.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_right_track_26.mux_l1_in_1__242 VGND VGND VPWR VPWR net242 sb_0__1_.mux_right_track_26.mux_l1_in_1__242/LO
+ sky130_fd_sc_hd__conb_1
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_14_0_prog_clk sb_0__1_.mem_right_track_16.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_18.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_14_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_3_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_right_track_8.mux_l2_in_1__259 VGND VGND VPWR VPWR net259 sb_0__1_.mux_right_track_8.mux_l2_in_1__259/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4__A1 net35 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_152_ net69 VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input64_A chany_top_in_0[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_top_track_28.mux_l2_in_1_ net265 net44 sb_0__1_.mem_top_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_83_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_2_0_prog_clk sb_0__1_.mem_right_track_30.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_30.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_17_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mux_top_track_2.mux_l1_in_2__A0 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__A1 net89 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_204_ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__clkbuf_1
X_135_ sb_0__1_.mux_right_track_4.out VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_top_track_0.mux_l1_in_0_ net118 net115 sb_0__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_bottom_track_7.mux_l1_in_3_ net231 right_width_0_height_0_subtile_2__pin_inpad_0_
+ sb_0__1_.mem_bottom_track_7.mem_out\[0\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mux_right_track_14.mux_l2_in_0__A0 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_18.mux_l1_in_0_ net91 net67 sb_0__1_.mem_right_track_18.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_0__1_.mux_right_track_10.mux_l2_in_1__233 VGND VGND VPWR VPWR net233 sb_0__1_.mux_right_track_10.mux_l2_in_1__233/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_60_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input27_A chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_4_2_0_prog_clk cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.ccff_tail
+ net98 VGND VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_118_ sb_0__1_.mux_right_track_38.out VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mux_right_track_20.mux_l1_in_0_ net87 net65 sb_0__1_.mem_right_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__1_.mux_bottom_track_53.mux_l2_in_0_ sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_0_X net120 VGND VGND VPWR VPWR
+ sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_11_0_prog_clk sb_0__1_.mem_top_track_0.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_2.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0_ sb_0__1_.mux_bottom_track_1.out
+ net54 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_76_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_8_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_right_track_32.mux_l2_in_0_ sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_32.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_29_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_0_0_prog_clk sb_0__1_.mem_right_track_36.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_36.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_15_0_prog_clk sb_0__1_.mem_right_track_2.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_4.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_20_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_right_track_2.mux_l1_in_2__A1 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_30.mux_l1_in_1__244 VGND VGND VPWR VPWR net244 sb_0__1_.mux_right_track_30.mux_l1_in_1__244/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_bottom_track_7.mux_l3_in_0_ sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_5_X
+ sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_4_X sb_0__1_.mem_bottom_track_11.ccff_head
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_1_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mux_bottom_track_53.mux_l1_in_1_ net230 net31 sb_0__1_.mem_bottom_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_input94_A gfpga_pad_io_soc_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_bottom_track_3.mux_l2_in_1__226 VGND VGND VPWR VPWR net226 sb_0__1_.mux_bottom_track_3.mux_l2_in_1__226/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_31_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_right_track_32.mux_l1_in_1_ net245 net56 sb_0__1_.mem_right_track_32.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_bottom_track_7.mux_l2_in_1_ sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X sb_0__1_.mem_bottom_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_22_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_top_track_4.mux_l1_in_0__A1 net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input1_A ccff_head VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_151_ net68 VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_2
XFILLER_77_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mux_right_track_22.mux_l2_in_0__A0 net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input57_A chany_bottom_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_top_track_28.mux_l2_in_0_ sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_top_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_53_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_2_0_prog_clk sb_0__1_.mem_right_track_28.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_30.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_0__1_.mux_top_track_28.mux_l1_in_0__A1 net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input111_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mux_top_track_2.mux_l1_in_2__A1 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_203_ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__clkbuf_1
X_134_ sb_0__1_.mux_right_track_6.out VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_2
Xsb_0__1_.mux_bottom_track_7.mux_l1_in_2_ right_width_0_height_0_subtile_0__pin_inpad_0_
+ net14 sb_0__1_.mem_bottom_track_7.mem_out\[0\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_bottom_track_11.mux_l1_in_3_ net276 right_width_0_height_0_subtile_3__pin_inpad_0_
+ sb_0__1_.mem_bottom_track_11.mem_out\[0\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_top_track_28.mux_l1_in_1_ net39 net4 sb_0__1_.mem_top_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_55_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_bottom_track_13.mux_l2_in_1__277 VGND VGND VPWR VPWR net277 sb_0__1_.mux_bottom_track_13.mux_l2_in_1__277/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_117_ sb_0__1_.mux_right_track_40.out VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_0__1_.mux_bottom_track_29.mux_l1_in_0__A0 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_0_0_prog_clk sb_0__1_.mem_right_track_36.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_36.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_4_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_right_track_8.mux_l3_in_0_ sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_4_X
+ sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_3_X sb_0__1_.mem_right_track_10.ccff_head
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_34_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input87_A chany_top_in_0[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_bottom_track_53.mux_l1_in_0_ net13 net65 sb_0__1_.mem_bottom_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_bottom_track_11.mux_l3_in_0_ sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_5_X
+ sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_4_X sb_0__1_.mem_bottom_track_11.ccff_tail
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_31_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_bottom_track_1.mux_l2_in_1__275 VGND VGND VPWR VPWR net275 sb_0__1_.mux_bottom_track_1.mux_l2_in_1__275/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_63_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_right_track_32.mux_l1_in_0_ net106 net86 sb_0__1_.mem_right_track_32.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_39_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_7_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_7_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_14_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_top_track_44.mux_l1_in_1__268 VGND VGND VPWR VPWR net268 sb_0__1_.mux_top_track_44.mux_l1_in_1__268/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_22_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_right_track_44.mux_l2_in_0_ net251 sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_right_track_44.ccff_tail VGND VGND VPWR VPWR sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_93_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_8.mux_l2_in_1_ net259 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_2_X
+ sb_0__1_.mem_right_track_8.mem_out\[1\] VGND VGND VPWR VPWR sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_bottom_track_7.mux_l2_in_0_ sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_bottom_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_36_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_bottom_track_11.mux_l2_in_1_ sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_3_X
+ sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_2_X sb_0__1_.mem_bottom_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xcby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_4_0_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[2\] net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
X_150_ net67 VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_1__A0 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input104_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mux_right_track_8.mux_l1_in_2_ net43 net111 sb_0__1_.mem_right_track_8.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
X_133_ sb_0__1_.mux_right_track_8.out VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_2
X_202_ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__clkbuf_1
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_bottom_track_7.mux_l1_in_1_ net6 net18 sb_0__1_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_73_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_bottom_track_11.mux_l1_in_2_ right_width_0_height_0_subtile_1__pin_inpad_0_
+ net25 sb_0__1_.mem_bottom_track_11.mem_out\[0\] VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__1_.mux_top_track_28.mux_l1_in_0_ net16 net117 sb_0__1_.mem_top_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_85_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_116_ net36 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_0__1_.mux_bottom_track_29.mux_l1_in_0__A1 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_3_0_prog_clk sb_0__1_.mem_right_track_34.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_right_track_36.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_4_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input32_A chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_0__1_.mux_right_track_30.mux_l1_in_1__A1 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_12_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_2.out sky130_fd_sc_hd__clkbuf_1
XFILLER_9_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1__A0 net81 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__1_.mux_right_track_8.mux_l2_in_0_ sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_right_track_8.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_3_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__1_.mux_bottom_track_11.mux_l2_in_0_ sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X sb_0__1_.mem_bottom_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_47_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_0_0_prog_clk
+ cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[1\] net98 VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_0__1_.mux_right_track_6.mux_l1_in_1__A1 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_18_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mux_right_track_22.mux_l2_in_1__240 VGND VGND VPWR VPWR net240 sb_0__1_.mux_right_track_22.mux_l2_in_1__240/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__1_.mux_right_track_44.mux_l1_in_0_ net40 net104 sb_0__1_.mem_right_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_3_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_right_track_8.mux_l1_in_1_ net108 net105 sb_0__1_.mem_right_track_8.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mux_bottom_track_37.mux_l1_in_0__A1 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_132_ sb_0__1_.mux_right_track_10.out VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_201_ cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__clkbuf_1
Xsb_0__1_.mux_right_track_56.mux_l2_in_0_ net257 sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__1_.mem_bottom_track_1.ccff_head VGND VGND VPWR VPWR sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_0__1_.mux_right_track_26.mux_l1_in_0__A0 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_bottom_track_7.mux_l1_in_0_ net89 net76 sb_0__1_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input62_A chany_bottom_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mux_bottom_track_7.mux_l1_in_3__231 VGND VGND VPWR VPWR net231 sb_0__1_.mux_bottom_track_7.mux_l1_in_3__231/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__1_.mux_bottom_track_11.mux_l1_in_1_ net7 net19 sb_0__1_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_64_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__211__A net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_115_ sb_0__1_.mux_right_track_44.out VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_0__1_.mux_right_track_18.mux_l1_in_0__A1 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_0__1_.mux_top_track_52.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_top_track_52.out sky130_fd_sc_hd__clkbuf_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3_ net272 net88 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__206__A net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input25_A chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_8_0_prog_clk sb_0__1_.mem_top_track_10.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_0__1_.mem_top_track_10.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_0_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__1_.mux_right_track_20.sky130_fd_sc_hd__buf_4_0_ sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_0__1_.mux_right_track_20.out sky130_fd_sc_hd__clkbuf_1
XFILLER_16_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
.ends

