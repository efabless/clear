magic
tech sky130A
magscale 1 2
timestamp 1625790302
<< locali >>
rect 5181 15351 5215 15521
rect 14197 11067 14231 11305
rect 6469 8279 6503 8449
rect 11529 8347 11563 8585
rect 9965 2499 9999 2601
<< viali >>
rect 2513 17289 2547 17323
rect 2881 17289 2915 17323
rect 3985 17289 4019 17323
rect 4721 17289 4755 17323
rect 5917 17289 5951 17323
rect 14197 17289 14231 17323
rect 14749 17289 14783 17323
rect 2053 17221 2087 17255
rect 3525 17221 3559 17255
rect 4261 17221 4295 17255
rect 4997 17221 5031 17255
rect 6561 17221 6595 17255
rect 7297 17221 7331 17255
rect 8033 17221 8067 17255
rect 8401 17221 8435 17255
rect 9229 17221 9263 17255
rect 3157 17153 3191 17187
rect 5365 17153 5399 17187
rect 6377 17153 6411 17187
rect 12265 17153 12299 17187
rect 13737 17153 13771 17187
rect 1409 17085 1443 17119
rect 1685 17085 1719 17119
rect 3709 17085 3743 17119
rect 6929 17085 6963 17119
rect 7665 17085 7699 17119
rect 7849 17085 7883 17119
rect 8585 17085 8619 17119
rect 10149 17085 10183 17119
rect 10517 17085 10551 17119
rect 10885 17085 10919 17119
rect 11253 17085 11287 17119
rect 11529 17085 11563 17119
rect 11989 17085 12023 17119
rect 13461 17085 13495 17119
rect 14013 17085 14047 17119
rect 15117 17085 15151 17119
rect 15485 17085 15519 17119
rect 2237 17017 2271 17051
rect 2605 17017 2639 17051
rect 2973 17017 3007 17051
rect 3341 17017 3375 17051
rect 4077 17017 4111 17051
rect 4445 17017 4479 17051
rect 4813 17017 4847 17051
rect 5181 17017 5215 17051
rect 5549 17017 5583 17051
rect 5825 17017 5859 17051
rect 6193 17017 6227 17051
rect 6745 17017 6779 17051
rect 7113 17017 7147 17051
rect 7481 17017 7515 17051
rect 8217 17017 8251 17051
rect 8769 17017 8803 17051
rect 8953 17017 8987 17051
rect 9413 17017 9447 17051
rect 12725 17017 12759 17051
rect 14657 17017 14691 17051
rect 14933 17017 14967 17051
rect 15301 17017 15335 17051
rect 9965 16949 9999 16983
rect 10333 16949 10367 16983
rect 10701 16949 10735 16983
rect 11069 16949 11103 16983
rect 11437 16949 11471 16983
rect 12081 16949 12115 16983
rect 12633 16949 12667 16983
rect 13921 16949 13955 16983
rect 1869 16745 1903 16779
rect 2881 16745 2915 16779
rect 3341 16745 3375 16779
rect 10241 16745 10275 16779
rect 10609 16745 10643 16779
rect 10977 16745 11011 16779
rect 11345 16745 11379 16779
rect 11805 16745 11839 16779
rect 13093 16745 13127 16779
rect 14105 16745 14139 16779
rect 1409 16677 1443 16711
rect 1961 16677 1995 16711
rect 2697 16677 2731 16711
rect 4997 16677 5031 16711
rect 5365 16677 5399 16711
rect 5733 16677 5767 16711
rect 12357 16677 12391 16711
rect 13461 16677 13495 16711
rect 14565 16677 14599 16711
rect 15301 16677 15335 16711
rect 1593 16609 1627 16643
rect 2145 16609 2179 16643
rect 2329 16609 2363 16643
rect 2513 16609 2547 16643
rect 3065 16609 3099 16643
rect 5181 16609 5215 16643
rect 5549 16609 5583 16643
rect 5917 16609 5951 16643
rect 12725 16609 12759 16643
rect 12909 16609 12943 16643
rect 14013 16609 14047 16643
rect 14933 16609 14967 16643
rect 15669 16609 15703 16643
rect 13645 16541 13679 16575
rect 3617 16473 3651 16507
rect 7113 16473 7147 16507
rect 12173 16473 12207 16507
rect 12541 16473 12575 16507
rect 13277 16473 13311 16507
rect 14749 16473 14783 16507
rect 15117 16473 15151 16507
rect 3249 16405 3283 16439
rect 3985 16405 4019 16439
rect 6745 16405 6779 16439
rect 14473 16405 14507 16439
rect 1501 16201 1535 16235
rect 5181 16201 5215 16235
rect 6745 16201 6779 16235
rect 7021 16201 7055 16235
rect 7297 16201 7331 16235
rect 8861 16201 8895 16235
rect 13645 16201 13679 16235
rect 14565 16201 14599 16235
rect 14749 16201 14783 16235
rect 14933 16201 14967 16235
rect 2053 16133 2087 16167
rect 6469 16133 6503 16167
rect 13829 16133 13863 16167
rect 2329 16065 2363 16099
rect 8033 16065 8067 16099
rect 1961 15997 1995 16031
rect 2237 15997 2271 16031
rect 5365 15997 5399 16031
rect 6653 15997 6687 16031
rect 6929 15997 6963 16031
rect 7205 15997 7239 16031
rect 7481 15997 7515 16031
rect 8677 15997 8711 16031
rect 15393 15997 15427 16031
rect 15577 15997 15611 16031
rect 1593 15929 1627 15963
rect 8217 15929 8251 15963
rect 15025 15929 15059 15963
rect 15209 15929 15243 15963
rect 2513 15861 2547 15895
rect 2789 15861 2823 15895
rect 4721 15861 4755 15895
rect 5549 15861 5583 15895
rect 7573 15861 7607 15895
rect 7757 15861 7791 15895
rect 8401 15861 8435 15895
rect 3893 15657 3927 15691
rect 4169 15657 4203 15691
rect 4721 15657 4755 15691
rect 5273 15657 5307 15691
rect 5549 15657 5583 15691
rect 6745 15657 6779 15691
rect 8033 15657 8067 15691
rect 8585 15657 8619 15691
rect 9137 15657 9171 15691
rect 9413 15657 9447 15691
rect 9689 15657 9723 15691
rect 9965 15657 9999 15691
rect 15393 15657 15427 15691
rect 1869 15589 1903 15623
rect 6101 15589 6135 15623
rect 7665 15589 7699 15623
rect 15485 15589 15519 15623
rect 1593 15521 1627 15555
rect 4077 15521 4111 15555
rect 4353 15521 4387 15555
rect 4629 15521 4663 15555
rect 4905 15521 4939 15555
rect 5181 15521 5215 15555
rect 5457 15521 5491 15555
rect 5733 15521 5767 15555
rect 6837 15521 6871 15555
rect 7573 15521 7607 15555
rect 8217 15521 8251 15555
rect 8493 15521 8527 15555
rect 8769 15521 8803 15555
rect 9321 15521 9355 15555
rect 9597 15521 9631 15555
rect 9873 15521 9907 15555
rect 10149 15521 10183 15555
rect 15025 15521 15059 15555
rect 1409 15385 1443 15419
rect 4445 15385 4479 15419
rect 5089 15385 5123 15419
rect 7021 15453 7055 15487
rect 7849 15453 7883 15487
rect 15209 15453 15243 15487
rect 6285 15385 6319 15419
rect 8309 15385 8343 15419
rect 8953 15385 8987 15419
rect 5181 15317 5215 15351
rect 5825 15317 5859 15351
rect 6377 15317 6411 15351
rect 7205 15317 7239 15351
rect 10333 15317 10367 15351
rect 5549 15113 5583 15147
rect 8125 15113 8159 15147
rect 8953 15113 8987 15147
rect 9321 15113 9355 15147
rect 5273 14977 5307 15011
rect 6193 14977 6227 15011
rect 7021 14977 7055 15011
rect 7849 14977 7883 15011
rect 8677 14977 8711 15011
rect 4537 14909 4571 14943
rect 5917 14909 5951 14943
rect 6009 14909 6043 14943
rect 7757 14909 7791 14943
rect 9137 14909 9171 14943
rect 6929 14841 6963 14875
rect 8585 14841 8619 14875
rect 4721 14773 4755 14807
rect 5089 14773 5123 14807
rect 5181 14773 5215 14807
rect 6469 14773 6503 14807
rect 6837 14773 6871 14807
rect 7297 14773 7331 14807
rect 7665 14773 7699 14807
rect 8493 14773 8527 14807
rect 9505 14773 9539 14807
rect 4629 14569 4663 14603
rect 4997 14569 5031 14603
rect 5457 14569 5491 14603
rect 4537 14501 4571 14535
rect 7052 14501 7086 14535
rect 7757 14501 7791 14535
rect 8493 14501 8527 14535
rect 9689 14501 9723 14535
rect 10149 14501 10183 14535
rect 1593 14433 1627 14467
rect 7849 14433 7883 14467
rect 8585 14433 8619 14467
rect 4353 14365 4387 14399
rect 5549 14365 5583 14399
rect 5641 14365 5675 14399
rect 7297 14365 7331 14399
rect 7941 14365 7975 14399
rect 8309 14365 8343 14399
rect 1409 14297 1443 14331
rect 9413 14297 9447 14331
rect 9597 14297 9631 14331
rect 9873 14297 9907 14331
rect 5089 14229 5123 14263
rect 5917 14229 5951 14263
rect 7389 14229 7423 14263
rect 8953 14229 8987 14263
rect 9229 14229 9263 14263
rect 2513 14025 2547 14059
rect 2789 14025 2823 14059
rect 8769 14025 8803 14059
rect 4077 13957 4111 13991
rect 6469 13957 6503 13991
rect 7941 13957 7975 13991
rect 4537 13889 4571 13923
rect 4721 13889 4755 13923
rect 8493 13889 8527 13923
rect 9229 13889 9263 13923
rect 9321 13889 9355 13923
rect 10241 13889 10275 13923
rect 2697 13821 2731 13855
rect 2973 13821 3007 13855
rect 4905 13821 4939 13855
rect 5161 13821 5195 13855
rect 7593 13821 7627 13855
rect 7849 13821 7883 13855
rect 10057 13821 10091 13855
rect 8309 13753 8343 13787
rect 4445 13685 4479 13719
rect 6285 13685 6319 13719
rect 8401 13685 8435 13719
rect 9137 13685 9171 13719
rect 9597 13685 9631 13719
rect 9965 13685 9999 13719
rect 10425 13685 10459 13719
rect 10609 13685 10643 13719
rect 2605 13481 2639 13515
rect 3433 13481 3467 13515
rect 3893 13481 3927 13515
rect 4537 13481 4571 13515
rect 8309 13481 8343 13515
rect 8861 13481 8895 13515
rect 9965 13481 9999 13515
rect 10425 13481 10459 13515
rect 1593 13413 1627 13447
rect 6592 13413 6626 13447
rect 7196 13413 7230 13447
rect 8585 13413 8619 13447
rect 1409 13345 1443 13379
rect 2789 13345 2823 13379
rect 3341 13345 3375 13379
rect 4077 13345 4111 13379
rect 4353 13345 4387 13379
rect 4997 13345 5031 13379
rect 9505 13345 9539 13379
rect 10333 13345 10367 13379
rect 10977 13345 11011 13379
rect 3525 13277 3559 13311
rect 5089 13277 5123 13311
rect 5273 13277 5307 13311
rect 6837 13277 6871 13311
rect 6929 13277 6963 13311
rect 9597 13277 9631 13311
rect 9689 13277 9723 13311
rect 10609 13277 10643 13311
rect 4629 13209 4663 13243
rect 9137 13209 9171 13243
rect 11345 13209 11379 13243
rect 2973 13141 3007 13175
rect 5457 13141 5491 13175
rect 10793 13141 10827 13175
rect 11161 13141 11195 13175
rect 2605 12937 2639 12971
rect 6285 12937 6319 12971
rect 7849 12937 7883 12971
rect 11437 12937 11471 12971
rect 2513 12869 2547 12903
rect 9321 12869 9355 12903
rect 10241 12869 10275 12903
rect 1961 12801 1995 12835
rect 3249 12801 3283 12835
rect 9965 12801 9999 12835
rect 10701 12801 10735 12835
rect 10885 12801 10919 12835
rect 11345 12801 11379 12835
rect 2145 12733 2179 12767
rect 2973 12733 3007 12767
rect 4813 12733 4847 12767
rect 4905 12733 4939 12767
rect 6469 12733 6503 12767
rect 7941 12733 7975 12767
rect 9781 12733 9815 12767
rect 11897 12733 11931 12767
rect 3065 12665 3099 12699
rect 4546 12665 4580 12699
rect 5150 12665 5184 12699
rect 6714 12665 6748 12699
rect 8186 12665 8220 12699
rect 9873 12665 9907 12699
rect 11805 12665 11839 12699
rect 2053 12597 2087 12631
rect 3433 12597 3467 12631
rect 9413 12597 9447 12631
rect 10609 12597 10643 12631
rect 11069 12597 11103 12631
rect 1869 12393 1903 12427
rect 3341 12393 3375 12427
rect 3709 12393 3743 12427
rect 4077 12393 4111 12427
rect 6009 12393 6043 12427
rect 6101 12393 6135 12427
rect 7573 12393 7607 12427
rect 10609 12393 10643 12427
rect 10977 12393 11011 12427
rect 11069 12393 11103 12427
rect 11805 12393 11839 12427
rect 12265 12393 12299 12427
rect 12725 12393 12759 12427
rect 13185 12393 13219 12427
rect 1409 12325 1443 12359
rect 1593 12325 1627 12359
rect 4537 12325 4571 12359
rect 9382 12325 9416 12359
rect 12633 12325 12667 12359
rect 2053 12257 2087 12291
rect 2513 12257 2547 12291
rect 4261 12257 4295 12291
rect 4896 12257 4930 12291
rect 7214 12257 7248 12291
rect 7481 12257 7515 12291
rect 8686 12257 8720 12291
rect 2329 12189 2363 12223
rect 2421 12189 2455 12223
rect 3065 12189 3099 12223
rect 3249 12189 3283 12223
rect 4629 12189 4663 12223
rect 8953 12189 8987 12223
rect 9137 12189 9171 12223
rect 11161 12189 11195 12223
rect 11897 12189 11931 12223
rect 12081 12189 12115 12223
rect 12817 12189 12851 12223
rect 2881 12121 2915 12155
rect 10517 12121 10551 12155
rect 11437 12053 11471 12087
rect 2421 11849 2455 11883
rect 3985 11849 4019 11883
rect 7941 11849 7975 11883
rect 11253 11849 11287 11883
rect 11713 11849 11747 11883
rect 12541 11849 12575 11883
rect 12725 11849 12759 11883
rect 13369 11849 13403 11883
rect 13093 11781 13127 11815
rect 1777 11713 1811 11747
rect 3065 11713 3099 11747
rect 3341 11713 3375 11747
rect 3525 11713 3559 11747
rect 4629 11713 4663 11747
rect 6469 11713 6503 11747
rect 9321 11713 9355 11747
rect 9965 11713 9999 11747
rect 10793 11713 10827 11747
rect 11345 11713 11379 11747
rect 12265 11713 12299 11747
rect 12909 11713 12943 11747
rect 2789 11645 2823 11679
rect 4905 11645 4939 11679
rect 5161 11645 5195 11679
rect 9054 11645 9088 11679
rect 9781 11645 9815 11679
rect 11069 11645 11103 11679
rect 1961 11577 1995 11611
rect 2881 11577 2915 11611
rect 4445 11577 4479 11611
rect 6714 11577 6748 11611
rect 10609 11577 10643 11611
rect 12081 11577 12115 11611
rect 1869 11509 1903 11543
rect 2329 11509 2363 11543
rect 3617 11509 3651 11543
rect 4077 11509 4111 11543
rect 4537 11509 4571 11543
rect 6285 11509 6319 11543
rect 7849 11509 7883 11543
rect 9413 11509 9447 11543
rect 9873 11509 9907 11543
rect 10241 11509 10275 11543
rect 10701 11509 10735 11543
rect 12173 11509 12207 11543
rect 1501 11305 1535 11339
rect 1869 11305 1903 11339
rect 3433 11305 3467 11339
rect 9137 11305 9171 11339
rect 9597 11305 9631 11339
rect 10333 11305 10367 11339
rect 11161 11305 11195 11339
rect 14197 11305 14231 11339
rect 14381 11305 14415 11339
rect 14749 11305 14783 11339
rect 14841 11305 14875 11339
rect 15301 11305 15335 11339
rect 1593 11237 1627 11271
rect 8042 11237 8076 11271
rect 11253 11237 11287 11271
rect 12817 11237 12851 11271
rect 12909 11237 12943 11271
rect 13829 11237 13863 11271
rect 2053 11169 2087 11203
rect 2513 11169 2547 11203
rect 3341 11169 3375 11203
rect 5109 11169 5143 11203
rect 6570 11169 6604 11203
rect 6837 11169 6871 11203
rect 8585 11169 8619 11203
rect 9505 11169 9539 11203
rect 10425 11169 10459 11203
rect 11989 11169 12023 11203
rect 2605 11101 2639 11135
rect 2789 11101 2823 11135
rect 3617 11101 3651 11135
rect 5365 11101 5399 11135
rect 8309 11101 8343 11135
rect 8861 11101 8895 11135
rect 9781 11101 9815 11135
rect 10609 11101 10643 11135
rect 11345 11101 11379 11135
rect 11713 11101 11747 11135
rect 11897 11101 11931 11135
rect 13001 11101 13035 11135
rect 13461 11101 13495 11135
rect 14933 11101 14967 11135
rect 2973 11033 3007 11067
rect 3985 11033 4019 11067
rect 5457 11033 5491 11067
rect 6929 11033 6963 11067
rect 12357 11033 12391 11067
rect 12449 11033 12483 11067
rect 13737 11033 13771 11067
rect 14105 11033 14139 11067
rect 14197 11033 14231 11067
rect 2145 10965 2179 10999
rect 9965 10965 9999 10999
rect 10793 10965 10827 10999
rect 13277 10965 13311 10999
rect 2513 10761 2547 10795
rect 3341 10761 3375 10795
rect 9413 10761 9447 10795
rect 10241 10761 10275 10795
rect 11069 10761 11103 10795
rect 11437 10761 11471 10795
rect 12541 10761 12575 10795
rect 14197 10761 14231 10795
rect 6285 10693 6319 10727
rect 9321 10693 9355 10727
rect 11253 10693 11287 10727
rect 1961 10625 1995 10659
rect 2789 10625 2823 10659
rect 2881 10625 2915 10659
rect 4905 10625 4939 10659
rect 9873 10625 9907 10659
rect 9965 10625 9999 10659
rect 10701 10625 10735 10659
rect 10885 10625 10919 10659
rect 11805 10625 11839 10659
rect 11989 10625 12023 10659
rect 13093 10625 13127 10659
rect 13461 10625 13495 10659
rect 14749 10625 14783 10659
rect 3433 10557 3467 10591
rect 6469 10557 6503 10591
rect 7941 10557 7975 10591
rect 10609 10557 10643 10591
rect 13737 10557 13771 10591
rect 14565 10557 14599 10591
rect 1593 10489 1627 10523
rect 2145 10489 2179 10523
rect 3700 10489 3734 10523
rect 5150 10489 5184 10523
rect 6714 10489 6748 10523
rect 8186 10489 8220 10523
rect 12081 10489 12115 10523
rect 12909 10489 12943 10523
rect 13645 10489 13679 10523
rect 15025 10489 15059 10523
rect 1501 10421 1535 10455
rect 2053 10421 2087 10455
rect 2973 10421 3007 10455
rect 4813 10421 4847 10455
rect 7849 10421 7883 10455
rect 9781 10421 9815 10455
rect 12449 10421 12483 10455
rect 13001 10421 13035 10455
rect 14105 10421 14139 10455
rect 14657 10421 14691 10455
rect 1869 10217 1903 10251
rect 2145 10217 2179 10251
rect 4353 10217 4387 10251
rect 8125 10217 8159 10251
rect 9137 10217 9171 10251
rect 9505 10217 9539 10251
rect 9597 10217 9631 10251
rect 10333 10217 10367 10251
rect 10701 10217 10735 10251
rect 11161 10217 11195 10251
rect 11621 10217 11655 10251
rect 11989 10217 12023 10251
rect 12449 10217 12483 10251
rect 12909 10217 12943 10251
rect 13277 10217 13311 10251
rect 13737 10217 13771 10251
rect 14841 10217 14875 10251
rect 4813 10149 4847 10183
rect 6898 10149 6932 10183
rect 8493 10149 8527 10183
rect 11253 10149 11287 10183
rect 12081 10149 12115 10183
rect 13645 10149 13679 10183
rect 2053 10081 2087 10115
rect 2513 10081 2547 10115
rect 3341 10081 3375 10115
rect 3433 10081 3467 10115
rect 4077 10081 4111 10115
rect 4721 10081 4755 10115
rect 5437 10081 5471 10115
rect 8585 10081 8619 10115
rect 12817 10081 12851 10115
rect 14105 10081 14139 10115
rect 14749 10081 14783 10115
rect 15485 10081 15519 10115
rect 2605 10013 2639 10047
rect 2789 10013 2823 10047
rect 3617 10013 3651 10047
rect 4997 10013 5031 10047
rect 5181 10013 5215 10047
rect 6653 10013 6687 10047
rect 8677 10013 8711 10047
rect 9781 10013 9815 10047
rect 10057 10013 10091 10047
rect 10241 10013 10275 10047
rect 11345 10013 11379 10047
rect 12173 10013 12207 10047
rect 13093 10013 13127 10047
rect 13829 10013 13863 10047
rect 14933 10013 14967 10047
rect 4261 9945 4295 9979
rect 8033 9945 8067 9979
rect 10793 9945 10827 9979
rect 14381 9945 14415 9979
rect 15669 9945 15703 9979
rect 1777 9877 1811 9911
rect 2973 9877 3007 9911
rect 3985 9877 4019 9911
rect 6561 9877 6595 9911
rect 15209 9877 15243 9911
rect 11529 9673 11563 9707
rect 11713 9673 11747 9707
rect 15209 9673 15243 9707
rect 2513 9605 2547 9639
rect 4813 9605 4847 9639
rect 6285 9605 6319 9639
rect 6469 9605 6503 9639
rect 9137 9605 9171 9639
rect 9321 9605 9355 9639
rect 11161 9605 11195 9639
rect 13369 9605 13403 9639
rect 1961 9537 1995 9571
rect 3249 9537 3283 9571
rect 3433 9537 3467 9571
rect 7021 9537 7055 9571
rect 7481 9537 7515 9571
rect 7757 9537 7791 9571
rect 12173 9537 12207 9571
rect 12357 9537 12391 9571
rect 12633 9537 12667 9571
rect 13921 9537 13955 9571
rect 14289 9537 14323 9571
rect 1409 9469 1443 9503
rect 2145 9469 2179 9503
rect 4905 9469 4939 9503
rect 5172 9469 5206 9503
rect 9413 9469 9447 9503
rect 11345 9469 11379 9503
rect 12081 9469 12115 9503
rect 12817 9469 12851 9503
rect 14565 9469 14599 9503
rect 15025 9469 15059 9503
rect 1593 9401 1627 9435
rect 2053 9401 2087 9435
rect 3700 9401 3734 9435
rect 8024 9401 8058 9435
rect 9658 9401 9692 9435
rect 11069 9401 11103 9435
rect 13829 9401 13863 9435
rect 15485 9401 15519 9435
rect 2605 9333 2639 9367
rect 2973 9333 3007 9367
rect 3065 9333 3099 9367
rect 6837 9333 6871 9367
rect 6929 9333 6963 9367
rect 7573 9333 7607 9367
rect 10793 9333 10827 9367
rect 12909 9333 12943 9367
rect 13277 9333 13311 9367
rect 13737 9333 13771 9367
rect 14473 9333 14507 9367
rect 14933 9333 14967 9367
rect 15301 9333 15335 9367
rect 1501 9129 1535 9163
rect 1869 9129 1903 9163
rect 2881 9129 2915 9163
rect 3341 9129 3375 9163
rect 3985 9129 4019 9163
rect 8861 9129 8895 9163
rect 10517 9129 10551 9163
rect 11345 9129 11379 9163
rect 11713 9129 11747 9163
rect 12173 9129 12207 9163
rect 13093 9129 13127 9163
rect 13553 9129 13587 9163
rect 14381 9129 14415 9163
rect 14749 9129 14783 9163
rect 5702 9061 5736 9095
rect 9382 9061 9416 9095
rect 1593 8993 1627 9027
rect 2053 8993 2087 9027
rect 2421 8993 2455 9027
rect 2513 8993 2547 9027
rect 3433 8993 3467 9027
rect 5109 8993 5143 9027
rect 8053 8993 8087 9027
rect 10977 8993 11011 9027
rect 11805 8993 11839 9027
rect 12633 8993 12667 9027
rect 13461 8993 13495 9027
rect 15393 8993 15427 9027
rect 2329 8925 2363 8959
rect 3617 8925 3651 8959
rect 5365 8925 5399 8959
rect 5457 8925 5491 8959
rect 8309 8925 8343 8959
rect 8585 8925 8619 8959
rect 9137 8925 9171 8959
rect 10701 8925 10735 8959
rect 10885 8925 10919 8959
rect 11529 8925 11563 8959
rect 12725 8925 12759 8959
rect 12909 8925 12943 8959
rect 13645 8925 13679 8959
rect 14841 8925 14875 8959
rect 14933 8925 14967 8959
rect 6837 8857 6871 8891
rect 12265 8857 12299 8891
rect 13921 8857 13955 8891
rect 15209 8857 15243 8891
rect 1777 8789 1811 8823
rect 2973 8789 3007 8823
rect 6929 8789 6963 8823
rect 14105 8789 14139 8823
rect 9873 8585 9907 8619
rect 11345 8585 11379 8619
rect 11529 8585 11563 8619
rect 11713 8585 11747 8619
rect 14933 8585 14967 8619
rect 2605 8517 2639 8551
rect 6285 8517 6319 8551
rect 8401 8517 8435 8551
rect 2237 8449 2271 8483
rect 2421 8449 2455 8483
rect 3249 8449 3283 8483
rect 3433 8449 3467 8483
rect 6469 8449 6503 8483
rect 9781 8449 9815 8483
rect 11253 8449 11287 8483
rect 2145 8381 2179 8415
rect 3700 8381 3734 8415
rect 4905 8381 4939 8415
rect 1409 8313 1443 8347
rect 1593 8313 1627 8347
rect 5172 8313 5206 8347
rect 12541 8517 12575 8551
rect 13369 8517 13403 8551
rect 15025 8517 15059 8551
rect 12265 8449 12299 8483
rect 13093 8449 13127 8483
rect 13921 8449 13955 8483
rect 14289 8449 14323 8483
rect 15209 8449 15243 8483
rect 12081 8381 12115 8415
rect 13001 8381 13035 8415
rect 13737 8381 13771 8415
rect 6561 8313 6595 8347
rect 8309 8313 8343 8347
rect 9536 8313 9570 8347
rect 10986 8313 11020 8347
rect 11529 8313 11563 8347
rect 12909 8313 12943 8347
rect 13829 8313 13863 8347
rect 14565 8313 14599 8347
rect 1777 8245 1811 8279
rect 2973 8245 3007 8279
rect 3065 8245 3099 8279
rect 4813 8245 4847 8279
rect 6469 8245 6503 8279
rect 12173 8245 12207 8279
rect 14473 8245 14507 8279
rect 1501 8041 1535 8075
rect 2881 8041 2915 8075
rect 3249 8041 3283 8075
rect 3893 8041 3927 8075
rect 7573 8041 7607 8075
rect 11805 8041 11839 8075
rect 11897 8041 11931 8075
rect 15117 8041 15151 8075
rect 1777 7973 1811 8007
rect 4169 7973 4203 8007
rect 10977 7973 11011 8007
rect 13461 7973 13495 8007
rect 14565 7973 14599 8007
rect 2053 7905 2087 7939
rect 2421 7905 2455 7939
rect 2513 7905 2547 7939
rect 3341 7905 3375 7939
rect 4077 7905 4111 7939
rect 4353 7905 4387 7939
rect 4885 7905 4919 7939
rect 7214 7905 7248 7939
rect 8686 7905 8720 7939
rect 8953 7905 8987 7939
rect 10250 7905 10284 7939
rect 12633 7905 12667 7939
rect 13553 7905 13587 7939
rect 14381 7905 14415 7939
rect 2329 7837 2363 7871
rect 3065 7837 3099 7871
rect 4629 7837 4663 7871
rect 7481 7837 7515 7871
rect 10517 7837 10551 7871
rect 11069 7837 11103 7871
rect 11161 7837 11195 7871
rect 11989 7837 12023 7871
rect 12725 7837 12759 7871
rect 12909 7837 12943 7871
rect 13645 7837 13679 7871
rect 12265 7769 12299 7803
rect 1869 7701 1903 7735
rect 3709 7701 3743 7735
rect 4537 7701 4571 7735
rect 6009 7701 6043 7735
rect 6101 7701 6135 7735
rect 9137 7701 9171 7735
rect 10609 7701 10643 7735
rect 11437 7701 11471 7735
rect 13093 7701 13127 7735
rect 14013 7701 14047 7735
rect 14197 7701 14231 7735
rect 14749 7701 14783 7735
rect 14933 7701 14967 7735
rect 3341 7497 3375 7531
rect 11437 7497 11471 7531
rect 13369 7497 13403 7531
rect 2513 7429 2547 7463
rect 6285 7429 6319 7463
rect 10793 7429 10827 7463
rect 11069 7429 11103 7463
rect 1409 7361 1443 7395
rect 1961 7361 1995 7395
rect 2789 7361 2823 7395
rect 9413 7361 9447 7395
rect 12173 7361 12207 7395
rect 12265 7361 12299 7395
rect 13093 7361 13127 7395
rect 13921 7361 13955 7395
rect 1593 7293 1627 7327
rect 2053 7293 2087 7327
rect 3433 7293 3467 7327
rect 4905 7293 4939 7327
rect 7849 7293 7883 7327
rect 7941 7293 7975 7327
rect 10885 7293 10919 7327
rect 11161 7293 11195 7327
rect 13737 7293 13771 7327
rect 14565 7293 14599 7327
rect 3700 7225 3734 7259
rect 5172 7225 5206 7259
rect 7582 7225 7616 7259
rect 8208 7225 8242 7259
rect 9680 7225 9714 7259
rect 2145 7157 2179 7191
rect 2881 7157 2915 7191
rect 2973 7157 3007 7191
rect 4813 7157 4847 7191
rect 6469 7157 6503 7191
rect 9321 7157 9355 7191
rect 11345 7157 11379 7191
rect 11713 7157 11747 7191
rect 12081 7157 12115 7191
rect 12541 7157 12575 7191
rect 12909 7157 12943 7191
rect 13001 7157 13035 7191
rect 13829 7157 13863 7191
rect 14197 7157 14231 7191
rect 14381 7157 14415 7191
rect 1593 6953 1627 6987
rect 4721 6953 4755 6987
rect 12265 6953 12299 6987
rect 13093 6953 13127 6987
rect 13553 6953 13587 6987
rect 13737 6953 13771 6987
rect 2513 6885 2547 6919
rect 3341 6885 3375 6919
rect 4813 6885 4847 6919
rect 8493 6885 8527 6919
rect 11437 6885 11471 6919
rect 11529 6885 11563 6919
rect 12357 6885 12391 6919
rect 14381 6885 14415 6919
rect 14565 6885 14599 6919
rect 1685 6817 1719 6851
rect 2053 6817 2087 6851
rect 4261 6817 4295 6851
rect 6294 6817 6328 6851
rect 6561 6817 6595 6851
rect 7766 6817 7800 6851
rect 8033 6817 8067 6851
rect 8585 6817 8619 6851
rect 9965 6817 9999 6851
rect 10609 6817 10643 6851
rect 10701 6817 10735 6851
rect 13185 6817 13219 6851
rect 2237 6749 2271 6783
rect 2421 6749 2455 6783
rect 3433 6749 3467 6783
rect 3617 6749 3651 6783
rect 4997 6749 5031 6783
rect 8677 6749 8711 6783
rect 9413 6749 9447 6783
rect 10793 6749 10827 6783
rect 11713 6749 11747 6783
rect 12449 6749 12483 6783
rect 13277 6749 13311 6783
rect 2973 6681 3007 6715
rect 4077 6681 4111 6715
rect 6653 6681 6687 6715
rect 11897 6681 11931 6715
rect 13921 6681 13955 6715
rect 1869 6613 1903 6647
rect 2881 6613 2915 6647
rect 3893 6613 3927 6647
rect 4353 6613 4387 6647
rect 5181 6613 5215 6647
rect 8125 6613 8159 6647
rect 10241 6613 10275 6647
rect 11069 6613 11103 6647
rect 12725 6613 12759 6647
rect 14197 6613 14231 6647
rect 14749 6613 14783 6647
rect 1501 6409 1535 6443
rect 2513 6409 2547 6443
rect 3433 6409 3467 6443
rect 4905 6409 4939 6443
rect 7849 6409 7883 6443
rect 9413 6341 9447 6375
rect 1961 6273 1995 6307
rect 2053 6273 2087 6307
rect 3249 6273 3283 6307
rect 11345 6273 11379 6307
rect 12357 6273 12391 6307
rect 13093 6273 13127 6307
rect 13921 6273 13955 6307
rect 14381 6273 14415 6307
rect 1593 6205 1627 6239
rect 4813 6205 4847 6239
rect 6285 6205 6319 6239
rect 6469 6205 6503 6239
rect 9321 6205 9355 6239
rect 10793 6205 10827 6239
rect 11069 6205 11103 6239
rect 13737 6205 13771 6239
rect 4568 6137 4602 6171
rect 6040 6137 6074 6171
rect 6714 6137 6748 6171
rect 9054 6137 9088 6171
rect 10526 6137 10560 6171
rect 11437 6137 11471 6171
rect 12173 6137 12207 6171
rect 12909 6137 12943 6171
rect 14197 6137 14231 6171
rect 2145 6069 2179 6103
rect 2605 6069 2639 6103
rect 2973 6069 3007 6103
rect 3065 6069 3099 6103
rect 7941 6069 7975 6103
rect 11713 6069 11747 6103
rect 12081 6069 12115 6103
rect 12541 6069 12575 6103
rect 13001 6069 13035 6103
rect 13369 6069 13403 6103
rect 13829 6069 13863 6103
rect 2881 5865 2915 5899
rect 3249 5865 3283 5899
rect 4077 5865 4111 5899
rect 5181 5865 5215 5899
rect 8677 5865 8711 5899
rect 10517 5865 10551 5899
rect 11897 5865 11931 5899
rect 12633 5865 12667 5899
rect 13369 5865 13403 5899
rect 1501 5797 1535 5831
rect 4813 5797 4847 5831
rect 9382 5797 9416 5831
rect 10977 5797 11011 5831
rect 11069 5797 11103 5831
rect 12725 5797 12759 5831
rect 13093 5797 13127 5831
rect 13553 5797 13587 5831
rect 13737 5797 13771 5831
rect 13921 5797 13955 5831
rect 2053 5729 2087 5763
rect 2513 5729 2547 5763
rect 3341 5729 3375 5763
rect 3893 5729 3927 5763
rect 5273 5729 5307 5763
rect 5540 5729 5574 5763
rect 7858 5729 7892 5763
rect 8585 5729 8619 5763
rect 9137 5729 9171 5763
rect 11805 5729 11839 5763
rect 2329 5661 2363 5695
rect 2421 5661 2455 5695
rect 3157 5661 3191 5695
rect 4353 5661 4387 5695
rect 4629 5661 4663 5695
rect 4721 5661 4755 5695
rect 8125 5661 8159 5695
rect 8769 5661 8803 5695
rect 11253 5661 11287 5695
rect 11989 5661 12023 5695
rect 12817 5661 12851 5695
rect 3709 5593 3743 5627
rect 6745 5593 6779 5627
rect 10609 5593 10643 5627
rect 11437 5593 11471 5627
rect 12265 5593 12299 5627
rect 1685 5525 1719 5559
rect 1869 5525 1903 5559
rect 6653 5525 6687 5559
rect 8217 5525 8251 5559
rect 14013 5525 14047 5559
rect 1501 5321 1535 5355
rect 3341 5321 3375 5355
rect 10241 5321 10275 5355
rect 12909 5321 12943 5355
rect 13277 5321 13311 5355
rect 3433 5253 3467 5287
rect 7941 5253 7975 5287
rect 13553 5253 13587 5287
rect 1961 5185 1995 5219
rect 2053 5185 2087 5219
rect 2789 5185 2823 5219
rect 4813 5185 4847 5219
rect 9873 5185 9907 5219
rect 9965 5185 9999 5219
rect 10793 5185 10827 5219
rect 11529 5185 11563 5219
rect 12265 5185 12299 5219
rect 1593 5117 1627 5151
rect 2973 5117 3007 5151
rect 6285 5117 6319 5151
rect 6469 5117 6503 5151
rect 9054 5117 9088 5151
rect 9321 5117 9355 5151
rect 9781 5117 9815 5151
rect 12081 5117 12115 5151
rect 12173 5117 12207 5151
rect 2145 5049 2179 5083
rect 4568 5049 4602 5083
rect 6040 5049 6074 5083
rect 6714 5049 6748 5083
rect 10609 5049 10643 5083
rect 10701 5049 10735 5083
rect 11069 5049 11103 5083
rect 11253 5049 11287 5083
rect 12633 5049 12667 5083
rect 2513 4981 2547 5015
rect 2881 4981 2915 5015
rect 4905 4981 4939 5015
rect 7849 4981 7883 5015
rect 9413 4981 9447 5015
rect 11713 4981 11747 5015
rect 12725 4981 12759 5015
rect 13093 4981 13127 5015
rect 13645 4981 13679 5015
rect 2145 4777 2179 4811
rect 2973 4777 3007 4811
rect 4813 4777 4847 4811
rect 4905 4777 4939 4811
rect 9597 4777 9631 4811
rect 10425 4777 10459 4811
rect 11713 4777 11747 4811
rect 13001 4777 13035 4811
rect 13461 4777 13495 4811
rect 14105 4777 14139 4811
rect 1593 4709 1627 4743
rect 10333 4709 10367 4743
rect 11069 4709 11103 4743
rect 12173 4709 12207 4743
rect 1777 4641 1811 4675
rect 2329 4641 2363 4675
rect 2605 4641 2639 4675
rect 2881 4641 2915 4675
rect 3341 4641 3375 4675
rect 4169 4641 4203 4675
rect 4445 4641 4479 4675
rect 6478 4641 6512 4675
rect 6745 4641 6779 4675
rect 7961 4641 7995 4675
rect 8769 4641 8803 4675
rect 9505 4641 9539 4675
rect 11161 4641 11195 4675
rect 11805 4641 11839 4675
rect 12541 4641 12575 4675
rect 13645 4641 13679 4675
rect 13829 4641 13863 4675
rect 3433 4573 3467 4607
rect 3617 4573 3651 4607
rect 4721 4573 4755 4607
rect 8217 4573 8251 4607
rect 8493 4573 8527 4607
rect 9689 4573 9723 4607
rect 10517 4573 10551 4607
rect 10885 4573 10919 4607
rect 2697 4505 2731 4539
rect 9137 4505 9171 4539
rect 9965 4505 9999 4539
rect 11529 4505 11563 4539
rect 11989 4505 12023 4539
rect 12725 4505 12759 4539
rect 13277 4505 13311 4539
rect 1501 4437 1535 4471
rect 1961 4437 1995 4471
rect 2421 4437 2455 4471
rect 3985 4437 4019 4471
rect 5273 4437 5307 4471
rect 5365 4437 5399 4471
rect 6837 4437 6871 4471
rect 8861 4437 8895 4471
rect 12449 4437 12483 4471
rect 13093 4437 13127 4471
rect 3893 4233 3927 4267
rect 4721 4233 4755 4267
rect 7849 4233 7883 4267
rect 7941 4233 7975 4267
rect 10425 4233 10459 4267
rect 12265 4233 12299 4267
rect 12541 4233 12575 4267
rect 12817 4233 12851 4267
rect 13553 4233 13587 4267
rect 14289 4233 14323 4267
rect 14473 4233 14507 4267
rect 2697 4165 2731 4199
rect 10977 4165 11011 4199
rect 11345 4165 11379 4199
rect 11989 4165 12023 4199
rect 13737 4165 13771 4199
rect 13921 4165 13955 4199
rect 14105 4165 14139 4199
rect 14657 4165 14691 4199
rect 3525 4097 3559 4131
rect 3709 4097 3743 4131
rect 4353 4097 4387 4131
rect 4537 4097 4571 4131
rect 5273 4097 5307 4131
rect 6101 4097 6135 4131
rect 8585 4097 8619 4131
rect 9321 4097 9355 4131
rect 10057 4097 10091 4131
rect 10149 4097 10183 4131
rect 13277 4097 13311 4131
rect 13461 4097 13495 4131
rect 1593 4029 1627 4063
rect 2237 4029 2271 4063
rect 2513 4029 2547 4063
rect 2789 4029 2823 4063
rect 6476 4029 6510 4063
rect 6725 4029 6759 4063
rect 8309 4029 8343 4063
rect 10609 4029 10643 4063
rect 10885 4029 10919 4063
rect 11153 4029 11187 4063
rect 12081 4029 12115 4063
rect 15485 4029 15519 4063
rect 1961 3961 1995 3995
rect 8401 3961 8435 3995
rect 9137 3961 9171 3995
rect 9965 3961 9999 3995
rect 12633 3961 12667 3995
rect 13001 3961 13035 3995
rect 1501 3893 1535 3927
rect 1869 3893 1903 3927
rect 2421 3893 2455 3927
rect 2973 3893 3007 3927
rect 3065 3893 3099 3927
rect 3433 3893 3467 3927
rect 4261 3893 4295 3927
rect 5089 3893 5123 3927
rect 5181 3893 5215 3927
rect 5549 3893 5583 3927
rect 5917 3893 5951 3927
rect 6009 3893 6043 3927
rect 8769 3893 8803 3927
rect 9229 3893 9263 3927
rect 9597 3893 9631 3927
rect 10701 3893 10735 3927
rect 11437 3893 11471 3927
rect 11713 3893 11747 3927
rect 15117 3893 15151 3927
rect 15301 3893 15335 3927
rect 15669 3893 15703 3927
rect 2145 3689 2179 3723
rect 3893 3689 3927 3723
rect 4353 3689 4387 3723
rect 4721 3689 4755 3723
rect 5181 3689 5215 3723
rect 5825 3689 5859 3723
rect 7021 3689 7055 3723
rect 7849 3689 7883 3723
rect 10701 3689 10735 3723
rect 11069 3689 11103 3723
rect 11713 3689 11747 3723
rect 15117 3689 15151 3723
rect 1961 3621 1995 3655
rect 8309 3621 8343 3655
rect 9597 3621 9631 3655
rect 11621 3621 11655 3655
rect 12173 3621 12207 3655
rect 13921 3621 13955 3655
rect 15485 3621 15519 3655
rect 1593 3553 1627 3587
rect 2329 3553 2363 3587
rect 2605 3553 2639 3587
rect 2881 3553 2915 3587
rect 3157 3553 3191 3587
rect 3433 3553 3467 3587
rect 3709 3553 3743 3587
rect 4261 3553 4295 3587
rect 5089 3553 5123 3587
rect 5733 3553 5767 3587
rect 6193 3553 6227 3587
rect 8493 3553 8527 3587
rect 9505 3553 9539 3587
rect 10149 3553 10183 3587
rect 10241 3553 10275 3587
rect 10517 3553 10551 3587
rect 10793 3553 10827 3587
rect 11244 3553 11278 3587
rect 11897 3553 11931 3587
rect 13369 3553 13403 3587
rect 13553 3553 13587 3587
rect 13829 3553 13863 3587
rect 14749 3553 14783 3587
rect 14841 3553 14875 3587
rect 15301 3553 15335 3587
rect 4537 3485 4571 3519
rect 5273 3485 5307 3519
rect 6285 3485 6319 3519
rect 6377 3485 6411 3519
rect 6745 3485 6779 3519
rect 6929 3485 6963 3519
rect 7941 3485 7975 3519
rect 8125 3485 8159 3519
rect 8677 3485 8711 3519
rect 9781 3485 9815 3519
rect 12909 3485 12943 3519
rect 1409 3417 1443 3451
rect 2697 3417 2731 3451
rect 3249 3417 3283 3451
rect 5549 3417 5583 3451
rect 7389 3417 7423 3451
rect 9965 3417 9999 3451
rect 11345 3417 11379 3451
rect 14105 3417 14139 3451
rect 14565 3417 14599 3451
rect 15025 3417 15059 3451
rect 15669 3417 15703 3451
rect 1869 3349 1903 3383
rect 2421 3349 2455 3383
rect 2973 3349 3007 3383
rect 3525 3349 3559 3383
rect 7481 3349 7515 3383
rect 9137 3349 9171 3383
rect 10425 3349 10459 3383
rect 10977 3349 11011 3383
rect 12449 3349 12483 3383
rect 12633 3349 12667 3383
rect 13093 3349 13127 3383
rect 13185 3349 13219 3383
rect 14473 3349 14507 3383
rect 4721 3145 4755 3179
rect 6469 3145 6503 3179
rect 7297 3145 7331 3179
rect 9045 3145 9079 3179
rect 10793 3145 10827 3179
rect 11897 3145 11931 3179
rect 12081 3145 12115 3179
rect 12449 3145 12483 3179
rect 14105 3145 14139 3179
rect 2145 3077 2179 3111
rect 3249 3077 3283 3111
rect 5549 3077 5583 3111
rect 11345 3077 11379 3111
rect 3617 3009 3651 3043
rect 5273 3009 5307 3043
rect 6193 3009 6227 3043
rect 6929 3009 6963 3043
rect 7021 3009 7055 3043
rect 7757 3009 7791 3043
rect 7849 3009 7883 3043
rect 8677 3009 8711 3043
rect 9321 3009 9355 3043
rect 12725 3009 12759 3043
rect 15209 3009 15243 3043
rect 1593 2941 1627 2975
rect 1961 2941 1995 2975
rect 2329 2941 2363 2975
rect 2697 2941 2731 2975
rect 3985 2941 4019 2975
rect 4169 2941 4203 2975
rect 4445 2941 4479 2975
rect 5917 2941 5951 2975
rect 6837 2941 6871 2975
rect 7665 2941 7699 2975
rect 8493 2941 8527 2975
rect 9137 2941 9171 2975
rect 9873 2941 9907 2975
rect 10149 2941 10183 2975
rect 10417 2941 10451 2975
rect 10525 2941 10559 2975
rect 10977 2941 11011 2975
rect 11253 2941 11287 2975
rect 11529 2941 11563 2975
rect 11713 2941 11747 2975
rect 12265 2941 12299 2975
rect 12633 2941 12667 2975
rect 13093 2941 13127 2975
rect 13553 2941 13587 2975
rect 14280 2941 14314 2975
rect 14389 2941 14423 2975
rect 14657 2941 14691 2975
rect 15117 2941 15151 2975
rect 1409 2873 1443 2907
rect 2881 2873 2915 2907
rect 3065 2873 3099 2907
rect 3433 2873 3467 2907
rect 3801 2873 3835 2907
rect 4629 2873 4663 2907
rect 5089 2873 5123 2907
rect 5181 2873 5215 2907
rect 9505 2873 9539 2907
rect 12909 2873 12943 2907
rect 13737 2873 13771 2907
rect 15485 2873 15519 2907
rect 15669 2873 15703 2907
rect 1869 2805 1903 2839
rect 2605 2805 2639 2839
rect 6009 2805 6043 2839
rect 8125 2805 8159 2839
rect 8585 2805 8619 2839
rect 9689 2805 9723 2839
rect 9965 2805 9999 2839
rect 10241 2805 10275 2839
rect 10701 2805 10735 2839
rect 11069 2805 11103 2839
rect 13277 2805 13311 2839
rect 13921 2805 13955 2839
rect 14565 2805 14599 2839
rect 14841 2805 14875 2839
rect 14933 2805 14967 2839
rect 5365 2601 5399 2635
rect 5641 2601 5675 2635
rect 6561 2601 6595 2635
rect 7021 2601 7055 2635
rect 7389 2601 7423 2635
rect 9689 2601 9723 2635
rect 9965 2601 9999 2635
rect 11529 2601 11563 2635
rect 12909 2601 12943 2635
rect 13277 2601 13311 2635
rect 14381 2601 14415 2635
rect 1593 2533 1627 2567
rect 4445 2533 4479 2567
rect 7757 2533 7791 2567
rect 7849 2533 7883 2567
rect 11345 2533 11379 2567
rect 12449 2533 12483 2567
rect 14749 2533 14783 2567
rect 15485 2533 15519 2567
rect 2053 2465 2087 2499
rect 2585 2465 2619 2499
rect 3893 2465 3927 2499
rect 4077 2465 4111 2499
rect 4813 2465 4847 2499
rect 5181 2465 5215 2499
rect 5549 2465 5583 2499
rect 6009 2465 6043 2499
rect 6929 2465 6963 2499
rect 8493 2465 8527 2499
rect 8861 2465 8895 2499
rect 9505 2465 9539 2499
rect 9873 2465 9907 2499
rect 9965 2465 9999 2499
rect 10241 2465 10275 2499
rect 10609 2465 10643 2499
rect 10977 2465 11011 2499
rect 11713 2465 11747 2499
rect 12081 2465 12115 2499
rect 13001 2465 13035 2499
rect 13369 2465 13403 2499
rect 13737 2465 13771 2499
rect 13921 2465 13955 2499
rect 14197 2465 14231 2499
rect 15117 2465 15151 2499
rect 2329 2397 2363 2431
rect 6101 2397 6135 2431
rect 6285 2397 6319 2431
rect 7205 2397 7239 2431
rect 7941 2397 7975 2431
rect 12633 2397 12667 2431
rect 14933 2397 14967 2431
rect 1409 2329 1443 2363
rect 1869 2329 1903 2363
rect 4261 2329 4295 2363
rect 4997 2329 5031 2363
rect 8953 2329 8987 2363
rect 10793 2329 10827 2363
rect 11897 2329 11931 2363
rect 13553 2329 13587 2363
rect 14105 2329 14139 2363
rect 15301 2329 15335 2363
rect 2145 2261 2179 2295
rect 3709 2261 3743 2295
rect 4721 2261 4755 2295
rect 8309 2261 8343 2295
rect 8677 2261 8711 2295
rect 9321 2261 9355 2295
rect 10149 2261 10183 2295
rect 10517 2261 10551 2295
rect 11253 2261 11287 2295
rect 12357 2261 12391 2295
rect 15577 2261 15611 2295
<< metal1 >>
rect 8386 17620 8392 17672
rect 8444 17660 8450 17672
rect 8846 17660 8852 17672
rect 8444 17632 8852 17660
rect 8444 17620 8450 17632
rect 8846 17620 8852 17632
rect 8904 17620 8910 17672
rect 1104 17434 16008 17456
rect 1104 17382 3480 17434
rect 3532 17382 3544 17434
rect 3596 17382 3608 17434
rect 3660 17382 3672 17434
rect 3724 17382 8478 17434
rect 8530 17382 8542 17434
rect 8594 17382 8606 17434
rect 8658 17382 8670 17434
rect 8722 17382 13475 17434
rect 13527 17382 13539 17434
rect 13591 17382 13603 17434
rect 13655 17382 13667 17434
rect 13719 17382 16008 17434
rect 1104 17360 16008 17382
rect 2501 17323 2559 17329
rect 2501 17289 2513 17323
rect 2547 17320 2559 17323
rect 2774 17320 2780 17332
rect 2547 17292 2780 17320
rect 2547 17289 2559 17292
rect 2501 17283 2559 17289
rect 2774 17280 2780 17292
rect 2832 17280 2838 17332
rect 2869 17323 2927 17329
rect 2869 17289 2881 17323
rect 2915 17289 2927 17323
rect 2869 17283 2927 17289
rect 2038 17252 2044 17264
rect 1999 17224 2044 17252
rect 2038 17212 2044 17224
rect 2096 17212 2102 17264
rect 2406 17212 2412 17264
rect 2464 17252 2470 17264
rect 2884 17252 2912 17283
rect 3142 17280 3148 17332
rect 3200 17320 3206 17332
rect 3973 17323 4031 17329
rect 3973 17320 3985 17323
rect 3200 17292 3985 17320
rect 3200 17280 3206 17292
rect 3973 17289 3985 17292
rect 4019 17289 4031 17323
rect 3973 17283 4031 17289
rect 4154 17280 4160 17332
rect 4212 17320 4218 17332
rect 4709 17323 4767 17329
rect 4709 17320 4721 17323
rect 4212 17292 4721 17320
rect 4212 17280 4218 17292
rect 4709 17289 4721 17292
rect 4755 17289 4767 17323
rect 4709 17283 4767 17289
rect 5905 17323 5963 17329
rect 5905 17289 5917 17323
rect 5951 17320 5963 17323
rect 9490 17320 9496 17332
rect 5951 17292 8524 17320
rect 5951 17289 5963 17292
rect 5905 17283 5963 17289
rect 3513 17255 3571 17261
rect 3513 17252 3525 17255
rect 2464 17224 2912 17252
rect 3252 17224 3525 17252
rect 2464 17212 2470 17224
rect 2774 17184 2780 17196
rect 2424 17156 2780 17184
rect 2424 17128 2452 17156
rect 2774 17144 2780 17156
rect 2832 17144 2838 17196
rect 2866 17144 2872 17196
rect 2924 17184 2930 17196
rect 3145 17187 3203 17193
rect 3145 17184 3157 17187
rect 2924 17156 3157 17184
rect 2924 17144 2930 17156
rect 3145 17153 3157 17156
rect 3191 17153 3203 17187
rect 3145 17147 3203 17153
rect 1394 17116 1400 17128
rect 1355 17088 1400 17116
rect 1394 17076 1400 17088
rect 1452 17076 1458 17128
rect 1673 17119 1731 17125
rect 1673 17085 1685 17119
rect 1719 17116 1731 17119
rect 2130 17116 2136 17128
rect 1719 17088 2136 17116
rect 1719 17085 1731 17088
rect 1673 17079 1731 17085
rect 2130 17076 2136 17088
rect 2188 17076 2194 17128
rect 2406 17076 2412 17128
rect 2464 17076 2470 17128
rect 3252 17116 3280 17224
rect 3513 17221 3525 17224
rect 3559 17221 3571 17255
rect 3513 17215 3571 17221
rect 3786 17212 3792 17264
rect 3844 17252 3850 17264
rect 4249 17255 4307 17261
rect 4249 17252 4261 17255
rect 3844 17224 4261 17252
rect 3844 17212 3850 17224
rect 4249 17221 4261 17224
rect 4295 17221 4307 17255
rect 4249 17215 4307 17221
rect 4338 17212 4344 17264
rect 4396 17252 4402 17264
rect 4985 17255 5043 17261
rect 4985 17252 4997 17255
rect 4396 17224 4997 17252
rect 4396 17212 4402 17224
rect 4985 17221 4997 17224
rect 5031 17221 5043 17255
rect 4985 17215 5043 17221
rect 6178 17212 6184 17264
rect 6236 17252 6242 17264
rect 6549 17255 6607 17261
rect 6549 17252 6561 17255
rect 6236 17224 6561 17252
rect 6236 17212 6242 17224
rect 6549 17221 6561 17224
rect 6595 17221 6607 17255
rect 6549 17215 6607 17221
rect 6914 17212 6920 17264
rect 6972 17252 6978 17264
rect 7285 17255 7343 17261
rect 7285 17252 7297 17255
rect 6972 17224 7297 17252
rect 6972 17212 6978 17224
rect 7285 17221 7297 17224
rect 7331 17221 7343 17255
rect 7285 17215 7343 17221
rect 7650 17212 7656 17264
rect 7708 17252 7714 17264
rect 8021 17255 8079 17261
rect 8021 17252 8033 17255
rect 7708 17224 8033 17252
rect 7708 17212 7714 17224
rect 8021 17221 8033 17224
rect 8067 17221 8079 17255
rect 8021 17215 8079 17221
rect 8294 17212 8300 17264
rect 8352 17252 8358 17264
rect 8389 17255 8447 17261
rect 8389 17252 8401 17255
rect 8352 17224 8401 17252
rect 8352 17212 8358 17224
rect 8389 17221 8401 17224
rect 8435 17221 8447 17255
rect 8496 17252 8524 17292
rect 8864 17292 9496 17320
rect 8864 17252 8892 17292
rect 9490 17280 9496 17292
rect 9548 17280 9554 17332
rect 13814 17280 13820 17332
rect 13872 17320 13878 17332
rect 14185 17323 14243 17329
rect 14185 17320 14197 17323
rect 13872 17292 14197 17320
rect 13872 17280 13878 17292
rect 14185 17289 14197 17292
rect 14231 17289 14243 17323
rect 14185 17283 14243 17289
rect 14642 17280 14648 17332
rect 14700 17320 14706 17332
rect 14737 17323 14795 17329
rect 14737 17320 14749 17323
rect 14700 17292 14749 17320
rect 14700 17280 14706 17292
rect 14737 17289 14749 17292
rect 14783 17289 14795 17323
rect 14737 17283 14795 17289
rect 8496 17224 8892 17252
rect 8389 17215 8447 17221
rect 8938 17212 8944 17264
rect 8996 17252 9002 17264
rect 9217 17255 9275 17261
rect 9217 17252 9229 17255
rect 8996 17224 9229 17252
rect 8996 17212 9002 17224
rect 9217 17221 9229 17224
rect 9263 17221 9275 17255
rect 9217 17215 9275 17221
rect 4154 17184 4160 17196
rect 2746 17088 3280 17116
rect 3344 17156 4160 17184
rect 2222 17048 2228 17060
rect 2183 17020 2228 17048
rect 2222 17008 2228 17020
rect 2280 17008 2286 17060
rect 2593 17051 2651 17057
rect 2593 17017 2605 17051
rect 2639 17017 2651 17051
rect 2593 17011 2651 17017
rect 2608 16980 2636 17011
rect 2746 16980 2774 17088
rect 2958 17048 2964 17060
rect 2919 17020 2964 17048
rect 2958 17008 2964 17020
rect 3016 17008 3022 17060
rect 3344 17057 3372 17156
rect 4154 17144 4160 17156
rect 4212 17144 4218 17196
rect 4614 17144 4620 17196
rect 4672 17184 4678 17196
rect 5353 17187 5411 17193
rect 5353 17184 5365 17187
rect 4672 17156 5365 17184
rect 4672 17144 4678 17156
rect 5353 17153 5365 17156
rect 5399 17153 5411 17187
rect 5353 17147 5411 17153
rect 6365 17187 6423 17193
rect 6365 17153 6377 17187
rect 6411 17184 6423 17187
rect 9030 17184 9036 17196
rect 6411 17156 9036 17184
rect 6411 17153 6423 17156
rect 6365 17147 6423 17153
rect 9030 17144 9036 17156
rect 9088 17144 9094 17196
rect 12253 17187 12311 17193
rect 12253 17184 12265 17187
rect 11532 17156 12265 17184
rect 3697 17119 3755 17125
rect 3697 17085 3709 17119
rect 3743 17116 3755 17119
rect 3786 17116 3792 17128
rect 3743 17088 3792 17116
rect 3743 17085 3755 17088
rect 3697 17079 3755 17085
rect 3786 17076 3792 17088
rect 3844 17076 3850 17128
rect 6546 17076 6552 17128
rect 6604 17116 6610 17128
rect 6917 17119 6975 17125
rect 6917 17116 6929 17119
rect 6604 17088 6929 17116
rect 6604 17076 6610 17088
rect 6917 17085 6929 17088
rect 6963 17085 6975 17119
rect 6917 17079 6975 17085
rect 7282 17076 7288 17128
rect 7340 17116 7346 17128
rect 7653 17119 7711 17125
rect 7653 17116 7665 17119
rect 7340 17088 7665 17116
rect 7340 17076 7346 17088
rect 7653 17085 7665 17088
rect 7699 17085 7711 17119
rect 7653 17079 7711 17085
rect 7837 17119 7895 17125
rect 7837 17085 7849 17119
rect 7883 17116 7895 17119
rect 8478 17116 8484 17128
rect 7883 17088 8484 17116
rect 7883 17085 7895 17088
rect 7837 17079 7895 17085
rect 8478 17076 8484 17088
rect 8536 17076 8542 17128
rect 8573 17119 8631 17125
rect 8573 17085 8585 17119
rect 8619 17116 8631 17119
rect 9122 17116 9128 17128
rect 8619 17088 9128 17116
rect 8619 17085 8631 17088
rect 8573 17079 8631 17085
rect 9122 17076 9128 17088
rect 9180 17076 9186 17128
rect 9858 17076 9864 17128
rect 9916 17116 9922 17128
rect 10137 17119 10195 17125
rect 10137 17116 10149 17119
rect 9916 17088 10149 17116
rect 9916 17076 9922 17088
rect 10137 17085 10149 17088
rect 10183 17085 10195 17119
rect 10137 17079 10195 17085
rect 10226 17076 10232 17128
rect 10284 17116 10290 17128
rect 10505 17119 10563 17125
rect 10505 17116 10517 17119
rect 10284 17088 10517 17116
rect 10284 17076 10290 17088
rect 10505 17085 10517 17088
rect 10551 17116 10563 17119
rect 10594 17116 10600 17128
rect 10551 17088 10600 17116
rect 10551 17085 10563 17088
rect 10505 17079 10563 17085
rect 10594 17076 10600 17088
rect 10652 17076 10658 17128
rect 10686 17076 10692 17128
rect 10744 17116 10750 17128
rect 10873 17119 10931 17125
rect 10873 17116 10885 17119
rect 10744 17088 10885 17116
rect 10744 17076 10750 17088
rect 10873 17085 10885 17088
rect 10919 17085 10931 17119
rect 10873 17079 10931 17085
rect 11054 17076 11060 17128
rect 11112 17116 11118 17128
rect 11241 17119 11299 17125
rect 11241 17116 11253 17119
rect 11112 17088 11253 17116
rect 11112 17076 11118 17088
rect 11241 17085 11253 17088
rect 11287 17116 11299 17119
rect 11330 17116 11336 17128
rect 11287 17088 11336 17116
rect 11287 17085 11299 17088
rect 11241 17079 11299 17085
rect 11330 17076 11336 17088
rect 11388 17076 11394 17128
rect 11422 17076 11428 17128
rect 11480 17116 11486 17128
rect 11532 17125 11560 17156
rect 12253 17153 12265 17156
rect 12299 17153 12311 17187
rect 12253 17147 12311 17153
rect 12894 17144 12900 17196
rect 12952 17184 12958 17196
rect 13725 17187 13783 17193
rect 13725 17184 13737 17187
rect 12952 17156 13737 17184
rect 12952 17144 12958 17156
rect 13725 17153 13737 17156
rect 13771 17153 13783 17187
rect 13725 17147 13783 17153
rect 14734 17144 14740 17196
rect 14792 17184 14798 17196
rect 14792 17156 15516 17184
rect 14792 17144 14798 17156
rect 11517 17119 11575 17125
rect 11517 17116 11529 17119
rect 11480 17088 11529 17116
rect 11480 17076 11486 17088
rect 11517 17085 11529 17088
rect 11563 17085 11575 17119
rect 11517 17079 11575 17085
rect 11790 17076 11796 17128
rect 11848 17116 11854 17128
rect 11977 17119 12035 17125
rect 11977 17116 11989 17119
rect 11848 17088 11989 17116
rect 11848 17076 11854 17088
rect 11977 17085 11989 17088
rect 12023 17085 12035 17119
rect 11977 17079 12035 17085
rect 13078 17076 13084 17128
rect 13136 17116 13142 17128
rect 13449 17119 13507 17125
rect 13449 17116 13461 17119
rect 13136 17088 13461 17116
rect 13136 17076 13142 17088
rect 13449 17085 13461 17088
rect 13495 17085 13507 17119
rect 13449 17079 13507 17085
rect 13814 17076 13820 17128
rect 13872 17116 13878 17128
rect 14001 17119 14059 17125
rect 14001 17116 14013 17119
rect 13872 17088 14013 17116
rect 13872 17076 13878 17088
rect 14001 17085 14013 17088
rect 14047 17085 14059 17119
rect 14001 17079 14059 17085
rect 14090 17076 14096 17128
rect 14148 17116 14154 17128
rect 14148 17088 14320 17116
rect 14148 17076 14154 17088
rect 3329 17051 3387 17057
rect 3329 17017 3341 17051
rect 3375 17017 3387 17051
rect 3329 17011 3387 17017
rect 4065 17051 4123 17057
rect 4065 17017 4077 17051
rect 4111 17048 4123 17051
rect 4246 17048 4252 17060
rect 4111 17020 4252 17048
rect 4111 17017 4123 17020
rect 4065 17011 4123 17017
rect 4246 17008 4252 17020
rect 4304 17008 4310 17060
rect 4430 17048 4436 17060
rect 4391 17020 4436 17048
rect 4430 17008 4436 17020
rect 4488 17008 4494 17060
rect 4798 17048 4804 17060
rect 4759 17020 4804 17048
rect 4798 17008 4804 17020
rect 4856 17008 4862 17060
rect 5166 17048 5172 17060
rect 5127 17020 5172 17048
rect 5166 17008 5172 17020
rect 5224 17008 5230 17060
rect 5534 17048 5540 17060
rect 5495 17020 5540 17048
rect 5534 17008 5540 17020
rect 5592 17008 5598 17060
rect 5810 17048 5816 17060
rect 5771 17020 5816 17048
rect 5810 17008 5816 17020
rect 5868 17008 5874 17060
rect 6181 17051 6239 17057
rect 6181 17017 6193 17051
rect 6227 17048 6239 17051
rect 6638 17048 6644 17060
rect 6227 17020 6644 17048
rect 6227 17017 6239 17020
rect 6181 17011 6239 17017
rect 6638 17008 6644 17020
rect 6696 17008 6702 17060
rect 6733 17051 6791 17057
rect 6733 17017 6745 17051
rect 6779 17017 6791 17051
rect 7098 17048 7104 17060
rect 7059 17020 7104 17048
rect 6733 17011 6791 17017
rect 2608 16952 2774 16980
rect 2866 16940 2872 16992
rect 2924 16980 2930 16992
rect 3234 16980 3240 16992
rect 2924 16952 3240 16980
rect 2924 16940 2930 16952
rect 3234 16940 3240 16952
rect 3292 16940 3298 16992
rect 6748 16980 6776 17011
rect 7098 17008 7104 17020
rect 7156 17008 7162 17060
rect 7469 17051 7527 17057
rect 7469 17017 7481 17051
rect 7515 17017 7527 17051
rect 7469 17011 7527 17017
rect 8205 17051 8263 17057
rect 8205 17017 8217 17051
rect 8251 17048 8263 17051
rect 8294 17048 8300 17060
rect 8251 17020 8300 17048
rect 8251 17017 8263 17020
rect 8205 17011 8263 17017
rect 7282 16980 7288 16992
rect 6748 16952 7288 16980
rect 7282 16940 7288 16952
rect 7340 16940 7346 16992
rect 7484 16980 7512 17011
rect 8294 17008 8300 17020
rect 8352 17008 8358 17060
rect 8754 17048 8760 17060
rect 8715 17020 8760 17048
rect 8754 17008 8760 17020
rect 8812 17008 8818 17060
rect 8938 17048 8944 17060
rect 8899 17020 8944 17048
rect 8938 17008 8944 17020
rect 8996 17008 9002 17060
rect 9398 17048 9404 17060
rect 9359 17020 9404 17048
rect 9398 17008 9404 17020
rect 9456 17008 9462 17060
rect 12713 17051 12771 17057
rect 12713 17017 12725 17051
rect 12759 17048 12771 17051
rect 12802 17048 12808 17060
rect 12759 17020 12808 17048
rect 12759 17017 12771 17020
rect 12713 17011 12771 17017
rect 12802 17008 12808 17020
rect 12860 17048 12866 17060
rect 14292 17048 14320 17088
rect 14366 17076 14372 17128
rect 14424 17116 14430 17128
rect 15488 17125 15516 17156
rect 15105 17119 15163 17125
rect 15105 17116 15117 17119
rect 14424 17088 15117 17116
rect 14424 17076 14430 17088
rect 15105 17085 15117 17088
rect 15151 17085 15163 17119
rect 15105 17079 15163 17085
rect 15473 17119 15531 17125
rect 15473 17085 15485 17119
rect 15519 17085 15531 17119
rect 15473 17079 15531 17085
rect 14645 17051 14703 17057
rect 14645 17048 14657 17051
rect 12860 17020 14228 17048
rect 14292 17020 14657 17048
rect 12860 17008 12866 17020
rect 8846 16980 8852 16992
rect 7484 16952 8852 16980
rect 8846 16940 8852 16952
rect 8904 16940 8910 16992
rect 9306 16940 9312 16992
rect 9364 16980 9370 16992
rect 9953 16983 10011 16989
rect 9953 16980 9965 16983
rect 9364 16952 9965 16980
rect 9364 16940 9370 16952
rect 9953 16949 9965 16952
rect 9999 16949 10011 16983
rect 9953 16943 10011 16949
rect 10226 16940 10232 16992
rect 10284 16980 10290 16992
rect 10321 16983 10379 16989
rect 10321 16980 10333 16983
rect 10284 16952 10333 16980
rect 10284 16940 10290 16952
rect 10321 16949 10333 16952
rect 10367 16949 10379 16983
rect 10321 16943 10379 16949
rect 10502 16940 10508 16992
rect 10560 16980 10566 16992
rect 10689 16983 10747 16989
rect 10689 16980 10701 16983
rect 10560 16952 10701 16980
rect 10560 16940 10566 16952
rect 10689 16949 10701 16952
rect 10735 16949 10747 16983
rect 10689 16943 10747 16949
rect 10778 16940 10784 16992
rect 10836 16980 10842 16992
rect 11057 16983 11115 16989
rect 11057 16980 11069 16983
rect 10836 16952 11069 16980
rect 10836 16940 10842 16952
rect 11057 16949 11069 16952
rect 11103 16949 11115 16983
rect 11057 16943 11115 16949
rect 11425 16983 11483 16989
rect 11425 16949 11437 16983
rect 11471 16980 11483 16983
rect 11882 16980 11888 16992
rect 11471 16952 11888 16980
rect 11471 16949 11483 16952
rect 11425 16943 11483 16949
rect 11882 16940 11888 16952
rect 11940 16940 11946 16992
rect 12066 16980 12072 16992
rect 12027 16952 12072 16980
rect 12066 16940 12072 16952
rect 12124 16940 12130 16992
rect 12618 16980 12624 16992
rect 12579 16952 12624 16980
rect 12618 16940 12624 16952
rect 12676 16940 12682 16992
rect 13909 16983 13967 16989
rect 13909 16949 13921 16983
rect 13955 16980 13967 16983
rect 14090 16980 14096 16992
rect 13955 16952 14096 16980
rect 13955 16949 13967 16952
rect 13909 16943 13967 16949
rect 14090 16940 14096 16952
rect 14148 16940 14154 16992
rect 14200 16980 14228 17020
rect 14645 17017 14657 17020
rect 14691 17017 14703 17051
rect 14645 17011 14703 17017
rect 14826 17008 14832 17060
rect 14884 17048 14890 17060
rect 14921 17051 14979 17057
rect 14921 17048 14933 17051
rect 14884 17020 14933 17048
rect 14884 17008 14890 17020
rect 14921 17017 14933 17020
rect 14967 17017 14979 17051
rect 15286 17048 15292 17060
rect 15247 17020 15292 17048
rect 14921 17011 14979 17017
rect 15286 17008 15292 17020
rect 15344 17008 15350 17060
rect 16574 16980 16580 16992
rect 14200 16952 16580 16980
rect 16574 16940 16580 16952
rect 16632 16940 16638 16992
rect 1104 16890 16008 16912
rect 1104 16838 5979 16890
rect 6031 16838 6043 16890
rect 6095 16838 6107 16890
rect 6159 16838 6171 16890
rect 6223 16838 10976 16890
rect 11028 16838 11040 16890
rect 11092 16838 11104 16890
rect 11156 16838 11168 16890
rect 11220 16838 16008 16890
rect 1104 16816 16008 16838
rect 566 16736 572 16788
rect 624 16776 630 16788
rect 1857 16779 1915 16785
rect 1857 16776 1869 16779
rect 624 16748 1869 16776
rect 624 16736 630 16748
rect 1857 16745 1869 16748
rect 1903 16745 1915 16779
rect 1857 16739 1915 16745
rect 2222 16736 2228 16788
rect 2280 16776 2286 16788
rect 2869 16779 2927 16785
rect 2869 16776 2881 16779
rect 2280 16748 2881 16776
rect 2280 16736 2286 16748
rect 2869 16745 2881 16748
rect 2915 16745 2927 16779
rect 2869 16739 2927 16745
rect 3234 16736 3240 16788
rect 3292 16776 3298 16788
rect 3329 16779 3387 16785
rect 3329 16776 3341 16779
rect 3292 16748 3341 16776
rect 3292 16736 3298 16748
rect 3329 16745 3341 16748
rect 3375 16745 3387 16779
rect 3329 16739 3387 16745
rect 5810 16736 5816 16788
rect 5868 16736 5874 16788
rect 6638 16736 6644 16788
rect 6696 16776 6702 16788
rect 9674 16776 9680 16788
rect 6696 16748 9680 16776
rect 6696 16736 6702 16748
rect 9674 16736 9680 16748
rect 9732 16736 9738 16788
rect 9858 16736 9864 16788
rect 9916 16776 9922 16788
rect 10229 16779 10287 16785
rect 10229 16776 10241 16779
rect 9916 16748 10241 16776
rect 9916 16736 9922 16748
rect 10229 16745 10241 16748
rect 10275 16745 10287 16779
rect 10594 16776 10600 16788
rect 10555 16748 10600 16776
rect 10229 16739 10287 16745
rect 10594 16736 10600 16748
rect 10652 16736 10658 16788
rect 10686 16736 10692 16788
rect 10744 16776 10750 16788
rect 10965 16779 11023 16785
rect 10965 16776 10977 16779
rect 10744 16748 10977 16776
rect 10744 16736 10750 16748
rect 10965 16745 10977 16748
rect 11011 16745 11023 16779
rect 11330 16776 11336 16788
rect 11291 16748 11336 16776
rect 10965 16739 11023 16745
rect 11330 16736 11336 16748
rect 11388 16736 11394 16788
rect 11790 16776 11796 16788
rect 11751 16748 11796 16776
rect 11790 16736 11796 16748
rect 11848 16736 11854 16788
rect 13081 16779 13139 16785
rect 13081 16776 13093 16779
rect 12544 16748 13093 16776
rect 198 16668 204 16720
rect 256 16708 262 16720
rect 1397 16711 1455 16717
rect 1397 16708 1409 16711
rect 256 16680 1409 16708
rect 256 16668 262 16680
rect 1397 16677 1409 16680
rect 1443 16677 1455 16711
rect 1949 16711 2007 16717
rect 1397 16671 1455 16677
rect 1504 16680 1808 16708
rect 1302 16600 1308 16652
rect 1360 16640 1366 16652
rect 1504 16640 1532 16680
rect 1360 16612 1532 16640
rect 1581 16643 1639 16649
rect 1360 16600 1366 16612
rect 1581 16609 1593 16643
rect 1627 16609 1639 16643
rect 1780 16640 1808 16680
rect 1949 16677 1961 16711
rect 1995 16708 2007 16711
rect 2685 16711 2743 16717
rect 1995 16680 2636 16708
rect 1995 16677 2007 16680
rect 1949 16671 2007 16677
rect 2133 16643 2191 16649
rect 2133 16640 2145 16643
rect 1780 16612 2145 16640
rect 1581 16603 1639 16609
rect 2133 16609 2145 16612
rect 2179 16609 2191 16643
rect 2133 16603 2191 16609
rect 2317 16643 2375 16649
rect 2317 16609 2329 16643
rect 2363 16640 2375 16643
rect 2406 16640 2412 16652
rect 2363 16612 2412 16640
rect 2363 16609 2375 16612
rect 2317 16603 2375 16609
rect 1596 16504 1624 16603
rect 2406 16600 2412 16612
rect 2464 16600 2470 16652
rect 2501 16643 2559 16649
rect 2501 16609 2513 16643
rect 2547 16609 2559 16643
rect 2608 16640 2636 16680
rect 2685 16677 2697 16711
rect 2731 16708 2743 16711
rect 4982 16708 4988 16720
rect 2731 16680 3648 16708
rect 4943 16680 4988 16708
rect 2731 16677 2743 16680
rect 2685 16671 2743 16677
rect 2866 16640 2872 16652
rect 2608 16612 2872 16640
rect 2501 16603 2559 16609
rect 1670 16532 1676 16584
rect 1728 16572 1734 16584
rect 2516 16572 2544 16603
rect 2866 16600 2872 16612
rect 2924 16600 2930 16652
rect 3053 16643 3111 16649
rect 3053 16609 3065 16643
rect 3099 16640 3111 16643
rect 3099 16612 3280 16640
rect 3099 16609 3111 16612
rect 3053 16603 3111 16609
rect 1728 16544 2544 16572
rect 1728 16532 1734 16544
rect 2038 16504 2044 16516
rect 1596 16476 2044 16504
rect 2038 16464 2044 16476
rect 2096 16464 2102 16516
rect 3252 16445 3280 16612
rect 3620 16513 3648 16680
rect 4982 16668 4988 16680
rect 5040 16668 5046 16720
rect 5350 16708 5356 16720
rect 5311 16680 5356 16708
rect 5350 16668 5356 16680
rect 5408 16668 5414 16720
rect 5718 16708 5724 16720
rect 5679 16680 5724 16708
rect 5718 16668 5724 16680
rect 5776 16668 5782 16720
rect 5828 16708 5856 16736
rect 9950 16708 9956 16720
rect 5828 16680 9956 16708
rect 9950 16668 9956 16680
rect 10008 16668 10014 16720
rect 12158 16668 12164 16720
rect 12216 16708 12222 16720
rect 12345 16711 12403 16717
rect 12345 16708 12357 16711
rect 12216 16680 12357 16708
rect 12216 16668 12222 16680
rect 12345 16677 12357 16680
rect 12391 16708 12403 16711
rect 12544 16708 12572 16748
rect 13081 16745 13093 16748
rect 13127 16745 13139 16779
rect 13081 16739 13139 16745
rect 13998 16736 14004 16788
rect 14056 16776 14062 16788
rect 14093 16779 14151 16785
rect 14093 16776 14105 16779
rect 14056 16748 14105 16776
rect 14056 16736 14062 16748
rect 14093 16745 14105 16748
rect 14139 16745 14151 16779
rect 16206 16776 16212 16788
rect 14093 16739 14151 16745
rect 14568 16748 16212 16776
rect 14568 16720 14596 16748
rect 16206 16736 16212 16748
rect 16264 16736 16270 16788
rect 12391 16680 12572 16708
rect 12391 16677 12403 16680
rect 12345 16671 12403 16677
rect 13354 16668 13360 16720
rect 13412 16708 13418 16720
rect 13449 16711 13507 16717
rect 13449 16708 13461 16711
rect 13412 16680 13461 16708
rect 13412 16668 13418 16680
rect 13449 16677 13461 16680
rect 13495 16677 13507 16711
rect 14550 16708 14556 16720
rect 14463 16680 14556 16708
rect 13449 16671 13507 16677
rect 14550 16668 14556 16680
rect 14608 16668 14614 16720
rect 15194 16668 15200 16720
rect 15252 16708 15258 16720
rect 15289 16711 15347 16717
rect 15289 16708 15301 16711
rect 15252 16680 15301 16708
rect 15252 16668 15258 16680
rect 15289 16677 15301 16680
rect 15335 16677 15347 16711
rect 15289 16671 15347 16677
rect 5169 16643 5227 16649
rect 5169 16609 5181 16643
rect 5215 16640 5227 16643
rect 5537 16643 5595 16649
rect 5215 16612 5488 16640
rect 5215 16609 5227 16612
rect 5169 16603 5227 16609
rect 5460 16572 5488 16612
rect 5537 16609 5549 16643
rect 5583 16640 5595 16643
rect 5810 16640 5816 16652
rect 5583 16612 5816 16640
rect 5583 16609 5595 16612
rect 5537 16603 5595 16609
rect 5810 16600 5816 16612
rect 5868 16600 5874 16652
rect 5905 16643 5963 16649
rect 5905 16609 5917 16643
rect 5951 16640 5963 16643
rect 7006 16640 7012 16652
rect 5951 16612 7012 16640
rect 5951 16609 5963 16612
rect 5905 16603 5963 16609
rect 7006 16600 7012 16612
rect 7064 16600 7070 16652
rect 8478 16600 8484 16652
rect 8536 16640 8542 16652
rect 9030 16640 9036 16652
rect 8536 16612 9036 16640
rect 8536 16600 8542 16612
rect 9030 16600 9036 16612
rect 9088 16600 9094 16652
rect 12526 16600 12532 16652
rect 12584 16640 12590 16652
rect 12713 16643 12771 16649
rect 12713 16640 12725 16643
rect 12584 16612 12725 16640
rect 12584 16600 12590 16612
rect 12713 16609 12725 16612
rect 12759 16609 12771 16643
rect 12713 16603 12771 16609
rect 6454 16572 6460 16584
rect 5460 16544 6460 16572
rect 6454 16532 6460 16544
rect 6512 16532 6518 16584
rect 9766 16572 9772 16584
rect 6564 16544 9772 16572
rect 3605 16507 3663 16513
rect 3605 16473 3617 16507
rect 3651 16504 3663 16507
rect 3878 16504 3884 16516
rect 3651 16476 3884 16504
rect 3651 16473 3663 16476
rect 3605 16467 3663 16473
rect 3878 16464 3884 16476
rect 3936 16464 3942 16516
rect 4522 16464 4528 16516
rect 4580 16504 4586 16516
rect 6564 16504 6592 16544
rect 9766 16532 9772 16544
rect 9824 16532 9830 16584
rect 12728 16572 12756 16603
rect 12802 16600 12808 16652
rect 12860 16640 12866 16652
rect 12897 16643 12955 16649
rect 12897 16640 12909 16643
rect 12860 16612 12909 16640
rect 12860 16600 12866 16612
rect 12897 16609 12909 16612
rect 12943 16609 12955 16643
rect 12897 16603 12955 16609
rect 14001 16643 14059 16649
rect 14001 16609 14013 16643
rect 14047 16640 14059 16643
rect 14366 16640 14372 16652
rect 14047 16612 14372 16640
rect 14047 16609 14059 16612
rect 14001 16603 14059 16609
rect 14366 16600 14372 16612
rect 14424 16600 14430 16652
rect 14921 16643 14979 16649
rect 14921 16609 14933 16643
rect 14967 16640 14979 16643
rect 15470 16640 15476 16652
rect 14967 16612 15476 16640
rect 14967 16609 14979 16612
rect 14921 16603 14979 16609
rect 15470 16600 15476 16612
rect 15528 16600 15534 16652
rect 15654 16640 15660 16652
rect 15615 16612 15660 16640
rect 15654 16600 15660 16612
rect 15712 16600 15718 16652
rect 13633 16575 13691 16581
rect 13633 16572 13645 16575
rect 12728 16544 13645 16572
rect 13633 16541 13645 16544
rect 13679 16541 13691 16575
rect 13633 16535 13691 16541
rect 4580 16476 6592 16504
rect 4580 16464 4586 16476
rect 6914 16464 6920 16516
rect 6972 16504 6978 16516
rect 7101 16507 7159 16513
rect 7101 16504 7113 16507
rect 6972 16476 7113 16504
rect 6972 16464 6978 16476
rect 7101 16473 7113 16476
rect 7147 16504 7159 16507
rect 12158 16504 12164 16516
rect 7147 16476 12020 16504
rect 12119 16476 12164 16504
rect 7147 16473 7159 16476
rect 7101 16467 7159 16473
rect 3237 16439 3295 16445
rect 3237 16405 3249 16439
rect 3283 16436 3295 16439
rect 3786 16436 3792 16448
rect 3283 16408 3792 16436
rect 3283 16405 3295 16408
rect 3237 16399 3295 16405
rect 3786 16396 3792 16408
rect 3844 16436 3850 16448
rect 3973 16439 4031 16445
rect 3973 16436 3985 16439
rect 3844 16408 3985 16436
rect 3844 16396 3850 16408
rect 3973 16405 3985 16408
rect 4019 16436 4031 16439
rect 5074 16436 5080 16448
rect 4019 16408 5080 16436
rect 4019 16405 4031 16408
rect 3973 16399 4031 16405
rect 5074 16396 5080 16408
rect 5132 16396 5138 16448
rect 6730 16436 6736 16448
rect 6691 16408 6736 16436
rect 6730 16396 6736 16408
rect 6788 16396 6794 16448
rect 7190 16396 7196 16448
rect 7248 16436 7254 16448
rect 9766 16436 9772 16448
rect 7248 16408 9772 16436
rect 7248 16396 7254 16408
rect 9766 16396 9772 16408
rect 9824 16396 9830 16448
rect 11992 16436 12020 16476
rect 12158 16464 12164 16476
rect 12216 16464 12222 16516
rect 12529 16507 12587 16513
rect 12529 16473 12541 16507
rect 12575 16504 12587 16507
rect 13262 16504 13268 16516
rect 12575 16476 13124 16504
rect 13223 16476 13268 16504
rect 12575 16473 12587 16476
rect 12529 16467 12587 16473
rect 12802 16436 12808 16448
rect 11992 16408 12808 16436
rect 12802 16396 12808 16408
rect 12860 16396 12866 16448
rect 13096 16436 13124 16476
rect 13262 16464 13268 16476
rect 13320 16464 13326 16516
rect 13906 16464 13912 16516
rect 13964 16504 13970 16516
rect 14737 16507 14795 16513
rect 14737 16504 14749 16507
rect 13964 16476 14749 16504
rect 13964 16464 13970 16476
rect 14737 16473 14749 16476
rect 14783 16473 14795 16507
rect 15102 16504 15108 16516
rect 15063 16476 15108 16504
rect 14737 16467 14795 16473
rect 15102 16464 15108 16476
rect 15160 16464 15166 16516
rect 13170 16436 13176 16448
rect 13096 16408 13176 16436
rect 13170 16396 13176 16408
rect 13228 16396 13234 16448
rect 14458 16436 14464 16448
rect 14419 16408 14464 16436
rect 14458 16396 14464 16408
rect 14516 16396 14522 16448
rect 1104 16346 16008 16368
rect 1104 16294 3480 16346
rect 3532 16294 3544 16346
rect 3596 16294 3608 16346
rect 3660 16294 3672 16346
rect 3724 16294 8478 16346
rect 8530 16294 8542 16346
rect 8594 16294 8606 16346
rect 8658 16294 8670 16346
rect 8722 16294 13475 16346
rect 13527 16294 13539 16346
rect 13591 16294 13603 16346
rect 13655 16294 13667 16346
rect 13719 16294 16008 16346
rect 1104 16272 16008 16294
rect 1486 16232 1492 16244
rect 1447 16204 1492 16232
rect 1486 16192 1492 16204
rect 1544 16192 1550 16244
rect 4798 16192 4804 16244
rect 4856 16232 4862 16244
rect 5169 16235 5227 16241
rect 5169 16232 5181 16235
rect 4856 16204 5181 16232
rect 4856 16192 4862 16204
rect 5169 16201 5181 16204
rect 5215 16201 5227 16235
rect 5169 16195 5227 16201
rect 5810 16192 5816 16244
rect 5868 16232 5874 16244
rect 6733 16235 6791 16241
rect 6733 16232 6745 16235
rect 5868 16204 6745 16232
rect 5868 16192 5874 16204
rect 6733 16201 6745 16204
rect 6779 16201 6791 16235
rect 7006 16232 7012 16244
rect 6967 16204 7012 16232
rect 6733 16195 6791 16201
rect 7006 16192 7012 16204
rect 7064 16192 7070 16244
rect 7282 16232 7288 16244
rect 7243 16204 7288 16232
rect 7282 16192 7288 16204
rect 7340 16192 7346 16244
rect 8849 16235 8907 16241
rect 8849 16201 8861 16235
rect 8895 16232 8907 16235
rect 8938 16232 8944 16244
rect 8895 16204 8944 16232
rect 8895 16201 8907 16204
rect 8849 16195 8907 16201
rect 8938 16192 8944 16204
rect 8996 16192 9002 16244
rect 13354 16192 13360 16244
rect 13412 16232 13418 16244
rect 13633 16235 13691 16241
rect 13633 16232 13645 16235
rect 13412 16204 13645 16232
rect 13412 16192 13418 16204
rect 13633 16201 13645 16204
rect 13679 16201 13691 16235
rect 14550 16232 14556 16244
rect 14511 16204 14556 16232
rect 13633 16195 13691 16201
rect 14550 16192 14556 16204
rect 14608 16192 14614 16244
rect 14734 16232 14740 16244
rect 14695 16204 14740 16232
rect 14734 16192 14740 16204
rect 14792 16192 14798 16244
rect 14918 16232 14924 16244
rect 14879 16204 14924 16232
rect 14918 16192 14924 16204
rect 14976 16192 14982 16244
rect 934 16124 940 16176
rect 992 16164 998 16176
rect 2041 16167 2099 16173
rect 2041 16164 2053 16167
rect 992 16136 2053 16164
rect 992 16124 998 16136
rect 2041 16133 2053 16136
rect 2087 16133 2099 16167
rect 6454 16164 6460 16176
rect 6415 16136 6460 16164
rect 2041 16127 2099 16133
rect 6454 16124 6460 16136
rect 6512 16124 6518 16176
rect 12894 16124 12900 16176
rect 12952 16164 12958 16176
rect 13817 16167 13875 16173
rect 13817 16164 13829 16167
rect 12952 16136 13829 16164
rect 12952 16124 12958 16136
rect 13817 16133 13829 16136
rect 13863 16133 13875 16167
rect 13817 16127 13875 16133
rect 2317 16099 2375 16105
rect 2317 16096 2329 16099
rect 1964 16068 2329 16096
rect 1964 16040 1992 16068
rect 2317 16065 2329 16068
rect 2363 16065 2375 16099
rect 8021 16099 8079 16105
rect 8021 16096 8033 16099
rect 2317 16059 2375 16065
rect 7208 16068 8033 16096
rect 1946 16028 1952 16040
rect 1907 16000 1952 16028
rect 1946 15988 1952 16000
rect 2004 15988 2010 16040
rect 2130 15988 2136 16040
rect 2188 16028 2194 16040
rect 2225 16031 2283 16037
rect 2225 16028 2237 16031
rect 2188 16000 2237 16028
rect 2188 15988 2194 16000
rect 2225 15997 2237 16000
rect 2271 15997 2283 16031
rect 2225 15991 2283 15997
rect 5353 16031 5411 16037
rect 5353 15997 5365 16031
rect 5399 16028 5411 16031
rect 5399 16000 5580 16028
rect 5399 15997 5411 16000
rect 5353 15991 5411 15997
rect 1581 15963 1639 15969
rect 1581 15929 1593 15963
rect 1627 15960 1639 15963
rect 3878 15960 3884 15972
rect 1627 15932 3884 15960
rect 1627 15929 1639 15932
rect 1581 15923 1639 15929
rect 3878 15920 3884 15932
rect 3936 15920 3942 15972
rect 2038 15852 2044 15904
rect 2096 15892 2102 15904
rect 2406 15892 2412 15904
rect 2096 15864 2412 15892
rect 2096 15852 2102 15864
rect 2406 15852 2412 15864
rect 2464 15892 2470 15904
rect 2501 15895 2559 15901
rect 2501 15892 2513 15895
rect 2464 15864 2513 15892
rect 2464 15852 2470 15864
rect 2501 15861 2513 15864
rect 2547 15861 2559 15895
rect 2501 15855 2559 15861
rect 2777 15895 2835 15901
rect 2777 15861 2789 15895
rect 2823 15892 2835 15895
rect 2866 15892 2872 15904
rect 2823 15864 2872 15892
rect 2823 15861 2835 15864
rect 2777 15855 2835 15861
rect 2866 15852 2872 15864
rect 2924 15852 2930 15904
rect 4706 15892 4712 15904
rect 4667 15864 4712 15892
rect 4706 15852 4712 15864
rect 4764 15852 4770 15904
rect 5552 15901 5580 16000
rect 6454 15988 6460 16040
rect 6512 16028 6518 16040
rect 6641 16031 6699 16037
rect 6641 16028 6653 16031
rect 6512 16000 6653 16028
rect 6512 15988 6518 16000
rect 6641 15997 6653 16000
rect 6687 16028 6699 16031
rect 6730 16028 6736 16040
rect 6687 16000 6736 16028
rect 6687 15997 6699 16000
rect 6641 15991 6699 15997
rect 6730 15988 6736 16000
rect 6788 15988 6794 16040
rect 6914 16028 6920 16040
rect 6875 16000 6920 16028
rect 6914 15988 6920 16000
rect 6972 15988 6978 16040
rect 7208 16037 7236 16068
rect 8021 16065 8033 16068
rect 8067 16096 8079 16099
rect 9214 16096 9220 16108
rect 8067 16068 9220 16096
rect 8067 16065 8079 16068
rect 8021 16059 8079 16065
rect 9214 16056 9220 16068
rect 9272 16056 9278 16108
rect 7193 16031 7251 16037
rect 7193 15997 7205 16031
rect 7239 15997 7251 16031
rect 7193 15991 7251 15997
rect 7469 16031 7527 16037
rect 7469 15997 7481 16031
rect 7515 16028 7527 16031
rect 8665 16031 8723 16037
rect 7515 16000 7696 16028
rect 7515 15997 7527 16000
rect 7469 15991 7527 15997
rect 5537 15895 5595 15901
rect 5537 15861 5549 15895
rect 5583 15892 5595 15895
rect 7282 15892 7288 15904
rect 5583 15864 7288 15892
rect 5583 15861 5595 15864
rect 5537 15855 5595 15861
rect 7282 15852 7288 15864
rect 7340 15852 7346 15904
rect 7558 15892 7564 15904
rect 7519 15864 7564 15892
rect 7558 15852 7564 15864
rect 7616 15852 7622 15904
rect 7668 15892 7696 16000
rect 8665 15997 8677 16031
rect 8711 16028 8723 16031
rect 9582 16028 9588 16040
rect 8711 16000 9588 16028
rect 8711 15997 8723 16000
rect 8665 15991 8723 15997
rect 9582 15988 9588 16000
rect 9640 15988 9646 16040
rect 11514 15988 11520 16040
rect 11572 16028 11578 16040
rect 15381 16031 15439 16037
rect 15381 16028 15393 16031
rect 11572 16000 15393 16028
rect 11572 15988 11578 16000
rect 15381 15997 15393 16000
rect 15427 15997 15439 16031
rect 15381 15991 15439 15997
rect 15565 16031 15623 16037
rect 15565 15997 15577 16031
rect 15611 16028 15623 16031
rect 15838 16028 15844 16040
rect 15611 16000 15844 16028
rect 15611 15997 15623 16000
rect 15565 15991 15623 15997
rect 15838 15988 15844 16000
rect 15896 15988 15902 16040
rect 8202 15960 8208 15972
rect 8115 15932 8208 15960
rect 8202 15920 8208 15932
rect 8260 15960 8266 15972
rect 9306 15960 9312 15972
rect 8260 15932 9312 15960
rect 8260 15920 8266 15932
rect 9306 15920 9312 15932
rect 9364 15920 9370 15972
rect 13814 15920 13820 15972
rect 13872 15960 13878 15972
rect 15013 15963 15071 15969
rect 15013 15960 15025 15963
rect 13872 15932 15025 15960
rect 13872 15920 13878 15932
rect 15013 15929 15025 15932
rect 15059 15929 15071 15963
rect 15013 15923 15071 15929
rect 15197 15963 15255 15969
rect 15197 15929 15209 15963
rect 15243 15960 15255 15963
rect 16942 15960 16948 15972
rect 15243 15932 16948 15960
rect 15243 15929 15255 15932
rect 15197 15923 15255 15929
rect 15396 15904 15424 15932
rect 16942 15920 16948 15932
rect 17000 15920 17006 15972
rect 7742 15892 7748 15904
rect 7668 15864 7748 15892
rect 7742 15852 7748 15864
rect 7800 15852 7806 15904
rect 7926 15852 7932 15904
rect 7984 15892 7990 15904
rect 8389 15895 8447 15901
rect 8389 15892 8401 15895
rect 7984 15864 8401 15892
rect 7984 15852 7990 15864
rect 8389 15861 8401 15864
rect 8435 15892 8447 15895
rect 9490 15892 9496 15904
rect 8435 15864 9496 15892
rect 8435 15861 8447 15864
rect 8389 15855 8447 15861
rect 9490 15852 9496 15864
rect 9548 15892 9554 15904
rect 10502 15892 10508 15904
rect 9548 15864 10508 15892
rect 9548 15852 9554 15864
rect 10502 15852 10508 15864
rect 10560 15852 10566 15904
rect 15378 15852 15384 15904
rect 15436 15852 15442 15904
rect 1104 15802 16008 15824
rect 1104 15750 5979 15802
rect 6031 15750 6043 15802
rect 6095 15750 6107 15802
rect 6159 15750 6171 15802
rect 6223 15750 10976 15802
rect 11028 15750 11040 15802
rect 11092 15750 11104 15802
rect 11156 15750 11168 15802
rect 11220 15750 16008 15802
rect 1104 15728 16008 15750
rect 2958 15648 2964 15700
rect 3016 15688 3022 15700
rect 3881 15691 3939 15697
rect 3881 15688 3893 15691
rect 3016 15660 3893 15688
rect 3016 15648 3022 15660
rect 3881 15657 3893 15660
rect 3927 15657 3939 15691
rect 4154 15688 4160 15700
rect 4115 15660 4160 15688
rect 3881 15651 3939 15657
rect 4154 15648 4160 15660
rect 4212 15648 4218 15700
rect 4430 15648 4436 15700
rect 4488 15688 4494 15700
rect 4709 15691 4767 15697
rect 4709 15688 4721 15691
rect 4488 15660 4721 15688
rect 4488 15648 4494 15660
rect 4709 15657 4721 15660
rect 4755 15657 4767 15691
rect 4709 15651 4767 15657
rect 5166 15648 5172 15700
rect 5224 15688 5230 15700
rect 5261 15691 5319 15697
rect 5261 15688 5273 15691
rect 5224 15660 5273 15688
rect 5224 15648 5230 15660
rect 5261 15657 5273 15660
rect 5307 15657 5319 15691
rect 5534 15688 5540 15700
rect 5495 15660 5540 15688
rect 5261 15651 5319 15657
rect 5534 15648 5540 15660
rect 5592 15648 5598 15700
rect 6730 15688 6736 15700
rect 6691 15660 6736 15688
rect 6730 15648 6736 15660
rect 6788 15648 6794 15700
rect 7098 15648 7104 15700
rect 7156 15688 7162 15700
rect 8021 15691 8079 15697
rect 8021 15688 8033 15691
rect 7156 15660 8033 15688
rect 7156 15648 7162 15660
rect 8021 15657 8033 15660
rect 8067 15657 8079 15691
rect 8021 15651 8079 15657
rect 8294 15648 8300 15700
rect 8352 15688 8358 15700
rect 8573 15691 8631 15697
rect 8573 15688 8585 15691
rect 8352 15660 8585 15688
rect 8352 15648 8358 15660
rect 8573 15657 8585 15660
rect 8619 15657 8631 15691
rect 9122 15688 9128 15700
rect 9083 15660 9128 15688
rect 8573 15651 8631 15657
rect 9122 15648 9128 15660
rect 9180 15648 9186 15700
rect 9398 15688 9404 15700
rect 9359 15660 9404 15688
rect 9398 15648 9404 15660
rect 9456 15648 9462 15700
rect 9674 15688 9680 15700
rect 9635 15660 9680 15688
rect 9674 15648 9680 15660
rect 9732 15648 9738 15700
rect 9950 15688 9956 15700
rect 9911 15660 9956 15688
rect 9950 15648 9956 15660
rect 10008 15648 10014 15700
rect 15381 15691 15439 15697
rect 15381 15657 15393 15691
rect 15427 15688 15439 15691
rect 15838 15688 15844 15700
rect 15427 15660 15844 15688
rect 15427 15657 15439 15660
rect 15381 15651 15439 15657
rect 15838 15648 15844 15660
rect 15896 15648 15902 15700
rect 1394 15580 1400 15632
rect 1452 15620 1458 15632
rect 1857 15623 1915 15629
rect 1857 15620 1869 15623
rect 1452 15592 1869 15620
rect 1452 15580 1458 15592
rect 1857 15589 1869 15592
rect 1903 15620 1915 15623
rect 4522 15620 4528 15632
rect 1903 15592 4528 15620
rect 1903 15589 1915 15592
rect 1857 15583 1915 15589
rect 4522 15580 4528 15592
rect 4580 15580 4586 15632
rect 6089 15623 6147 15629
rect 6089 15620 6101 15623
rect 5460 15592 6101 15620
rect 1581 15555 1639 15561
rect 1581 15521 1593 15555
rect 1627 15552 1639 15555
rect 2774 15552 2780 15564
rect 1627 15524 2780 15552
rect 1627 15521 1639 15524
rect 1581 15515 1639 15521
rect 2774 15512 2780 15524
rect 2832 15512 2838 15564
rect 4065 15555 4123 15561
rect 4065 15521 4077 15555
rect 4111 15521 4123 15555
rect 4338 15552 4344 15564
rect 4299 15524 4344 15552
rect 4065 15515 4123 15521
rect 4080 15484 4108 15515
rect 4338 15512 4344 15524
rect 4396 15512 4402 15564
rect 4617 15555 4675 15561
rect 4617 15521 4629 15555
rect 4663 15552 4675 15555
rect 4706 15552 4712 15564
rect 4663 15524 4712 15552
rect 4663 15521 4675 15524
rect 4617 15515 4675 15521
rect 4632 15484 4660 15515
rect 4706 15512 4712 15524
rect 4764 15512 4770 15564
rect 5460 15561 5488 15592
rect 6089 15589 6101 15592
rect 6135 15620 6147 15623
rect 7190 15620 7196 15632
rect 6135 15592 7196 15620
rect 6135 15589 6147 15592
rect 6089 15583 6147 15589
rect 7190 15580 7196 15592
rect 7248 15580 7254 15632
rect 7653 15623 7711 15629
rect 7653 15589 7665 15623
rect 7699 15620 7711 15623
rect 7926 15620 7932 15632
rect 7699 15592 7932 15620
rect 7699 15589 7711 15592
rect 7653 15583 7711 15589
rect 7926 15580 7932 15592
rect 7984 15580 7990 15632
rect 11422 15620 11428 15632
rect 8312 15592 8800 15620
rect 8312 15564 8340 15592
rect 4893 15555 4951 15561
rect 4893 15521 4905 15555
rect 4939 15552 4951 15555
rect 5169 15555 5227 15561
rect 5169 15552 5181 15555
rect 4939 15524 5181 15552
rect 4939 15521 4951 15524
rect 4893 15515 4951 15521
rect 5169 15521 5181 15524
rect 5215 15521 5227 15555
rect 5169 15515 5227 15521
rect 5445 15555 5503 15561
rect 5445 15521 5457 15555
rect 5491 15521 5503 15555
rect 5445 15515 5503 15521
rect 5721 15555 5779 15561
rect 5721 15521 5733 15555
rect 5767 15552 5779 15555
rect 5994 15552 6000 15564
rect 5767 15524 6000 15552
rect 5767 15521 5779 15524
rect 5721 15515 5779 15521
rect 5994 15512 6000 15524
rect 6052 15512 6058 15564
rect 6178 15512 6184 15564
rect 6236 15552 6242 15564
rect 6825 15555 6883 15561
rect 6825 15552 6837 15555
rect 6236 15524 6837 15552
rect 6236 15512 6242 15524
rect 6825 15521 6837 15524
rect 6871 15552 6883 15555
rect 7466 15552 7472 15564
rect 6871 15524 7472 15552
rect 6871 15521 6883 15524
rect 6825 15515 6883 15521
rect 7466 15512 7472 15524
rect 7524 15512 7530 15564
rect 7561 15555 7619 15561
rect 7561 15521 7573 15555
rect 7607 15552 7619 15555
rect 7742 15552 7748 15564
rect 7607 15524 7748 15552
rect 7607 15521 7619 15524
rect 7561 15515 7619 15521
rect 5902 15484 5908 15496
rect 4080 15456 4568 15484
rect 4632 15456 5908 15484
rect 1394 15416 1400 15428
rect 1355 15388 1400 15416
rect 1394 15376 1400 15388
rect 1452 15376 1458 15428
rect 4246 15376 4252 15428
rect 4304 15416 4310 15428
rect 4433 15419 4491 15425
rect 4433 15416 4445 15419
rect 4304 15388 4445 15416
rect 4304 15376 4310 15388
rect 4433 15385 4445 15388
rect 4479 15385 4491 15419
rect 4540 15416 4568 15456
rect 5902 15444 5908 15456
rect 5960 15484 5966 15496
rect 7006 15484 7012 15496
rect 5960 15456 6316 15484
rect 6967 15456 7012 15484
rect 5960 15444 5966 15456
rect 5077 15419 5135 15425
rect 5077 15416 5089 15419
rect 4540 15388 5089 15416
rect 4433 15379 4491 15385
rect 5077 15385 5089 15388
rect 5123 15416 5135 15419
rect 6086 15416 6092 15428
rect 5123 15388 6092 15416
rect 5123 15385 5135 15388
rect 5077 15379 5135 15385
rect 6086 15376 6092 15388
rect 6144 15376 6150 15428
rect 6288 15425 6316 15456
rect 7006 15444 7012 15456
rect 7064 15444 7070 15496
rect 6273 15419 6331 15425
rect 6273 15385 6285 15419
rect 6319 15416 6331 15419
rect 6730 15416 6736 15428
rect 6319 15388 6736 15416
rect 6319 15385 6331 15388
rect 6273 15379 6331 15385
rect 6730 15376 6736 15388
rect 6788 15376 6794 15428
rect 5169 15351 5227 15357
rect 5169 15317 5181 15351
rect 5215 15348 5227 15351
rect 5810 15348 5816 15360
rect 5215 15320 5816 15348
rect 5215 15317 5227 15320
rect 5169 15311 5227 15317
rect 5810 15308 5816 15320
rect 5868 15308 5874 15360
rect 6362 15348 6368 15360
rect 6323 15320 6368 15348
rect 6362 15308 6368 15320
rect 6420 15308 6426 15360
rect 6914 15308 6920 15360
rect 6972 15348 6978 15360
rect 7193 15351 7251 15357
rect 7193 15348 7205 15351
rect 6972 15320 7205 15348
rect 6972 15308 6978 15320
rect 7193 15317 7205 15320
rect 7239 15317 7251 15351
rect 7576 15348 7604 15515
rect 7742 15512 7748 15524
rect 7800 15512 7806 15564
rect 8202 15552 8208 15564
rect 8163 15524 8208 15552
rect 8202 15512 8208 15524
rect 8260 15512 8266 15564
rect 8294 15512 8300 15564
rect 8352 15512 8358 15564
rect 8481 15555 8539 15561
rect 8481 15521 8493 15555
rect 8527 15552 8539 15555
rect 8662 15552 8668 15564
rect 8527 15524 8668 15552
rect 8527 15521 8539 15524
rect 8481 15515 8539 15521
rect 8662 15512 8668 15524
rect 8720 15512 8726 15564
rect 8772 15561 8800 15592
rect 9324 15592 11428 15620
rect 9324 15561 9352 15592
rect 11422 15580 11428 15592
rect 11480 15580 11486 15632
rect 15194 15580 15200 15632
rect 15252 15620 15258 15632
rect 15473 15623 15531 15629
rect 15473 15620 15485 15623
rect 15252 15592 15485 15620
rect 15252 15580 15258 15592
rect 15473 15589 15485 15592
rect 15519 15589 15531 15623
rect 15473 15583 15531 15589
rect 8757 15555 8815 15561
rect 8757 15521 8769 15555
rect 8803 15521 8815 15555
rect 8757 15515 8815 15521
rect 9309 15555 9367 15561
rect 9309 15521 9321 15555
rect 9355 15521 9367 15555
rect 9309 15515 9367 15521
rect 9585 15555 9643 15561
rect 9585 15521 9597 15555
rect 9631 15521 9643 15555
rect 9858 15552 9864 15564
rect 9819 15524 9864 15552
rect 9585 15515 9643 15521
rect 7650 15444 7656 15496
rect 7708 15484 7714 15496
rect 7837 15487 7895 15493
rect 7837 15484 7849 15487
rect 7708 15456 7849 15484
rect 7708 15444 7714 15456
rect 7837 15453 7849 15456
rect 7883 15484 7895 15487
rect 8018 15484 8024 15496
rect 7883 15456 8024 15484
rect 7883 15453 7895 15456
rect 7837 15447 7895 15453
rect 8018 15444 8024 15456
rect 8076 15444 8082 15496
rect 8846 15484 8852 15496
rect 8312 15456 8852 15484
rect 8312 15425 8340 15456
rect 8846 15444 8852 15456
rect 8904 15444 8910 15496
rect 9214 15444 9220 15496
rect 9272 15484 9278 15496
rect 9490 15484 9496 15496
rect 9272 15456 9496 15484
rect 9272 15444 9278 15456
rect 9490 15444 9496 15456
rect 9548 15444 9554 15496
rect 9600 15484 9628 15515
rect 9858 15512 9864 15524
rect 9916 15512 9922 15564
rect 10134 15552 10140 15564
rect 10095 15524 10140 15552
rect 10134 15512 10140 15524
rect 10192 15512 10198 15564
rect 15013 15555 15071 15561
rect 15013 15521 15025 15555
rect 15059 15552 15071 15555
rect 15378 15552 15384 15564
rect 15059 15524 15384 15552
rect 15059 15521 15071 15524
rect 15013 15515 15071 15521
rect 15378 15512 15384 15524
rect 15436 15512 15442 15564
rect 11790 15484 11796 15496
rect 9600 15456 11796 15484
rect 11790 15444 11796 15456
rect 11848 15444 11854 15496
rect 15197 15487 15255 15493
rect 15197 15453 15209 15487
rect 15243 15484 15255 15487
rect 15470 15484 15476 15496
rect 15243 15456 15476 15484
rect 15243 15453 15255 15456
rect 15197 15447 15255 15453
rect 15470 15444 15476 15456
rect 15528 15444 15534 15496
rect 8297 15419 8355 15425
rect 8297 15385 8309 15419
rect 8343 15385 8355 15419
rect 8297 15379 8355 15385
rect 8941 15419 8999 15425
rect 8941 15385 8953 15419
rect 8987 15416 8999 15419
rect 12802 15416 12808 15428
rect 8987 15388 12808 15416
rect 8987 15385 8999 15388
rect 8941 15379 8999 15385
rect 8956 15348 8984 15379
rect 12802 15376 12808 15388
rect 12860 15376 12866 15428
rect 7576 15320 8984 15348
rect 7193 15311 7251 15317
rect 9858 15308 9864 15360
rect 9916 15348 9922 15360
rect 10321 15351 10379 15357
rect 10321 15348 10333 15351
rect 9916 15320 10333 15348
rect 9916 15308 9922 15320
rect 10321 15317 10333 15320
rect 10367 15348 10379 15351
rect 10686 15348 10692 15360
rect 10367 15320 10692 15348
rect 10367 15317 10379 15320
rect 10321 15311 10379 15317
rect 10686 15308 10692 15320
rect 10744 15308 10750 15360
rect 1104 15258 16008 15280
rect 1104 15206 3480 15258
rect 3532 15206 3544 15258
rect 3596 15206 3608 15258
rect 3660 15206 3672 15258
rect 3724 15206 8478 15258
rect 8530 15206 8542 15258
rect 8594 15206 8606 15258
rect 8658 15206 8670 15258
rect 8722 15206 13475 15258
rect 13527 15206 13539 15258
rect 13591 15206 13603 15258
rect 13655 15206 13667 15258
rect 13719 15206 16008 15258
rect 1104 15184 16008 15206
rect 3326 15104 3332 15156
rect 3384 15144 3390 15156
rect 5537 15147 5595 15153
rect 5537 15144 5549 15147
rect 3384 15116 5549 15144
rect 3384 15104 3390 15116
rect 5537 15113 5549 15116
rect 5583 15113 5595 15147
rect 5537 15107 5595 15113
rect 7190 15104 7196 15156
rect 7248 15144 7254 15156
rect 8113 15147 8171 15153
rect 8113 15144 8125 15147
rect 7248 15116 8125 15144
rect 7248 15104 7254 15116
rect 8113 15113 8125 15116
rect 8159 15113 8171 15147
rect 8113 15107 8171 15113
rect 8941 15147 8999 15153
rect 8941 15113 8953 15147
rect 8987 15144 8999 15147
rect 9030 15144 9036 15156
rect 8987 15116 9036 15144
rect 8987 15113 8999 15116
rect 8941 15107 8999 15113
rect 9030 15104 9036 15116
rect 9088 15104 9094 15156
rect 9122 15104 9128 15156
rect 9180 15144 9186 15156
rect 9309 15147 9367 15153
rect 9309 15144 9321 15147
rect 9180 15116 9321 15144
rect 9180 15104 9186 15116
rect 9309 15113 9321 15116
rect 9355 15144 9367 15147
rect 9858 15144 9864 15156
rect 9355 15116 9864 15144
rect 9355 15113 9367 15116
rect 9309 15107 9367 15113
rect 9858 15104 9864 15116
rect 9916 15104 9922 15156
rect 7650 15076 7656 15088
rect 6196 15048 7656 15076
rect 5074 14968 5080 15020
rect 5132 15008 5138 15020
rect 6196 15017 6224 15048
rect 7650 15036 7656 15048
rect 7708 15036 7714 15088
rect 10042 15076 10048 15088
rect 7944 15048 10048 15076
rect 5261 15011 5319 15017
rect 5261 15008 5273 15011
rect 5132 14980 5273 15008
rect 5132 14968 5138 14980
rect 5261 14977 5273 14980
rect 5307 14977 5319 15011
rect 5261 14971 5319 14977
rect 6181 15011 6239 15017
rect 6181 14977 6193 15011
rect 6227 14977 6239 15011
rect 6181 14971 6239 14977
rect 6822 14968 6828 15020
rect 6880 15008 6886 15020
rect 7009 15011 7067 15017
rect 7009 15008 7021 15011
rect 6880 14980 7021 15008
rect 6880 14968 6886 14980
rect 7009 14977 7021 14980
rect 7055 15008 7067 15011
rect 7837 15011 7895 15017
rect 7837 15008 7849 15011
rect 7055 14980 7849 15008
rect 7055 14977 7067 14980
rect 7009 14971 7067 14977
rect 7837 14977 7849 14980
rect 7883 14977 7895 15011
rect 7837 14971 7895 14977
rect 4338 14900 4344 14952
rect 4396 14940 4402 14952
rect 4525 14943 4583 14949
rect 4525 14940 4537 14943
rect 4396 14912 4537 14940
rect 4396 14900 4402 14912
rect 4525 14909 4537 14912
rect 4571 14940 4583 14943
rect 5902 14940 5908 14952
rect 4571 14912 5534 14940
rect 5863 14912 5908 14940
rect 4571 14909 4583 14912
rect 4525 14903 4583 14909
rect 5506 14872 5534 14912
rect 5902 14900 5908 14912
rect 5960 14900 5966 14952
rect 5997 14943 6055 14949
rect 5997 14909 6009 14943
rect 6043 14940 6055 14943
rect 6362 14940 6368 14952
rect 6043 14912 6368 14940
rect 6043 14909 6055 14912
rect 5997 14903 6055 14909
rect 6362 14900 6368 14912
rect 6420 14900 6426 14952
rect 7745 14943 7803 14949
rect 6472 14912 7696 14940
rect 6472 14872 6500 14912
rect 4172 14844 4752 14872
rect 5506 14844 6500 14872
rect 2682 14764 2688 14816
rect 2740 14804 2746 14816
rect 4172 14804 4200 14844
rect 4724 14813 4752 14844
rect 6546 14832 6552 14884
rect 6604 14872 6610 14884
rect 6917 14875 6975 14881
rect 6917 14872 6929 14875
rect 6604 14844 6929 14872
rect 6604 14832 6610 14844
rect 6917 14841 6929 14844
rect 6963 14841 6975 14875
rect 7466 14872 7472 14884
rect 6917 14835 6975 14841
rect 7024 14844 7472 14872
rect 2740 14776 4200 14804
rect 4709 14807 4767 14813
rect 2740 14764 2746 14776
rect 4709 14773 4721 14807
rect 4755 14773 4767 14807
rect 4709 14767 4767 14773
rect 4982 14764 4988 14816
rect 5040 14804 5046 14816
rect 5077 14807 5135 14813
rect 5077 14804 5089 14807
rect 5040 14776 5089 14804
rect 5040 14764 5046 14776
rect 5077 14773 5089 14776
rect 5123 14773 5135 14807
rect 5077 14767 5135 14773
rect 5169 14807 5227 14813
rect 5169 14773 5181 14807
rect 5215 14804 5227 14807
rect 5258 14804 5264 14816
rect 5215 14776 5264 14804
rect 5215 14773 5227 14776
rect 5169 14767 5227 14773
rect 5258 14764 5264 14776
rect 5316 14764 5322 14816
rect 5718 14764 5724 14816
rect 5776 14804 5782 14816
rect 6457 14807 6515 14813
rect 6457 14804 6469 14807
rect 5776 14776 6469 14804
rect 5776 14764 5782 14776
rect 6457 14773 6469 14776
rect 6503 14773 6515 14807
rect 6457 14767 6515 14773
rect 6825 14807 6883 14813
rect 6825 14773 6837 14807
rect 6871 14804 6883 14807
rect 7024 14804 7052 14844
rect 7466 14832 7472 14844
rect 7524 14832 7530 14884
rect 7668 14872 7696 14912
rect 7745 14909 7757 14943
rect 7791 14940 7803 14943
rect 7944 14940 7972 15048
rect 10042 15036 10048 15048
rect 10100 15036 10106 15088
rect 8018 14968 8024 15020
rect 8076 15008 8082 15020
rect 8662 15008 8668 15020
rect 8076 14980 8668 15008
rect 8076 14968 8082 14980
rect 8662 14968 8668 14980
rect 8720 14968 8726 15020
rect 8754 14968 8760 15020
rect 8812 15008 8818 15020
rect 8812 14980 12434 15008
rect 8812 14968 8818 14980
rect 7791 14912 7972 14940
rect 9125 14943 9183 14949
rect 7791 14909 7803 14912
rect 7745 14903 7803 14909
rect 9125 14909 9137 14943
rect 9171 14940 9183 14943
rect 12250 14940 12256 14952
rect 9171 14912 12256 14940
rect 9171 14909 9183 14912
rect 9125 14903 9183 14909
rect 12250 14900 12256 14912
rect 12308 14900 12314 14952
rect 8386 14872 8392 14884
rect 7668 14844 8392 14872
rect 8386 14832 8392 14844
rect 8444 14832 8450 14884
rect 8573 14875 8631 14881
rect 8573 14841 8585 14875
rect 8619 14872 8631 14875
rect 12406 14872 12434 14980
rect 14366 14872 14372 14884
rect 8619 14844 9536 14872
rect 12406 14844 14372 14872
rect 8619 14841 8631 14844
rect 8573 14835 8631 14841
rect 6871 14776 7052 14804
rect 6871 14773 6883 14776
rect 6825 14767 6883 14773
rect 7098 14764 7104 14816
rect 7156 14804 7162 14816
rect 7285 14807 7343 14813
rect 7285 14804 7297 14807
rect 7156 14776 7297 14804
rect 7156 14764 7162 14776
rect 7285 14773 7297 14776
rect 7331 14773 7343 14807
rect 7285 14767 7343 14773
rect 7653 14807 7711 14813
rect 7653 14773 7665 14807
rect 7699 14804 7711 14807
rect 7742 14804 7748 14816
rect 7699 14776 7748 14804
rect 7699 14773 7711 14776
rect 7653 14767 7711 14773
rect 7742 14764 7748 14776
rect 7800 14764 7806 14816
rect 8481 14807 8539 14813
rect 8481 14773 8493 14807
rect 8527 14804 8539 14807
rect 9122 14804 9128 14816
rect 8527 14776 9128 14804
rect 8527 14773 8539 14776
rect 8481 14767 8539 14773
rect 9122 14764 9128 14776
rect 9180 14764 9186 14816
rect 9508 14813 9536 14844
rect 14366 14832 14372 14844
rect 14424 14832 14430 14884
rect 9493 14807 9551 14813
rect 9493 14773 9505 14807
rect 9539 14804 9551 14807
rect 14090 14804 14096 14816
rect 9539 14776 14096 14804
rect 9539 14773 9551 14776
rect 9493 14767 9551 14773
rect 14090 14764 14096 14776
rect 14148 14804 14154 14816
rect 14550 14804 14556 14816
rect 14148 14776 14556 14804
rect 14148 14764 14154 14776
rect 14550 14764 14556 14776
rect 14608 14764 14614 14816
rect 1104 14714 16008 14736
rect 1104 14662 5979 14714
rect 6031 14662 6043 14714
rect 6095 14662 6107 14714
rect 6159 14662 6171 14714
rect 6223 14662 10976 14714
rect 11028 14662 11040 14714
rect 11092 14662 11104 14714
rect 11156 14662 11168 14714
rect 11220 14662 16008 14714
rect 1104 14640 16008 14662
rect 4614 14600 4620 14612
rect 4575 14572 4620 14600
rect 4614 14560 4620 14572
rect 4672 14560 4678 14612
rect 4982 14600 4988 14612
rect 4943 14572 4988 14600
rect 4982 14560 4988 14572
rect 5040 14560 5046 14612
rect 5445 14603 5503 14609
rect 5445 14569 5457 14603
rect 5491 14600 5503 14603
rect 9858 14600 9864 14612
rect 5491 14572 8616 14600
rect 5491 14569 5503 14572
rect 5445 14563 5503 14569
rect 4525 14535 4583 14541
rect 4525 14501 4537 14535
rect 4571 14532 4583 14535
rect 7040 14535 7098 14541
rect 4571 14504 6960 14532
rect 4571 14501 4583 14504
rect 4525 14495 4583 14501
rect 1581 14467 1639 14473
rect 1581 14433 1593 14467
rect 1627 14464 1639 14467
rect 2498 14464 2504 14476
rect 1627 14436 2504 14464
rect 1627 14433 1639 14436
rect 1581 14427 1639 14433
rect 2498 14424 2504 14436
rect 2556 14424 2562 14476
rect 4062 14424 4068 14476
rect 4120 14464 4126 14476
rect 6546 14464 6552 14476
rect 4120 14436 6552 14464
rect 4120 14424 4126 14436
rect 6546 14424 6552 14436
rect 6604 14424 6610 14476
rect 6932 14464 6960 14504
rect 7040 14501 7052 14535
rect 7086 14532 7098 14535
rect 7650 14532 7656 14544
rect 7086 14504 7656 14532
rect 7086 14501 7098 14504
rect 7040 14495 7098 14501
rect 7650 14492 7656 14504
rect 7708 14492 7714 14544
rect 7745 14535 7803 14541
rect 7745 14501 7757 14535
rect 7791 14532 7803 14535
rect 7926 14532 7932 14544
rect 7791 14504 7932 14532
rect 7791 14501 7803 14504
rect 7745 14495 7803 14501
rect 7926 14492 7932 14504
rect 7984 14492 7990 14544
rect 8386 14492 8392 14544
rect 8444 14532 8450 14544
rect 8481 14535 8539 14541
rect 8481 14532 8493 14535
rect 8444 14504 8493 14532
rect 8444 14492 8450 14504
rect 8481 14501 8493 14504
rect 8527 14501 8539 14535
rect 8588 14532 8616 14572
rect 8864 14572 9864 14600
rect 8864 14532 8892 14572
rect 9858 14560 9864 14572
rect 9916 14560 9922 14612
rect 8588 14504 8892 14532
rect 8481 14495 8539 14501
rect 7837 14467 7895 14473
rect 6932 14436 7795 14464
rect 3786 14356 3792 14408
rect 3844 14396 3850 14408
rect 4341 14399 4399 14405
rect 4341 14396 4353 14399
rect 3844 14368 4353 14396
rect 3844 14356 3850 14368
rect 4341 14365 4353 14368
rect 4387 14365 4399 14399
rect 5534 14396 5540 14408
rect 5495 14368 5540 14396
rect 4341 14359 4399 14365
rect 5534 14356 5540 14368
rect 5592 14356 5598 14408
rect 5629 14399 5687 14405
rect 5629 14365 5641 14399
rect 5675 14365 5687 14399
rect 5629 14359 5687 14365
rect 7285 14399 7343 14405
rect 7285 14365 7297 14399
rect 7331 14396 7343 14399
rect 7650 14396 7656 14408
rect 7331 14368 7656 14396
rect 7331 14365 7343 14368
rect 7285 14359 7343 14365
rect 1394 14328 1400 14340
rect 1355 14300 1400 14328
rect 1394 14288 1400 14300
rect 1452 14288 1458 14340
rect 4614 14288 4620 14340
rect 4672 14328 4678 14340
rect 5644 14328 5672 14359
rect 7650 14356 7656 14368
rect 7708 14356 7714 14408
rect 6270 14328 6276 14340
rect 4672 14300 6276 14328
rect 4672 14288 4678 14300
rect 6270 14288 6276 14300
rect 6328 14288 6334 14340
rect 4522 14220 4528 14272
rect 4580 14260 4586 14272
rect 5077 14263 5135 14269
rect 5077 14260 5089 14263
rect 4580 14232 5089 14260
rect 4580 14220 4586 14232
rect 5077 14229 5089 14232
rect 5123 14229 5135 14263
rect 5902 14260 5908 14272
rect 5863 14232 5908 14260
rect 5077 14223 5135 14229
rect 5902 14220 5908 14232
rect 5960 14220 5966 14272
rect 7374 14260 7380 14272
rect 7335 14232 7380 14260
rect 7374 14220 7380 14232
rect 7432 14220 7438 14272
rect 7767 14260 7795 14436
rect 7837 14433 7849 14467
rect 7883 14433 7895 14467
rect 7837 14427 7895 14433
rect 7852 14340 7880 14427
rect 7929 14399 7987 14405
rect 7929 14365 7941 14399
rect 7975 14365 7987 14399
rect 7929 14359 7987 14365
rect 7834 14288 7840 14340
rect 7892 14288 7898 14340
rect 7944 14328 7972 14359
rect 8018 14356 8024 14408
rect 8076 14396 8082 14408
rect 8297 14399 8355 14405
rect 8297 14396 8309 14399
rect 8076 14368 8309 14396
rect 8076 14356 8082 14368
rect 8297 14365 8309 14368
rect 8343 14365 8355 14399
rect 8297 14359 8355 14365
rect 8110 14328 8116 14340
rect 7944 14300 8116 14328
rect 8110 14288 8116 14300
rect 8168 14288 8174 14340
rect 8496 14328 8524 14495
rect 8938 14492 8944 14544
rect 8996 14532 9002 14544
rect 9306 14532 9312 14544
rect 8996 14504 9312 14532
rect 8996 14492 9002 14504
rect 9306 14492 9312 14504
rect 9364 14532 9370 14544
rect 9677 14535 9735 14541
rect 9677 14532 9689 14535
rect 9364 14504 9689 14532
rect 9364 14492 9370 14504
rect 9677 14501 9689 14504
rect 9723 14501 9735 14535
rect 9677 14495 9735 14501
rect 10137 14535 10195 14541
rect 10137 14501 10149 14535
rect 10183 14532 10195 14535
rect 10502 14532 10508 14544
rect 10183 14504 10508 14532
rect 10183 14501 10195 14504
rect 10137 14495 10195 14501
rect 10502 14492 10508 14504
rect 10560 14492 10566 14544
rect 8573 14467 8631 14473
rect 8573 14433 8585 14467
rect 8619 14464 8631 14467
rect 8619 14436 10088 14464
rect 8619 14433 8631 14436
rect 8573 14427 8631 14433
rect 8662 14356 8668 14408
rect 8720 14396 8726 14408
rect 9950 14396 9956 14408
rect 8720 14368 9956 14396
rect 8720 14356 8726 14368
rect 9950 14356 9956 14368
rect 10008 14356 10014 14408
rect 9398 14328 9404 14340
rect 8496 14300 9404 14328
rect 9398 14288 9404 14300
rect 9456 14288 9462 14340
rect 9585 14331 9643 14337
rect 9585 14297 9597 14331
rect 9631 14328 9643 14331
rect 9674 14328 9680 14340
rect 9631 14300 9680 14328
rect 9631 14297 9643 14300
rect 9585 14291 9643 14297
rect 9674 14288 9680 14300
rect 9732 14288 9738 14340
rect 9861 14331 9919 14337
rect 9861 14297 9873 14331
rect 9907 14328 9919 14331
rect 10060 14328 10088 14436
rect 10226 14328 10232 14340
rect 9907 14300 10232 14328
rect 9907 14297 9919 14300
rect 9861 14291 9919 14297
rect 10226 14288 10232 14300
rect 10284 14328 10290 14340
rect 10870 14328 10876 14340
rect 10284 14300 10876 14328
rect 10284 14288 10290 14300
rect 10870 14288 10876 14300
rect 10928 14288 10934 14340
rect 8202 14260 8208 14272
rect 7767 14232 8208 14260
rect 8202 14220 8208 14232
rect 8260 14220 8266 14272
rect 8941 14263 8999 14269
rect 8941 14229 8953 14263
rect 8987 14260 8999 14263
rect 9030 14260 9036 14272
rect 8987 14232 9036 14260
rect 8987 14229 8999 14232
rect 8941 14223 8999 14229
rect 9030 14220 9036 14232
rect 9088 14220 9094 14272
rect 9217 14263 9275 14269
rect 9217 14229 9229 14263
rect 9263 14260 9275 14263
rect 9306 14260 9312 14272
rect 9263 14232 9312 14260
rect 9263 14229 9275 14232
rect 9217 14223 9275 14229
rect 9306 14220 9312 14232
rect 9364 14220 9370 14272
rect 10042 14220 10048 14272
rect 10100 14260 10106 14272
rect 10502 14260 10508 14272
rect 10100 14232 10508 14260
rect 10100 14220 10106 14232
rect 10502 14220 10508 14232
rect 10560 14220 10566 14272
rect 1104 14170 16008 14192
rect 1104 14118 3480 14170
rect 3532 14118 3544 14170
rect 3596 14118 3608 14170
rect 3660 14118 3672 14170
rect 3724 14118 8478 14170
rect 8530 14118 8542 14170
rect 8594 14118 8606 14170
rect 8658 14118 8670 14170
rect 8722 14118 13475 14170
rect 13527 14118 13539 14170
rect 13591 14118 13603 14170
rect 13655 14118 13667 14170
rect 13719 14118 16008 14170
rect 1104 14096 16008 14118
rect 2498 14056 2504 14068
rect 2459 14028 2504 14056
rect 2498 14016 2504 14028
rect 2556 14016 2562 14068
rect 2774 14016 2780 14068
rect 2832 14056 2838 14068
rect 2832 14028 2877 14056
rect 2832 14016 2838 14028
rect 5534 14016 5540 14068
rect 5592 14056 5598 14068
rect 8757 14059 8815 14065
rect 8757 14056 8769 14059
rect 5592 14028 8769 14056
rect 5592 14016 5598 14028
rect 8757 14025 8769 14028
rect 8803 14025 8815 14059
rect 8757 14019 8815 14025
rect 9490 14016 9496 14068
rect 9548 14056 9554 14068
rect 11330 14056 11336 14068
rect 9548 14028 11336 14056
rect 9548 14016 9554 14028
rect 11330 14016 11336 14028
rect 11388 14016 11394 14068
rect 4065 13991 4123 13997
rect 4065 13988 4077 13991
rect 2746 13960 4077 13988
rect 2746 13920 2774 13960
rect 4065 13957 4077 13960
rect 4111 13957 4123 13991
rect 4065 13951 4123 13957
rect 4356 13960 4936 13988
rect 2700 13892 2774 13920
rect 2700 13861 2728 13892
rect 3510 13880 3516 13932
rect 3568 13920 3574 13932
rect 4356 13920 4384 13960
rect 4522 13920 4528 13932
rect 3568 13892 4384 13920
rect 4483 13892 4528 13920
rect 3568 13880 3574 13892
rect 4522 13880 4528 13892
rect 4580 13880 4586 13932
rect 4706 13920 4712 13932
rect 4667 13892 4712 13920
rect 4706 13880 4712 13892
rect 4764 13880 4770 13932
rect 4908 13920 4936 13960
rect 6270 13948 6276 14000
rect 6328 13988 6334 14000
rect 6457 13991 6515 13997
rect 6457 13988 6469 13991
rect 6328 13960 6469 13988
rect 6328 13948 6334 13960
rect 6457 13957 6469 13960
rect 6503 13957 6515 13991
rect 7926 13988 7932 14000
rect 7887 13960 7932 13988
rect 6457 13951 6515 13957
rect 7926 13948 7932 13960
rect 7984 13948 7990 14000
rect 8202 13948 8208 14000
rect 8260 13988 8266 14000
rect 14182 13988 14188 14000
rect 8260 13960 14188 13988
rect 8260 13948 8266 13960
rect 14182 13948 14188 13960
rect 14240 13948 14246 14000
rect 4908 13892 5028 13920
rect 2685 13855 2743 13861
rect 2685 13821 2697 13855
rect 2731 13821 2743 13855
rect 2958 13852 2964 13864
rect 2919 13824 2964 13852
rect 2685 13815 2743 13821
rect 2958 13812 2964 13824
rect 3016 13812 3022 13864
rect 4890 13852 4896 13864
rect 4851 13824 4896 13852
rect 4890 13812 4896 13824
rect 4948 13812 4954 13864
rect 5000 13852 5028 13892
rect 6012 13892 6868 13920
rect 5149 13855 5207 13861
rect 5149 13852 5161 13855
rect 5000 13824 5161 13852
rect 5149 13821 5161 13824
rect 5195 13852 5207 13855
rect 5902 13852 5908 13864
rect 5195 13824 5908 13852
rect 5195 13821 5207 13824
rect 5149 13815 5207 13821
rect 5902 13812 5908 13824
rect 5960 13812 5966 13864
rect 2774 13744 2780 13796
rect 2832 13784 2838 13796
rect 6012 13784 6040 13892
rect 6270 13812 6276 13864
rect 6328 13852 6334 13864
rect 6730 13852 6736 13864
rect 6328 13824 6736 13852
rect 6328 13812 6334 13824
rect 6730 13812 6736 13824
rect 6788 13812 6794 13864
rect 6840 13852 6868 13892
rect 8110 13880 8116 13932
rect 8168 13920 8174 13932
rect 8481 13923 8539 13929
rect 8481 13920 8493 13923
rect 8168 13892 8493 13920
rect 8168 13880 8174 13892
rect 8481 13889 8493 13892
rect 8527 13889 8539 13923
rect 8481 13883 8539 13889
rect 9030 13880 9036 13932
rect 9088 13920 9094 13932
rect 9217 13923 9275 13929
rect 9217 13920 9229 13923
rect 9088 13892 9229 13920
rect 9088 13880 9094 13892
rect 9217 13889 9229 13892
rect 9263 13889 9275 13923
rect 9217 13883 9275 13889
rect 9309 13923 9367 13929
rect 9309 13889 9321 13923
rect 9355 13920 9367 13923
rect 10229 13923 10287 13929
rect 10229 13920 10241 13923
rect 9355 13892 10241 13920
rect 9355 13889 9367 13892
rect 9309 13883 9367 13889
rect 10229 13889 10241 13892
rect 10275 13920 10287 13923
rect 12342 13920 12348 13932
rect 10275 13892 12348 13920
rect 10275 13889 10287 13892
rect 10229 13883 10287 13889
rect 7098 13852 7104 13864
rect 6840 13824 7104 13852
rect 7098 13812 7104 13824
rect 7156 13812 7162 13864
rect 7581 13855 7639 13861
rect 7581 13821 7593 13855
rect 7627 13821 7639 13855
rect 7834 13852 7840 13864
rect 7795 13824 7840 13852
rect 7581 13815 7639 13821
rect 2832 13756 6040 13784
rect 7596 13784 7624 13815
rect 7834 13812 7840 13824
rect 7892 13812 7898 13864
rect 8386 13852 8392 13864
rect 8128 13824 8392 13852
rect 8128 13784 8156 13824
rect 8386 13812 8392 13824
rect 8444 13852 8450 13864
rect 9324 13852 9352 13883
rect 12342 13880 12348 13892
rect 12400 13880 12406 13932
rect 10045 13855 10103 13861
rect 8444 13824 9352 13852
rect 9508 13824 9674 13852
rect 8444 13812 8450 13824
rect 7596 13756 8156 13784
rect 2832 13744 2838 13756
rect 8202 13744 8208 13796
rect 8260 13784 8266 13796
rect 8297 13787 8355 13793
rect 8297 13784 8309 13787
rect 8260 13756 8309 13784
rect 8260 13744 8266 13756
rect 8297 13753 8309 13756
rect 8343 13784 8355 13787
rect 8343 13756 8616 13784
rect 8343 13753 8355 13756
rect 8297 13747 8355 13753
rect 2498 13676 2504 13728
rect 2556 13716 2562 13728
rect 4433 13719 4491 13725
rect 4433 13716 4445 13719
rect 2556 13688 4445 13716
rect 2556 13676 2562 13688
rect 4433 13685 4445 13688
rect 4479 13685 4491 13719
rect 4433 13679 4491 13685
rect 5626 13676 5632 13728
rect 5684 13716 5690 13728
rect 6273 13719 6331 13725
rect 6273 13716 6285 13719
rect 5684 13688 6285 13716
rect 5684 13676 5690 13688
rect 6273 13685 6285 13688
rect 6319 13685 6331 13719
rect 6273 13679 6331 13685
rect 7558 13676 7564 13728
rect 7616 13716 7622 13728
rect 8389 13719 8447 13725
rect 8389 13716 8401 13719
rect 7616 13688 8401 13716
rect 7616 13676 7622 13688
rect 8389 13685 8401 13688
rect 8435 13716 8447 13719
rect 8478 13716 8484 13728
rect 8435 13688 8484 13716
rect 8435 13685 8447 13688
rect 8389 13679 8447 13685
rect 8478 13676 8484 13688
rect 8536 13676 8542 13728
rect 8588 13716 8616 13756
rect 8662 13744 8668 13796
rect 8720 13784 8726 13796
rect 9508 13784 9536 13824
rect 8720 13756 9536 13784
rect 9646 13784 9674 13824
rect 10045 13821 10057 13855
rect 10091 13852 10103 13855
rect 14274 13852 14280 13864
rect 10091 13824 14280 13852
rect 10091 13821 10103 13824
rect 10045 13815 10103 13821
rect 14274 13812 14280 13824
rect 14332 13852 14338 13864
rect 14458 13852 14464 13864
rect 14332 13824 14464 13852
rect 14332 13812 14338 13824
rect 14458 13812 14464 13824
rect 14516 13812 14522 13864
rect 11698 13784 11704 13796
rect 9646 13756 11704 13784
rect 8720 13744 8726 13756
rect 11698 13744 11704 13756
rect 11756 13744 11762 13796
rect 8938 13716 8944 13728
rect 8588 13688 8944 13716
rect 8938 13676 8944 13688
rect 8996 13676 9002 13728
rect 9122 13716 9128 13728
rect 9083 13688 9128 13716
rect 9122 13676 9128 13688
rect 9180 13676 9186 13728
rect 9306 13676 9312 13728
rect 9364 13716 9370 13728
rect 9585 13719 9643 13725
rect 9585 13716 9597 13719
rect 9364 13688 9597 13716
rect 9364 13676 9370 13688
rect 9585 13685 9597 13688
rect 9631 13685 9643 13719
rect 9585 13679 9643 13685
rect 9674 13676 9680 13728
rect 9732 13716 9738 13728
rect 9953 13719 10011 13725
rect 9953 13716 9965 13719
rect 9732 13688 9965 13716
rect 9732 13676 9738 13688
rect 9953 13685 9965 13688
rect 9999 13685 10011 13719
rect 10410 13716 10416 13728
rect 10371 13688 10416 13716
rect 9953 13679 10011 13685
rect 10410 13676 10416 13688
rect 10468 13676 10474 13728
rect 10502 13676 10508 13728
rect 10560 13716 10566 13728
rect 10597 13719 10655 13725
rect 10597 13716 10609 13719
rect 10560 13688 10609 13716
rect 10560 13676 10566 13688
rect 10597 13685 10609 13688
rect 10643 13685 10655 13719
rect 10597 13679 10655 13685
rect 14458 13676 14464 13728
rect 14516 13716 14522 13728
rect 14826 13716 14832 13728
rect 14516 13688 14832 13716
rect 14516 13676 14522 13688
rect 14826 13676 14832 13688
rect 14884 13676 14890 13728
rect 1104 13626 16008 13648
rect 1104 13574 5979 13626
rect 6031 13574 6043 13626
rect 6095 13574 6107 13626
rect 6159 13574 6171 13626
rect 6223 13574 10976 13626
rect 11028 13574 11040 13626
rect 11092 13574 11104 13626
rect 11156 13574 11168 13626
rect 11220 13574 16008 13626
rect 1104 13552 16008 13574
rect 2593 13515 2651 13521
rect 2593 13481 2605 13515
rect 2639 13481 2651 13515
rect 3418 13512 3424 13524
rect 3379 13484 3424 13512
rect 2593 13475 2651 13481
rect 1581 13447 1639 13453
rect 1581 13413 1593 13447
rect 1627 13444 1639 13447
rect 2608 13444 2636 13475
rect 3418 13472 3424 13484
rect 3476 13472 3482 13524
rect 3878 13512 3884 13524
rect 3839 13484 3884 13512
rect 3878 13472 3884 13484
rect 3936 13472 3942 13524
rect 4525 13515 4583 13521
rect 4525 13481 4537 13515
rect 4571 13512 4583 13515
rect 4890 13512 4896 13524
rect 4571 13484 4896 13512
rect 4571 13481 4583 13484
rect 4525 13475 4583 13481
rect 4890 13472 4896 13484
rect 4948 13472 4954 13524
rect 8297 13515 8355 13521
rect 6472 13484 8248 13512
rect 6472 13444 6500 13484
rect 1627 13416 2636 13444
rect 4080 13416 6500 13444
rect 6580 13447 6638 13453
rect 1627 13413 1639 13416
rect 1581 13407 1639 13413
rect 1394 13376 1400 13388
rect 1355 13348 1400 13376
rect 1394 13336 1400 13348
rect 1452 13336 1458 13388
rect 2590 13336 2596 13388
rect 2648 13376 2654 13388
rect 4080 13385 4108 13416
rect 6580 13413 6592 13447
rect 6626 13444 6638 13447
rect 6822 13444 6828 13456
rect 6626 13416 6828 13444
rect 6626 13413 6638 13416
rect 6580 13407 6638 13413
rect 6822 13404 6828 13416
rect 6880 13404 6886 13456
rect 7190 13453 7196 13456
rect 7184 13407 7196 13453
rect 7248 13444 7254 13456
rect 8018 13444 8024 13456
rect 7248 13416 8024 13444
rect 7190 13404 7196 13407
rect 7248 13404 7254 13416
rect 8018 13404 8024 13416
rect 8076 13404 8082 13456
rect 8220 13444 8248 13484
rect 8297 13481 8309 13515
rect 8343 13512 8355 13515
rect 8386 13512 8392 13524
rect 8343 13484 8392 13512
rect 8343 13481 8355 13484
rect 8297 13475 8355 13481
rect 8386 13472 8392 13484
rect 8444 13472 8450 13524
rect 8662 13512 8668 13524
rect 8496 13484 8668 13512
rect 8496 13444 8524 13484
rect 8662 13472 8668 13484
rect 8720 13472 8726 13524
rect 8849 13515 8907 13521
rect 8849 13481 8861 13515
rect 8895 13512 8907 13515
rect 9030 13512 9036 13524
rect 8895 13484 9036 13512
rect 8895 13481 8907 13484
rect 8849 13475 8907 13481
rect 9030 13472 9036 13484
rect 9088 13472 9094 13524
rect 9858 13472 9864 13524
rect 9916 13512 9922 13524
rect 9953 13515 10011 13521
rect 9953 13512 9965 13515
rect 9916 13484 9965 13512
rect 9916 13472 9922 13484
rect 9953 13481 9965 13484
rect 9999 13481 10011 13515
rect 9953 13475 10011 13481
rect 10226 13472 10232 13524
rect 10284 13512 10290 13524
rect 10413 13515 10471 13521
rect 10413 13512 10425 13515
rect 10284 13484 10425 13512
rect 10284 13472 10290 13484
rect 10413 13481 10425 13484
rect 10459 13512 10471 13515
rect 10778 13512 10784 13524
rect 10459 13484 10784 13512
rect 10459 13481 10471 13484
rect 10413 13475 10471 13481
rect 10778 13472 10784 13484
rect 10836 13512 10842 13524
rect 11606 13512 11612 13524
rect 10836 13484 11612 13512
rect 10836 13472 10842 13484
rect 11606 13472 11612 13484
rect 11664 13472 11670 13524
rect 8220 13416 8524 13444
rect 8573 13447 8631 13453
rect 8573 13413 8585 13447
rect 8619 13444 8631 13447
rect 8938 13444 8944 13456
rect 8619 13416 8944 13444
rect 8619 13413 8631 13416
rect 8573 13407 8631 13413
rect 8938 13404 8944 13416
rect 8996 13404 9002 13456
rect 9398 13404 9404 13456
rect 9456 13444 9462 13456
rect 9582 13444 9588 13456
rect 9456 13416 9588 13444
rect 9456 13404 9462 13416
rect 9582 13404 9588 13416
rect 9640 13404 9646 13456
rect 11054 13444 11060 13456
rect 10888 13416 11060 13444
rect 2777 13379 2835 13385
rect 2777 13376 2789 13379
rect 2648 13348 2789 13376
rect 2648 13336 2654 13348
rect 2777 13345 2789 13348
rect 2823 13345 2835 13379
rect 2777 13339 2835 13345
rect 3329 13379 3387 13385
rect 3329 13345 3341 13379
rect 3375 13376 3387 13379
rect 4065 13379 4123 13385
rect 3375 13348 4016 13376
rect 3375 13345 3387 13348
rect 3329 13339 3387 13345
rect 3050 13268 3056 13320
rect 3108 13308 3114 13320
rect 3510 13308 3516 13320
rect 3108 13280 3516 13308
rect 3108 13268 3114 13280
rect 3510 13268 3516 13280
rect 3568 13268 3574 13320
rect 2130 13132 2136 13184
rect 2188 13172 2194 13184
rect 2961 13175 3019 13181
rect 2961 13172 2973 13175
rect 2188 13144 2973 13172
rect 2188 13132 2194 13144
rect 2961 13141 2973 13144
rect 3007 13141 3019 13175
rect 3988 13172 4016 13348
rect 4065 13345 4077 13379
rect 4111 13345 4123 13379
rect 4065 13339 4123 13345
rect 4341 13379 4399 13385
rect 4341 13345 4353 13379
rect 4387 13376 4399 13379
rect 4614 13376 4620 13388
rect 4387 13348 4620 13376
rect 4387 13345 4399 13348
rect 4341 13339 4399 13345
rect 4614 13336 4620 13348
rect 4672 13336 4678 13388
rect 4985 13379 5043 13385
rect 4985 13345 4997 13379
rect 5031 13376 5043 13379
rect 5031 13348 7972 13376
rect 5031 13345 5043 13348
rect 4985 13339 5043 13345
rect 4246 13268 4252 13320
rect 4304 13308 4310 13320
rect 5077 13311 5135 13317
rect 5077 13308 5089 13311
rect 4304 13280 5089 13308
rect 4304 13268 4310 13280
rect 5077 13277 5089 13280
rect 5123 13277 5135 13311
rect 5077 13271 5135 13277
rect 5261 13311 5319 13317
rect 5261 13277 5273 13311
rect 5307 13308 5319 13311
rect 5810 13308 5816 13320
rect 5307 13280 5816 13308
rect 5307 13277 5319 13280
rect 5261 13271 5319 13277
rect 5810 13268 5816 13280
rect 5868 13268 5874 13320
rect 6825 13311 6883 13317
rect 6825 13277 6837 13311
rect 6871 13308 6883 13311
rect 6917 13311 6975 13317
rect 6917 13308 6929 13311
rect 6871 13280 6929 13308
rect 6871 13277 6883 13280
rect 6825 13271 6883 13277
rect 6917 13277 6929 13280
rect 6963 13277 6975 13311
rect 6917 13271 6975 13277
rect 4154 13200 4160 13252
rect 4212 13240 4218 13252
rect 4617 13243 4675 13249
rect 4617 13240 4629 13243
rect 4212 13212 4629 13240
rect 4212 13200 4218 13212
rect 4617 13209 4629 13212
rect 4663 13209 4675 13243
rect 4617 13203 4675 13209
rect 4982 13172 4988 13184
rect 3988 13144 4988 13172
rect 2961 13135 3019 13141
rect 4982 13132 4988 13144
rect 5040 13132 5046 13184
rect 5442 13172 5448 13184
rect 5403 13144 5448 13172
rect 5442 13132 5448 13144
rect 5500 13132 5506 13184
rect 6932 13172 6960 13271
rect 7650 13172 7656 13184
rect 6932 13144 7656 13172
rect 7650 13132 7656 13144
rect 7708 13172 7714 13184
rect 7834 13172 7840 13184
rect 7708 13144 7840 13172
rect 7708 13132 7714 13144
rect 7834 13132 7840 13144
rect 7892 13132 7898 13184
rect 7944 13172 7972 13348
rect 8846 13336 8852 13388
rect 8904 13376 8910 13388
rect 9493 13379 9551 13385
rect 9493 13376 9505 13379
rect 8904 13348 9505 13376
rect 8904 13336 8910 13348
rect 9493 13345 9505 13348
rect 9539 13376 9551 13379
rect 9766 13376 9772 13388
rect 9539 13348 9772 13376
rect 9539 13345 9551 13348
rect 9493 13339 9551 13345
rect 9766 13336 9772 13348
rect 9824 13336 9830 13388
rect 10321 13379 10379 13385
rect 10321 13345 10333 13379
rect 10367 13376 10379 13379
rect 10888 13376 10916 13416
rect 11054 13404 11060 13416
rect 11112 13404 11118 13456
rect 10367 13348 10916 13376
rect 10965 13379 11023 13385
rect 10367 13345 10379 13348
rect 10321 13339 10379 13345
rect 10965 13345 10977 13379
rect 11011 13376 11023 13379
rect 11330 13376 11336 13388
rect 11011 13348 11336 13376
rect 11011 13345 11023 13348
rect 10965 13339 11023 13345
rect 11330 13336 11336 13348
rect 11388 13336 11394 13388
rect 8864 13280 9352 13308
rect 8864 13252 8892 13280
rect 8846 13200 8852 13252
rect 8904 13200 8910 13252
rect 9122 13240 9128 13252
rect 9083 13212 9128 13240
rect 9122 13200 9128 13212
rect 9180 13200 9186 13252
rect 9324 13240 9352 13280
rect 9398 13268 9404 13320
rect 9456 13308 9462 13320
rect 9585 13311 9643 13317
rect 9585 13308 9597 13311
rect 9456 13280 9597 13308
rect 9456 13268 9462 13280
rect 9585 13277 9597 13280
rect 9631 13277 9643 13311
rect 9585 13271 9643 13277
rect 9677 13311 9735 13317
rect 9677 13277 9689 13311
rect 9723 13277 9735 13311
rect 10597 13311 10655 13317
rect 9677 13271 9735 13277
rect 9968 13280 10548 13308
rect 9692 13240 9720 13271
rect 9858 13240 9864 13252
rect 9324 13212 9864 13240
rect 9858 13200 9864 13212
rect 9916 13200 9922 13252
rect 9968 13172 9996 13280
rect 10520 13252 10548 13280
rect 10597 13277 10609 13311
rect 10643 13308 10655 13311
rect 12342 13308 12348 13320
rect 10643 13280 12348 13308
rect 10643 13277 10655 13280
rect 10597 13271 10655 13277
rect 12342 13268 12348 13280
rect 12400 13268 12406 13320
rect 10502 13200 10508 13252
rect 10560 13200 10566 13252
rect 11333 13243 11391 13249
rect 11333 13209 11345 13243
rect 11379 13240 11391 13243
rect 11606 13240 11612 13252
rect 11379 13212 11612 13240
rect 11379 13209 11391 13212
rect 11333 13203 11391 13209
rect 11606 13200 11612 13212
rect 11664 13200 11670 13252
rect 7944 13144 9996 13172
rect 10042 13132 10048 13184
rect 10100 13172 10106 13184
rect 10781 13175 10839 13181
rect 10781 13172 10793 13175
rect 10100 13144 10793 13172
rect 10100 13132 10106 13144
rect 10781 13141 10793 13144
rect 10827 13141 10839 13175
rect 11146 13172 11152 13184
rect 11107 13144 11152 13172
rect 10781 13135 10839 13141
rect 11146 13132 11152 13144
rect 11204 13132 11210 13184
rect 11238 13132 11244 13184
rect 11296 13172 11302 13184
rect 11422 13172 11428 13184
rect 11296 13144 11428 13172
rect 11296 13132 11302 13144
rect 11422 13132 11428 13144
rect 11480 13132 11486 13184
rect 1104 13082 16008 13104
rect 1104 13030 3480 13082
rect 3532 13030 3544 13082
rect 3596 13030 3608 13082
rect 3660 13030 3672 13082
rect 3724 13030 8478 13082
rect 8530 13030 8542 13082
rect 8594 13030 8606 13082
rect 8658 13030 8670 13082
rect 8722 13030 13475 13082
rect 13527 13030 13539 13082
rect 13591 13030 13603 13082
rect 13655 13030 13667 13082
rect 13719 13030 16008 13082
rect 1104 13008 16008 13030
rect 2590 12968 2596 12980
rect 2551 12940 2596 12968
rect 2590 12928 2596 12940
rect 2648 12928 2654 12980
rect 5626 12968 5632 12980
rect 3160 12940 5632 12968
rect 2501 12903 2559 12909
rect 2501 12869 2513 12903
rect 2547 12900 2559 12903
rect 2958 12900 2964 12912
rect 2547 12872 2964 12900
rect 2547 12869 2559 12872
rect 2501 12863 2559 12869
rect 2958 12860 2964 12872
rect 3016 12860 3022 12912
rect 1949 12835 2007 12841
rect 1949 12801 1961 12835
rect 1995 12832 2007 12835
rect 3160 12832 3188 12940
rect 5626 12928 5632 12940
rect 5684 12928 5690 12980
rect 6273 12971 6331 12977
rect 6273 12937 6285 12971
rect 6319 12968 6331 12971
rect 7190 12968 7196 12980
rect 6319 12940 7196 12968
rect 6319 12937 6331 12940
rect 6273 12931 6331 12937
rect 7190 12928 7196 12940
rect 7248 12928 7254 12980
rect 7837 12971 7895 12977
rect 7837 12937 7849 12971
rect 7883 12968 7895 12971
rect 8110 12968 8116 12980
rect 7883 12940 8116 12968
rect 7883 12937 7895 12940
rect 7837 12931 7895 12937
rect 8110 12928 8116 12940
rect 8168 12968 8174 12980
rect 8168 12940 9085 12968
rect 8168 12928 8174 12940
rect 9057 12844 9085 12940
rect 9674 12928 9680 12980
rect 9732 12968 9738 12980
rect 10042 12968 10048 12980
rect 9732 12940 10048 12968
rect 9732 12928 9738 12940
rect 10042 12928 10048 12940
rect 10100 12928 10106 12980
rect 11422 12968 11428 12980
rect 11383 12940 11428 12968
rect 11422 12928 11428 12940
rect 11480 12928 11486 12980
rect 9122 12860 9128 12912
rect 9180 12900 9186 12912
rect 9309 12903 9367 12909
rect 9309 12900 9321 12903
rect 9180 12872 9321 12900
rect 9180 12860 9186 12872
rect 9309 12869 9321 12872
rect 9355 12869 9367 12903
rect 9309 12863 9367 12869
rect 10229 12903 10287 12909
rect 10229 12869 10241 12903
rect 10275 12900 10287 12903
rect 10594 12900 10600 12912
rect 10275 12872 10600 12900
rect 10275 12869 10287 12872
rect 10229 12863 10287 12869
rect 10594 12860 10600 12872
rect 10652 12860 10658 12912
rect 14458 12900 14464 12912
rect 10704 12872 14464 12900
rect 1995 12804 3188 12832
rect 3237 12835 3295 12841
rect 1995 12801 2007 12804
rect 1949 12795 2007 12801
rect 3237 12801 3249 12835
rect 3283 12801 3295 12835
rect 9030 12832 9036 12844
rect 8952 12804 9036 12832
rect 3237 12795 3295 12801
rect 2130 12764 2136 12776
rect 2091 12736 2136 12764
rect 2130 12724 2136 12736
rect 2188 12724 2194 12776
rect 2774 12724 2780 12776
rect 2832 12764 2838 12776
rect 2961 12767 3019 12773
rect 2961 12764 2973 12767
rect 2832 12736 2973 12764
rect 2832 12724 2838 12736
rect 2961 12733 2973 12736
rect 3007 12733 3019 12767
rect 3252 12764 3280 12795
rect 9030 12792 9036 12804
rect 9088 12832 9094 12844
rect 10704 12841 10732 12872
rect 14458 12860 14464 12872
rect 14516 12860 14522 12912
rect 9953 12835 10011 12841
rect 9953 12832 9965 12835
rect 9088 12804 9965 12832
rect 9088 12792 9094 12804
rect 9953 12801 9965 12804
rect 9999 12801 10011 12835
rect 9953 12795 10011 12801
rect 10689 12835 10747 12841
rect 10689 12801 10701 12835
rect 10735 12801 10747 12835
rect 10870 12832 10876 12844
rect 10831 12804 10876 12832
rect 10689 12795 10747 12801
rect 10870 12792 10876 12804
rect 10928 12792 10934 12844
rect 11333 12835 11391 12841
rect 11333 12801 11345 12835
rect 11379 12832 11391 12835
rect 11606 12832 11612 12844
rect 11379 12804 11612 12832
rect 11379 12801 11391 12804
rect 11333 12795 11391 12801
rect 11606 12792 11612 12804
rect 11664 12832 11670 12844
rect 12434 12832 12440 12844
rect 11664 12804 12440 12832
rect 11664 12792 11670 12804
rect 12434 12792 12440 12804
rect 12492 12792 12498 12844
rect 4801 12767 4859 12773
rect 3252 12736 4660 12764
rect 2961 12727 3019 12733
rect 3053 12699 3111 12705
rect 3053 12665 3065 12699
rect 3099 12696 3111 12699
rect 3510 12696 3516 12708
rect 3099 12668 3516 12696
rect 3099 12665 3111 12668
rect 3053 12659 3111 12665
rect 3510 12656 3516 12668
rect 3568 12656 3574 12708
rect 3602 12656 3608 12708
rect 3660 12696 3666 12708
rect 4062 12696 4068 12708
rect 3660 12668 4068 12696
rect 3660 12656 3666 12668
rect 4062 12656 4068 12668
rect 4120 12656 4126 12708
rect 4522 12696 4528 12708
rect 4580 12705 4586 12708
rect 4492 12668 4528 12696
rect 4522 12656 4528 12668
rect 4580 12659 4592 12705
rect 4632 12696 4660 12736
rect 4801 12733 4813 12767
rect 4847 12764 4859 12767
rect 4890 12764 4896 12776
rect 4847 12736 4896 12764
rect 4847 12733 4859 12736
rect 4801 12727 4859 12733
rect 4890 12724 4896 12736
rect 4948 12724 4954 12776
rect 6454 12764 6460 12776
rect 6367 12736 6460 12764
rect 6454 12724 6460 12736
rect 6512 12764 6518 12776
rect 7650 12764 7656 12776
rect 6512 12736 7656 12764
rect 6512 12724 6518 12736
rect 7650 12724 7656 12736
rect 7708 12764 7714 12776
rect 7834 12764 7840 12776
rect 7708 12736 7840 12764
rect 7708 12724 7714 12736
rect 7834 12724 7840 12736
rect 7892 12764 7898 12776
rect 7929 12767 7987 12773
rect 7929 12764 7941 12767
rect 7892 12736 7941 12764
rect 7892 12724 7898 12736
rect 7929 12733 7941 12736
rect 7975 12764 7987 12767
rect 9674 12764 9680 12776
rect 7975 12736 9680 12764
rect 7975 12733 7987 12736
rect 7929 12727 7987 12733
rect 9674 12724 9680 12736
rect 9732 12724 9738 12776
rect 9766 12724 9772 12776
rect 9824 12764 9830 12776
rect 10410 12764 10416 12776
rect 9824 12736 10416 12764
rect 9824 12724 9830 12736
rect 10410 12724 10416 12736
rect 10468 12764 10474 12776
rect 11885 12767 11943 12773
rect 11885 12764 11897 12767
rect 10468 12736 11897 12764
rect 10468 12724 10474 12736
rect 11885 12733 11897 12736
rect 11931 12764 11943 12767
rect 12158 12764 12164 12776
rect 11931 12736 12164 12764
rect 11931 12733 11943 12736
rect 11885 12727 11943 12733
rect 12158 12724 12164 12736
rect 12216 12724 12222 12776
rect 12250 12724 12256 12776
rect 12308 12764 12314 12776
rect 14090 12764 14096 12776
rect 12308 12736 14096 12764
rect 12308 12724 12314 12736
rect 14090 12724 14096 12736
rect 14148 12724 14154 12776
rect 5138 12699 5196 12705
rect 5138 12696 5150 12699
rect 4632 12668 5150 12696
rect 5138 12665 5150 12668
rect 5184 12696 5196 12699
rect 5442 12696 5448 12708
rect 5184 12668 5448 12696
rect 5184 12665 5196 12668
rect 5138 12659 5196 12665
rect 4580 12656 4586 12659
rect 5442 12656 5448 12668
rect 5500 12656 5506 12708
rect 5810 12656 5816 12708
rect 5868 12696 5874 12708
rect 6702 12699 6760 12705
rect 6702 12696 6714 12699
rect 5868 12668 6714 12696
rect 5868 12656 5874 12668
rect 6702 12665 6714 12668
rect 6748 12665 6760 12699
rect 6702 12659 6760 12665
rect 8018 12656 8024 12708
rect 8076 12696 8082 12708
rect 8174 12699 8232 12705
rect 8174 12696 8186 12699
rect 8076 12668 8186 12696
rect 8076 12656 8082 12668
rect 8174 12665 8186 12668
rect 8220 12665 8232 12699
rect 8174 12659 8232 12665
rect 8754 12656 8760 12708
rect 8812 12696 8818 12708
rect 8938 12696 8944 12708
rect 8812 12668 8944 12696
rect 8812 12656 8818 12668
rect 8938 12656 8944 12668
rect 8996 12656 9002 12708
rect 9858 12696 9864 12708
rect 9232 12668 9536 12696
rect 9819 12668 9864 12696
rect 2038 12628 2044 12640
rect 1999 12600 2044 12628
rect 2038 12588 2044 12600
rect 2096 12588 2102 12640
rect 3421 12631 3479 12637
rect 3421 12597 3433 12631
rect 3467 12628 3479 12631
rect 4706 12628 4712 12640
rect 3467 12600 4712 12628
rect 3467 12597 3479 12600
rect 3421 12591 3479 12597
rect 4706 12588 4712 12600
rect 4764 12588 4770 12640
rect 4982 12588 4988 12640
rect 5040 12628 5046 12640
rect 9232 12628 9260 12668
rect 5040 12600 9260 12628
rect 5040 12588 5046 12600
rect 9306 12588 9312 12640
rect 9364 12628 9370 12640
rect 9401 12631 9459 12637
rect 9401 12628 9413 12631
rect 9364 12600 9413 12628
rect 9364 12588 9370 12600
rect 9401 12597 9413 12600
rect 9447 12597 9459 12631
rect 9508 12628 9536 12668
rect 9858 12656 9864 12668
rect 9916 12656 9922 12708
rect 10428 12668 11192 12696
rect 10428 12628 10456 12668
rect 10594 12628 10600 12640
rect 9508 12600 10456 12628
rect 10555 12600 10600 12628
rect 9401 12591 9459 12597
rect 10594 12588 10600 12600
rect 10652 12588 10658 12640
rect 10778 12588 10784 12640
rect 10836 12628 10842 12640
rect 11057 12631 11115 12637
rect 11057 12628 11069 12631
rect 10836 12600 11069 12628
rect 10836 12588 10842 12600
rect 11057 12597 11069 12600
rect 11103 12597 11115 12631
rect 11164 12628 11192 12668
rect 11238 12656 11244 12708
rect 11296 12696 11302 12708
rect 11514 12696 11520 12708
rect 11296 12668 11520 12696
rect 11296 12656 11302 12668
rect 11514 12656 11520 12668
rect 11572 12656 11578 12708
rect 11793 12699 11851 12705
rect 11793 12665 11805 12699
rect 11839 12696 11851 12699
rect 11974 12696 11980 12708
rect 11839 12668 11980 12696
rect 11839 12665 11851 12668
rect 11793 12659 11851 12665
rect 11974 12656 11980 12668
rect 12032 12656 12038 12708
rect 12250 12628 12256 12640
rect 11164 12600 12256 12628
rect 11057 12591 11115 12597
rect 12250 12588 12256 12600
rect 12308 12588 12314 12640
rect 1104 12538 16008 12560
rect 1104 12486 5979 12538
rect 6031 12486 6043 12538
rect 6095 12486 6107 12538
rect 6159 12486 6171 12538
rect 6223 12486 10976 12538
rect 11028 12486 11040 12538
rect 11092 12486 11104 12538
rect 11156 12486 11168 12538
rect 11220 12486 16008 12538
rect 1104 12464 16008 12486
rect 1857 12427 1915 12433
rect 1857 12393 1869 12427
rect 1903 12393 1915 12427
rect 3329 12427 3387 12433
rect 1857 12387 1915 12393
rect 2056 12396 3096 12424
rect 1394 12356 1400 12368
rect 1355 12328 1400 12356
rect 1394 12316 1400 12328
rect 1452 12316 1458 12368
rect 1581 12359 1639 12365
rect 1581 12325 1593 12359
rect 1627 12356 1639 12359
rect 1872 12356 1900 12387
rect 1627 12328 1900 12356
rect 1627 12325 1639 12328
rect 1581 12319 1639 12325
rect 2056 12297 2084 12396
rect 3068 12356 3096 12396
rect 3329 12393 3341 12427
rect 3375 12424 3387 12427
rect 3602 12424 3608 12436
rect 3375 12396 3608 12424
rect 3375 12393 3387 12396
rect 3329 12387 3387 12393
rect 3602 12384 3608 12396
rect 3660 12384 3666 12436
rect 3697 12427 3755 12433
rect 3697 12393 3709 12427
rect 3743 12424 3755 12427
rect 3878 12424 3884 12436
rect 3743 12396 3884 12424
rect 3743 12393 3755 12396
rect 3697 12387 3755 12393
rect 3878 12384 3884 12396
rect 3936 12384 3942 12436
rect 4062 12424 4068 12436
rect 4023 12396 4068 12424
rect 4062 12384 4068 12396
rect 4120 12384 4126 12436
rect 4430 12384 4436 12436
rect 4488 12424 4494 12436
rect 5258 12424 5264 12436
rect 4488 12396 5264 12424
rect 4488 12384 4494 12396
rect 5258 12384 5264 12396
rect 5316 12384 5322 12436
rect 5810 12384 5816 12436
rect 5868 12424 5874 12436
rect 5997 12427 6055 12433
rect 5997 12424 6009 12427
rect 5868 12396 6009 12424
rect 5868 12384 5874 12396
rect 5997 12393 6009 12396
rect 6043 12393 6055 12427
rect 5997 12387 6055 12393
rect 6089 12427 6147 12433
rect 6089 12393 6101 12427
rect 6135 12424 6147 12427
rect 6730 12424 6736 12436
rect 6135 12396 6736 12424
rect 6135 12393 6147 12396
rect 6089 12387 6147 12393
rect 4154 12356 4160 12368
rect 3068 12328 4160 12356
rect 4154 12316 4160 12328
rect 4212 12316 4218 12368
rect 4525 12359 4583 12365
rect 4525 12325 4537 12359
rect 4571 12356 4583 12359
rect 5902 12356 5908 12368
rect 4571 12328 5908 12356
rect 4571 12325 4583 12328
rect 4525 12319 4583 12325
rect 5902 12316 5908 12328
rect 5960 12316 5966 12368
rect 2041 12291 2099 12297
rect 2041 12257 2053 12291
rect 2087 12257 2099 12291
rect 2041 12251 2099 12257
rect 2501 12291 2559 12297
rect 2501 12257 2513 12291
rect 2547 12288 2559 12291
rect 3142 12288 3148 12300
rect 2547 12260 3148 12288
rect 2547 12257 2559 12260
rect 2501 12251 2559 12257
rect 3142 12248 3148 12260
rect 3200 12248 3206 12300
rect 4249 12291 4307 12297
rect 4249 12257 4261 12291
rect 4295 12288 4307 12291
rect 4884 12291 4942 12297
rect 4884 12288 4896 12291
rect 4295 12260 4384 12288
rect 4295 12257 4307 12260
rect 4249 12251 4307 12257
rect 4356 12232 4384 12260
rect 4448 12260 4896 12288
rect 2314 12220 2320 12232
rect 2275 12192 2320 12220
rect 2314 12180 2320 12192
rect 2372 12180 2378 12232
rect 2406 12180 2412 12232
rect 2464 12220 2470 12232
rect 3053 12223 3111 12229
rect 2464 12192 2509 12220
rect 2464 12180 2470 12192
rect 3053 12189 3065 12223
rect 3099 12189 3111 12223
rect 3234 12220 3240 12232
rect 3195 12192 3240 12220
rect 3053 12183 3111 12189
rect 2590 12112 2596 12164
rect 2648 12152 2654 12164
rect 2869 12155 2927 12161
rect 2869 12152 2881 12155
rect 2648 12124 2881 12152
rect 2648 12112 2654 12124
rect 2869 12121 2881 12124
rect 2915 12121 2927 12155
rect 2869 12115 2927 12121
rect 3068 12084 3096 12183
rect 3234 12180 3240 12192
rect 3292 12180 3298 12232
rect 4338 12180 4344 12232
rect 4396 12180 4402 12232
rect 3142 12112 3148 12164
rect 3200 12152 3206 12164
rect 4448 12152 4476 12260
rect 4884 12257 4896 12260
rect 4930 12288 4942 12291
rect 6104 12288 6132 12387
rect 6730 12384 6736 12396
rect 6788 12384 6794 12436
rect 6822 12384 6828 12436
rect 6880 12424 6886 12436
rect 7561 12427 7619 12433
rect 7561 12424 7573 12427
rect 6880 12396 7573 12424
rect 6880 12384 6886 12396
rect 7561 12393 7573 12396
rect 7607 12393 7619 12427
rect 7561 12387 7619 12393
rect 7742 12384 7748 12436
rect 7800 12424 7806 12436
rect 10597 12427 10655 12433
rect 10597 12424 10609 12427
rect 7800 12396 10609 12424
rect 7800 12384 7806 12396
rect 10597 12393 10609 12396
rect 10643 12393 10655 12427
rect 10597 12387 10655 12393
rect 10686 12384 10692 12436
rect 10744 12424 10750 12436
rect 10965 12427 11023 12433
rect 10965 12424 10977 12427
rect 10744 12396 10977 12424
rect 10744 12384 10750 12396
rect 10965 12393 10977 12396
rect 11011 12393 11023 12427
rect 10965 12387 11023 12393
rect 11057 12427 11115 12433
rect 11057 12393 11069 12427
rect 11103 12424 11115 12427
rect 11422 12424 11428 12436
rect 11103 12396 11428 12424
rect 11103 12393 11115 12396
rect 11057 12387 11115 12393
rect 11422 12384 11428 12396
rect 11480 12384 11486 12436
rect 11790 12424 11796 12436
rect 11751 12396 11796 12424
rect 11790 12384 11796 12396
rect 11848 12384 11854 12436
rect 12250 12424 12256 12436
rect 12211 12396 12256 12424
rect 12250 12384 12256 12396
rect 12308 12384 12314 12436
rect 12710 12424 12716 12436
rect 12671 12396 12716 12424
rect 12710 12384 12716 12396
rect 12768 12424 12774 12436
rect 12986 12424 12992 12436
rect 12768 12396 12992 12424
rect 12768 12384 12774 12396
rect 12986 12384 12992 12396
rect 13044 12384 13050 12436
rect 13173 12427 13231 12433
rect 13173 12393 13185 12427
rect 13219 12424 13231 12427
rect 13262 12424 13268 12436
rect 13219 12396 13268 12424
rect 13219 12393 13231 12396
rect 13173 12387 13231 12393
rect 13262 12384 13268 12396
rect 13320 12384 13326 12436
rect 4930 12260 6132 12288
rect 6472 12328 9260 12356
rect 4930 12257 4942 12260
rect 4884 12251 4942 12257
rect 4522 12180 4528 12232
rect 4580 12220 4586 12232
rect 4617 12223 4675 12229
rect 4617 12220 4629 12223
rect 4580 12192 4629 12220
rect 4580 12180 4586 12192
rect 4617 12189 4629 12192
rect 4663 12189 4675 12223
rect 4617 12183 4675 12189
rect 5902 12180 5908 12232
rect 5960 12220 5966 12232
rect 6472 12220 6500 12328
rect 7190 12288 7196 12300
rect 7248 12297 7254 12300
rect 7160 12260 7196 12288
rect 7190 12248 7196 12260
rect 7248 12251 7260 12297
rect 7469 12291 7527 12297
rect 7469 12257 7481 12291
rect 7515 12288 7527 12291
rect 7650 12288 7656 12300
rect 7515 12260 7656 12288
rect 7515 12257 7527 12260
rect 7469 12251 7527 12257
rect 7248 12248 7254 12251
rect 7650 12248 7656 12260
rect 7708 12248 7714 12300
rect 8674 12291 8732 12297
rect 8674 12288 8686 12291
rect 7944 12260 8686 12288
rect 5960 12192 6500 12220
rect 5960 12180 5966 12192
rect 3200 12124 4476 12152
rect 3200 12112 3206 12124
rect 7944 12096 7972 12260
rect 8674 12257 8686 12260
rect 8720 12288 8732 12291
rect 8846 12288 8852 12300
rect 8720 12260 8852 12288
rect 8720 12257 8732 12260
rect 8674 12251 8732 12257
rect 8846 12248 8852 12260
rect 8904 12248 8910 12300
rect 9232 12288 9260 12328
rect 9306 12316 9312 12368
rect 9364 12365 9370 12368
rect 9364 12359 9428 12365
rect 9364 12325 9382 12359
rect 9416 12325 9428 12359
rect 12621 12359 12679 12365
rect 12621 12356 12633 12359
rect 9364 12319 9428 12325
rect 9646 12328 12633 12356
rect 9364 12316 9370 12319
rect 9646 12288 9674 12328
rect 12621 12325 12633 12328
rect 12667 12325 12679 12359
rect 12621 12319 12679 12325
rect 9232 12260 9674 12288
rect 9950 12248 9956 12300
rect 10008 12288 10014 12300
rect 10008 12260 10456 12288
rect 10008 12248 10014 12260
rect 8941 12223 8999 12229
rect 8941 12189 8953 12223
rect 8987 12220 8999 12223
rect 9125 12223 9183 12229
rect 9125 12220 9137 12223
rect 8987 12192 9137 12220
rect 8987 12189 8999 12192
rect 8941 12183 8999 12189
rect 9125 12189 9137 12192
rect 9171 12189 9183 12223
rect 9125 12183 9183 12189
rect 7926 12084 7932 12096
rect 3068 12056 7932 12084
rect 7926 12044 7932 12056
rect 7984 12044 7990 12096
rect 9140 12084 9168 12183
rect 10428 12152 10456 12260
rect 10962 12180 10968 12232
rect 11020 12220 11026 12232
rect 11149 12223 11207 12229
rect 11149 12220 11161 12223
rect 11020 12192 11161 12220
rect 11020 12180 11026 12192
rect 11149 12189 11161 12192
rect 11195 12189 11207 12223
rect 11149 12183 11207 12189
rect 11790 12180 11796 12232
rect 11848 12220 11854 12232
rect 11885 12223 11943 12229
rect 11885 12220 11897 12223
rect 11848 12192 11897 12220
rect 11848 12180 11854 12192
rect 11885 12189 11897 12192
rect 11931 12189 11943 12223
rect 11885 12183 11943 12189
rect 12069 12223 12127 12229
rect 12069 12189 12081 12223
rect 12115 12220 12127 12223
rect 12342 12220 12348 12232
rect 12115 12192 12348 12220
rect 12115 12189 12127 12192
rect 12069 12183 12127 12189
rect 12342 12180 12348 12192
rect 12400 12180 12406 12232
rect 12805 12223 12863 12229
rect 12805 12189 12817 12223
rect 12851 12189 12863 12223
rect 12805 12183 12863 12189
rect 10505 12155 10563 12161
rect 10505 12152 10517 12155
rect 10428 12124 10517 12152
rect 10505 12121 10517 12124
rect 10551 12152 10563 12155
rect 12820 12152 12848 12183
rect 10551 12124 12848 12152
rect 10551 12121 10563 12124
rect 10505 12115 10563 12121
rect 9306 12084 9312 12096
rect 9140 12056 9312 12084
rect 9306 12044 9312 12056
rect 9364 12044 9370 12096
rect 9490 12044 9496 12096
rect 9548 12084 9554 12096
rect 11238 12084 11244 12096
rect 9548 12056 11244 12084
rect 9548 12044 9554 12056
rect 11238 12044 11244 12056
rect 11296 12044 11302 12096
rect 11422 12084 11428 12096
rect 11383 12056 11428 12084
rect 11422 12044 11428 12056
rect 11480 12044 11486 12096
rect 11790 12044 11796 12096
rect 11848 12084 11854 12096
rect 12066 12084 12072 12096
rect 11848 12056 12072 12084
rect 11848 12044 11854 12056
rect 12066 12044 12072 12056
rect 12124 12084 12130 12096
rect 13354 12084 13360 12096
rect 12124 12056 13360 12084
rect 12124 12044 12130 12056
rect 13354 12044 13360 12056
rect 13412 12044 13418 12096
rect 13998 12044 14004 12096
rect 14056 12084 14062 12096
rect 14642 12084 14648 12096
rect 14056 12056 14648 12084
rect 14056 12044 14062 12056
rect 14642 12044 14648 12056
rect 14700 12044 14706 12096
rect 1104 11994 16008 12016
rect 1104 11942 3480 11994
rect 3532 11942 3544 11994
rect 3596 11942 3608 11994
rect 3660 11942 3672 11994
rect 3724 11942 8478 11994
rect 8530 11942 8542 11994
rect 8594 11942 8606 11994
rect 8658 11942 8670 11994
rect 8722 11942 13475 11994
rect 13527 11942 13539 11994
rect 13591 11942 13603 11994
rect 13655 11942 13667 11994
rect 13719 11942 16008 11994
rect 1104 11920 16008 11942
rect 2038 11840 2044 11892
rect 2096 11880 2102 11892
rect 2409 11883 2467 11889
rect 2409 11880 2421 11883
rect 2096 11852 2421 11880
rect 2096 11840 2102 11852
rect 2409 11849 2421 11852
rect 2455 11849 2467 11883
rect 3786 11880 3792 11892
rect 2409 11843 2467 11849
rect 2884 11852 3792 11880
rect 1765 11747 1823 11753
rect 1765 11713 1777 11747
rect 1811 11744 1823 11747
rect 2884 11744 2912 11852
rect 3786 11840 3792 11852
rect 3844 11840 3850 11892
rect 3970 11880 3976 11892
rect 3931 11852 3976 11880
rect 3970 11840 3976 11852
rect 4028 11840 4034 11892
rect 7926 11880 7932 11892
rect 7887 11852 7932 11880
rect 7926 11840 7932 11852
rect 7984 11840 7990 11892
rect 11241 11883 11299 11889
rect 11241 11849 11253 11883
rect 11287 11880 11299 11883
rect 11330 11880 11336 11892
rect 11287 11852 11336 11880
rect 11287 11849 11299 11852
rect 11241 11843 11299 11849
rect 11330 11840 11336 11852
rect 11388 11840 11394 11892
rect 11698 11880 11704 11892
rect 11659 11852 11704 11880
rect 11698 11840 11704 11852
rect 11756 11840 11762 11892
rect 12526 11880 12532 11892
rect 12487 11852 12532 11880
rect 12526 11840 12532 11852
rect 12584 11880 12590 11892
rect 12713 11883 12771 11889
rect 12713 11880 12725 11883
rect 12584 11852 12725 11880
rect 12584 11840 12590 11852
rect 12713 11849 12725 11852
rect 12759 11849 12771 11883
rect 13354 11880 13360 11892
rect 13315 11852 13360 11880
rect 12713 11843 12771 11849
rect 13354 11840 13360 11852
rect 13412 11840 13418 11892
rect 4798 11812 4804 11824
rect 4448 11784 4804 11812
rect 3050 11744 3056 11756
rect 1811 11716 2912 11744
rect 3011 11716 3056 11744
rect 1811 11713 1823 11716
rect 1765 11707 1823 11713
rect 3050 11704 3056 11716
rect 3108 11704 3114 11756
rect 3142 11704 3148 11756
rect 3200 11744 3206 11756
rect 3329 11747 3387 11753
rect 3329 11744 3341 11747
rect 3200 11716 3341 11744
rect 3200 11704 3206 11716
rect 3329 11713 3341 11716
rect 3375 11713 3387 11747
rect 3329 11707 3387 11713
rect 3513 11747 3571 11753
rect 3513 11713 3525 11747
rect 3559 11744 3571 11747
rect 4338 11744 4344 11756
rect 3559 11716 4344 11744
rect 3559 11713 3571 11716
rect 3513 11707 3571 11713
rect 4338 11704 4344 11716
rect 4396 11704 4402 11756
rect 2777 11679 2835 11685
rect 2777 11645 2789 11679
rect 2823 11676 2835 11679
rect 4448 11676 4476 11784
rect 4798 11772 4804 11784
rect 4856 11772 4862 11824
rect 10226 11812 10232 11824
rect 9784 11784 10232 11812
rect 4614 11744 4620 11756
rect 4575 11716 4620 11744
rect 4614 11704 4620 11716
rect 4672 11744 4678 11756
rect 6454 11744 6460 11756
rect 4672 11716 5028 11744
rect 6415 11716 6460 11744
rect 4672 11704 4678 11716
rect 2823 11648 4476 11676
rect 2823 11645 2835 11648
rect 2777 11639 2835 11645
rect 4522 11636 4528 11688
rect 4580 11676 4586 11688
rect 4890 11676 4896 11688
rect 4580 11648 4896 11676
rect 4580 11636 4586 11648
rect 4890 11636 4896 11648
rect 4948 11636 4954 11688
rect 5000 11676 5028 11716
rect 6454 11704 6460 11716
rect 6512 11704 6518 11756
rect 9306 11744 9312 11756
rect 9219 11716 9312 11744
rect 9306 11704 9312 11716
rect 9364 11744 9370 11756
rect 9674 11744 9680 11756
rect 9364 11716 9680 11744
rect 9364 11704 9370 11716
rect 9674 11704 9680 11716
rect 9732 11704 9738 11756
rect 5149 11679 5207 11685
rect 5149 11676 5161 11679
rect 5000 11648 5161 11676
rect 5149 11645 5161 11648
rect 5195 11645 5207 11679
rect 5149 11639 5207 11645
rect 5442 11636 5448 11688
rect 5500 11676 5506 11688
rect 8294 11676 8300 11688
rect 5500 11648 8300 11676
rect 5500 11636 5506 11648
rect 8294 11636 8300 11648
rect 8352 11636 8358 11688
rect 9030 11636 9036 11688
rect 9088 11685 9094 11688
rect 9784 11685 9812 11784
rect 10226 11772 10232 11784
rect 10284 11772 10290 11824
rect 11974 11812 11980 11824
rect 10612 11784 10824 11812
rect 10612 11756 10640 11784
rect 9953 11747 10011 11753
rect 9953 11713 9965 11747
rect 9999 11744 10011 11747
rect 10594 11744 10600 11756
rect 9999 11716 10600 11744
rect 9999 11713 10011 11716
rect 9953 11707 10011 11713
rect 9088 11676 9100 11685
rect 9769 11679 9827 11685
rect 9088 11648 9133 11676
rect 9088 11639 9100 11648
rect 9769 11645 9781 11679
rect 9815 11645 9827 11679
rect 9769 11639 9827 11645
rect 9088 11636 9094 11639
rect 1946 11608 1952 11620
rect 1907 11580 1952 11608
rect 1946 11568 1952 11580
rect 2004 11568 2010 11620
rect 2869 11611 2927 11617
rect 2332 11580 2774 11608
rect 1857 11543 1915 11549
rect 1857 11509 1869 11543
rect 1903 11540 1915 11543
rect 2222 11540 2228 11552
rect 1903 11512 2228 11540
rect 1903 11509 1915 11512
rect 1857 11503 1915 11509
rect 2222 11500 2228 11512
rect 2280 11500 2286 11552
rect 2332 11549 2360 11580
rect 2317 11543 2375 11549
rect 2317 11509 2329 11543
rect 2363 11509 2375 11543
rect 2746 11540 2774 11580
rect 2869 11577 2881 11611
rect 2915 11608 2927 11611
rect 3326 11608 3332 11620
rect 2915 11580 3332 11608
rect 2915 11577 2927 11580
rect 2869 11571 2927 11577
rect 3326 11568 3332 11580
rect 3384 11568 3390 11620
rect 4338 11608 4344 11620
rect 3436 11580 4344 11608
rect 3436 11540 3464 11580
rect 4338 11568 4344 11580
rect 4396 11568 4402 11620
rect 4433 11611 4491 11617
rect 4433 11577 4445 11611
rect 4479 11608 4491 11611
rect 5810 11608 5816 11620
rect 4479 11580 5816 11608
rect 4479 11577 4491 11580
rect 4433 11571 4491 11577
rect 5810 11568 5816 11580
rect 5868 11568 5874 11620
rect 6702 11611 6760 11617
rect 6702 11608 6714 11611
rect 6288 11580 6714 11608
rect 2746 11512 3464 11540
rect 2317 11503 2375 11509
rect 3602 11500 3608 11552
rect 3660 11540 3666 11552
rect 3660 11512 3705 11540
rect 3660 11500 3666 11512
rect 4062 11500 4068 11552
rect 4120 11540 4126 11552
rect 4120 11512 4165 11540
rect 4120 11500 4126 11512
rect 4522 11500 4528 11552
rect 4580 11540 4586 11552
rect 4580 11512 4625 11540
rect 4580 11500 4586 11512
rect 4798 11500 4804 11552
rect 4856 11540 4862 11552
rect 6288 11549 6316 11580
rect 6702 11577 6714 11580
rect 6748 11577 6760 11611
rect 9968 11608 9996 11707
rect 10594 11704 10600 11716
rect 10652 11704 10658 11756
rect 10796 11753 10824 11784
rect 10989 11784 11980 11812
rect 10781 11747 10839 11753
rect 10781 11713 10793 11747
rect 10827 11713 10839 11747
rect 10781 11707 10839 11713
rect 6702 11571 6760 11577
rect 7852 11580 9996 11608
rect 10597 11611 10655 11617
rect 7852 11552 7880 11580
rect 10597 11577 10609 11611
rect 10643 11608 10655 11611
rect 10989 11608 11017 11784
rect 11974 11772 11980 11784
rect 12032 11772 12038 11824
rect 12434 11772 12440 11824
rect 12492 11812 12498 11824
rect 12986 11812 12992 11824
rect 12492 11784 12992 11812
rect 12492 11772 12498 11784
rect 12986 11772 12992 11784
rect 13044 11812 13050 11824
rect 13081 11815 13139 11821
rect 13081 11812 13093 11815
rect 13044 11784 13093 11812
rect 13044 11772 13050 11784
rect 13081 11781 13093 11784
rect 13127 11781 13139 11815
rect 13081 11775 13139 11781
rect 11238 11704 11244 11756
rect 11296 11744 11302 11756
rect 11333 11747 11391 11753
rect 11333 11744 11345 11747
rect 11296 11716 11345 11744
rect 11296 11704 11302 11716
rect 11333 11713 11345 11716
rect 11379 11744 11391 11747
rect 11379 11716 11468 11744
rect 11379 11713 11391 11716
rect 11333 11707 11391 11713
rect 11440 11688 11468 11716
rect 11606 11704 11612 11756
rect 11664 11744 11670 11756
rect 12253 11747 12311 11753
rect 12253 11744 12265 11747
rect 11664 11716 12265 11744
rect 11664 11704 11670 11716
rect 12253 11713 12265 11716
rect 12299 11713 12311 11747
rect 12253 11707 12311 11713
rect 12710 11704 12716 11756
rect 12768 11744 12774 11756
rect 12897 11747 12955 11753
rect 12897 11744 12909 11747
rect 12768 11716 12909 11744
rect 12768 11704 12774 11716
rect 12897 11713 12909 11716
rect 12943 11744 12955 11747
rect 13998 11744 14004 11756
rect 12943 11716 14004 11744
rect 12943 11713 12955 11716
rect 12897 11707 12955 11713
rect 13998 11704 14004 11716
rect 14056 11704 14062 11756
rect 11054 11636 11060 11688
rect 11112 11676 11118 11688
rect 11112 11648 11157 11676
rect 11112 11636 11118 11648
rect 11422 11636 11428 11688
rect 11480 11636 11486 11688
rect 14734 11676 14740 11688
rect 11532 11648 14740 11676
rect 10643 11580 11017 11608
rect 10643 11577 10655 11580
rect 10597 11571 10655 11577
rect 6273 11543 6331 11549
rect 6273 11540 6285 11543
rect 4856 11512 6285 11540
rect 4856 11500 4862 11512
rect 6273 11509 6285 11512
rect 6319 11509 6331 11543
rect 7834 11540 7840 11552
rect 7795 11512 7840 11540
rect 6273 11503 6331 11509
rect 7834 11500 7840 11512
rect 7892 11500 7898 11552
rect 8386 11500 8392 11552
rect 8444 11540 8450 11552
rect 8846 11540 8852 11552
rect 8444 11512 8852 11540
rect 8444 11500 8450 11512
rect 8846 11500 8852 11512
rect 8904 11500 8910 11552
rect 9398 11540 9404 11552
rect 9359 11512 9404 11540
rect 9398 11500 9404 11512
rect 9456 11500 9462 11552
rect 9490 11500 9496 11552
rect 9548 11540 9554 11552
rect 9861 11543 9919 11549
rect 9861 11540 9873 11543
rect 9548 11512 9873 11540
rect 9548 11500 9554 11512
rect 9861 11509 9873 11512
rect 9907 11509 9919 11543
rect 10226 11540 10232 11552
rect 10187 11512 10232 11540
rect 9861 11503 9919 11509
rect 10226 11500 10232 11512
rect 10284 11500 10290 11552
rect 10686 11540 10692 11552
rect 10647 11512 10692 11540
rect 10686 11500 10692 11512
rect 10744 11500 10750 11552
rect 10870 11500 10876 11552
rect 10928 11540 10934 11552
rect 11532 11540 11560 11648
rect 14734 11636 14740 11648
rect 14792 11636 14798 11688
rect 12069 11611 12127 11617
rect 12069 11577 12081 11611
rect 12115 11608 12127 11611
rect 12618 11608 12624 11620
rect 12115 11580 12624 11608
rect 12115 11577 12127 11580
rect 12069 11571 12127 11577
rect 12618 11568 12624 11580
rect 12676 11568 12682 11620
rect 13170 11568 13176 11620
rect 13228 11608 13234 11620
rect 14642 11608 14648 11620
rect 13228 11580 14648 11608
rect 13228 11568 13234 11580
rect 14642 11568 14648 11580
rect 14700 11568 14706 11620
rect 10928 11512 11560 11540
rect 10928 11500 10934 11512
rect 11698 11500 11704 11552
rect 11756 11540 11762 11552
rect 12161 11543 12219 11549
rect 12161 11540 12173 11543
rect 11756 11512 12173 11540
rect 11756 11500 11762 11512
rect 12161 11509 12173 11512
rect 12207 11509 12219 11543
rect 12161 11503 12219 11509
rect 13078 11500 13084 11552
rect 13136 11540 13142 11552
rect 14458 11540 14464 11552
rect 13136 11512 14464 11540
rect 13136 11500 13142 11512
rect 14458 11500 14464 11512
rect 14516 11500 14522 11552
rect 1104 11450 16008 11472
rect 1104 11398 5979 11450
rect 6031 11398 6043 11450
rect 6095 11398 6107 11450
rect 6159 11398 6171 11450
rect 6223 11398 10976 11450
rect 11028 11398 11040 11450
rect 11092 11398 11104 11450
rect 11156 11398 11168 11450
rect 11220 11398 16008 11450
rect 1104 11376 16008 11398
rect 1486 11336 1492 11348
rect 1447 11308 1492 11336
rect 1486 11296 1492 11308
rect 1544 11296 1550 11348
rect 1857 11339 1915 11345
rect 1857 11305 1869 11339
rect 1903 11305 1915 11339
rect 1857 11299 1915 11305
rect 3421 11339 3479 11345
rect 3421 11305 3433 11339
rect 3467 11336 3479 11339
rect 4062 11336 4068 11348
rect 3467 11308 4068 11336
rect 3467 11305 3479 11308
rect 3421 11299 3479 11305
rect 1581 11271 1639 11277
rect 1581 11237 1593 11271
rect 1627 11268 1639 11271
rect 1872 11268 1900 11299
rect 4062 11296 4068 11308
rect 4120 11296 4126 11348
rect 4154 11296 4160 11348
rect 4212 11336 4218 11348
rect 9125 11339 9183 11345
rect 9125 11336 9137 11339
rect 4212 11308 9137 11336
rect 4212 11296 4218 11308
rect 9125 11305 9137 11308
rect 9171 11305 9183 11339
rect 9125 11299 9183 11305
rect 9490 11296 9496 11348
rect 9548 11336 9554 11348
rect 9585 11339 9643 11345
rect 9585 11336 9597 11339
rect 9548 11308 9597 11336
rect 9548 11296 9554 11308
rect 9585 11305 9597 11308
rect 9631 11305 9643 11339
rect 9585 11299 9643 11305
rect 10321 11339 10379 11345
rect 10321 11305 10333 11339
rect 10367 11336 10379 11339
rect 10778 11336 10784 11348
rect 10367 11308 10784 11336
rect 10367 11305 10379 11308
rect 10321 11299 10379 11305
rect 10778 11296 10784 11308
rect 10836 11336 10842 11348
rect 11149 11339 11207 11345
rect 10836 11308 11008 11336
rect 10836 11296 10842 11308
rect 10980 11280 11008 11308
rect 11149 11305 11161 11339
rect 11195 11336 11207 11339
rect 11514 11336 11520 11348
rect 11195 11308 11520 11336
rect 11195 11305 11207 11308
rect 11149 11299 11207 11305
rect 11514 11296 11520 11308
rect 11572 11296 11578 11348
rect 11974 11296 11980 11348
rect 12032 11336 12038 11348
rect 14185 11339 14243 11345
rect 14185 11336 14197 11339
rect 12032 11308 14197 11336
rect 12032 11296 12038 11308
rect 14185 11305 14197 11308
rect 14231 11305 14243 11339
rect 14366 11336 14372 11348
rect 14327 11308 14372 11336
rect 14185 11299 14243 11305
rect 14366 11296 14372 11308
rect 14424 11296 14430 11348
rect 14734 11336 14740 11348
rect 14695 11308 14740 11336
rect 14734 11296 14740 11308
rect 14792 11296 14798 11348
rect 14829 11339 14887 11345
rect 14829 11305 14841 11339
rect 14875 11336 14887 11339
rect 15286 11336 15292 11348
rect 14875 11308 15292 11336
rect 14875 11305 14887 11308
rect 14829 11299 14887 11305
rect 15286 11296 15292 11308
rect 15344 11296 15350 11348
rect 1627 11240 1900 11268
rect 1627 11237 1639 11240
rect 1581 11231 1639 11237
rect 3602 11228 3608 11280
rect 3660 11268 3666 11280
rect 3660 11240 5856 11268
rect 3660 11228 3666 11240
rect 2041 11203 2099 11209
rect 2041 11169 2053 11203
rect 2087 11169 2099 11203
rect 2498 11200 2504 11212
rect 2459 11172 2504 11200
rect 2041 11163 2099 11169
rect 2056 11064 2084 11163
rect 2498 11160 2504 11172
rect 2556 11160 2562 11212
rect 3326 11200 3332 11212
rect 3287 11172 3332 11200
rect 3326 11160 3332 11172
rect 3384 11160 3390 11212
rect 4798 11200 4804 11212
rect 3620 11172 4804 11200
rect 2590 11132 2596 11144
rect 2551 11104 2596 11132
rect 2590 11092 2596 11104
rect 2648 11092 2654 11144
rect 3620 11141 3648 11172
rect 4798 11160 4804 11172
rect 4856 11160 4862 11212
rect 5097 11203 5155 11209
rect 5097 11169 5109 11203
rect 5143 11200 5155 11203
rect 5258 11200 5264 11212
rect 5143 11172 5264 11200
rect 5143 11169 5155 11172
rect 5097 11163 5155 11169
rect 5258 11160 5264 11172
rect 5316 11160 5322 11212
rect 2777 11135 2835 11141
rect 2777 11101 2789 11135
rect 2823 11132 2835 11135
rect 3605 11135 3663 11141
rect 2823 11104 3556 11132
rect 2823 11101 2835 11104
rect 2777 11095 2835 11101
rect 2961 11067 3019 11073
rect 2961 11064 2973 11067
rect 2056 11036 2973 11064
rect 2961 11033 2973 11036
rect 3007 11033 3019 11067
rect 2961 11027 3019 11033
rect 2130 10996 2136 11008
rect 2091 10968 2136 10996
rect 2130 10956 2136 10968
rect 2188 10956 2194 11008
rect 3528 10996 3556 11104
rect 3605 11101 3617 11135
rect 3651 11101 3663 11135
rect 3605 11095 3663 11101
rect 5353 11135 5411 11141
rect 5353 11101 5365 11135
rect 5399 11132 5411 11135
rect 5534 11132 5540 11144
rect 5399 11104 5540 11132
rect 5399 11101 5411 11104
rect 5353 11095 5411 11101
rect 5534 11092 5540 11104
rect 5592 11092 5598 11144
rect 3786 11024 3792 11076
rect 3844 11064 3850 11076
rect 3973 11067 4031 11073
rect 3973 11064 3985 11067
rect 3844 11036 3985 11064
rect 3844 11024 3850 11036
rect 3973 11033 3985 11036
rect 4019 11033 4031 11067
rect 3973 11027 4031 11033
rect 5445 11067 5503 11073
rect 5445 11033 5457 11067
rect 5491 11033 5503 11067
rect 5828 11064 5856 11240
rect 6454 11228 6460 11280
rect 6512 11268 6518 11280
rect 6512 11240 6868 11268
rect 6512 11228 6518 11240
rect 6270 11160 6276 11212
rect 6328 11200 6334 11212
rect 6840 11209 6868 11240
rect 7834 11228 7840 11280
rect 7892 11268 7898 11280
rect 8030 11271 8088 11277
rect 8030 11268 8042 11271
rect 7892 11240 8042 11268
rect 7892 11228 7898 11240
rect 8030 11237 8042 11240
rect 8076 11237 8088 11271
rect 8030 11231 8088 11237
rect 8202 11228 8208 11280
rect 8260 11268 8266 11280
rect 9950 11268 9956 11280
rect 8260 11240 9956 11268
rect 8260 11228 8266 11240
rect 9950 11228 9956 11240
rect 10008 11228 10014 11280
rect 10686 11228 10692 11280
rect 10744 11268 10750 11280
rect 10870 11268 10876 11280
rect 10744 11240 10876 11268
rect 10744 11228 10750 11240
rect 10870 11228 10876 11240
rect 10928 11228 10934 11280
rect 10962 11228 10968 11280
rect 11020 11228 11026 11280
rect 11241 11271 11299 11277
rect 11241 11237 11253 11271
rect 11287 11268 11299 11271
rect 11287 11240 12112 11268
rect 11287 11237 11299 11240
rect 11241 11231 11299 11237
rect 6558 11203 6616 11209
rect 6558 11200 6570 11203
rect 6328 11172 6570 11200
rect 6328 11160 6334 11172
rect 6558 11169 6570 11172
rect 6604 11169 6616 11203
rect 6558 11163 6616 11169
rect 6825 11203 6883 11209
rect 6825 11169 6837 11203
rect 6871 11169 6883 11203
rect 8573 11203 8631 11209
rect 6825 11163 6883 11169
rect 7300 11172 8524 11200
rect 7300 11132 7328 11172
rect 6840 11104 7328 11132
rect 8297 11135 8355 11141
rect 5828 11036 5948 11064
rect 5445 11027 5503 11033
rect 4430 10996 4436 11008
rect 3528 10968 4436 10996
rect 4430 10956 4436 10968
rect 4488 10956 4494 11008
rect 4614 10956 4620 11008
rect 4672 10996 4678 11008
rect 5460 10996 5488 11027
rect 4672 10968 5488 10996
rect 5920 10996 5948 11036
rect 6840 10996 6868 11104
rect 8297 11101 8309 11135
rect 8343 11101 8355 11135
rect 8297 11095 8355 11101
rect 6917 11067 6975 11073
rect 6917 11033 6929 11067
rect 6963 11064 6975 11067
rect 7190 11064 7196 11076
rect 6963 11036 7196 11064
rect 6963 11033 6975 11036
rect 6917 11027 6975 11033
rect 7190 11024 7196 11036
rect 7248 11024 7254 11076
rect 5920 10968 6868 10996
rect 4672 10956 4678 10968
rect 7926 10956 7932 11008
rect 7984 10996 7990 11008
rect 8312 10996 8340 11095
rect 7984 10968 8340 10996
rect 8496 10996 8524 11172
rect 8573 11169 8585 11203
rect 8619 11200 8631 11203
rect 9493 11203 9551 11209
rect 9493 11200 9505 11203
rect 8619 11172 9505 11200
rect 8619 11169 8631 11172
rect 8573 11163 8631 11169
rect 9493 11169 9505 11172
rect 9539 11169 9551 11203
rect 9493 11163 9551 11169
rect 9582 11160 9588 11212
rect 9640 11200 9646 11212
rect 10413 11203 10471 11209
rect 10413 11200 10425 11203
rect 9640 11172 10425 11200
rect 9640 11160 9646 11172
rect 10413 11169 10425 11172
rect 10459 11200 10471 11203
rect 11054 11200 11060 11212
rect 10459 11172 11060 11200
rect 10459 11169 10471 11172
rect 10413 11163 10471 11169
rect 11054 11160 11060 11172
rect 11112 11160 11118 11212
rect 11974 11200 11980 11212
rect 11935 11172 11980 11200
rect 11974 11160 11980 11172
rect 12032 11160 12038 11212
rect 8849 11135 8907 11141
rect 8849 11101 8861 11135
rect 8895 11132 8907 11135
rect 9766 11132 9772 11144
rect 8895 11104 9674 11132
rect 9727 11104 9772 11132
rect 8895 11101 8907 11104
rect 8849 11095 8907 11101
rect 9646 11064 9674 11104
rect 9766 11092 9772 11104
rect 9824 11092 9830 11144
rect 10594 11132 10600 11144
rect 10555 11104 10600 11132
rect 10594 11092 10600 11104
rect 10652 11092 10658 11144
rect 10870 11092 10876 11144
rect 10928 11132 10934 11144
rect 11333 11135 11391 11141
rect 11333 11132 11345 11135
rect 10928 11104 11345 11132
rect 10928 11092 10934 11104
rect 11333 11101 11345 11104
rect 11379 11101 11391 11135
rect 11333 11095 11391 11101
rect 11514 11092 11520 11144
rect 11572 11132 11578 11144
rect 11701 11135 11759 11141
rect 11701 11132 11713 11135
rect 11572 11104 11713 11132
rect 11572 11092 11578 11104
rect 11701 11101 11713 11104
rect 11747 11101 11759 11135
rect 11882 11132 11888 11144
rect 11843 11104 11888 11132
rect 11701 11095 11759 11101
rect 11882 11092 11888 11104
rect 11940 11092 11946 11144
rect 12084 11132 12112 11240
rect 12250 11228 12256 11280
rect 12308 11268 12314 11280
rect 12308 11240 12480 11268
rect 12308 11228 12314 11240
rect 12452 11200 12480 11240
rect 12526 11228 12532 11280
rect 12584 11268 12590 11280
rect 12805 11271 12863 11277
rect 12805 11268 12817 11271
rect 12584 11240 12817 11268
rect 12584 11228 12590 11240
rect 12805 11237 12817 11240
rect 12851 11237 12863 11271
rect 12805 11231 12863 11237
rect 12897 11271 12955 11277
rect 12897 11237 12909 11271
rect 12943 11268 12955 11271
rect 12986 11268 12992 11280
rect 12943 11240 12992 11268
rect 12943 11237 12955 11240
rect 12897 11231 12955 11237
rect 12986 11228 12992 11240
rect 13044 11268 13050 11280
rect 13170 11268 13176 11280
rect 13044 11240 13176 11268
rect 13044 11228 13050 11240
rect 13170 11228 13176 11240
rect 13228 11268 13234 11280
rect 13817 11271 13875 11277
rect 13817 11268 13829 11271
rect 13228 11240 13829 11268
rect 13228 11228 13234 11240
rect 13817 11237 13829 11240
rect 13863 11237 13875 11271
rect 13817 11231 13875 11237
rect 14734 11200 14740 11212
rect 12452 11172 14740 11200
rect 12710 11132 12716 11144
rect 12084 11104 12716 11132
rect 12710 11092 12716 11104
rect 12768 11092 12774 11144
rect 13004 11141 13032 11172
rect 14734 11160 14740 11172
rect 14792 11200 14798 11212
rect 14792 11172 14964 11200
rect 14792 11160 14798 11172
rect 12989 11135 13047 11141
rect 12989 11101 13001 11135
rect 13035 11101 13047 11135
rect 12989 11095 13047 11101
rect 13262 11092 13268 11144
rect 13320 11132 13326 11144
rect 14936 11141 14964 11172
rect 13449 11135 13507 11141
rect 13449 11132 13461 11135
rect 13320 11104 13461 11132
rect 13320 11092 13326 11104
rect 13449 11101 13461 11104
rect 13495 11101 13507 11135
rect 13449 11095 13507 11101
rect 14921 11135 14979 11141
rect 14921 11101 14933 11135
rect 14967 11101 14979 11135
rect 14921 11095 14979 11101
rect 10318 11064 10324 11076
rect 9646 11036 10324 11064
rect 10318 11024 10324 11036
rect 10376 11024 10382 11076
rect 12158 11024 12164 11076
rect 12216 11064 12222 11076
rect 12345 11067 12403 11073
rect 12345 11064 12357 11067
rect 12216 11036 12357 11064
rect 12216 11024 12222 11036
rect 12345 11033 12357 11036
rect 12391 11033 12403 11067
rect 12345 11027 12403 11033
rect 12434 11024 12440 11076
rect 12492 11064 12498 11076
rect 12492 11036 12537 11064
rect 12492 11024 12498 11036
rect 9490 10996 9496 11008
rect 8496 10968 9496 10996
rect 7984 10956 7990 10968
rect 9490 10956 9496 10968
rect 9548 10956 9554 11008
rect 9582 10956 9588 11008
rect 9640 10996 9646 11008
rect 9766 10996 9772 11008
rect 9640 10968 9772 10996
rect 9640 10956 9646 10968
rect 9766 10956 9772 10968
rect 9824 10956 9830 11008
rect 9950 10996 9956 11008
rect 9911 10968 9956 10996
rect 9950 10956 9956 10968
rect 10008 10956 10014 11008
rect 10778 10996 10784 11008
rect 10739 10968 10784 10996
rect 10778 10956 10784 10968
rect 10836 10956 10842 11008
rect 11606 10956 11612 11008
rect 11664 10996 11670 11008
rect 13265 10999 13323 11005
rect 13265 10996 13277 10999
rect 11664 10968 13277 10996
rect 11664 10956 11670 10968
rect 13265 10965 13277 10968
rect 13311 10996 13323 10999
rect 13354 10996 13360 11008
rect 13311 10968 13360 10996
rect 13311 10965 13323 10968
rect 13265 10959 13323 10965
rect 13354 10956 13360 10968
rect 13412 10956 13418 11008
rect 13464 10996 13492 11095
rect 13725 11067 13783 11073
rect 13725 11033 13737 11067
rect 13771 11064 13783 11067
rect 13998 11064 14004 11076
rect 13771 11036 14004 11064
rect 13771 11033 13783 11036
rect 13725 11027 13783 11033
rect 13998 11024 14004 11036
rect 14056 11024 14062 11076
rect 14093 11067 14151 11073
rect 14093 11033 14105 11067
rect 14139 11064 14151 11067
rect 14185 11067 14243 11073
rect 14185 11064 14197 11067
rect 14139 11036 14197 11064
rect 14139 11033 14151 11036
rect 14093 11027 14151 11033
rect 14185 11033 14197 11036
rect 14231 11064 14243 11067
rect 14550 11064 14556 11076
rect 14231 11036 14556 11064
rect 14231 11033 14243 11036
rect 14185 11027 14243 11033
rect 14550 11024 14556 11036
rect 14608 11024 14614 11076
rect 15102 10996 15108 11008
rect 13464 10968 15108 10996
rect 15102 10956 15108 10968
rect 15160 10956 15166 11008
rect 1104 10906 16008 10928
rect 1104 10854 3480 10906
rect 3532 10854 3544 10906
rect 3596 10854 3608 10906
rect 3660 10854 3672 10906
rect 3724 10854 8478 10906
rect 8530 10854 8542 10906
rect 8594 10854 8606 10906
rect 8658 10854 8670 10906
rect 8722 10854 13475 10906
rect 13527 10854 13539 10906
rect 13591 10854 13603 10906
rect 13655 10854 13667 10906
rect 13719 10854 16008 10906
rect 1104 10832 16008 10854
rect 2501 10795 2559 10801
rect 2501 10761 2513 10795
rect 2547 10792 2559 10795
rect 2590 10792 2596 10804
rect 2547 10764 2596 10792
rect 2547 10761 2559 10764
rect 2501 10755 2559 10761
rect 2590 10752 2596 10764
rect 2648 10752 2654 10804
rect 3326 10792 3332 10804
rect 3287 10764 3332 10792
rect 3326 10752 3332 10764
rect 3384 10752 3390 10804
rect 9401 10795 9459 10801
rect 9401 10792 9413 10795
rect 3436 10764 9413 10792
rect 1949 10659 2007 10665
rect 1949 10625 1961 10659
rect 1995 10656 2007 10659
rect 2682 10656 2688 10668
rect 1995 10628 2688 10656
rect 1995 10625 2007 10628
rect 1949 10619 2007 10625
rect 2682 10616 2688 10628
rect 2740 10616 2746 10668
rect 2777 10659 2835 10665
rect 2777 10625 2789 10659
rect 2823 10625 2835 10659
rect 2777 10619 2835 10625
rect 2869 10659 2927 10665
rect 2869 10625 2881 10659
rect 2915 10656 2927 10659
rect 3436 10656 3464 10764
rect 9401 10761 9413 10764
rect 9447 10761 9459 10795
rect 9401 10755 9459 10761
rect 9490 10752 9496 10804
rect 9548 10792 9554 10804
rect 10229 10795 10287 10801
rect 10229 10792 10241 10795
rect 9548 10764 10241 10792
rect 9548 10752 9554 10764
rect 10229 10761 10241 10764
rect 10275 10761 10287 10795
rect 10229 10755 10287 10761
rect 10686 10752 10692 10804
rect 10744 10792 10750 10804
rect 11054 10792 11060 10804
rect 10744 10764 11060 10792
rect 10744 10752 10750 10764
rect 11054 10752 11060 10764
rect 11112 10752 11118 10804
rect 11422 10792 11428 10804
rect 11383 10764 11428 10792
rect 11422 10752 11428 10764
rect 11480 10792 11486 10804
rect 12066 10792 12072 10804
rect 11480 10764 12072 10792
rect 11480 10752 11486 10764
rect 12066 10752 12072 10764
rect 12124 10752 12130 10804
rect 12529 10795 12587 10801
rect 12529 10761 12541 10795
rect 12575 10792 12587 10795
rect 12618 10792 12624 10804
rect 12575 10764 12624 10792
rect 12575 10761 12587 10764
rect 12529 10755 12587 10761
rect 12618 10752 12624 10764
rect 12676 10752 12682 10804
rect 12802 10752 12808 10804
rect 12860 10792 12866 10804
rect 13078 10792 13084 10804
rect 12860 10764 13084 10792
rect 12860 10752 12866 10764
rect 13078 10752 13084 10764
rect 13136 10752 13142 10804
rect 14182 10792 14188 10804
rect 14143 10764 14188 10792
rect 14182 10752 14188 10764
rect 14240 10752 14246 10804
rect 6273 10727 6331 10733
rect 6273 10693 6285 10727
rect 6319 10693 6331 10727
rect 9306 10724 9312 10736
rect 9267 10696 9312 10724
rect 6273 10687 6331 10693
rect 4890 10656 4896 10668
rect 2915 10628 3464 10656
rect 4851 10628 4896 10656
rect 2915 10625 2927 10628
rect 2869 10619 2927 10625
rect 2792 10588 2820 10619
rect 4890 10616 4896 10628
rect 4948 10616 4954 10668
rect 5902 10616 5908 10668
rect 5960 10656 5966 10668
rect 6288 10656 6316 10687
rect 9306 10684 9312 10696
rect 9364 10684 9370 10736
rect 9766 10724 9772 10736
rect 9416 10696 9772 10724
rect 5960 10628 6601 10656
rect 5960 10616 5966 10628
rect 2792 10560 3372 10588
rect 1581 10523 1639 10529
rect 1581 10489 1593 10523
rect 1627 10520 1639 10523
rect 1854 10520 1860 10532
rect 1627 10492 1860 10520
rect 1627 10489 1639 10492
rect 1581 10483 1639 10489
rect 1854 10480 1860 10492
rect 1912 10480 1918 10532
rect 2133 10523 2191 10529
rect 2133 10489 2145 10523
rect 2179 10520 2191 10523
rect 3234 10520 3240 10532
rect 2179 10492 3240 10520
rect 2179 10489 2191 10492
rect 2133 10483 2191 10489
rect 3234 10480 3240 10492
rect 3292 10480 3298 10532
rect 3344 10520 3372 10560
rect 3418 10548 3424 10600
rect 3476 10588 3482 10600
rect 4614 10588 4620 10600
rect 3476 10560 3521 10588
rect 3620 10560 4620 10588
rect 3476 10548 3482 10560
rect 3620 10520 3648 10560
rect 4614 10548 4620 10560
rect 4672 10548 4678 10600
rect 4798 10548 4804 10600
rect 4856 10588 4862 10600
rect 4856 10560 5304 10588
rect 4856 10548 4862 10560
rect 3344 10492 3648 10520
rect 3688 10523 3746 10529
rect 3688 10489 3700 10523
rect 3734 10520 3746 10523
rect 3786 10520 3792 10532
rect 3734 10492 3792 10520
rect 3734 10489 3746 10492
rect 3688 10483 3746 10489
rect 3786 10480 3792 10492
rect 3844 10480 3850 10532
rect 3970 10480 3976 10532
rect 4028 10520 4034 10532
rect 4430 10520 4436 10532
rect 4028 10492 4436 10520
rect 4028 10480 4034 10492
rect 4430 10480 4436 10492
rect 4488 10520 4494 10532
rect 5138 10523 5196 10529
rect 5138 10520 5150 10523
rect 4488 10492 5150 10520
rect 4488 10480 4494 10492
rect 5138 10489 5150 10492
rect 5184 10489 5196 10523
rect 5276 10520 5304 10560
rect 5534 10548 5540 10600
rect 5592 10588 5598 10600
rect 6457 10591 6515 10597
rect 6457 10588 6469 10591
rect 5592 10560 6469 10588
rect 5592 10548 5598 10560
rect 6457 10557 6469 10560
rect 6503 10557 6515 10591
rect 6573 10588 6601 10628
rect 7484 10628 8055 10656
rect 7484 10588 7512 10628
rect 7926 10588 7932 10600
rect 6573 10560 7512 10588
rect 7887 10560 7932 10588
rect 6457 10551 6515 10557
rect 7926 10548 7932 10560
rect 7984 10548 7990 10600
rect 8027 10588 8055 10628
rect 9122 10616 9128 10668
rect 9180 10656 9186 10668
rect 9416 10656 9444 10696
rect 9766 10684 9772 10696
rect 9824 10684 9830 10736
rect 10594 10684 10600 10736
rect 10652 10724 10658 10736
rect 10652 10696 11017 10724
rect 10652 10684 10658 10696
rect 9180 10628 9444 10656
rect 9180 10616 9186 10628
rect 9674 10616 9680 10668
rect 9732 10656 9738 10668
rect 9861 10659 9919 10665
rect 9861 10656 9873 10659
rect 9732 10628 9873 10656
rect 9732 10616 9738 10628
rect 9861 10625 9873 10628
rect 9907 10625 9919 10659
rect 9861 10619 9919 10625
rect 9953 10659 10011 10665
rect 9953 10625 9965 10659
rect 9999 10625 10011 10659
rect 9953 10619 10011 10625
rect 8027 10560 8340 10588
rect 5902 10520 5908 10532
rect 5276 10492 5908 10520
rect 5138 10483 5196 10489
rect 5902 10480 5908 10492
rect 5960 10480 5966 10532
rect 6546 10480 6552 10532
rect 6604 10520 6610 10532
rect 6702 10523 6760 10529
rect 6702 10520 6714 10523
rect 6604 10492 6714 10520
rect 6604 10480 6610 10492
rect 6702 10489 6714 10492
rect 6748 10489 6760 10523
rect 6702 10483 6760 10489
rect 8018 10480 8024 10532
rect 8076 10520 8082 10532
rect 8174 10523 8232 10529
rect 8174 10520 8186 10523
rect 8076 10492 8186 10520
rect 8076 10480 8082 10492
rect 8174 10489 8186 10492
rect 8220 10489 8232 10523
rect 8312 10520 8340 10560
rect 8662 10548 8668 10600
rect 8720 10588 8726 10600
rect 9582 10588 9588 10600
rect 8720 10560 9588 10588
rect 8720 10548 8726 10560
rect 9582 10548 9588 10560
rect 9640 10588 9646 10600
rect 9968 10588 9996 10619
rect 10226 10616 10232 10668
rect 10284 10656 10290 10668
rect 10689 10659 10747 10665
rect 10689 10656 10701 10659
rect 10284 10628 10701 10656
rect 10284 10616 10290 10628
rect 10689 10625 10701 10628
rect 10735 10625 10747 10659
rect 10870 10656 10876 10668
rect 10831 10628 10876 10656
rect 10689 10619 10747 10625
rect 10870 10616 10876 10628
rect 10928 10616 10934 10668
rect 9640 10560 9996 10588
rect 9640 10548 9646 10560
rect 10410 10548 10416 10600
rect 10468 10588 10474 10600
rect 10597 10591 10655 10597
rect 10597 10588 10609 10591
rect 10468 10560 10609 10588
rect 10468 10548 10474 10560
rect 10597 10557 10609 10560
rect 10643 10557 10655 10591
rect 10989 10588 11017 10696
rect 11072 10656 11100 10752
rect 11238 10724 11244 10736
rect 11199 10696 11244 10724
rect 11238 10684 11244 10696
rect 11296 10724 11302 10736
rect 11296 10696 12020 10724
rect 11296 10684 11302 10696
rect 11606 10656 11612 10668
rect 11072 10628 11612 10656
rect 11606 10616 11612 10628
rect 11664 10616 11670 10668
rect 11992 10665 12020 10696
rect 12894 10684 12900 10736
rect 12952 10724 12958 10736
rect 13906 10724 13912 10736
rect 12952 10696 13912 10724
rect 12952 10684 12958 10696
rect 13906 10684 13912 10696
rect 13964 10684 13970 10736
rect 11793 10659 11851 10665
rect 11793 10625 11805 10659
rect 11839 10625 11851 10659
rect 11793 10619 11851 10625
rect 11977 10659 12035 10665
rect 11977 10625 11989 10659
rect 12023 10625 12035 10659
rect 11977 10619 12035 10625
rect 11808 10588 11836 10619
rect 12618 10616 12624 10668
rect 12676 10656 12682 10668
rect 13081 10659 13139 10665
rect 13081 10656 13093 10659
rect 12676 10628 13093 10656
rect 12676 10616 12682 10628
rect 13081 10625 13093 10628
rect 13127 10625 13139 10659
rect 13081 10619 13139 10625
rect 13449 10659 13507 10665
rect 13449 10625 13461 10659
rect 13495 10625 13507 10659
rect 14734 10656 14740 10668
rect 14695 10628 14740 10656
rect 13449 10619 13507 10625
rect 13464 10588 13492 10619
rect 14734 10616 14740 10628
rect 14792 10616 14798 10668
rect 10989 10560 11836 10588
rect 11900 10560 13492 10588
rect 13725 10591 13783 10597
rect 10597 10551 10655 10557
rect 11900 10520 11928 10560
rect 13725 10557 13737 10591
rect 13771 10588 13783 10591
rect 13998 10588 14004 10600
rect 13771 10560 14004 10588
rect 13771 10557 13783 10560
rect 13725 10551 13783 10557
rect 13998 10548 14004 10560
rect 14056 10548 14062 10600
rect 14090 10548 14096 10600
rect 14148 10588 14154 10600
rect 14553 10591 14611 10597
rect 14553 10588 14565 10591
rect 14148 10560 14565 10588
rect 14148 10548 14154 10560
rect 14553 10557 14565 10560
rect 14599 10557 14611 10591
rect 14553 10551 14611 10557
rect 8312 10492 11928 10520
rect 12069 10523 12127 10529
rect 8174 10483 8232 10489
rect 12069 10489 12081 10523
rect 12115 10520 12127 10523
rect 12250 10520 12256 10532
rect 12115 10492 12256 10520
rect 12115 10489 12127 10492
rect 12069 10483 12127 10489
rect 1486 10452 1492 10464
rect 1447 10424 1492 10452
rect 1486 10412 1492 10424
rect 1544 10412 1550 10464
rect 2038 10452 2044 10464
rect 1999 10424 2044 10452
rect 2038 10412 2044 10424
rect 2096 10412 2102 10464
rect 2961 10455 3019 10461
rect 2961 10421 2973 10455
rect 3007 10452 3019 10455
rect 4154 10452 4160 10464
rect 3007 10424 4160 10452
rect 3007 10421 3019 10424
rect 2961 10415 3019 10421
rect 4154 10412 4160 10424
rect 4212 10412 4218 10464
rect 4801 10455 4859 10461
rect 4801 10421 4813 10455
rect 4847 10452 4859 10455
rect 4982 10452 4988 10464
rect 4847 10424 4988 10452
rect 4847 10421 4859 10424
rect 4801 10415 4859 10421
rect 4982 10412 4988 10424
rect 5040 10412 5046 10464
rect 6270 10412 6276 10464
rect 6328 10452 6334 10464
rect 7837 10455 7895 10461
rect 7837 10452 7849 10455
rect 6328 10424 7849 10452
rect 6328 10412 6334 10424
rect 7837 10421 7849 10424
rect 7883 10452 7895 10455
rect 8662 10452 8668 10464
rect 7883 10424 8668 10452
rect 7883 10421 7895 10424
rect 7837 10415 7895 10421
rect 8662 10412 8668 10424
rect 8720 10412 8726 10464
rect 8846 10412 8852 10464
rect 8904 10452 8910 10464
rect 9769 10455 9827 10461
rect 9769 10452 9781 10455
rect 8904 10424 9781 10452
rect 8904 10412 8910 10424
rect 9769 10421 9781 10424
rect 9815 10421 9827 10455
rect 9769 10415 9827 10421
rect 10318 10412 10324 10464
rect 10376 10452 10382 10464
rect 12084 10452 12112 10483
rect 12250 10480 12256 10492
rect 12308 10480 12314 10532
rect 12897 10523 12955 10529
rect 12897 10489 12909 10523
rect 12943 10520 12955 10523
rect 13262 10520 13268 10532
rect 12943 10492 13268 10520
rect 12943 10489 12955 10492
rect 12897 10483 12955 10489
rect 13262 10480 13268 10492
rect 13320 10480 13326 10532
rect 13354 10480 13360 10532
rect 13412 10520 13418 10532
rect 13633 10523 13691 10529
rect 13633 10520 13645 10523
rect 13412 10492 13645 10520
rect 13412 10480 13418 10492
rect 13633 10489 13645 10492
rect 13679 10489 13691 10523
rect 15013 10523 15071 10529
rect 15013 10520 15025 10523
rect 13633 10483 13691 10489
rect 13740 10492 15025 10520
rect 13740 10464 13768 10492
rect 15013 10489 15025 10492
rect 15059 10489 15071 10523
rect 15013 10483 15071 10489
rect 10376 10424 12112 10452
rect 10376 10412 10382 10424
rect 12434 10412 12440 10464
rect 12492 10452 12498 10464
rect 12492 10424 12537 10452
rect 12492 10412 12498 10424
rect 12802 10412 12808 10464
rect 12860 10452 12866 10464
rect 12989 10455 13047 10461
rect 12989 10452 13001 10455
rect 12860 10424 13001 10452
rect 12860 10412 12866 10424
rect 12989 10421 13001 10424
rect 13035 10421 13047 10455
rect 12989 10415 13047 10421
rect 13722 10412 13728 10464
rect 13780 10412 13786 10464
rect 14090 10452 14096 10464
rect 14051 10424 14096 10452
rect 14090 10412 14096 10424
rect 14148 10412 14154 10464
rect 14550 10412 14556 10464
rect 14608 10452 14614 10464
rect 14645 10455 14703 10461
rect 14645 10452 14657 10455
rect 14608 10424 14657 10452
rect 14608 10412 14614 10424
rect 14645 10421 14657 10424
rect 14691 10421 14703 10455
rect 14645 10415 14703 10421
rect 1104 10362 16008 10384
rect 1104 10310 5979 10362
rect 6031 10310 6043 10362
rect 6095 10310 6107 10362
rect 6159 10310 6171 10362
rect 6223 10310 10976 10362
rect 11028 10310 11040 10362
rect 11092 10310 11104 10362
rect 11156 10310 11168 10362
rect 11220 10310 16008 10362
rect 1104 10288 16008 10310
rect 1854 10248 1860 10260
rect 1815 10220 1860 10248
rect 1854 10208 1860 10220
rect 1912 10208 1918 10260
rect 2038 10208 2044 10260
rect 2096 10248 2102 10260
rect 2133 10251 2191 10257
rect 2133 10248 2145 10251
rect 2096 10220 2145 10248
rect 2096 10208 2102 10220
rect 2133 10217 2145 10220
rect 2179 10217 2191 10251
rect 4341 10251 4399 10257
rect 2133 10211 2191 10217
rect 2792 10220 4292 10248
rect 2041 10115 2099 10121
rect 2041 10081 2053 10115
rect 2087 10112 2099 10115
rect 2406 10112 2412 10124
rect 2087 10084 2412 10112
rect 2087 10081 2099 10084
rect 2041 10075 2099 10081
rect 2406 10072 2412 10084
rect 2464 10072 2470 10124
rect 2501 10115 2559 10121
rect 2501 10081 2513 10115
rect 2547 10112 2559 10115
rect 2682 10112 2688 10124
rect 2547 10084 2688 10112
rect 2547 10081 2559 10084
rect 2501 10075 2559 10081
rect 2682 10072 2688 10084
rect 2740 10072 2746 10124
rect 2590 10044 2596 10056
rect 2551 10016 2596 10044
rect 2590 10004 2596 10016
rect 2648 10004 2654 10056
rect 2792 10053 2820 10220
rect 4264 10180 4292 10220
rect 4341 10217 4353 10251
rect 4387 10248 4399 10251
rect 4522 10248 4528 10260
rect 4387 10220 4528 10248
rect 4387 10217 4399 10220
rect 4341 10211 4399 10217
rect 4522 10208 4528 10220
rect 4580 10208 4586 10260
rect 4614 10208 4620 10260
rect 4672 10248 4678 10260
rect 5258 10248 5264 10260
rect 4672 10220 5264 10248
rect 4672 10208 4678 10220
rect 5258 10208 5264 10220
rect 5316 10208 5322 10260
rect 5626 10208 5632 10260
rect 5684 10248 5690 10260
rect 8113 10251 8171 10257
rect 8113 10248 8125 10251
rect 5684 10220 6592 10248
rect 5684 10208 5690 10220
rect 4430 10180 4436 10192
rect 4264 10152 4436 10180
rect 4430 10140 4436 10152
rect 4488 10140 4494 10192
rect 4801 10183 4859 10189
rect 4801 10149 4813 10183
rect 4847 10180 4859 10183
rect 6454 10180 6460 10192
rect 4847 10152 6460 10180
rect 4847 10149 4859 10152
rect 4801 10143 4859 10149
rect 6454 10140 6460 10152
rect 6512 10140 6518 10192
rect 6564 10180 6592 10220
rect 7024 10220 8125 10248
rect 6886 10183 6944 10189
rect 6886 10180 6898 10183
rect 6564 10152 6898 10180
rect 6886 10149 6898 10152
rect 6932 10149 6944 10183
rect 6886 10143 6944 10149
rect 3142 10072 3148 10124
rect 3200 10112 3206 10124
rect 3329 10115 3387 10121
rect 3329 10112 3341 10115
rect 3200 10084 3341 10112
rect 3200 10072 3206 10084
rect 3329 10081 3341 10084
rect 3375 10081 3387 10115
rect 3329 10075 3387 10081
rect 3421 10115 3479 10121
rect 3421 10081 3433 10115
rect 3467 10112 3479 10115
rect 3694 10112 3700 10124
rect 3467 10084 3700 10112
rect 3467 10081 3479 10084
rect 3421 10075 3479 10081
rect 3694 10072 3700 10084
rect 3752 10072 3758 10124
rect 3878 10072 3884 10124
rect 3936 10112 3942 10124
rect 4065 10115 4123 10121
rect 4065 10112 4077 10115
rect 3936 10084 4077 10112
rect 3936 10072 3942 10084
rect 4065 10081 4077 10084
rect 4111 10081 4123 10115
rect 4065 10075 4123 10081
rect 4522 10072 4528 10124
rect 4580 10112 4586 10124
rect 4709 10115 4767 10121
rect 4709 10112 4721 10115
rect 4580 10084 4721 10112
rect 4580 10072 4586 10084
rect 4709 10081 4721 10084
rect 4755 10081 4767 10115
rect 4709 10075 4767 10081
rect 5074 10072 5080 10124
rect 5132 10112 5138 10124
rect 5425 10115 5483 10121
rect 5425 10112 5437 10115
rect 5132 10084 5437 10112
rect 5132 10072 5138 10084
rect 5425 10081 5437 10084
rect 5471 10081 5483 10115
rect 5425 10075 5483 10081
rect 5810 10072 5816 10124
rect 5868 10112 5874 10124
rect 7024 10112 7052 10220
rect 8113 10217 8125 10220
rect 8159 10217 8171 10251
rect 8113 10211 8171 10217
rect 8294 10208 8300 10260
rect 8352 10248 8358 10260
rect 9125 10251 9183 10257
rect 9125 10248 9137 10251
rect 8352 10220 9137 10248
rect 8352 10208 8358 10220
rect 9125 10217 9137 10220
rect 9171 10217 9183 10251
rect 9125 10211 9183 10217
rect 9398 10208 9404 10260
rect 9456 10248 9462 10260
rect 9493 10251 9551 10257
rect 9493 10248 9505 10251
rect 9456 10220 9505 10248
rect 9456 10208 9462 10220
rect 9493 10217 9505 10220
rect 9539 10217 9551 10251
rect 9493 10211 9551 10217
rect 9585 10251 9643 10257
rect 9585 10217 9597 10251
rect 9631 10248 9643 10251
rect 9950 10248 9956 10260
rect 9631 10220 9956 10248
rect 9631 10217 9643 10220
rect 9585 10211 9643 10217
rect 9950 10208 9956 10220
rect 10008 10208 10014 10260
rect 10226 10208 10232 10260
rect 10284 10248 10290 10260
rect 10321 10251 10379 10257
rect 10321 10248 10333 10251
rect 10284 10220 10333 10248
rect 10284 10208 10290 10220
rect 10321 10217 10333 10220
rect 10367 10217 10379 10251
rect 10321 10211 10379 10217
rect 10689 10251 10747 10257
rect 10689 10217 10701 10251
rect 10735 10248 10747 10251
rect 11149 10251 11207 10257
rect 11149 10248 11161 10251
rect 10735 10220 11161 10248
rect 10735 10217 10747 10220
rect 10689 10211 10747 10217
rect 11149 10217 11161 10220
rect 11195 10217 11207 10251
rect 11149 10211 11207 10217
rect 11609 10251 11667 10257
rect 11609 10217 11621 10251
rect 11655 10248 11667 10251
rect 11977 10251 12035 10257
rect 11655 10220 11836 10248
rect 11655 10217 11667 10220
rect 11609 10211 11667 10217
rect 8481 10183 8539 10189
rect 8481 10149 8493 10183
rect 8527 10180 8539 10183
rect 8938 10180 8944 10192
rect 8527 10152 8944 10180
rect 8527 10149 8539 10152
rect 8481 10143 8539 10149
rect 8938 10140 8944 10152
rect 8996 10140 9002 10192
rect 9030 10140 9036 10192
rect 9088 10180 9094 10192
rect 9088 10152 10548 10180
rect 9088 10140 9094 10152
rect 5868 10084 7052 10112
rect 8573 10115 8631 10121
rect 5868 10072 5874 10084
rect 8573 10081 8585 10115
rect 8619 10112 8631 10115
rect 8619 10084 8800 10112
rect 8619 10081 8631 10084
rect 8573 10075 8631 10081
rect 2777 10047 2835 10053
rect 2777 10013 2789 10047
rect 2823 10013 2835 10047
rect 2777 10007 2835 10013
rect 2866 10004 2872 10056
rect 2924 10044 2930 10056
rect 3050 10044 3056 10056
rect 2924 10016 3056 10044
rect 2924 10004 2930 10016
rect 3050 10004 3056 10016
rect 3108 10004 3114 10056
rect 3605 10047 3663 10053
rect 3605 10013 3617 10047
rect 3651 10044 3663 10047
rect 4154 10044 4160 10056
rect 3651 10016 4160 10044
rect 3651 10013 3663 10016
rect 3605 10007 3663 10013
rect 4154 10004 4160 10016
rect 4212 10004 4218 10056
rect 4985 10047 5043 10053
rect 4985 10013 4997 10047
rect 5031 10013 5043 10047
rect 5166 10044 5172 10056
rect 5127 10016 5172 10044
rect 4985 10007 5043 10013
rect 1578 9936 1584 9988
rect 1636 9976 1642 9988
rect 4249 9979 4307 9985
rect 4249 9976 4261 9979
rect 1636 9948 3096 9976
rect 1636 9936 1642 9948
rect 1762 9908 1768 9920
rect 1723 9880 1768 9908
rect 1762 9868 1768 9880
rect 1820 9868 1826 9920
rect 2866 9868 2872 9920
rect 2924 9908 2930 9920
rect 2961 9911 3019 9917
rect 2961 9908 2973 9911
rect 2924 9880 2973 9908
rect 2924 9868 2930 9880
rect 2961 9877 2973 9880
rect 3007 9877 3019 9911
rect 3068 9908 3096 9948
rect 3896 9948 4261 9976
rect 3896 9908 3924 9948
rect 4249 9945 4261 9948
rect 4295 9976 4307 9979
rect 4706 9976 4712 9988
rect 4295 9948 4712 9976
rect 4295 9945 4307 9948
rect 4249 9939 4307 9945
rect 4706 9936 4712 9948
rect 4764 9936 4770 9988
rect 3068 9880 3924 9908
rect 3973 9911 4031 9917
rect 2961 9871 3019 9877
rect 3973 9877 3985 9911
rect 4019 9908 4031 9911
rect 4522 9908 4528 9920
rect 4019 9880 4528 9908
rect 4019 9877 4031 9880
rect 3973 9871 4031 9877
rect 4522 9868 4528 9880
rect 4580 9868 4586 9920
rect 5000 9908 5028 10007
rect 5166 10004 5172 10016
rect 5224 10004 5230 10056
rect 6641 10047 6699 10053
rect 6641 10013 6653 10047
rect 6687 10013 6699 10047
rect 8662 10044 8668 10056
rect 8623 10016 8668 10044
rect 6641 10007 6699 10013
rect 6270 9908 6276 9920
rect 5000 9880 6276 9908
rect 6270 9868 6276 9880
rect 6328 9868 6334 9920
rect 6546 9908 6552 9920
rect 6507 9880 6552 9908
rect 6546 9868 6552 9880
rect 6604 9868 6610 9920
rect 6656 9908 6684 10007
rect 8662 10004 8668 10016
rect 8720 10004 8726 10056
rect 8772 10044 8800 10084
rect 8846 10072 8852 10124
rect 8904 10112 8910 10124
rect 10410 10112 10416 10124
rect 8904 10084 9674 10112
rect 8904 10072 8910 10084
rect 9122 10044 9128 10056
rect 8772 10016 9128 10044
rect 9122 10004 9128 10016
rect 9180 10004 9186 10056
rect 9646 10044 9674 10084
rect 10060 10084 10416 10112
rect 10060 10053 10088 10084
rect 10410 10072 10416 10084
rect 10468 10072 10474 10124
rect 9769 10047 9827 10053
rect 9769 10044 9781 10047
rect 9646 10016 9781 10044
rect 9769 10013 9781 10016
rect 9815 10044 9827 10047
rect 10045 10047 10103 10053
rect 10045 10044 10057 10047
rect 9815 10016 10057 10044
rect 9815 10013 9827 10016
rect 9769 10007 9827 10013
rect 10045 10013 10057 10016
rect 10091 10013 10103 10047
rect 10045 10007 10103 10013
rect 10134 10004 10140 10056
rect 10192 10044 10198 10056
rect 10229 10047 10287 10053
rect 10229 10044 10241 10047
rect 10192 10016 10241 10044
rect 10192 10004 10198 10016
rect 10229 10013 10241 10016
rect 10275 10013 10287 10047
rect 10520 10044 10548 10152
rect 10778 10140 10784 10192
rect 10836 10180 10842 10192
rect 11241 10183 11299 10189
rect 11241 10180 11253 10183
rect 10836 10152 11253 10180
rect 10836 10140 10842 10152
rect 11241 10149 11253 10152
rect 11287 10149 11299 10183
rect 11241 10143 11299 10149
rect 11054 10072 11060 10124
rect 11112 10112 11118 10124
rect 11808 10112 11836 10220
rect 11977 10217 11989 10251
rect 12023 10248 12035 10251
rect 12250 10248 12256 10260
rect 12023 10220 12256 10248
rect 12023 10217 12035 10220
rect 11977 10211 12035 10217
rect 12250 10208 12256 10220
rect 12308 10208 12314 10260
rect 12437 10251 12495 10257
rect 12437 10217 12449 10251
rect 12483 10217 12495 10251
rect 12437 10211 12495 10217
rect 12066 10180 12072 10192
rect 12027 10152 12072 10180
rect 12066 10140 12072 10152
rect 12124 10140 12130 10192
rect 11974 10112 11980 10124
rect 11112 10084 11468 10112
rect 11808 10084 11980 10112
rect 11112 10072 11118 10084
rect 11333 10047 11391 10053
rect 11333 10044 11345 10047
rect 10520 10016 11345 10044
rect 10229 10007 10287 10013
rect 11333 10013 11345 10016
rect 11379 10013 11391 10047
rect 11440 10044 11468 10084
rect 11974 10072 11980 10084
rect 12032 10072 12038 10124
rect 12342 10072 12348 10124
rect 12400 10112 12406 10124
rect 12452 10112 12480 10211
rect 12526 10208 12532 10260
rect 12584 10248 12590 10260
rect 12897 10251 12955 10257
rect 12897 10248 12909 10251
rect 12584 10220 12909 10248
rect 12584 10208 12590 10220
rect 12897 10217 12909 10220
rect 12943 10217 12955 10251
rect 13262 10248 13268 10260
rect 13223 10220 13268 10248
rect 12897 10211 12955 10217
rect 13262 10208 13268 10220
rect 13320 10208 13326 10260
rect 13725 10251 13783 10257
rect 13725 10217 13737 10251
rect 13771 10248 13783 10251
rect 13814 10248 13820 10260
rect 13771 10220 13820 10248
rect 13771 10217 13783 10220
rect 13725 10211 13783 10217
rect 13814 10208 13820 10220
rect 13872 10208 13878 10260
rect 14090 10208 14096 10260
rect 14148 10248 14154 10260
rect 14829 10251 14887 10257
rect 14829 10248 14841 10251
rect 14148 10220 14841 10248
rect 14148 10208 14154 10220
rect 14829 10217 14841 10220
rect 14875 10217 14887 10251
rect 14829 10211 14887 10217
rect 13633 10183 13691 10189
rect 13633 10180 13645 10183
rect 12912 10152 13645 10180
rect 12400 10084 12480 10112
rect 12805 10115 12863 10121
rect 12400 10072 12406 10084
rect 12805 10081 12817 10115
rect 12851 10081 12863 10115
rect 12805 10075 12863 10081
rect 12161 10047 12219 10053
rect 12161 10044 12173 10047
rect 11440 10016 12173 10044
rect 11333 10007 11391 10013
rect 12161 10013 12173 10016
rect 12207 10013 12219 10047
rect 12161 10007 12219 10013
rect 12434 10004 12440 10056
rect 12492 10044 12498 10056
rect 12820 10044 12848 10075
rect 12492 10016 12848 10044
rect 12492 10004 12498 10016
rect 8018 9976 8024 9988
rect 7979 9948 8024 9976
rect 8018 9936 8024 9948
rect 8076 9976 8082 9988
rect 8076 9948 10456 9976
rect 8076 9936 8082 9948
rect 7926 9908 7932 9920
rect 6656 9880 7932 9908
rect 7926 9868 7932 9880
rect 7984 9868 7990 9920
rect 9030 9868 9036 9920
rect 9088 9908 9094 9920
rect 9306 9908 9312 9920
rect 9088 9880 9312 9908
rect 9088 9868 9094 9880
rect 9306 9868 9312 9880
rect 9364 9868 9370 9920
rect 9674 9868 9680 9920
rect 9732 9908 9738 9920
rect 10042 9908 10048 9920
rect 9732 9880 10048 9908
rect 9732 9868 9738 9880
rect 10042 9868 10048 9880
rect 10100 9868 10106 9920
rect 10428 9908 10456 9948
rect 10502 9936 10508 9988
rect 10560 9976 10566 9988
rect 10781 9979 10839 9985
rect 10781 9976 10793 9979
rect 10560 9948 10793 9976
rect 10560 9936 10566 9948
rect 10781 9945 10793 9948
rect 10827 9945 10839 9979
rect 10781 9939 10839 9945
rect 11238 9936 11244 9988
rect 11296 9976 11302 9988
rect 12710 9976 12716 9988
rect 11296 9948 12716 9976
rect 11296 9936 11302 9948
rect 12710 9936 12716 9948
rect 12768 9936 12774 9988
rect 10594 9908 10600 9920
rect 10428 9880 10600 9908
rect 10594 9868 10600 9880
rect 10652 9908 10658 9920
rect 11054 9908 11060 9920
rect 10652 9880 11060 9908
rect 10652 9868 10658 9880
rect 11054 9868 11060 9880
rect 11112 9868 11118 9920
rect 11146 9868 11152 9920
rect 11204 9908 11210 9920
rect 12912 9908 12940 10152
rect 13633 10149 13645 10152
rect 13679 10149 13691 10183
rect 14274 10180 14280 10192
rect 13633 10143 13691 10149
rect 13740 10152 14280 10180
rect 13262 10072 13268 10124
rect 13320 10112 13326 10124
rect 13740 10112 13768 10152
rect 14274 10140 14280 10152
rect 14332 10140 14338 10192
rect 13320 10084 13768 10112
rect 13320 10072 13326 10084
rect 13906 10072 13912 10124
rect 13964 10112 13970 10124
rect 14093 10115 14151 10121
rect 14093 10112 14105 10115
rect 13964 10084 14105 10112
rect 13964 10072 13970 10084
rect 14093 10081 14105 10084
rect 14139 10112 14151 10115
rect 14182 10112 14188 10124
rect 14139 10084 14188 10112
rect 14139 10081 14151 10084
rect 14093 10075 14151 10081
rect 14182 10072 14188 10084
rect 14240 10112 14246 10124
rect 14737 10115 14795 10121
rect 14737 10112 14749 10115
rect 14240 10084 14749 10112
rect 14240 10072 14246 10084
rect 14737 10081 14749 10084
rect 14783 10081 14795 10115
rect 15470 10112 15476 10124
rect 15431 10084 15476 10112
rect 14737 10075 14795 10081
rect 15470 10072 15476 10084
rect 15528 10072 15534 10124
rect 13081 10047 13139 10053
rect 13081 10013 13093 10047
rect 13127 10044 13139 10047
rect 13446 10044 13452 10056
rect 13127 10016 13452 10044
rect 13127 10013 13139 10016
rect 13081 10007 13139 10013
rect 13446 10004 13452 10016
rect 13504 10044 13510 10056
rect 13817 10047 13875 10053
rect 13817 10044 13829 10047
rect 13504 10016 13829 10044
rect 13504 10004 13510 10016
rect 13817 10013 13829 10016
rect 13863 10013 13875 10047
rect 13817 10007 13875 10013
rect 14826 10004 14832 10056
rect 14884 10044 14890 10056
rect 14921 10047 14979 10053
rect 14921 10044 14933 10047
rect 14884 10016 14933 10044
rect 14884 10004 14890 10016
rect 14921 10013 14933 10016
rect 14967 10013 14979 10047
rect 14921 10007 14979 10013
rect 14366 9976 14372 9988
rect 14327 9948 14372 9976
rect 14366 9936 14372 9948
rect 14424 9936 14430 9988
rect 15654 9976 15660 9988
rect 15615 9948 15660 9976
rect 15654 9936 15660 9948
rect 15712 9936 15718 9988
rect 11204 9880 12940 9908
rect 11204 9868 11210 9880
rect 13998 9868 14004 9920
rect 14056 9908 14062 9920
rect 15197 9911 15255 9917
rect 15197 9908 15209 9911
rect 14056 9880 15209 9908
rect 14056 9868 14062 9880
rect 15197 9877 15209 9880
rect 15243 9877 15255 9911
rect 15197 9871 15255 9877
rect 1104 9818 16008 9840
rect 1104 9766 3480 9818
rect 3532 9766 3544 9818
rect 3596 9766 3608 9818
rect 3660 9766 3672 9818
rect 3724 9766 8478 9818
rect 8530 9766 8542 9818
rect 8594 9766 8606 9818
rect 8658 9766 8670 9818
rect 8722 9766 13475 9818
rect 13527 9766 13539 9818
rect 13591 9766 13603 9818
rect 13655 9766 13667 9818
rect 13719 9766 16008 9818
rect 1104 9744 16008 9766
rect 2424 9676 2912 9704
rect 2222 9596 2228 9648
rect 2280 9636 2286 9648
rect 2424 9636 2452 9676
rect 2280 9608 2452 9636
rect 2501 9639 2559 9645
rect 2280 9596 2286 9608
rect 2501 9605 2513 9639
rect 2547 9636 2559 9639
rect 2774 9636 2780 9648
rect 2547 9608 2780 9636
rect 2547 9605 2559 9608
rect 2501 9599 2559 9605
rect 2774 9596 2780 9608
rect 2832 9596 2838 9648
rect 2884 9636 2912 9676
rect 3234 9664 3240 9716
rect 3292 9704 3298 9716
rect 11238 9704 11244 9716
rect 3292 9676 11244 9704
rect 3292 9664 3298 9676
rect 11238 9664 11244 9676
rect 11296 9664 11302 9716
rect 11517 9707 11575 9713
rect 11517 9673 11529 9707
rect 11563 9704 11575 9707
rect 11606 9704 11612 9716
rect 11563 9676 11612 9704
rect 11563 9673 11575 9676
rect 11517 9667 11575 9673
rect 11606 9664 11612 9676
rect 11664 9664 11670 9716
rect 11698 9664 11704 9716
rect 11756 9704 11762 9716
rect 11756 9676 11801 9704
rect 11756 9664 11762 9676
rect 11974 9664 11980 9716
rect 12032 9704 12038 9716
rect 12894 9704 12900 9716
rect 12032 9676 12900 9704
rect 12032 9664 12038 9676
rect 12894 9664 12900 9676
rect 12952 9664 12958 9716
rect 15197 9707 15255 9713
rect 13280 9676 13952 9704
rect 3326 9636 3332 9648
rect 2884 9608 3332 9636
rect 3326 9596 3332 9608
rect 3384 9636 3390 9648
rect 3384 9608 3464 9636
rect 3384 9596 3390 9608
rect 1949 9571 2007 9577
rect 1949 9537 1961 9571
rect 1995 9568 2007 9571
rect 2314 9568 2320 9580
rect 1995 9540 2320 9568
rect 1995 9537 2007 9540
rect 1949 9531 2007 9537
rect 2314 9528 2320 9540
rect 2372 9528 2378 9580
rect 2866 9528 2872 9580
rect 2924 9528 2930 9580
rect 3234 9568 3240 9580
rect 3195 9540 3240 9568
rect 3234 9528 3240 9540
rect 3292 9528 3298 9580
rect 3436 9577 3464 9608
rect 4614 9596 4620 9648
rect 4672 9636 4678 9648
rect 4801 9639 4859 9645
rect 4801 9636 4813 9639
rect 4672 9608 4813 9636
rect 4672 9596 4678 9608
rect 4801 9605 4813 9608
rect 4847 9605 4859 9639
rect 6270 9636 6276 9648
rect 6231 9608 6276 9636
rect 4801 9599 4859 9605
rect 6270 9596 6276 9608
rect 6328 9596 6334 9648
rect 6454 9636 6460 9648
rect 6415 9608 6460 9636
rect 6454 9596 6460 9608
rect 6512 9596 6518 9648
rect 7650 9636 7656 9648
rect 7484 9608 7656 9636
rect 3421 9571 3479 9577
rect 3421 9537 3433 9571
rect 3467 9537 3479 9571
rect 3421 9531 3479 9537
rect 1394 9500 1400 9512
rect 1355 9472 1400 9500
rect 1394 9460 1400 9472
rect 1452 9460 1458 9512
rect 2133 9503 2191 9509
rect 2133 9469 2145 9503
rect 2179 9500 2191 9503
rect 2884 9500 2912 9528
rect 2179 9472 2912 9500
rect 3436 9500 3464 9531
rect 4430 9528 4436 9580
rect 4488 9568 4494 9580
rect 4488 9540 5028 9568
rect 4488 9528 4494 9540
rect 4890 9500 4896 9512
rect 3436 9472 4896 9500
rect 2179 9469 2191 9472
rect 2133 9463 2191 9469
rect 4890 9460 4896 9472
rect 4948 9460 4954 9512
rect 5000 9500 5028 9540
rect 6546 9528 6552 9580
rect 6604 9568 6610 9580
rect 7484 9577 7512 9608
rect 7650 9596 7656 9608
rect 7708 9596 7714 9648
rect 9125 9639 9183 9645
rect 9125 9605 9137 9639
rect 9171 9605 9183 9639
rect 9125 9599 9183 9605
rect 9309 9639 9367 9645
rect 9309 9605 9321 9639
rect 9355 9636 9367 9639
rect 9398 9636 9404 9648
rect 9355 9608 9404 9636
rect 9355 9605 9367 9608
rect 9309 9599 9367 9605
rect 7009 9571 7067 9577
rect 7009 9568 7021 9571
rect 6604 9540 7021 9568
rect 6604 9528 6610 9540
rect 7009 9537 7021 9540
rect 7055 9537 7067 9571
rect 7009 9531 7067 9537
rect 7469 9571 7527 9577
rect 7469 9537 7481 9571
rect 7515 9537 7527 9571
rect 7469 9531 7527 9537
rect 7745 9571 7803 9577
rect 7745 9537 7757 9571
rect 7791 9568 7803 9571
rect 9140 9568 9168 9599
rect 9398 9596 9404 9608
rect 9456 9596 9462 9648
rect 10502 9596 10508 9648
rect 10560 9636 10566 9648
rect 11149 9639 11207 9645
rect 11149 9636 11161 9639
rect 10560 9608 11161 9636
rect 10560 9596 10566 9608
rect 11149 9605 11161 9608
rect 11195 9605 11207 9639
rect 13280 9636 13308 9676
rect 11149 9599 11207 9605
rect 11256 9608 12388 9636
rect 11256 9568 11284 9608
rect 12360 9580 12388 9608
rect 12452 9608 13308 9636
rect 13357 9639 13415 9645
rect 12158 9568 12164 9580
rect 7791 9540 7880 9568
rect 9140 9540 9536 9568
rect 7791 9537 7803 9540
rect 7745 9531 7803 9537
rect 7852 9512 7880 9540
rect 5160 9503 5218 9509
rect 5160 9500 5172 9503
rect 5000 9472 5172 9500
rect 5160 9469 5172 9472
rect 5206 9500 5218 9503
rect 5206 9472 5396 9500
rect 5206 9469 5218 9472
rect 5160 9463 5218 9469
rect 1581 9435 1639 9441
rect 1581 9401 1593 9435
rect 1627 9432 1639 9435
rect 1854 9432 1860 9444
rect 1627 9404 1860 9432
rect 1627 9401 1639 9404
rect 1581 9395 1639 9401
rect 1854 9392 1860 9404
rect 1912 9392 1918 9444
rect 2041 9435 2099 9441
rect 2041 9401 2053 9435
rect 2087 9432 2099 9435
rect 3688 9435 3746 9441
rect 2087 9404 2636 9432
rect 2087 9401 2099 9404
rect 2041 9395 2099 9401
rect 2608 9373 2636 9404
rect 3688 9401 3700 9435
rect 3734 9432 3746 9435
rect 3734 9404 4200 9432
rect 3734 9401 3746 9404
rect 3688 9395 3746 9401
rect 2593 9367 2651 9373
rect 2593 9333 2605 9367
rect 2639 9333 2651 9367
rect 2958 9364 2964 9376
rect 2919 9336 2964 9364
rect 2593 9327 2651 9333
rect 2958 9324 2964 9336
rect 3016 9324 3022 9376
rect 3050 9324 3056 9376
rect 3108 9364 3114 9376
rect 4172 9364 4200 9404
rect 4246 9392 4252 9444
rect 4304 9432 4310 9444
rect 5368 9432 5396 9472
rect 7300 9472 7788 9500
rect 7300 9432 7328 9472
rect 4304 9404 5304 9432
rect 5368 9404 7328 9432
rect 4304 9392 4310 9404
rect 4798 9364 4804 9376
rect 3108 9336 3153 9364
rect 4172 9336 4804 9364
rect 3108 9324 3114 9336
rect 4798 9324 4804 9336
rect 4856 9324 4862 9376
rect 5276 9364 5304 9404
rect 5442 9364 5448 9376
rect 5276 9336 5448 9364
rect 5442 9324 5448 9336
rect 5500 9324 5506 9376
rect 5534 9324 5540 9376
rect 5592 9364 5598 9376
rect 6822 9364 6828 9376
rect 5592 9336 6828 9364
rect 5592 9324 5598 9336
rect 6822 9324 6828 9336
rect 6880 9324 6886 9376
rect 6917 9367 6975 9373
rect 6917 9333 6929 9367
rect 6963 9364 6975 9367
rect 7466 9364 7472 9376
rect 6963 9336 7472 9364
rect 6963 9333 6975 9336
rect 6917 9327 6975 9333
rect 7466 9324 7472 9336
rect 7524 9364 7530 9376
rect 7561 9367 7619 9373
rect 7561 9364 7573 9367
rect 7524 9336 7573 9364
rect 7524 9324 7530 9336
rect 7561 9333 7573 9336
rect 7607 9333 7619 9367
rect 7760 9364 7788 9472
rect 7834 9460 7840 9512
rect 7892 9500 7898 9512
rect 9122 9500 9128 9512
rect 7892 9472 9128 9500
rect 7892 9460 7898 9472
rect 9122 9460 9128 9472
rect 9180 9500 9186 9512
rect 9401 9503 9459 9509
rect 9401 9500 9413 9503
rect 9180 9472 9413 9500
rect 9180 9460 9186 9472
rect 9401 9469 9413 9472
rect 9447 9469 9459 9503
rect 9401 9463 9459 9469
rect 9508 9500 9536 9540
rect 10980 9540 11284 9568
rect 11532 9540 12020 9568
rect 12119 9540 12164 9568
rect 10980 9500 11008 9540
rect 9508 9472 11008 9500
rect 8012 9435 8070 9441
rect 8012 9401 8024 9435
rect 8058 9432 8070 9435
rect 9030 9432 9036 9444
rect 8058 9404 9036 9432
rect 8058 9401 8070 9404
rect 8012 9395 8070 9401
rect 9030 9392 9036 9404
rect 9088 9392 9094 9444
rect 9306 9392 9312 9444
rect 9364 9432 9370 9444
rect 9508 9432 9536 9472
rect 11146 9460 11152 9512
rect 11204 9460 11210 9512
rect 11330 9500 11336 9512
rect 11291 9472 11336 9500
rect 11330 9460 11336 9472
rect 11388 9460 11394 9512
rect 9364 9404 9536 9432
rect 9364 9392 9370 9404
rect 9582 9392 9588 9444
rect 9640 9441 9646 9444
rect 9640 9435 9704 9441
rect 9640 9401 9658 9435
rect 9692 9401 9704 9435
rect 9640 9395 9704 9401
rect 9640 9392 9646 9395
rect 9766 9392 9772 9444
rect 9824 9432 9830 9444
rect 10962 9432 10968 9444
rect 9824 9404 10968 9432
rect 9824 9392 9830 9404
rect 10962 9392 10968 9404
rect 11020 9392 11026 9444
rect 11057 9435 11115 9441
rect 11057 9401 11069 9435
rect 11103 9432 11115 9435
rect 11164 9432 11192 9460
rect 11103 9404 11192 9432
rect 11103 9401 11115 9404
rect 11057 9395 11115 9401
rect 10781 9367 10839 9373
rect 10781 9364 10793 9367
rect 7760 9336 10793 9364
rect 7561 9327 7619 9333
rect 10781 9333 10793 9336
rect 10827 9364 10839 9367
rect 11532 9364 11560 9540
rect 11992 9432 12020 9540
rect 12158 9528 12164 9540
rect 12216 9528 12222 9580
rect 12342 9568 12348 9580
rect 12303 9540 12348 9568
rect 12342 9528 12348 9540
rect 12400 9528 12406 9580
rect 12069 9503 12127 9509
rect 12069 9469 12081 9503
rect 12115 9500 12127 9503
rect 12250 9500 12256 9512
rect 12115 9472 12256 9500
rect 12115 9469 12127 9472
rect 12069 9463 12127 9469
rect 12250 9460 12256 9472
rect 12308 9460 12314 9512
rect 12452 9432 12480 9608
rect 13357 9605 13369 9639
rect 13403 9605 13415 9639
rect 13357 9599 13415 9605
rect 12526 9528 12532 9580
rect 12584 9568 12590 9580
rect 12621 9571 12679 9577
rect 12621 9568 12633 9571
rect 12584 9540 12633 9568
rect 12584 9528 12590 9540
rect 12621 9537 12633 9540
rect 12667 9537 12679 9571
rect 12621 9531 12679 9537
rect 12710 9528 12716 9580
rect 12768 9568 12774 9580
rect 13372 9568 13400 9599
rect 13924 9577 13952 9676
rect 15197 9673 15209 9707
rect 15243 9704 15255 9707
rect 15470 9704 15476 9716
rect 15243 9676 15476 9704
rect 15243 9673 15255 9676
rect 15197 9667 15255 9673
rect 15470 9664 15476 9676
rect 15528 9664 15534 9716
rect 12768 9540 13400 9568
rect 13909 9571 13967 9577
rect 12768 9528 12774 9540
rect 13909 9537 13921 9571
rect 13955 9568 13967 9571
rect 14274 9568 14280 9580
rect 13955 9540 14280 9568
rect 13955 9537 13967 9540
rect 13909 9531 13967 9537
rect 14274 9528 14280 9540
rect 14332 9528 14338 9580
rect 12802 9500 12808 9512
rect 12763 9472 12808 9500
rect 12802 9460 12808 9472
rect 12860 9460 12866 9512
rect 14553 9503 14611 9509
rect 14553 9500 14565 9503
rect 13096 9472 14565 9500
rect 13096 9432 13124 9472
rect 14553 9469 14565 9472
rect 14599 9469 14611 9503
rect 14553 9463 14611 9469
rect 15013 9503 15071 9509
rect 15013 9469 15025 9503
rect 15059 9500 15071 9503
rect 15102 9500 15108 9512
rect 15059 9472 15108 9500
rect 15059 9469 15071 9472
rect 15013 9463 15071 9469
rect 15102 9460 15108 9472
rect 15160 9460 15166 9512
rect 13817 9435 13875 9441
rect 13817 9432 13829 9435
rect 11992 9404 12480 9432
rect 12544 9404 13124 9432
rect 13280 9404 13829 9432
rect 10827 9336 11560 9364
rect 10827 9333 10839 9336
rect 10781 9327 10839 9333
rect 11882 9324 11888 9376
rect 11940 9364 11946 9376
rect 12544 9364 12572 9404
rect 11940 9336 12572 9364
rect 11940 9324 11946 9336
rect 12894 9324 12900 9376
rect 12952 9364 12958 9376
rect 13280 9373 13308 9404
rect 13817 9401 13829 9404
rect 13863 9401 13875 9435
rect 15470 9432 15476 9444
rect 15431 9404 15476 9432
rect 13817 9395 13875 9401
rect 15470 9392 15476 9404
rect 15528 9392 15534 9444
rect 13265 9367 13323 9373
rect 12952 9336 12997 9364
rect 12952 9324 12958 9336
rect 13265 9333 13277 9367
rect 13311 9333 13323 9367
rect 13722 9364 13728 9376
rect 13683 9336 13728 9364
rect 13265 9327 13323 9333
rect 13722 9324 13728 9336
rect 13780 9324 13786 9376
rect 14458 9364 14464 9376
rect 14419 9336 14464 9364
rect 14458 9324 14464 9336
rect 14516 9324 14522 9376
rect 14734 9324 14740 9376
rect 14792 9364 14798 9376
rect 14921 9367 14979 9373
rect 14921 9364 14933 9367
rect 14792 9336 14933 9364
rect 14792 9324 14798 9336
rect 14921 9333 14933 9336
rect 14967 9333 14979 9367
rect 14921 9327 14979 9333
rect 15102 9324 15108 9376
rect 15160 9364 15166 9376
rect 15289 9367 15347 9373
rect 15289 9364 15301 9367
rect 15160 9336 15301 9364
rect 15160 9324 15166 9336
rect 15289 9333 15301 9336
rect 15335 9333 15347 9367
rect 15289 9327 15347 9333
rect 1104 9274 16008 9296
rect 1104 9222 5979 9274
rect 6031 9222 6043 9274
rect 6095 9222 6107 9274
rect 6159 9222 6171 9274
rect 6223 9222 10976 9274
rect 11028 9222 11040 9274
rect 11092 9222 11104 9274
rect 11156 9222 11168 9274
rect 11220 9222 16008 9274
rect 1104 9200 16008 9222
rect 1486 9160 1492 9172
rect 1447 9132 1492 9160
rect 1486 9120 1492 9132
rect 1544 9120 1550 9172
rect 1854 9160 1860 9172
rect 1815 9132 1860 9160
rect 1854 9120 1860 9132
rect 1912 9120 1918 9172
rect 2869 9163 2927 9169
rect 2869 9129 2881 9163
rect 2915 9160 2927 9163
rect 3050 9160 3056 9172
rect 2915 9132 3056 9160
rect 2915 9129 2927 9132
rect 2869 9123 2927 9129
rect 3050 9120 3056 9132
rect 3108 9120 3114 9172
rect 3329 9163 3387 9169
rect 3329 9129 3341 9163
rect 3375 9160 3387 9163
rect 3602 9160 3608 9172
rect 3375 9132 3608 9160
rect 3375 9129 3387 9132
rect 3329 9123 3387 9129
rect 3602 9120 3608 9132
rect 3660 9120 3666 9172
rect 3970 9160 3976 9172
rect 3931 9132 3976 9160
rect 3970 9120 3976 9132
rect 4028 9120 4034 9172
rect 8849 9163 8907 9169
rect 4908 9132 8800 9160
rect 2958 9052 2964 9104
rect 3016 9092 3022 9104
rect 4908 9092 4936 9132
rect 3016 9064 4936 9092
rect 3016 9052 3022 9064
rect 4982 9052 4988 9104
rect 5040 9092 5046 9104
rect 5690 9095 5748 9101
rect 5690 9092 5702 9095
rect 5040 9064 5702 9092
rect 5040 9052 5046 9064
rect 5690 9061 5702 9064
rect 5736 9061 5748 9095
rect 5690 9055 5748 9061
rect 6270 9052 6276 9104
rect 6328 9092 6334 9104
rect 7926 9092 7932 9104
rect 6328 9064 7932 9092
rect 6328 9052 6334 9064
rect 7926 9052 7932 9064
rect 7984 9052 7990 9104
rect 1578 9024 1584 9036
rect 1539 8996 1584 9024
rect 1578 8984 1584 8996
rect 1636 8984 1642 9036
rect 2041 9027 2099 9033
rect 2041 8993 2053 9027
rect 2087 9024 2099 9027
rect 2130 9024 2136 9036
rect 2087 8996 2136 9024
rect 2087 8993 2099 8996
rect 2041 8987 2099 8993
rect 2130 8984 2136 8996
rect 2188 8984 2194 9036
rect 2406 9024 2412 9036
rect 2367 8996 2412 9024
rect 2406 8984 2412 8996
rect 2464 8984 2470 9036
rect 2498 8984 2504 9036
rect 2556 9024 2562 9036
rect 3421 9027 3479 9033
rect 2556 8996 2601 9024
rect 2556 8984 2562 8996
rect 3421 8993 3433 9027
rect 3467 9024 3479 9027
rect 4062 9024 4068 9036
rect 3467 8996 4068 9024
rect 3467 8993 3479 8996
rect 3421 8987 3479 8993
rect 4062 8984 4068 8996
rect 4120 8984 4126 9036
rect 4338 8984 4344 9036
rect 4396 9024 4402 9036
rect 5097 9027 5155 9033
rect 5097 9024 5109 9027
rect 4396 8996 5109 9024
rect 4396 8984 4402 8996
rect 5097 8993 5109 8996
rect 5143 9024 5155 9027
rect 6288 9024 6316 9052
rect 8041 9027 8099 9033
rect 8041 9024 8053 9027
rect 5143 8996 6316 9024
rect 7300 8996 8053 9024
rect 5143 8993 5155 8996
rect 5097 8987 5155 8993
rect 2317 8959 2375 8965
rect 2317 8925 2329 8959
rect 2363 8925 2375 8959
rect 2317 8919 2375 8925
rect 3605 8959 3663 8965
rect 3605 8925 3617 8959
rect 3651 8956 3663 8959
rect 4154 8956 4160 8968
rect 3651 8928 4160 8956
rect 3651 8925 3663 8928
rect 3605 8919 3663 8925
rect 2332 8888 2360 8919
rect 2332 8860 3188 8888
rect 1765 8823 1823 8829
rect 1765 8789 1777 8823
rect 1811 8820 1823 8823
rect 1854 8820 1860 8832
rect 1811 8792 1860 8820
rect 1811 8789 1823 8792
rect 1765 8783 1823 8789
rect 1854 8780 1860 8792
rect 1912 8780 1918 8832
rect 2130 8780 2136 8832
rect 2188 8820 2194 8832
rect 2961 8823 3019 8829
rect 2961 8820 2973 8823
rect 2188 8792 2973 8820
rect 2188 8780 2194 8792
rect 2961 8789 2973 8792
rect 3007 8789 3019 8823
rect 3160 8820 3188 8860
rect 3234 8848 3240 8900
rect 3292 8888 3298 8900
rect 3620 8888 3648 8919
rect 4154 8916 4160 8928
rect 4212 8916 4218 8968
rect 5350 8956 5356 8968
rect 5311 8928 5356 8956
rect 5350 8916 5356 8928
rect 5408 8956 5414 8968
rect 5445 8959 5503 8965
rect 5445 8956 5457 8959
rect 5408 8928 5457 8956
rect 5408 8916 5414 8928
rect 5445 8925 5457 8928
rect 5491 8925 5503 8959
rect 5445 8919 5503 8925
rect 4338 8888 4344 8900
rect 3292 8860 3648 8888
rect 4080 8860 4344 8888
rect 3292 8848 3298 8860
rect 4080 8820 4108 8860
rect 4338 8848 4344 8860
rect 4396 8848 4402 8900
rect 6825 8891 6883 8897
rect 6825 8857 6837 8891
rect 6871 8888 6883 8891
rect 7300 8888 7328 8996
rect 8041 8993 8053 8996
rect 8087 9024 8099 9027
rect 8202 9024 8208 9036
rect 8087 8996 8208 9024
rect 8087 8993 8099 8996
rect 8041 8987 8099 8993
rect 8202 8984 8208 8996
rect 8260 8984 8266 9036
rect 8772 9024 8800 9132
rect 8849 9129 8861 9163
rect 8895 9160 8907 9163
rect 9766 9160 9772 9172
rect 8895 9132 9772 9160
rect 8895 9129 8907 9132
rect 8849 9123 8907 9129
rect 9766 9120 9772 9132
rect 9824 9120 9830 9172
rect 10505 9163 10563 9169
rect 10505 9129 10517 9163
rect 10551 9160 10563 9163
rect 10778 9160 10784 9172
rect 10551 9132 10784 9160
rect 10551 9129 10563 9132
rect 10505 9123 10563 9129
rect 10778 9120 10784 9132
rect 10836 9160 10842 9172
rect 11330 9160 11336 9172
rect 10836 9132 11192 9160
rect 11291 9132 11336 9160
rect 10836 9120 10842 9132
rect 9306 9052 9312 9104
rect 9364 9101 9370 9104
rect 9364 9095 9428 9101
rect 9364 9061 9382 9095
rect 9416 9061 9428 9095
rect 9364 9055 9428 9061
rect 9364 9052 9370 9055
rect 9490 9052 9496 9104
rect 9548 9092 9554 9104
rect 11054 9092 11060 9104
rect 9548 9064 11060 9092
rect 9548 9052 9554 9064
rect 11054 9052 11060 9064
rect 11112 9052 11118 9104
rect 8772 8996 10180 9024
rect 8297 8959 8355 8965
rect 8297 8925 8309 8959
rect 8343 8925 8355 8959
rect 8297 8919 8355 8925
rect 8573 8959 8631 8965
rect 8573 8925 8585 8959
rect 8619 8956 8631 8959
rect 9030 8956 9036 8968
rect 8619 8928 9036 8956
rect 8619 8925 8631 8928
rect 8573 8919 8631 8925
rect 6871 8860 7328 8888
rect 6871 8857 6883 8860
rect 6825 8851 6883 8857
rect 3160 8792 4108 8820
rect 2961 8783 3019 8789
rect 4154 8780 4160 8832
rect 4212 8820 4218 8832
rect 5166 8820 5172 8832
rect 4212 8792 5172 8820
rect 4212 8780 4218 8792
rect 5166 8780 5172 8792
rect 5224 8780 5230 8832
rect 6914 8820 6920 8832
rect 6875 8792 6920 8820
rect 6914 8780 6920 8792
rect 6972 8780 6978 8832
rect 7926 8780 7932 8832
rect 7984 8820 7990 8832
rect 8312 8820 8340 8919
rect 9030 8916 9036 8928
rect 9088 8916 9094 8968
rect 9122 8916 9128 8968
rect 9180 8956 9186 8968
rect 9180 8928 9225 8956
rect 9180 8916 9186 8928
rect 10152 8888 10180 8996
rect 10502 8984 10508 9036
rect 10560 9024 10566 9036
rect 10962 9024 10968 9036
rect 10560 8996 10824 9024
rect 10923 8996 10968 9024
rect 10560 8984 10566 8996
rect 10594 8916 10600 8968
rect 10652 8956 10658 8968
rect 10689 8959 10747 8965
rect 10689 8956 10701 8959
rect 10652 8928 10701 8956
rect 10652 8916 10658 8928
rect 10689 8925 10701 8928
rect 10735 8925 10747 8959
rect 10796 8956 10824 8996
rect 10962 8984 10968 8996
rect 11020 8984 11026 9036
rect 11164 9024 11192 9132
rect 11330 9120 11336 9132
rect 11388 9120 11394 9172
rect 11701 9163 11759 9169
rect 11440 9132 11652 9160
rect 11238 9052 11244 9104
rect 11296 9092 11302 9104
rect 11440 9092 11468 9132
rect 11296 9064 11468 9092
rect 11624 9092 11652 9132
rect 11701 9129 11713 9163
rect 11747 9160 11759 9163
rect 11974 9160 11980 9172
rect 11747 9132 11980 9160
rect 11747 9129 11759 9132
rect 11701 9123 11759 9129
rect 11974 9120 11980 9132
rect 12032 9120 12038 9172
rect 12161 9163 12219 9169
rect 12161 9129 12173 9163
rect 12207 9160 12219 9163
rect 12618 9160 12624 9172
rect 12207 9132 12624 9160
rect 12207 9129 12219 9132
rect 12161 9123 12219 9129
rect 12618 9120 12624 9132
rect 12676 9120 12682 9172
rect 12802 9120 12808 9172
rect 12860 9160 12866 9172
rect 13081 9163 13139 9169
rect 13081 9160 13093 9163
rect 12860 9132 13093 9160
rect 12860 9120 12866 9132
rect 13081 9129 13093 9132
rect 13127 9129 13139 9163
rect 13081 9123 13139 9129
rect 13446 9120 13452 9172
rect 13504 9160 13510 9172
rect 13541 9163 13599 9169
rect 13541 9160 13553 9163
rect 13504 9132 13553 9160
rect 13504 9120 13510 9132
rect 13541 9129 13553 9132
rect 13587 9129 13599 9163
rect 13541 9123 13599 9129
rect 13906 9120 13912 9172
rect 13964 9160 13970 9172
rect 14369 9163 14427 9169
rect 14369 9160 14381 9163
rect 13964 9132 14381 9160
rect 13964 9120 13970 9132
rect 14369 9129 14381 9132
rect 14415 9129 14427 9163
rect 14734 9160 14740 9172
rect 14695 9132 14740 9160
rect 14369 9123 14427 9129
rect 14734 9120 14740 9132
rect 14792 9120 14798 9172
rect 11624 9064 14964 9092
rect 11296 9052 11302 9064
rect 11164 8996 11652 9024
rect 10873 8959 10931 8965
rect 10873 8956 10885 8959
rect 10796 8928 10885 8956
rect 10689 8919 10747 8925
rect 10873 8925 10885 8928
rect 10919 8956 10931 8959
rect 11330 8956 11336 8968
rect 10919 8928 11336 8956
rect 10919 8925 10931 8928
rect 10873 8919 10931 8925
rect 11330 8916 11336 8928
rect 11388 8916 11394 8968
rect 11514 8956 11520 8968
rect 11475 8928 11520 8956
rect 11514 8916 11520 8928
rect 11572 8916 11578 8968
rect 11624 8956 11652 8996
rect 11698 8984 11704 9036
rect 11756 9024 11762 9036
rect 11793 9027 11851 9033
rect 11793 9024 11805 9027
rect 11756 8996 11805 9024
rect 11756 8984 11762 8996
rect 11793 8993 11805 8996
rect 11839 8993 11851 9027
rect 11793 8987 11851 8993
rect 11882 8984 11888 9036
rect 11940 9024 11946 9036
rect 12621 9027 12679 9033
rect 12621 9024 12633 9027
rect 11940 8996 12633 9024
rect 11940 8984 11946 8996
rect 12621 8993 12633 8996
rect 12667 8993 12679 9027
rect 12621 8987 12679 8993
rect 13449 9027 13507 9033
rect 13449 8993 13461 9027
rect 13495 9024 13507 9027
rect 13495 8996 14320 9024
rect 13495 8993 13507 8996
rect 13449 8987 13507 8993
rect 12342 8956 12348 8968
rect 11624 8928 12348 8956
rect 12342 8916 12348 8928
rect 12400 8916 12406 8968
rect 12710 8916 12716 8968
rect 12768 8956 12774 8968
rect 12894 8956 12900 8968
rect 12768 8928 12813 8956
rect 12855 8928 12900 8956
rect 12768 8916 12774 8928
rect 12894 8916 12900 8928
rect 12952 8916 12958 8968
rect 13354 8916 13360 8968
rect 13412 8956 13418 8968
rect 13633 8959 13691 8965
rect 13633 8956 13645 8959
rect 13412 8928 13645 8956
rect 13412 8916 13418 8928
rect 13633 8925 13645 8928
rect 13679 8956 13691 8959
rect 13814 8956 13820 8968
rect 13679 8928 13820 8956
rect 13679 8925 13691 8928
rect 13633 8919 13691 8925
rect 13814 8916 13820 8928
rect 13872 8916 13878 8968
rect 12253 8891 12311 8897
rect 12253 8888 12265 8891
rect 10152 8860 12265 8888
rect 12253 8857 12265 8860
rect 12299 8857 12311 8891
rect 12253 8851 12311 8857
rect 12986 8848 12992 8900
rect 13044 8888 13050 8900
rect 13446 8888 13452 8900
rect 13044 8860 13452 8888
rect 13044 8848 13050 8860
rect 13446 8848 13452 8860
rect 13504 8888 13510 8900
rect 13909 8891 13967 8897
rect 13909 8888 13921 8891
rect 13504 8860 13921 8888
rect 13504 8848 13510 8860
rect 13909 8857 13921 8860
rect 13955 8857 13967 8891
rect 14292 8888 14320 8996
rect 14826 8956 14832 8968
rect 14787 8928 14832 8956
rect 14826 8916 14832 8928
rect 14884 8916 14890 8968
rect 14936 8965 14964 9064
rect 15194 8984 15200 9036
rect 15252 9024 15258 9036
rect 15381 9027 15439 9033
rect 15381 9024 15393 9027
rect 15252 8996 15393 9024
rect 15252 8984 15258 8996
rect 15381 8993 15393 8996
rect 15427 8993 15439 9027
rect 15381 8987 15439 8993
rect 14921 8959 14979 8965
rect 14921 8925 14933 8959
rect 14967 8925 14979 8959
rect 14921 8919 14979 8925
rect 14366 8888 14372 8900
rect 14279 8860 14372 8888
rect 13909 8851 13967 8857
rect 14366 8848 14372 8860
rect 14424 8888 14430 8900
rect 15197 8891 15255 8897
rect 15197 8888 15209 8891
rect 14424 8860 15209 8888
rect 14424 8848 14430 8860
rect 15197 8857 15209 8860
rect 15243 8857 15255 8891
rect 15197 8851 15255 8857
rect 7984 8792 8340 8820
rect 7984 8780 7990 8792
rect 8846 8780 8852 8832
rect 8904 8820 8910 8832
rect 9490 8820 9496 8832
rect 8904 8792 9496 8820
rect 8904 8780 8910 8792
rect 9490 8780 9496 8792
rect 9548 8820 9554 8832
rect 12526 8820 12532 8832
rect 9548 8792 12532 8820
rect 9548 8780 9554 8792
rect 12526 8780 12532 8792
rect 12584 8820 12590 8832
rect 13354 8820 13360 8832
rect 12584 8792 13360 8820
rect 12584 8780 12590 8792
rect 13354 8780 13360 8792
rect 13412 8780 13418 8832
rect 14090 8820 14096 8832
rect 14051 8792 14096 8820
rect 14090 8780 14096 8792
rect 14148 8780 14154 8832
rect 1104 8730 16008 8752
rect 1104 8678 3480 8730
rect 3532 8678 3544 8730
rect 3596 8678 3608 8730
rect 3660 8678 3672 8730
rect 3724 8678 8478 8730
rect 8530 8678 8542 8730
rect 8594 8678 8606 8730
rect 8658 8678 8670 8730
rect 8722 8678 13475 8730
rect 13527 8678 13539 8730
rect 13591 8678 13603 8730
rect 13655 8678 13667 8730
rect 13719 8678 16008 8730
rect 1104 8656 16008 8678
rect 1854 8576 1860 8628
rect 1912 8616 1918 8628
rect 2222 8616 2228 8628
rect 1912 8588 2228 8616
rect 1912 8576 1918 8588
rect 2222 8576 2228 8588
rect 2280 8616 2286 8628
rect 9861 8619 9919 8625
rect 9861 8616 9873 8619
rect 2280 8588 3464 8616
rect 2280 8576 2286 8588
rect 2593 8551 2651 8557
rect 2593 8548 2605 8551
rect 2240 8520 2605 8548
rect 2240 8489 2268 8520
rect 2593 8517 2605 8520
rect 2639 8517 2651 8551
rect 3326 8548 3332 8560
rect 2593 8511 2651 8517
rect 2746 8520 3332 8548
rect 2225 8483 2283 8489
rect 2225 8449 2237 8483
rect 2271 8449 2283 8483
rect 2225 8443 2283 8449
rect 2409 8483 2467 8489
rect 2409 8449 2421 8483
rect 2455 8480 2467 8483
rect 2746 8480 2774 8520
rect 3326 8508 3332 8520
rect 3384 8508 3390 8560
rect 3234 8480 3240 8492
rect 2455 8452 2774 8480
rect 3195 8452 3240 8480
rect 2455 8449 2467 8452
rect 2409 8443 2467 8449
rect 3234 8440 3240 8452
rect 3292 8440 3298 8492
rect 3436 8489 3464 8588
rect 4816 8588 9873 8616
rect 3421 8483 3479 8489
rect 3421 8449 3433 8483
rect 3467 8449 3479 8483
rect 3421 8443 3479 8449
rect 2130 8412 2136 8424
rect 2091 8384 2136 8412
rect 2130 8372 2136 8384
rect 2188 8372 2194 8424
rect 2314 8372 2320 8424
rect 2372 8412 2378 8424
rect 3688 8415 3746 8421
rect 3688 8412 3700 8415
rect 2372 8384 3700 8412
rect 2372 8372 2378 8384
rect 3688 8381 3700 8384
rect 3734 8412 3746 8415
rect 4816 8412 4844 8588
rect 9861 8585 9873 8588
rect 9907 8585 9919 8619
rect 10502 8616 10508 8628
rect 9861 8579 9919 8585
rect 10336 8588 10508 8616
rect 6273 8551 6331 8557
rect 6273 8517 6285 8551
rect 6319 8548 6331 8551
rect 6319 8520 6408 8548
rect 6319 8517 6331 8520
rect 6273 8511 6331 8517
rect 3734 8384 4844 8412
rect 3734 8381 3746 8384
rect 3688 8375 3746 8381
rect 4890 8372 4896 8424
rect 4948 8412 4954 8424
rect 6380 8412 6408 8520
rect 6546 8508 6552 8560
rect 6604 8548 6610 8560
rect 8386 8548 8392 8560
rect 6604 8520 8392 8548
rect 6604 8508 6610 8520
rect 8386 8508 8392 8520
rect 8444 8508 8450 8560
rect 10336 8548 10364 8588
rect 10502 8576 10508 8588
rect 10560 8576 10566 8628
rect 10594 8576 10600 8628
rect 10652 8616 10658 8628
rect 10652 8588 11284 8616
rect 10652 8576 10658 8588
rect 9784 8520 10364 8548
rect 9784 8492 9812 8520
rect 11256 8492 11284 8588
rect 11330 8576 11336 8628
rect 11388 8616 11394 8628
rect 11517 8619 11575 8625
rect 11517 8616 11529 8619
rect 11388 8588 11529 8616
rect 11388 8576 11394 8588
rect 11517 8585 11529 8588
rect 11563 8585 11575 8619
rect 11517 8579 11575 8585
rect 11701 8619 11759 8625
rect 11701 8585 11713 8619
rect 11747 8616 11759 8619
rect 12158 8616 12164 8628
rect 11747 8588 12164 8616
rect 11747 8585 11759 8588
rect 11701 8579 11759 8585
rect 12158 8576 12164 8588
rect 12216 8576 12222 8628
rect 12342 8576 12348 8628
rect 12400 8616 12406 8628
rect 13906 8616 13912 8628
rect 12400 8588 13912 8616
rect 12400 8576 12406 8588
rect 13906 8576 13912 8588
rect 13964 8576 13970 8628
rect 14826 8576 14832 8628
rect 14884 8616 14890 8628
rect 14921 8619 14979 8625
rect 14921 8616 14933 8619
rect 14884 8588 14933 8616
rect 14884 8576 14890 8588
rect 14921 8585 14933 8588
rect 14967 8585 14979 8619
rect 14921 8579 14979 8585
rect 12526 8548 12532 8560
rect 12487 8520 12532 8548
rect 12526 8508 12532 8520
rect 12584 8508 12590 8560
rect 13354 8548 13360 8560
rect 13315 8520 13360 8548
rect 13354 8508 13360 8520
rect 13412 8508 13418 8560
rect 13538 8508 13544 8560
rect 13596 8548 13602 8560
rect 15013 8551 15071 8557
rect 15013 8548 15025 8551
rect 13596 8520 15025 8548
rect 13596 8508 13602 8520
rect 15013 8517 15025 8520
rect 15059 8517 15071 8551
rect 15013 8511 15071 8517
rect 6457 8483 6515 8489
rect 6457 8449 6469 8483
rect 6503 8480 6515 8483
rect 8754 8480 8760 8492
rect 6503 8452 8760 8480
rect 6503 8449 6515 8452
rect 6457 8443 6515 8449
rect 8754 8440 8760 8452
rect 8812 8440 8818 8492
rect 9766 8480 9772 8492
rect 9727 8452 9772 8480
rect 9766 8440 9772 8452
rect 9824 8440 9830 8492
rect 11238 8480 11244 8492
rect 11199 8452 11244 8480
rect 11238 8440 11244 8452
rect 11296 8440 11302 8492
rect 12253 8483 12311 8489
rect 12253 8480 12265 8483
rect 11348 8452 12265 8480
rect 9674 8412 9680 8424
rect 4948 8384 4993 8412
rect 5092 8384 9680 8412
rect 4948 8372 4954 8384
rect 1394 8344 1400 8356
rect 1355 8316 1400 8344
rect 1394 8304 1400 8316
rect 1452 8304 1458 8356
rect 1581 8347 1639 8353
rect 1581 8313 1593 8347
rect 1627 8344 1639 8347
rect 3510 8344 3516 8356
rect 1627 8316 3516 8344
rect 1627 8313 1639 8316
rect 1581 8307 1639 8313
rect 3510 8304 3516 8316
rect 3568 8304 3574 8356
rect 5092 8344 5120 8384
rect 9674 8372 9680 8384
rect 9732 8372 9738 8424
rect 11348 8412 11376 8452
rect 12253 8449 12265 8452
rect 12299 8480 12311 8483
rect 12434 8480 12440 8492
rect 12299 8452 12440 8480
rect 12299 8449 12311 8452
rect 12253 8443 12311 8449
rect 12434 8440 12440 8452
rect 12492 8440 12498 8492
rect 12894 8480 12900 8492
rect 12544 8452 12900 8480
rect 12544 8424 12572 8452
rect 12894 8440 12900 8452
rect 12952 8480 12958 8492
rect 13081 8483 13139 8489
rect 13081 8480 13093 8483
rect 12952 8452 13093 8480
rect 12952 8440 12958 8452
rect 13081 8449 13093 8452
rect 13127 8480 13139 8483
rect 13630 8480 13636 8492
rect 13127 8452 13636 8480
rect 13127 8449 13139 8452
rect 13081 8443 13139 8449
rect 13630 8440 13636 8452
rect 13688 8440 13694 8492
rect 13814 8440 13820 8492
rect 13872 8480 13878 8492
rect 13909 8483 13967 8489
rect 13909 8480 13921 8483
rect 13872 8452 13921 8480
rect 13872 8440 13878 8452
rect 13909 8449 13921 8452
rect 13955 8449 13967 8483
rect 14274 8480 14280 8492
rect 14235 8452 14280 8480
rect 13909 8443 13967 8449
rect 14274 8440 14280 8452
rect 14332 8440 14338 8492
rect 15194 8480 15200 8492
rect 15155 8452 15200 8480
rect 15194 8440 15200 8452
rect 15252 8440 15258 8492
rect 11974 8412 11980 8424
rect 10428 8384 11376 8412
rect 11440 8384 11980 8412
rect 10428 8356 10456 8384
rect 5166 8353 5172 8356
rect 3620 8316 5120 8344
rect 1765 8279 1823 8285
rect 1765 8245 1777 8279
rect 1811 8276 1823 8279
rect 2038 8276 2044 8288
rect 1811 8248 2044 8276
rect 1811 8245 1823 8248
rect 1765 8239 1823 8245
rect 2038 8236 2044 8248
rect 2096 8236 2102 8288
rect 2958 8276 2964 8288
rect 2919 8248 2964 8276
rect 2958 8236 2964 8248
rect 3016 8236 3022 8288
rect 3050 8236 3056 8288
rect 3108 8276 3114 8288
rect 3108 8248 3153 8276
rect 3108 8236 3114 8248
rect 3326 8236 3332 8288
rect 3384 8276 3390 8288
rect 3620 8276 3648 8316
rect 5160 8307 5172 8353
rect 5224 8344 5230 8356
rect 5224 8316 5260 8344
rect 5166 8304 5172 8307
rect 5224 8304 5230 8316
rect 5442 8304 5448 8356
rect 5500 8344 5506 8356
rect 6549 8347 6607 8353
rect 6549 8344 6561 8347
rect 5500 8316 6561 8344
rect 5500 8304 5506 8316
rect 6549 8313 6561 8316
rect 6595 8313 6607 8347
rect 6549 8307 6607 8313
rect 8297 8347 8355 8353
rect 8297 8313 8309 8347
rect 8343 8344 8355 8347
rect 9306 8344 9312 8356
rect 8343 8316 9312 8344
rect 8343 8313 8355 8316
rect 8297 8307 8355 8313
rect 9306 8304 9312 8316
rect 9364 8304 9370 8356
rect 9524 8347 9582 8353
rect 9524 8313 9536 8347
rect 9570 8344 9582 8347
rect 10410 8344 10416 8356
rect 9570 8316 10416 8344
rect 9570 8313 9582 8316
rect 9524 8307 9582 8313
rect 10410 8304 10416 8316
rect 10468 8304 10474 8356
rect 10870 8304 10876 8356
rect 10928 8344 10934 8356
rect 10974 8347 11032 8353
rect 10974 8344 10986 8347
rect 10928 8316 10986 8344
rect 10928 8304 10934 8316
rect 10974 8313 10986 8316
rect 11020 8313 11032 8347
rect 10974 8307 11032 8313
rect 11146 8304 11152 8356
rect 11204 8344 11210 8356
rect 11440 8344 11468 8384
rect 11974 8372 11980 8384
rect 12032 8412 12038 8424
rect 12069 8415 12127 8421
rect 12069 8412 12081 8415
rect 12032 8384 12081 8412
rect 12032 8372 12038 8384
rect 12069 8381 12081 8384
rect 12115 8381 12127 8415
rect 12069 8375 12127 8381
rect 12158 8372 12164 8424
rect 12216 8412 12222 8424
rect 12216 8384 12296 8412
rect 12216 8372 12222 8384
rect 11204 8316 11468 8344
rect 11517 8347 11575 8353
rect 11204 8304 11210 8316
rect 11517 8313 11529 8347
rect 11563 8344 11575 8347
rect 11698 8344 11704 8356
rect 11563 8316 11704 8344
rect 11563 8313 11575 8316
rect 11517 8307 11575 8313
rect 11698 8304 11704 8316
rect 11756 8344 11762 8356
rect 12268 8344 12296 8384
rect 12526 8372 12532 8424
rect 12584 8372 12590 8424
rect 12618 8372 12624 8424
rect 12676 8412 12682 8424
rect 12989 8415 13047 8421
rect 12989 8412 13001 8415
rect 12676 8384 13001 8412
rect 12676 8372 12682 8384
rect 12989 8381 13001 8384
rect 13035 8412 13047 8415
rect 13538 8412 13544 8424
rect 13035 8384 13544 8412
rect 13035 8381 13047 8384
rect 12989 8375 13047 8381
rect 13538 8372 13544 8384
rect 13596 8372 13602 8424
rect 13725 8415 13783 8421
rect 13725 8381 13737 8415
rect 13771 8412 13783 8415
rect 13998 8412 14004 8424
rect 13771 8384 14004 8412
rect 13771 8381 13783 8384
rect 13725 8375 13783 8381
rect 13998 8372 14004 8384
rect 14056 8372 14062 8424
rect 12897 8347 12955 8353
rect 12897 8344 12909 8347
rect 11756 8316 12204 8344
rect 12268 8316 12909 8344
rect 11756 8304 11762 8316
rect 3384 8248 3648 8276
rect 3384 8236 3390 8248
rect 3694 8236 3700 8288
rect 3752 8276 3758 8288
rect 4522 8276 4528 8288
rect 3752 8248 4528 8276
rect 3752 8236 3758 8248
rect 4522 8236 4528 8248
rect 4580 8236 4586 8288
rect 4801 8279 4859 8285
rect 4801 8245 4813 8279
rect 4847 8276 4859 8279
rect 6457 8279 6515 8285
rect 6457 8276 6469 8279
rect 4847 8248 6469 8276
rect 4847 8245 4859 8248
rect 4801 8239 4859 8245
rect 6457 8245 6469 8248
rect 6503 8245 6515 8279
rect 6457 8239 6515 8245
rect 6638 8236 6644 8288
rect 6696 8276 6702 8288
rect 8110 8276 8116 8288
rect 6696 8248 8116 8276
rect 6696 8236 6702 8248
rect 8110 8236 8116 8248
rect 8168 8236 8174 8288
rect 8662 8236 8668 8288
rect 8720 8276 8726 8288
rect 11974 8276 11980 8288
rect 8720 8248 11980 8276
rect 8720 8236 8726 8248
rect 11974 8236 11980 8248
rect 12032 8236 12038 8288
rect 12176 8285 12204 8316
rect 12897 8313 12909 8316
rect 12943 8313 12955 8347
rect 12897 8307 12955 8313
rect 13446 8304 13452 8356
rect 13504 8344 13510 8356
rect 13817 8347 13875 8353
rect 13817 8344 13829 8347
rect 13504 8316 13829 8344
rect 13504 8304 13510 8316
rect 13817 8313 13829 8316
rect 13863 8344 13875 8347
rect 14090 8344 14096 8356
rect 13863 8316 14096 8344
rect 13863 8313 13875 8316
rect 13817 8307 13875 8313
rect 14090 8304 14096 8316
rect 14148 8304 14154 8356
rect 14274 8304 14280 8356
rect 14332 8344 14338 8356
rect 14553 8347 14611 8353
rect 14553 8344 14565 8347
rect 14332 8316 14565 8344
rect 14332 8304 14338 8316
rect 14553 8313 14565 8316
rect 14599 8313 14611 8347
rect 14553 8307 14611 8313
rect 12161 8279 12219 8285
rect 12161 8245 12173 8279
rect 12207 8245 12219 8279
rect 12161 8239 12219 8245
rect 12342 8236 12348 8288
rect 12400 8276 12406 8288
rect 13262 8276 13268 8288
rect 12400 8248 13268 8276
rect 12400 8236 12406 8248
rect 13262 8236 13268 8248
rect 13320 8276 13326 8288
rect 13722 8276 13728 8288
rect 13320 8248 13728 8276
rect 13320 8236 13326 8248
rect 13722 8236 13728 8248
rect 13780 8236 13786 8288
rect 14461 8279 14519 8285
rect 14461 8245 14473 8279
rect 14507 8276 14519 8279
rect 14826 8276 14832 8288
rect 14507 8248 14832 8276
rect 14507 8245 14519 8248
rect 14461 8239 14519 8245
rect 14826 8236 14832 8248
rect 14884 8236 14890 8288
rect 1104 8186 16008 8208
rect 1104 8134 5979 8186
rect 6031 8134 6043 8186
rect 6095 8134 6107 8186
rect 6159 8134 6171 8186
rect 6223 8134 10976 8186
rect 11028 8134 11040 8186
rect 11092 8134 11104 8186
rect 11156 8134 11168 8186
rect 11220 8134 16008 8186
rect 1104 8112 16008 8134
rect 1486 8072 1492 8084
rect 1447 8044 1492 8072
rect 1486 8032 1492 8044
rect 1544 8032 1550 8084
rect 1854 8032 1860 8084
rect 1912 8072 1918 8084
rect 2682 8072 2688 8084
rect 1912 8044 2688 8072
rect 1912 8032 1918 8044
rect 2682 8032 2688 8044
rect 2740 8032 2746 8084
rect 2869 8075 2927 8081
rect 2869 8041 2881 8075
rect 2915 8072 2927 8075
rect 3050 8072 3056 8084
rect 2915 8044 3056 8072
rect 2915 8041 2927 8044
rect 2869 8035 2927 8041
rect 3050 8032 3056 8044
rect 3108 8032 3114 8084
rect 3234 8072 3240 8084
rect 3195 8044 3240 8072
rect 3234 8032 3240 8044
rect 3292 8032 3298 8084
rect 3510 8032 3516 8084
rect 3568 8072 3574 8084
rect 3881 8075 3939 8081
rect 3881 8072 3893 8075
rect 3568 8044 3893 8072
rect 3568 8032 3574 8044
rect 3881 8041 3893 8044
rect 3927 8041 3939 8075
rect 5074 8072 5080 8084
rect 3881 8035 3939 8041
rect 4172 8044 5080 8072
rect 1578 7964 1584 8016
rect 1636 8004 1642 8016
rect 1765 8007 1823 8013
rect 1765 8004 1777 8007
rect 1636 7976 1777 8004
rect 1636 7964 1642 7976
rect 1765 7973 1777 7976
rect 1811 8004 1823 8007
rect 1811 7976 2544 8004
rect 1811 7973 1823 7976
rect 1765 7967 1823 7973
rect 2038 7936 2044 7948
rect 1999 7908 2044 7936
rect 2038 7896 2044 7908
rect 2096 7896 2102 7948
rect 2406 7936 2412 7948
rect 2367 7908 2412 7936
rect 2406 7896 2412 7908
rect 2464 7896 2470 7948
rect 2516 7945 2544 7976
rect 2774 7964 2780 8016
rect 2832 8004 2838 8016
rect 2832 7976 3832 8004
rect 2832 7964 2838 7976
rect 2501 7939 2559 7945
rect 2501 7905 2513 7939
rect 2547 7936 2559 7939
rect 2958 7936 2964 7948
rect 2547 7908 2964 7936
rect 2547 7905 2559 7908
rect 2501 7899 2559 7905
rect 2958 7896 2964 7908
rect 3016 7896 3022 7948
rect 3329 7939 3387 7945
rect 3329 7905 3341 7939
rect 3375 7936 3387 7939
rect 3602 7936 3608 7948
rect 3375 7908 3608 7936
rect 3375 7905 3387 7908
rect 3329 7899 3387 7905
rect 3602 7896 3608 7908
rect 3660 7896 3666 7948
rect 3804 7936 3832 7976
rect 3970 7964 3976 8016
rect 4028 8004 4034 8016
rect 4172 8013 4200 8044
rect 5074 8032 5080 8044
rect 5132 8032 5138 8084
rect 5166 8032 5172 8084
rect 5224 8072 5230 8084
rect 7561 8075 7619 8081
rect 7561 8072 7573 8075
rect 5224 8044 7573 8072
rect 5224 8032 5230 8044
rect 7561 8041 7573 8044
rect 7607 8041 7619 8075
rect 7561 8035 7619 8041
rect 8294 8032 8300 8084
rect 8352 8072 8358 8084
rect 8846 8072 8852 8084
rect 8352 8044 8852 8072
rect 8352 8032 8358 8044
rect 8846 8032 8852 8044
rect 8904 8032 8910 8084
rect 9398 8072 9404 8084
rect 8956 8044 9404 8072
rect 4157 8007 4215 8013
rect 4157 8004 4169 8007
rect 4028 7976 4169 8004
rect 4028 7964 4034 7976
rect 4157 7973 4169 7976
rect 4203 7973 4215 8007
rect 6914 8004 6920 8016
rect 4157 7967 4215 7973
rect 4264 7976 6920 8004
rect 4065 7939 4123 7945
rect 4065 7936 4077 7939
rect 3804 7908 4077 7936
rect 4065 7905 4077 7908
rect 4111 7905 4123 7939
rect 4065 7899 4123 7905
rect 2317 7871 2375 7877
rect 2317 7837 2329 7871
rect 2363 7837 2375 7871
rect 2317 7831 2375 7837
rect 2332 7800 2360 7831
rect 2682 7828 2688 7880
rect 2740 7868 2746 7880
rect 3050 7868 3056 7880
rect 2740 7840 3056 7868
rect 2740 7828 2746 7840
rect 3050 7828 3056 7840
rect 3108 7828 3114 7880
rect 4264 7868 4292 7976
rect 6914 7964 6920 7976
rect 6972 8004 6978 8016
rect 6972 7976 7972 8004
rect 6972 7964 6978 7976
rect 4341 7939 4399 7945
rect 4341 7905 4353 7939
rect 4387 7905 4399 7939
rect 4873 7939 4931 7945
rect 4873 7936 4885 7939
rect 4341 7899 4399 7905
rect 4540 7908 4885 7936
rect 3528 7840 4292 7868
rect 3528 7800 3556 7840
rect 4356 7812 4384 7899
rect 4540 7880 4568 7908
rect 4873 7905 4885 7908
rect 4919 7905 4931 7939
rect 4873 7899 4931 7905
rect 5718 7896 5724 7948
rect 5776 7936 5782 7948
rect 7202 7939 7260 7945
rect 7202 7936 7214 7939
rect 5776 7908 7214 7936
rect 5776 7896 5782 7908
rect 7202 7905 7214 7908
rect 7248 7936 7260 7939
rect 7834 7936 7840 7948
rect 7248 7908 7840 7936
rect 7248 7905 7260 7908
rect 7202 7899 7260 7905
rect 7834 7896 7840 7908
rect 7892 7896 7898 7948
rect 7944 7936 7972 7976
rect 8386 7964 8392 8016
rect 8444 8004 8450 8016
rect 8444 7976 8892 8004
rect 8444 7964 8450 7976
rect 8662 7936 8668 7948
rect 8720 7945 8726 7948
rect 7944 7908 8668 7936
rect 8662 7896 8668 7908
rect 8720 7899 8732 7945
rect 8720 7896 8726 7899
rect 4522 7828 4528 7880
rect 4580 7828 4586 7880
rect 4617 7871 4675 7877
rect 4617 7837 4629 7871
rect 4663 7837 4675 7871
rect 4617 7831 4675 7837
rect 2332 7772 3556 7800
rect 3602 7760 3608 7812
rect 3660 7800 3666 7812
rect 3660 7772 4108 7800
rect 3660 7760 3666 7772
rect 4080 7744 4108 7772
rect 4338 7760 4344 7812
rect 4396 7760 4402 7812
rect 1762 7692 1768 7744
rect 1820 7732 1826 7744
rect 1857 7735 1915 7741
rect 1857 7732 1869 7735
rect 1820 7704 1869 7732
rect 1820 7692 1826 7704
rect 1857 7701 1869 7704
rect 1903 7701 1915 7735
rect 1857 7695 1915 7701
rect 3697 7735 3755 7741
rect 3697 7701 3709 7735
rect 3743 7732 3755 7735
rect 3878 7732 3884 7744
rect 3743 7704 3884 7732
rect 3743 7701 3755 7704
rect 3697 7695 3755 7701
rect 3878 7692 3884 7704
rect 3936 7692 3942 7744
rect 4062 7692 4068 7744
rect 4120 7692 4126 7744
rect 4525 7735 4583 7741
rect 4525 7701 4537 7735
rect 4571 7732 4583 7735
rect 4632 7732 4660 7831
rect 5810 7828 5816 7880
rect 5868 7868 5874 7880
rect 7469 7871 7527 7877
rect 5868 7840 6224 7868
rect 5868 7828 5874 7840
rect 5626 7760 5632 7812
rect 5684 7800 5690 7812
rect 6196 7800 6224 7840
rect 7469 7837 7481 7871
rect 7515 7868 7527 7871
rect 7926 7868 7932 7880
rect 7515 7840 7932 7868
rect 7515 7837 7527 7840
rect 7469 7831 7527 7837
rect 7926 7828 7932 7840
rect 7984 7828 7990 7880
rect 8864 7868 8892 7976
rect 8956 7945 8984 8044
rect 9398 8032 9404 8044
rect 9456 8072 9462 8084
rect 10594 8072 10600 8084
rect 9456 8044 10600 8072
rect 9456 8032 9462 8044
rect 10594 8032 10600 8044
rect 10652 8032 10658 8084
rect 11790 8072 11796 8084
rect 10796 8044 11100 8072
rect 11751 8044 11796 8072
rect 9030 7964 9036 8016
rect 9088 8004 9094 8016
rect 10796 8004 10824 8044
rect 10962 8004 10968 8016
rect 9088 7976 10824 8004
rect 10923 7976 10968 8004
rect 9088 7964 9094 7976
rect 10962 7964 10968 7976
rect 11020 7964 11026 8016
rect 11072 8004 11100 8044
rect 11790 8032 11796 8044
rect 11848 8032 11854 8084
rect 11885 8075 11943 8081
rect 11885 8041 11897 8075
rect 11931 8072 11943 8075
rect 12250 8072 12256 8084
rect 11931 8044 12256 8072
rect 11931 8041 11943 8044
rect 11885 8035 11943 8041
rect 12250 8032 12256 8044
rect 12308 8032 12314 8084
rect 12342 8032 12348 8084
rect 12400 8072 12406 8084
rect 15105 8075 15163 8081
rect 15105 8072 15117 8075
rect 12400 8044 15117 8072
rect 12400 8032 12406 8044
rect 15105 8041 15117 8044
rect 15151 8041 15163 8075
rect 15105 8035 15163 8041
rect 13449 8007 13507 8013
rect 13449 8004 13461 8007
rect 11072 7976 13461 8004
rect 13449 7973 13461 7976
rect 13495 7973 13507 8007
rect 13449 7967 13507 7973
rect 13722 7964 13728 8016
rect 13780 8004 13786 8016
rect 14553 8007 14611 8013
rect 14553 8004 14565 8007
rect 13780 7976 14565 8004
rect 13780 7964 13786 7976
rect 14553 7973 14565 7976
rect 14599 8004 14611 8007
rect 15010 8004 15016 8016
rect 14599 7976 15016 8004
rect 14599 7973 14611 7976
rect 14553 7967 14611 7973
rect 15010 7964 15016 7976
rect 15068 7964 15074 8016
rect 8941 7939 8999 7945
rect 8941 7905 8953 7939
rect 8987 7905 8999 7939
rect 10238 7939 10296 7945
rect 10238 7936 10250 7939
rect 8941 7899 8999 7905
rect 9048 7908 10250 7936
rect 9048 7868 9076 7908
rect 10238 7905 10250 7908
rect 10284 7936 10296 7939
rect 12526 7936 12532 7948
rect 10284 7908 12532 7936
rect 10284 7905 10296 7908
rect 10238 7899 10296 7905
rect 12526 7896 12532 7908
rect 12584 7896 12590 7948
rect 12621 7939 12679 7945
rect 12621 7905 12633 7939
rect 12667 7936 12679 7939
rect 13078 7936 13084 7948
rect 12667 7908 13084 7936
rect 12667 7905 12679 7908
rect 12621 7899 12679 7905
rect 10502 7868 10508 7880
rect 8864 7840 9076 7868
rect 10463 7840 10508 7868
rect 10502 7828 10508 7840
rect 10560 7828 10566 7880
rect 10778 7828 10784 7880
rect 10836 7868 10842 7880
rect 11057 7871 11115 7877
rect 11057 7868 11069 7871
rect 10836 7840 11069 7868
rect 10836 7828 10842 7840
rect 11057 7837 11069 7840
rect 11103 7837 11115 7871
rect 11057 7831 11115 7837
rect 10870 7800 10876 7812
rect 5684 7772 6132 7800
rect 6196 7772 6592 7800
rect 5684 7760 5690 7772
rect 4890 7732 4896 7744
rect 4571 7704 4896 7732
rect 4571 7701 4583 7704
rect 4525 7695 4583 7701
rect 4890 7692 4896 7704
rect 4948 7692 4954 7744
rect 5994 7732 6000 7744
rect 5955 7704 6000 7732
rect 5994 7692 6000 7704
rect 6052 7692 6058 7744
rect 6104 7741 6132 7772
rect 6089 7735 6147 7741
rect 6089 7701 6101 7735
rect 6135 7732 6147 7735
rect 6454 7732 6460 7744
rect 6135 7704 6460 7732
rect 6135 7701 6147 7704
rect 6089 7695 6147 7701
rect 6454 7692 6460 7704
rect 6512 7692 6518 7744
rect 6564 7732 6592 7772
rect 10520 7772 10876 7800
rect 6822 7732 6828 7744
rect 6564 7704 6828 7732
rect 6822 7692 6828 7704
rect 6880 7692 6886 7744
rect 7190 7692 7196 7744
rect 7248 7732 7254 7744
rect 9125 7735 9183 7741
rect 9125 7732 9137 7735
rect 7248 7704 9137 7732
rect 7248 7692 7254 7704
rect 9125 7701 9137 7704
rect 9171 7732 9183 7735
rect 10520 7732 10548 7772
rect 10870 7760 10876 7772
rect 10928 7760 10934 7812
rect 11072 7800 11100 7831
rect 11146 7828 11152 7880
rect 11204 7868 11210 7880
rect 11974 7868 11980 7880
rect 11204 7840 11249 7868
rect 11935 7840 11980 7868
rect 11204 7828 11210 7840
rect 11974 7828 11980 7840
rect 12032 7828 12038 7880
rect 12434 7828 12440 7880
rect 12492 7868 12498 7880
rect 12636 7868 12664 7899
rect 13078 7896 13084 7908
rect 13136 7896 13142 7948
rect 13170 7896 13176 7948
rect 13228 7936 13234 7948
rect 13541 7939 13599 7945
rect 13541 7936 13553 7939
rect 13228 7908 13553 7936
rect 13228 7896 13234 7908
rect 13541 7905 13553 7908
rect 13587 7936 13599 7939
rect 13814 7936 13820 7948
rect 13587 7908 13820 7936
rect 13587 7905 13599 7908
rect 13541 7899 13599 7905
rect 13814 7896 13820 7908
rect 13872 7896 13878 7948
rect 14182 7896 14188 7948
rect 14240 7936 14246 7948
rect 14369 7939 14427 7945
rect 14369 7936 14381 7939
rect 14240 7908 14381 7936
rect 14240 7896 14246 7908
rect 14369 7905 14381 7908
rect 14415 7905 14427 7939
rect 14369 7899 14427 7905
rect 12492 7840 12664 7868
rect 12713 7871 12771 7877
rect 12492 7828 12498 7840
rect 12713 7837 12725 7871
rect 12759 7837 12771 7871
rect 12894 7868 12900 7880
rect 12855 7840 12900 7868
rect 12713 7831 12771 7837
rect 12250 7800 12256 7812
rect 11072 7772 11560 7800
rect 12211 7772 12256 7800
rect 9171 7704 10548 7732
rect 9171 7701 9183 7704
rect 9125 7695 9183 7701
rect 10594 7692 10600 7744
rect 10652 7732 10658 7744
rect 10652 7704 10697 7732
rect 10652 7692 10658 7704
rect 10778 7692 10784 7744
rect 10836 7732 10842 7744
rect 11238 7732 11244 7744
rect 10836 7704 11244 7732
rect 10836 7692 10842 7704
rect 11238 7692 11244 7704
rect 11296 7692 11302 7744
rect 11422 7732 11428 7744
rect 11383 7704 11428 7732
rect 11422 7692 11428 7704
rect 11480 7692 11486 7744
rect 11532 7732 11560 7772
rect 12250 7760 12256 7772
rect 12308 7760 12314 7812
rect 12728 7800 12756 7831
rect 12894 7828 12900 7840
rect 12952 7828 12958 7880
rect 13630 7868 13636 7880
rect 13591 7840 13636 7868
rect 13630 7828 13636 7840
rect 13688 7828 13694 7880
rect 14090 7800 14096 7812
rect 12728 7772 14096 7800
rect 14090 7760 14096 7772
rect 14148 7800 14154 7812
rect 14200 7800 14228 7896
rect 14148 7772 14228 7800
rect 14148 7760 14154 7772
rect 12342 7732 12348 7744
rect 11532 7704 12348 7732
rect 12342 7692 12348 7704
rect 12400 7692 12406 7744
rect 12526 7692 12532 7744
rect 12584 7732 12590 7744
rect 12986 7732 12992 7744
rect 12584 7704 12992 7732
rect 12584 7692 12590 7704
rect 12986 7692 12992 7704
rect 13044 7692 13050 7744
rect 13078 7692 13084 7744
rect 13136 7732 13142 7744
rect 14001 7735 14059 7741
rect 13136 7704 13181 7732
rect 13136 7692 13142 7704
rect 14001 7701 14013 7735
rect 14047 7732 14059 7735
rect 14182 7732 14188 7744
rect 14047 7704 14188 7732
rect 14047 7701 14059 7704
rect 14001 7695 14059 7701
rect 14182 7692 14188 7704
rect 14240 7692 14246 7744
rect 14734 7732 14740 7744
rect 14695 7704 14740 7732
rect 14734 7692 14740 7704
rect 14792 7692 14798 7744
rect 14918 7732 14924 7744
rect 14879 7704 14924 7732
rect 14918 7692 14924 7704
rect 14976 7692 14982 7744
rect 1104 7642 16008 7664
rect 1104 7590 3480 7642
rect 3532 7590 3544 7642
rect 3596 7590 3608 7642
rect 3660 7590 3672 7642
rect 3724 7590 8478 7642
rect 8530 7590 8542 7642
rect 8594 7590 8606 7642
rect 8658 7590 8670 7642
rect 8722 7590 13475 7642
rect 13527 7590 13539 7642
rect 13591 7590 13603 7642
rect 13655 7590 13667 7642
rect 13719 7590 16008 7642
rect 1104 7568 16008 7590
rect 3234 7488 3240 7540
rect 3292 7528 3298 7540
rect 3329 7531 3387 7537
rect 3329 7528 3341 7531
rect 3292 7500 3341 7528
rect 3292 7488 3298 7500
rect 3329 7497 3341 7500
rect 3375 7497 3387 7531
rect 10594 7528 10600 7540
rect 3329 7491 3387 7497
rect 3436 7500 10600 7528
rect 2501 7463 2559 7469
rect 2501 7429 2513 7463
rect 2547 7460 2559 7463
rect 3142 7460 3148 7472
rect 2547 7432 3148 7460
rect 2547 7429 2559 7432
rect 2501 7423 2559 7429
rect 3142 7420 3148 7432
rect 3200 7420 3206 7472
rect 1394 7392 1400 7404
rect 1355 7364 1400 7392
rect 1394 7352 1400 7364
rect 1452 7352 1458 7404
rect 1949 7395 2007 7401
rect 1949 7361 1961 7395
rect 1995 7392 2007 7395
rect 2682 7392 2688 7404
rect 1995 7364 2688 7392
rect 1995 7361 2007 7364
rect 1949 7355 2007 7361
rect 2682 7352 2688 7364
rect 2740 7352 2746 7404
rect 2777 7395 2835 7401
rect 2777 7361 2789 7395
rect 2823 7392 2835 7395
rect 2958 7392 2964 7404
rect 2823 7364 2964 7392
rect 2823 7361 2835 7364
rect 2777 7355 2835 7361
rect 2958 7352 2964 7364
rect 3016 7352 3022 7404
rect 3436 7392 3464 7500
rect 10594 7488 10600 7500
rect 10652 7488 10658 7540
rect 10870 7488 10876 7540
rect 10928 7528 10934 7540
rect 11425 7531 11483 7537
rect 11425 7528 11437 7531
rect 10928 7500 11437 7528
rect 10928 7488 10934 7500
rect 6273 7463 6331 7469
rect 6273 7460 6285 7463
rect 3344 7364 3464 7392
rect 5920 7432 6285 7460
rect 1581 7327 1639 7333
rect 1581 7293 1593 7327
rect 1627 7324 1639 7327
rect 1762 7324 1768 7336
rect 1627 7296 1768 7324
rect 1627 7293 1639 7296
rect 1581 7287 1639 7293
rect 1762 7284 1768 7296
rect 1820 7284 1826 7336
rect 2041 7327 2099 7333
rect 2041 7293 2053 7327
rect 2087 7324 2099 7327
rect 3344 7324 3372 7364
rect 2087 7296 3372 7324
rect 3421 7327 3479 7333
rect 2087 7293 2099 7296
rect 2041 7287 2099 7293
rect 3421 7293 3433 7327
rect 3467 7324 3479 7327
rect 4890 7324 4896 7336
rect 3467 7296 4896 7324
rect 3467 7293 3479 7296
rect 3421 7287 3479 7293
rect 4890 7284 4896 7296
rect 4948 7284 4954 7336
rect 5000 7296 5304 7324
rect 1670 7216 1676 7268
rect 1728 7256 1734 7268
rect 1728 7228 3004 7256
rect 1728 7216 1734 7228
rect 2130 7188 2136 7200
rect 2091 7160 2136 7188
rect 2130 7148 2136 7160
rect 2188 7148 2194 7200
rect 2866 7188 2872 7200
rect 2827 7160 2872 7188
rect 2866 7148 2872 7160
rect 2924 7148 2930 7200
rect 2976 7197 3004 7228
rect 3050 7216 3056 7268
rect 3108 7256 3114 7268
rect 3688 7259 3746 7265
rect 3688 7256 3700 7259
rect 3108 7228 3700 7256
rect 3108 7216 3114 7228
rect 3688 7225 3700 7228
rect 3734 7256 3746 7259
rect 5000 7256 5028 7296
rect 3734 7228 5028 7256
rect 5160 7259 5218 7265
rect 3734 7225 3746 7228
rect 3688 7219 3746 7225
rect 5160 7225 5172 7259
rect 5206 7225 5218 7259
rect 5276 7256 5304 7296
rect 5442 7284 5448 7336
rect 5500 7324 5506 7336
rect 5920 7324 5948 7432
rect 6273 7429 6285 7432
rect 6319 7460 6331 7463
rect 6362 7460 6368 7472
rect 6319 7432 6368 7460
rect 6319 7429 6331 7432
rect 6273 7423 6331 7429
rect 6362 7420 6368 7432
rect 6420 7420 6426 7472
rect 10410 7420 10416 7472
rect 10468 7460 10474 7472
rect 10781 7463 10839 7469
rect 10781 7460 10793 7463
rect 10468 7432 10793 7460
rect 10468 7420 10474 7432
rect 10781 7429 10793 7432
rect 10827 7429 10839 7463
rect 10781 7423 10839 7429
rect 11057 7463 11115 7469
rect 11057 7429 11069 7463
rect 11103 7429 11115 7463
rect 11057 7423 11115 7429
rect 9398 7392 9404 7404
rect 9359 7364 9404 7392
rect 9398 7352 9404 7364
rect 9456 7352 9462 7404
rect 10502 7352 10508 7404
rect 10560 7392 10566 7404
rect 10962 7392 10968 7404
rect 10560 7364 10968 7392
rect 10560 7352 10566 7364
rect 10962 7352 10968 7364
rect 11020 7352 11026 7404
rect 5500 7296 5948 7324
rect 5500 7284 5506 7296
rect 5994 7284 6000 7336
rect 6052 7324 6058 7336
rect 7837 7327 7895 7333
rect 6052 7296 7696 7324
rect 6052 7284 6058 7296
rect 7558 7256 7564 7268
rect 7616 7265 7622 7268
rect 5276 7228 7420 7256
rect 7528 7228 7564 7256
rect 5160 7219 5218 7225
rect 2961 7191 3019 7197
rect 2961 7157 2973 7191
rect 3007 7188 3019 7191
rect 4154 7188 4160 7200
rect 3007 7160 4160 7188
rect 3007 7157 3019 7160
rect 2961 7151 3019 7157
rect 4154 7148 4160 7160
rect 4212 7148 4218 7200
rect 4801 7191 4859 7197
rect 4801 7157 4813 7191
rect 4847 7188 4859 7191
rect 4982 7188 4988 7200
rect 4847 7160 4988 7188
rect 4847 7157 4859 7160
rect 4801 7151 4859 7157
rect 4982 7148 4988 7160
rect 5040 7148 5046 7200
rect 5074 7148 5080 7200
rect 5132 7188 5138 7200
rect 5175 7188 5203 7219
rect 5626 7188 5632 7200
rect 5132 7160 5632 7188
rect 5132 7148 5138 7160
rect 5626 7148 5632 7160
rect 5684 7148 5690 7200
rect 5810 7148 5816 7200
rect 5868 7188 5874 7200
rect 6457 7191 6515 7197
rect 6457 7188 6469 7191
rect 5868 7160 6469 7188
rect 5868 7148 5874 7160
rect 6457 7157 6469 7160
rect 6503 7157 6515 7191
rect 7392 7188 7420 7228
rect 7558 7216 7564 7228
rect 7616 7219 7628 7265
rect 7668 7256 7696 7296
rect 7837 7293 7849 7327
rect 7883 7324 7895 7327
rect 7926 7324 7932 7336
rect 7883 7296 7932 7324
rect 7883 7293 7895 7296
rect 7837 7287 7895 7293
rect 7926 7284 7932 7296
rect 7984 7324 7990 7336
rect 9416 7324 9444 7352
rect 10778 7324 10784 7336
rect 7984 7296 9444 7324
rect 9600 7296 10784 7324
rect 7984 7284 7990 7296
rect 8196 7259 8254 7265
rect 8196 7256 8208 7259
rect 7668 7228 8208 7256
rect 8196 7225 8208 7228
rect 8242 7256 8254 7259
rect 9600 7256 9628 7296
rect 10778 7284 10784 7296
rect 10836 7284 10842 7336
rect 10870 7284 10876 7336
rect 10928 7324 10934 7336
rect 11072 7324 11100 7423
rect 11164 7392 11192 7500
rect 11425 7497 11437 7500
rect 11471 7528 11483 7531
rect 12526 7528 12532 7540
rect 11471 7500 12532 7528
rect 11471 7497 11483 7500
rect 11425 7491 11483 7497
rect 12526 7488 12532 7500
rect 12584 7488 12590 7540
rect 12710 7488 12716 7540
rect 12768 7528 12774 7540
rect 13357 7531 13415 7537
rect 13357 7528 13369 7531
rect 12768 7500 13369 7528
rect 12768 7488 12774 7500
rect 13357 7497 13369 7500
rect 13403 7497 13415 7531
rect 13357 7491 13415 7497
rect 13998 7488 14004 7540
rect 14056 7528 14062 7540
rect 14274 7528 14280 7540
rect 14056 7500 14280 7528
rect 14056 7488 14062 7500
rect 14274 7488 14280 7500
rect 14332 7528 14338 7540
rect 14734 7528 14740 7540
rect 14332 7500 14740 7528
rect 14332 7488 14338 7500
rect 14734 7488 14740 7500
rect 14792 7488 14798 7540
rect 11238 7420 11244 7472
rect 11296 7460 11302 7472
rect 12986 7460 12992 7472
rect 11296 7432 12992 7460
rect 11296 7420 11302 7432
rect 12986 7420 12992 7432
rect 13044 7420 13050 7472
rect 12161 7395 12219 7401
rect 12161 7392 12173 7395
rect 11164 7364 12173 7392
rect 12161 7361 12173 7364
rect 12207 7361 12219 7395
rect 12161 7355 12219 7361
rect 12253 7395 12311 7401
rect 12253 7361 12265 7395
rect 12299 7361 12311 7395
rect 13078 7392 13084 7404
rect 13039 7364 13084 7392
rect 12253 7355 12311 7361
rect 11149 7327 11207 7333
rect 11149 7324 11161 7327
rect 10928 7296 10973 7324
rect 11072 7296 11161 7324
rect 10928 7284 10934 7296
rect 11149 7293 11161 7296
rect 11195 7324 11207 7327
rect 11330 7324 11336 7336
rect 11195 7296 11336 7324
rect 11195 7293 11207 7296
rect 11149 7287 11207 7293
rect 11330 7284 11336 7296
rect 11388 7284 11394 7336
rect 11974 7284 11980 7336
rect 12032 7324 12038 7336
rect 12268 7324 12296 7355
rect 13078 7352 13084 7364
rect 13136 7352 13142 7404
rect 13909 7395 13967 7401
rect 13909 7392 13921 7395
rect 13188 7364 13921 7392
rect 12032 7296 12296 7324
rect 12032 7284 12038 7296
rect 12894 7284 12900 7336
rect 12952 7324 12958 7336
rect 13188 7324 13216 7364
rect 13909 7361 13921 7364
rect 13955 7361 13967 7395
rect 13909 7355 13967 7361
rect 12952 7296 13216 7324
rect 13725 7327 13783 7333
rect 12952 7284 12958 7296
rect 13725 7293 13737 7327
rect 13771 7324 13783 7327
rect 13998 7324 14004 7336
rect 13771 7296 14004 7324
rect 13771 7293 13783 7296
rect 13725 7287 13783 7293
rect 13998 7284 14004 7296
rect 14056 7324 14062 7336
rect 14553 7327 14611 7333
rect 14553 7324 14565 7327
rect 14056 7296 14565 7324
rect 14056 7284 14062 7296
rect 14553 7293 14565 7296
rect 14599 7324 14611 7327
rect 14642 7324 14648 7336
rect 14599 7296 14648 7324
rect 14599 7293 14611 7296
rect 14553 7287 14611 7293
rect 14642 7284 14648 7296
rect 14700 7284 14706 7336
rect 9674 7265 9680 7268
rect 8242 7228 9628 7256
rect 8242 7225 8254 7228
rect 8196 7219 8254 7225
rect 9668 7219 9680 7265
rect 9732 7256 9738 7268
rect 9732 7228 9768 7256
rect 7616 7216 7622 7219
rect 9674 7216 9680 7219
rect 9732 7216 9738 7228
rect 10042 7216 10048 7268
rect 10100 7256 10106 7268
rect 12618 7256 12624 7268
rect 10100 7228 12624 7256
rect 10100 7216 10106 7228
rect 12618 7216 12624 7228
rect 12676 7216 12682 7268
rect 14458 7256 14464 7268
rect 13004 7228 14464 7256
rect 13004 7200 13032 7228
rect 14458 7216 14464 7228
rect 14516 7216 14522 7268
rect 9214 7188 9220 7200
rect 7392 7160 9220 7188
rect 6457 7151 6515 7157
rect 9214 7148 9220 7160
rect 9272 7148 9278 7200
rect 9306 7148 9312 7200
rect 9364 7188 9370 7200
rect 10318 7188 10324 7200
rect 9364 7160 10324 7188
rect 9364 7148 9370 7160
rect 10318 7148 10324 7160
rect 10376 7148 10382 7200
rect 11333 7191 11391 7197
rect 11333 7157 11345 7191
rect 11379 7188 11391 7191
rect 11422 7188 11428 7200
rect 11379 7160 11428 7188
rect 11379 7157 11391 7160
rect 11333 7151 11391 7157
rect 11422 7148 11428 7160
rect 11480 7148 11486 7200
rect 11698 7188 11704 7200
rect 11659 7160 11704 7188
rect 11698 7148 11704 7160
rect 11756 7148 11762 7200
rect 12069 7191 12127 7197
rect 12069 7157 12081 7191
rect 12115 7188 12127 7191
rect 12158 7188 12164 7200
rect 12115 7160 12164 7188
rect 12115 7157 12127 7160
rect 12069 7151 12127 7157
rect 12158 7148 12164 7160
rect 12216 7148 12222 7200
rect 12342 7148 12348 7200
rect 12400 7188 12406 7200
rect 12529 7191 12587 7197
rect 12529 7188 12541 7191
rect 12400 7160 12541 7188
rect 12400 7148 12406 7160
rect 12529 7157 12541 7160
rect 12575 7157 12587 7191
rect 12894 7188 12900 7200
rect 12855 7160 12900 7188
rect 12529 7151 12587 7157
rect 12894 7148 12900 7160
rect 12952 7148 12958 7200
rect 12986 7148 12992 7200
rect 13044 7188 13050 7200
rect 13814 7188 13820 7200
rect 13044 7160 13089 7188
rect 13775 7160 13820 7188
rect 13044 7148 13050 7160
rect 13814 7148 13820 7160
rect 13872 7188 13878 7200
rect 14185 7191 14243 7197
rect 14185 7188 14197 7191
rect 13872 7160 14197 7188
rect 13872 7148 13878 7160
rect 14185 7157 14197 7160
rect 14231 7157 14243 7191
rect 14366 7188 14372 7200
rect 14327 7160 14372 7188
rect 14185 7151 14243 7157
rect 14366 7148 14372 7160
rect 14424 7148 14430 7200
rect 1104 7098 16008 7120
rect 1104 7046 5979 7098
rect 6031 7046 6043 7098
rect 6095 7046 6107 7098
rect 6159 7046 6171 7098
rect 6223 7046 10976 7098
rect 11028 7046 11040 7098
rect 11092 7046 11104 7098
rect 11156 7046 11168 7098
rect 11220 7046 16008 7098
rect 1104 7024 16008 7046
rect 1581 6987 1639 6993
rect 1581 6953 1593 6987
rect 1627 6984 1639 6987
rect 1670 6984 1676 6996
rect 1627 6956 1676 6984
rect 1627 6953 1639 6956
rect 1581 6947 1639 6953
rect 1670 6944 1676 6956
rect 1728 6944 1734 6996
rect 2590 6984 2596 6996
rect 2332 6956 2596 6984
rect 1486 6876 1492 6928
rect 1544 6916 1550 6928
rect 2332 6916 2360 6956
rect 2590 6944 2596 6956
rect 2648 6984 2654 6996
rect 2648 6956 2820 6984
rect 2648 6944 2654 6956
rect 2498 6916 2504 6928
rect 1544 6888 2360 6916
rect 2459 6888 2504 6916
rect 1544 6876 1550 6888
rect 2498 6876 2504 6888
rect 2556 6876 2562 6928
rect 2792 6916 2820 6956
rect 2958 6944 2964 6996
rect 3016 6984 3022 6996
rect 3016 6956 4384 6984
rect 3016 6944 3022 6956
rect 3329 6919 3387 6925
rect 3329 6916 3341 6919
rect 2792 6888 3341 6916
rect 3329 6885 3341 6888
rect 3375 6885 3387 6919
rect 3329 6879 3387 6885
rect 1578 6808 1584 6860
rect 1636 6848 1642 6860
rect 1673 6851 1731 6857
rect 1673 6848 1685 6851
rect 1636 6820 1685 6848
rect 1636 6808 1642 6820
rect 1673 6817 1685 6820
rect 1719 6817 1731 6851
rect 1673 6811 1731 6817
rect 2041 6851 2099 6857
rect 2041 6817 2053 6851
rect 2087 6848 2099 6851
rect 2314 6848 2320 6860
rect 2087 6820 2320 6848
rect 2087 6817 2099 6820
rect 2041 6811 2099 6817
rect 2314 6808 2320 6820
rect 2372 6808 2378 6860
rect 4246 6848 4252 6860
rect 4207 6820 4252 6848
rect 4246 6808 4252 6820
rect 4304 6808 4310 6860
rect 2222 6780 2228 6792
rect 2183 6752 2228 6780
rect 2222 6740 2228 6752
rect 2280 6740 2286 6792
rect 2406 6780 2412 6792
rect 2367 6752 2412 6780
rect 2406 6740 2412 6752
rect 2464 6740 2470 6792
rect 3421 6783 3479 6789
rect 3421 6749 3433 6783
rect 3467 6749 3479 6783
rect 3602 6780 3608 6792
rect 3563 6752 3608 6780
rect 3421 6743 3479 6749
rect 2961 6715 3019 6721
rect 2961 6712 2973 6715
rect 2746 6684 2973 6712
rect 1854 6644 1860 6656
rect 1815 6616 1860 6644
rect 1854 6604 1860 6616
rect 1912 6604 1918 6656
rect 2038 6604 2044 6656
rect 2096 6644 2102 6656
rect 2746 6644 2774 6684
rect 2961 6681 2973 6684
rect 3007 6681 3019 6715
rect 2961 6675 3019 6681
rect 2866 6644 2872 6656
rect 2096 6616 2774 6644
rect 2827 6616 2872 6644
rect 2096 6604 2102 6616
rect 2866 6604 2872 6616
rect 2924 6604 2930 6656
rect 3050 6604 3056 6656
rect 3108 6644 3114 6656
rect 3436 6644 3464 6743
rect 3602 6740 3608 6752
rect 3660 6740 3666 6792
rect 4356 6780 4384 6956
rect 4706 6944 4712 6996
rect 4764 6984 4770 6996
rect 8386 6984 8392 6996
rect 4764 6956 4809 6984
rect 4908 6956 8392 6984
rect 4764 6944 4770 6956
rect 4798 6916 4804 6928
rect 4759 6888 4804 6916
rect 4798 6876 4804 6888
rect 4856 6876 4862 6928
rect 4908 6848 4936 6956
rect 8386 6944 8392 6956
rect 8444 6944 8450 6996
rect 8754 6944 8760 6996
rect 8812 6984 8818 6996
rect 11974 6984 11980 6996
rect 8812 6956 11980 6984
rect 8812 6944 8818 6956
rect 11974 6944 11980 6956
rect 12032 6944 12038 6996
rect 12250 6984 12256 6996
rect 12211 6956 12256 6984
rect 12250 6944 12256 6956
rect 12308 6944 12314 6996
rect 12710 6944 12716 6996
rect 12768 6984 12774 6996
rect 13081 6987 13139 6993
rect 13081 6984 13093 6987
rect 12768 6956 13093 6984
rect 12768 6944 12774 6956
rect 13081 6953 13093 6956
rect 13127 6984 13139 6987
rect 13170 6984 13176 6996
rect 13127 6956 13176 6984
rect 13127 6953 13139 6956
rect 13081 6947 13139 6953
rect 13170 6944 13176 6956
rect 13228 6984 13234 6996
rect 13541 6987 13599 6993
rect 13541 6984 13553 6987
rect 13228 6956 13553 6984
rect 13228 6944 13234 6956
rect 13541 6953 13553 6956
rect 13587 6953 13599 6987
rect 13541 6947 13599 6953
rect 13725 6987 13783 6993
rect 13725 6953 13737 6987
rect 13771 6984 13783 6987
rect 14090 6984 14096 6996
rect 13771 6956 14096 6984
rect 13771 6953 13783 6956
rect 13725 6947 13783 6953
rect 14090 6944 14096 6956
rect 14148 6944 14154 6996
rect 5258 6876 5264 6928
rect 5316 6916 5322 6928
rect 6086 6916 6092 6928
rect 5316 6888 6092 6916
rect 5316 6876 5322 6888
rect 6086 6876 6092 6888
rect 6144 6876 6150 6928
rect 6454 6876 6460 6928
rect 6512 6916 6518 6928
rect 7558 6916 7564 6928
rect 6512 6888 7564 6916
rect 6512 6876 6518 6888
rect 7558 6876 7564 6888
rect 7616 6876 7622 6928
rect 7926 6916 7932 6928
rect 7668 6888 7932 6916
rect 4816 6820 4936 6848
rect 4816 6780 4844 6820
rect 5718 6808 5724 6860
rect 5776 6848 5782 6860
rect 6282 6851 6340 6857
rect 6282 6848 6294 6851
rect 5776 6820 6294 6848
rect 5776 6808 5782 6820
rect 6282 6817 6294 6820
rect 6328 6817 6340 6851
rect 6282 6811 6340 6817
rect 6549 6851 6607 6857
rect 6549 6817 6561 6851
rect 6595 6848 6607 6851
rect 7668 6848 7696 6888
rect 7926 6876 7932 6888
rect 7984 6916 7990 6928
rect 7984 6888 8064 6916
rect 7984 6876 7990 6888
rect 6595 6820 7696 6848
rect 6595 6817 6607 6820
rect 6549 6811 6607 6817
rect 7742 6808 7748 6860
rect 7800 6857 7806 6860
rect 8036 6857 8064 6888
rect 8202 6876 8208 6928
rect 8260 6916 8266 6928
rect 8481 6919 8539 6925
rect 8481 6916 8493 6919
rect 8260 6888 8493 6916
rect 8260 6876 8266 6888
rect 8481 6885 8493 6888
rect 8527 6916 8539 6919
rect 8527 6888 8800 6916
rect 8527 6885 8539 6888
rect 8481 6879 8539 6885
rect 7800 6848 7812 6857
rect 8021 6851 8079 6857
rect 7800 6820 7992 6848
rect 7800 6811 7812 6820
rect 7800 6808 7806 6811
rect 4356 6752 4844 6780
rect 4985 6783 5043 6789
rect 4985 6749 4997 6783
rect 5031 6780 5043 6783
rect 5534 6780 5540 6792
rect 5031 6752 5540 6780
rect 5031 6749 5043 6752
rect 4985 6743 5043 6749
rect 5534 6740 5540 6752
rect 5592 6740 5598 6792
rect 7964 6780 7992 6820
rect 8021 6817 8033 6851
rect 8067 6817 8079 6851
rect 8021 6811 8079 6817
rect 8110 6808 8116 6860
rect 8168 6848 8174 6860
rect 8573 6851 8631 6857
rect 8573 6848 8585 6851
rect 8168 6820 8585 6848
rect 8168 6808 8174 6820
rect 8573 6817 8585 6820
rect 8619 6817 8631 6851
rect 8772 6848 8800 6888
rect 8846 6876 8852 6928
rect 8904 6916 8910 6928
rect 9306 6916 9312 6928
rect 8904 6888 9312 6916
rect 8904 6876 8910 6888
rect 9306 6876 9312 6888
rect 9364 6876 9370 6928
rect 10042 6916 10048 6928
rect 9600 6888 10048 6916
rect 9600 6848 9628 6888
rect 10042 6876 10048 6888
rect 10100 6916 10106 6928
rect 11425 6919 11483 6925
rect 11425 6916 11437 6919
rect 10100 6888 11437 6916
rect 10100 6876 10106 6888
rect 11425 6885 11437 6888
rect 11471 6885 11483 6919
rect 11425 6879 11483 6885
rect 11517 6919 11575 6925
rect 11517 6885 11529 6919
rect 11563 6916 11575 6919
rect 11606 6916 11612 6928
rect 11563 6888 11612 6916
rect 11563 6885 11575 6888
rect 11517 6879 11575 6885
rect 11606 6876 11612 6888
rect 11664 6876 11670 6928
rect 11790 6876 11796 6928
rect 11848 6916 11854 6928
rect 12342 6916 12348 6928
rect 11848 6888 12204 6916
rect 12303 6888 12348 6916
rect 11848 6876 11854 6888
rect 8772 6820 9628 6848
rect 8573 6811 8631 6817
rect 9858 6808 9864 6860
rect 9916 6848 9922 6860
rect 9953 6851 10011 6857
rect 9953 6848 9965 6851
rect 9916 6820 9965 6848
rect 9916 6808 9922 6820
rect 9953 6817 9965 6820
rect 9999 6848 10011 6851
rect 10410 6848 10416 6860
rect 9999 6820 10416 6848
rect 9999 6817 10011 6820
rect 9953 6811 10011 6817
rect 10410 6808 10416 6820
rect 10468 6808 10474 6860
rect 10502 6808 10508 6860
rect 10560 6848 10566 6860
rect 10597 6851 10655 6857
rect 10597 6848 10609 6851
rect 10560 6820 10609 6848
rect 10560 6808 10566 6820
rect 10597 6817 10609 6820
rect 10643 6817 10655 6851
rect 10597 6811 10655 6817
rect 10689 6851 10747 6857
rect 10689 6817 10701 6851
rect 10735 6848 10747 6851
rect 11146 6848 11152 6860
rect 10735 6820 11152 6848
rect 10735 6817 10747 6820
rect 10689 6811 10747 6817
rect 11146 6808 11152 6820
rect 11204 6808 11210 6860
rect 11624 6848 11652 6876
rect 11974 6848 11980 6860
rect 11624 6820 11980 6848
rect 11974 6808 11980 6820
rect 12032 6808 12038 6860
rect 12176 6848 12204 6888
rect 12342 6876 12348 6888
rect 12400 6916 12406 6928
rect 14369 6919 14427 6925
rect 14369 6916 14381 6919
rect 12400 6888 14381 6916
rect 12400 6876 12406 6888
rect 14369 6885 14381 6888
rect 14415 6916 14427 6919
rect 14553 6919 14611 6925
rect 14553 6916 14565 6919
rect 14415 6888 14565 6916
rect 14415 6885 14427 6888
rect 14369 6879 14427 6885
rect 14553 6885 14565 6888
rect 14599 6916 14611 6919
rect 14918 6916 14924 6928
rect 14599 6888 14924 6916
rect 14599 6885 14611 6888
rect 14553 6879 14611 6885
rect 14918 6876 14924 6888
rect 14976 6876 14982 6928
rect 12802 6848 12808 6860
rect 12176 6820 12808 6848
rect 12802 6808 12808 6820
rect 12860 6808 12866 6860
rect 13173 6851 13231 6857
rect 13173 6817 13185 6851
rect 13219 6848 13231 6851
rect 13219 6820 13400 6848
rect 13219 6817 13231 6820
rect 13173 6811 13231 6817
rect 8202 6780 8208 6792
rect 7964 6752 8208 6780
rect 8202 6740 8208 6752
rect 8260 6740 8266 6792
rect 8665 6783 8723 6789
rect 8665 6749 8677 6783
rect 8711 6749 8723 6783
rect 8665 6743 8723 6749
rect 3970 6712 3976 6724
rect 3896 6684 3976 6712
rect 3896 6653 3924 6684
rect 3970 6672 3976 6684
rect 4028 6672 4034 6724
rect 4062 6672 4068 6724
rect 4120 6712 4126 6724
rect 4120 6684 4165 6712
rect 4120 6672 4126 6684
rect 4706 6672 4712 6724
rect 4764 6712 4770 6724
rect 6641 6715 6699 6721
rect 4764 6684 5672 6712
rect 4764 6672 4770 6684
rect 3881 6647 3939 6653
rect 3881 6644 3893 6647
rect 3108 6616 3893 6644
rect 3108 6604 3114 6616
rect 3881 6613 3893 6616
rect 3927 6613 3939 6647
rect 3881 6607 3939 6613
rect 4246 6604 4252 6656
rect 4304 6644 4310 6656
rect 4341 6647 4399 6653
rect 4341 6644 4353 6647
rect 4304 6616 4353 6644
rect 4304 6604 4310 6616
rect 4341 6613 4353 6616
rect 4387 6613 4399 6647
rect 4341 6607 4399 6613
rect 4522 6604 4528 6656
rect 4580 6644 4586 6656
rect 5169 6647 5227 6653
rect 5169 6644 5181 6647
rect 4580 6616 5181 6644
rect 4580 6604 4586 6616
rect 5169 6613 5181 6616
rect 5215 6613 5227 6647
rect 5644 6644 5672 6684
rect 6641 6681 6653 6715
rect 6687 6712 6699 6715
rect 6730 6712 6736 6724
rect 6687 6684 6736 6712
rect 6687 6681 6699 6684
rect 6641 6675 6699 6681
rect 6730 6672 6736 6684
rect 6788 6672 6794 6724
rect 8018 6672 8024 6724
rect 8076 6712 8082 6724
rect 8680 6712 8708 6743
rect 8846 6740 8852 6792
rect 8904 6780 8910 6792
rect 8904 6752 9345 6780
rect 8904 6740 8910 6752
rect 9030 6712 9036 6724
rect 8076 6684 9036 6712
rect 8076 6672 8082 6684
rect 9030 6672 9036 6684
rect 9088 6672 9094 6724
rect 9317 6712 9345 6752
rect 9398 6740 9404 6792
rect 9456 6780 9462 6792
rect 10781 6783 10839 6789
rect 10781 6780 10793 6783
rect 9456 6752 9501 6780
rect 9539 6752 10793 6780
rect 9456 6740 9462 6752
rect 9539 6712 9567 6752
rect 10781 6749 10793 6752
rect 10827 6780 10839 6783
rect 11514 6780 11520 6792
rect 10827 6752 11520 6780
rect 10827 6749 10839 6752
rect 10781 6743 10839 6749
rect 11514 6740 11520 6752
rect 11572 6740 11578 6792
rect 11698 6780 11704 6792
rect 11659 6752 11704 6780
rect 11698 6740 11704 6752
rect 11756 6740 11762 6792
rect 11790 6740 11796 6792
rect 11848 6780 11854 6792
rect 12437 6783 12495 6789
rect 12437 6780 12449 6783
rect 11848 6752 12449 6780
rect 11848 6740 11854 6752
rect 12437 6749 12449 6752
rect 12483 6780 12495 6783
rect 12618 6780 12624 6792
rect 12483 6752 12624 6780
rect 12483 6749 12495 6752
rect 12437 6743 12495 6749
rect 12618 6740 12624 6752
rect 12676 6740 12682 6792
rect 13262 6780 13268 6792
rect 13223 6752 13268 6780
rect 13262 6740 13268 6752
rect 13320 6740 13326 6792
rect 13372 6780 13400 6820
rect 13372 6752 14228 6780
rect 9317 6684 9567 6712
rect 9674 6672 9680 6724
rect 9732 6712 9738 6724
rect 11885 6715 11943 6721
rect 11885 6712 11897 6715
rect 9732 6684 11897 6712
rect 9732 6672 9738 6684
rect 11885 6681 11897 6684
rect 11931 6681 11943 6715
rect 11885 6675 11943 6681
rect 12250 6672 12256 6724
rect 12308 6712 12314 6724
rect 13909 6715 13967 6721
rect 13909 6712 13921 6715
rect 12308 6684 13921 6712
rect 12308 6672 12314 6684
rect 13909 6681 13921 6684
rect 13955 6681 13967 6715
rect 13909 6675 13967 6681
rect 7006 6644 7012 6656
rect 5644 6616 7012 6644
rect 5169 6607 5227 6613
rect 7006 6604 7012 6616
rect 7064 6604 7070 6656
rect 7098 6604 7104 6656
rect 7156 6644 7162 6656
rect 8113 6647 8171 6653
rect 8113 6644 8125 6647
rect 7156 6616 8125 6644
rect 7156 6604 7162 6616
rect 8113 6613 8125 6616
rect 8159 6613 8171 6647
rect 8113 6607 8171 6613
rect 8202 6604 8208 6656
rect 8260 6644 8266 6656
rect 10229 6647 10287 6653
rect 10229 6644 10241 6647
rect 8260 6616 10241 6644
rect 8260 6604 8266 6616
rect 10229 6613 10241 6616
rect 10275 6613 10287 6647
rect 10229 6607 10287 6613
rect 10410 6604 10416 6656
rect 10468 6644 10474 6656
rect 10870 6644 10876 6656
rect 10468 6616 10876 6644
rect 10468 6604 10474 6616
rect 10870 6604 10876 6616
rect 10928 6604 10934 6656
rect 11054 6644 11060 6656
rect 11015 6616 11060 6644
rect 11054 6604 11060 6616
rect 11112 6604 11118 6656
rect 11146 6604 11152 6656
rect 11204 6644 11210 6656
rect 14200 6653 14228 6752
rect 12713 6647 12771 6653
rect 12713 6644 12725 6647
rect 11204 6616 12725 6644
rect 11204 6604 11210 6616
rect 12713 6613 12725 6616
rect 12759 6613 12771 6647
rect 12713 6607 12771 6613
rect 14185 6647 14243 6653
rect 14185 6613 14197 6647
rect 14231 6644 14243 6647
rect 14274 6644 14280 6656
rect 14231 6616 14280 6644
rect 14231 6613 14243 6616
rect 14185 6607 14243 6613
rect 14274 6604 14280 6616
rect 14332 6604 14338 6656
rect 14734 6644 14740 6656
rect 14695 6616 14740 6644
rect 14734 6604 14740 6616
rect 14792 6604 14798 6656
rect 1104 6554 16008 6576
rect 1104 6502 3480 6554
rect 3532 6502 3544 6554
rect 3596 6502 3608 6554
rect 3660 6502 3672 6554
rect 3724 6502 8478 6554
rect 8530 6502 8542 6554
rect 8594 6502 8606 6554
rect 8658 6502 8670 6554
rect 8722 6502 13475 6554
rect 13527 6502 13539 6554
rect 13591 6502 13603 6554
rect 13655 6502 13667 6554
rect 13719 6502 16008 6554
rect 1104 6480 16008 6502
rect 1486 6440 1492 6452
rect 1447 6412 1492 6440
rect 1486 6400 1492 6412
rect 1544 6400 1550 6452
rect 2406 6400 2412 6452
rect 2464 6440 2470 6452
rect 2501 6443 2559 6449
rect 2501 6440 2513 6443
rect 2464 6412 2513 6440
rect 2464 6400 2470 6412
rect 2501 6409 2513 6412
rect 2547 6409 2559 6443
rect 2501 6403 2559 6409
rect 3421 6443 3479 6449
rect 3421 6409 3433 6443
rect 3467 6440 3479 6443
rect 3786 6440 3792 6452
rect 3467 6412 3792 6440
rect 3467 6409 3479 6412
rect 3421 6403 3479 6409
rect 3786 6400 3792 6412
rect 3844 6440 3850 6452
rect 4430 6440 4436 6452
rect 3844 6412 4436 6440
rect 3844 6400 3850 6412
rect 4430 6400 4436 6412
rect 4488 6400 4494 6452
rect 4893 6443 4951 6449
rect 4893 6409 4905 6443
rect 4939 6440 4951 6443
rect 5258 6440 5264 6452
rect 4939 6412 5264 6440
rect 4939 6409 4951 6412
rect 4893 6403 4951 6409
rect 5258 6400 5264 6412
rect 5316 6400 5322 6452
rect 5534 6400 5540 6452
rect 5592 6440 5598 6452
rect 7837 6443 7895 6449
rect 7837 6440 7849 6443
rect 5592 6412 7849 6440
rect 5592 6400 5598 6412
rect 7837 6409 7849 6412
rect 7883 6440 7895 6443
rect 8018 6440 8024 6452
rect 7883 6412 8024 6440
rect 7883 6409 7895 6412
rect 7837 6403 7895 6409
rect 8018 6400 8024 6412
rect 8076 6400 8082 6452
rect 8294 6400 8300 6452
rect 8352 6440 8358 6452
rect 10042 6440 10048 6452
rect 8352 6412 10048 6440
rect 8352 6400 8358 6412
rect 10042 6400 10048 6412
rect 10100 6400 10106 6452
rect 10410 6400 10416 6452
rect 10468 6440 10474 6452
rect 11790 6440 11796 6452
rect 10468 6412 11796 6440
rect 10468 6400 10474 6412
rect 11790 6400 11796 6412
rect 11848 6400 11854 6452
rect 12986 6440 12992 6452
rect 12268 6412 12992 6440
rect 2222 6332 2228 6384
rect 2280 6372 2286 6384
rect 3602 6372 3608 6384
rect 2280 6344 3608 6372
rect 2280 6332 2286 6344
rect 3602 6332 3608 6344
rect 3660 6332 3666 6384
rect 5074 6332 5080 6384
rect 5132 6332 5138 6384
rect 9398 6332 9404 6384
rect 9456 6372 9462 6384
rect 9456 6344 9501 6372
rect 9456 6332 9462 6344
rect 10778 6332 10784 6384
rect 10836 6332 10842 6384
rect 10870 6332 10876 6384
rect 10928 6372 10934 6384
rect 11882 6372 11888 6384
rect 10928 6344 11888 6372
rect 10928 6332 10934 6344
rect 11882 6332 11888 6344
rect 11940 6332 11946 6384
rect 1949 6307 2007 6313
rect 1949 6273 1961 6307
rect 1995 6273 2007 6307
rect 1949 6267 2007 6273
rect 1581 6239 1639 6245
rect 1581 6205 1593 6239
rect 1627 6236 1639 6239
rect 1854 6236 1860 6248
rect 1627 6208 1860 6236
rect 1627 6205 1639 6208
rect 1581 6199 1639 6205
rect 1854 6196 1860 6208
rect 1912 6196 1918 6248
rect 1964 6236 1992 6267
rect 2038 6264 2044 6316
rect 2096 6304 2102 6316
rect 2096 6276 2141 6304
rect 2096 6264 2102 6276
rect 2314 6264 2320 6316
rect 2372 6304 2378 6316
rect 2682 6304 2688 6316
rect 2372 6276 2688 6304
rect 2372 6264 2378 6276
rect 2682 6264 2688 6276
rect 2740 6264 2746 6316
rect 3237 6307 3295 6313
rect 3237 6273 3249 6307
rect 3283 6304 3295 6307
rect 3326 6304 3332 6316
rect 3283 6276 3332 6304
rect 3283 6273 3295 6276
rect 3237 6267 3295 6273
rect 3326 6264 3332 6276
rect 3384 6264 3390 6316
rect 5092 6304 5120 6332
rect 10796 6304 10824 6332
rect 11146 6304 11152 6316
rect 4724 6276 5120 6304
rect 6196 6276 6601 6304
rect 10796 6276 11152 6304
rect 4724 6236 4752 6276
rect 1964 6208 4752 6236
rect 4801 6239 4859 6245
rect 4801 6205 4813 6239
rect 4847 6236 4859 6239
rect 4890 6236 4896 6248
rect 4847 6208 4896 6236
rect 4847 6205 4859 6208
rect 4801 6199 4859 6205
rect 4890 6196 4896 6208
rect 4948 6236 4954 6248
rect 5074 6236 5080 6248
rect 4948 6208 5080 6236
rect 4948 6196 4954 6208
rect 5074 6196 5080 6208
rect 5132 6196 5138 6248
rect 6196 6236 6224 6276
rect 5828 6208 6224 6236
rect 6273 6239 6331 6245
rect 5828 6180 5856 6208
rect 6273 6205 6285 6239
rect 6319 6236 6331 6239
rect 6454 6236 6460 6248
rect 6319 6208 6460 6236
rect 6319 6205 6331 6208
rect 6273 6199 6331 6205
rect 6454 6196 6460 6208
rect 6512 6196 6518 6248
rect 6573 6236 6601 6276
rect 11146 6264 11152 6276
rect 11204 6264 11210 6316
rect 11333 6307 11391 6313
rect 11333 6273 11345 6307
rect 11379 6304 11391 6307
rect 12268 6304 12296 6412
rect 12986 6400 12992 6412
rect 13044 6400 13050 6452
rect 12618 6332 12624 6384
rect 12676 6372 12682 6384
rect 12676 6344 13952 6372
rect 12676 6332 12682 6344
rect 11379 6276 12296 6304
rect 12345 6307 12403 6313
rect 11379 6273 11391 6276
rect 11333 6267 11391 6273
rect 12345 6273 12357 6307
rect 12391 6304 12403 6307
rect 12710 6304 12716 6316
rect 12391 6276 12716 6304
rect 12391 6273 12403 6276
rect 12345 6267 12403 6273
rect 12710 6264 12716 6276
rect 12768 6264 12774 6316
rect 13078 6304 13084 6316
rect 13039 6276 13084 6304
rect 13078 6264 13084 6276
rect 13136 6264 13142 6316
rect 13924 6313 13952 6344
rect 13909 6307 13967 6313
rect 13909 6273 13921 6307
rect 13955 6273 13967 6307
rect 14366 6304 14372 6316
rect 14327 6276 14372 6304
rect 13909 6267 13967 6273
rect 14366 6264 14372 6276
rect 14424 6264 14430 6316
rect 8754 6236 8760 6248
rect 6573 6208 8760 6236
rect 8754 6196 8760 6208
rect 8812 6196 8818 6248
rect 9214 6196 9220 6248
rect 9272 6236 9278 6248
rect 9309 6239 9367 6245
rect 9309 6236 9321 6239
rect 9272 6208 9321 6236
rect 9272 6196 9278 6208
rect 9309 6205 9321 6208
rect 9355 6236 9367 6239
rect 10781 6239 10839 6245
rect 10781 6236 10793 6239
rect 9355 6208 10793 6236
rect 9355 6205 9367 6208
rect 9309 6199 9367 6205
rect 10781 6205 10793 6208
rect 10827 6236 10839 6239
rect 11057 6239 11115 6245
rect 10827 6208 10916 6236
rect 10827 6205 10839 6208
rect 10781 6199 10839 6205
rect 4556 6171 4614 6177
rect 4556 6168 4568 6171
rect 3620 6140 4568 6168
rect 3620 6112 3648 6140
rect 4556 6137 4568 6140
rect 4602 6168 4614 6171
rect 5442 6168 5448 6180
rect 4602 6140 5448 6168
rect 4602 6137 4614 6140
rect 4556 6131 4614 6137
rect 5442 6128 5448 6140
rect 5500 6128 5506 6180
rect 5810 6128 5816 6180
rect 5868 6128 5874 6180
rect 6028 6171 6086 6177
rect 6028 6137 6040 6171
rect 6074 6168 6086 6171
rect 6362 6168 6368 6180
rect 6074 6140 6368 6168
rect 6074 6137 6086 6140
rect 6028 6131 6086 6137
rect 6362 6128 6368 6140
rect 6420 6128 6426 6180
rect 6546 6128 6552 6180
rect 6604 6168 6610 6180
rect 6702 6171 6760 6177
rect 6702 6168 6714 6171
rect 6604 6140 6714 6168
rect 6604 6128 6610 6140
rect 6702 6137 6714 6140
rect 6748 6137 6760 6171
rect 6702 6131 6760 6137
rect 7006 6128 7012 6180
rect 7064 6168 7070 6180
rect 8294 6168 8300 6180
rect 7064 6140 8300 6168
rect 7064 6128 7070 6140
rect 8294 6128 8300 6140
rect 8352 6128 8358 6180
rect 8846 6128 8852 6180
rect 8904 6168 8910 6180
rect 9042 6171 9100 6177
rect 9042 6168 9054 6171
rect 8904 6140 9054 6168
rect 8904 6128 8910 6140
rect 9042 6137 9054 6140
rect 9088 6137 9100 6171
rect 9042 6131 9100 6137
rect 9674 6128 9680 6180
rect 9732 6168 9738 6180
rect 10226 6168 10232 6180
rect 9732 6140 10232 6168
rect 9732 6128 9738 6140
rect 10226 6128 10232 6140
rect 10284 6128 10290 6180
rect 10318 6128 10324 6180
rect 10376 6168 10382 6180
rect 10514 6171 10572 6177
rect 10514 6168 10526 6171
rect 10376 6140 10526 6168
rect 10376 6128 10382 6140
rect 10514 6137 10526 6140
rect 10560 6137 10572 6171
rect 10514 6131 10572 6137
rect 10888 6112 10916 6208
rect 11057 6205 11069 6239
rect 11103 6236 11115 6239
rect 12618 6236 12624 6248
rect 11103 6208 12624 6236
rect 11103 6205 11115 6208
rect 11057 6199 11115 6205
rect 12618 6196 12624 6208
rect 12676 6196 12682 6248
rect 12986 6196 12992 6248
rect 13044 6236 13050 6248
rect 13725 6239 13783 6245
rect 13725 6236 13737 6239
rect 13044 6208 13737 6236
rect 13044 6196 13050 6208
rect 13725 6205 13737 6208
rect 13771 6205 13783 6239
rect 13725 6199 13783 6205
rect 10962 6128 10968 6180
rect 11020 6168 11026 6180
rect 11422 6168 11428 6180
rect 11020 6140 11428 6168
rect 11020 6128 11026 6140
rect 11422 6128 11428 6140
rect 11480 6128 11486 6180
rect 11974 6128 11980 6180
rect 12032 6168 12038 6180
rect 12161 6171 12219 6177
rect 12161 6168 12173 6171
rect 12032 6140 12173 6168
rect 12032 6128 12038 6140
rect 12161 6137 12173 6140
rect 12207 6137 12219 6171
rect 12161 6131 12219 6137
rect 12897 6171 12955 6177
rect 12897 6137 12909 6171
rect 12943 6168 12955 6171
rect 13538 6168 13544 6180
rect 12943 6140 13544 6168
rect 12943 6137 12955 6140
rect 12897 6131 12955 6137
rect 13538 6128 13544 6140
rect 13596 6128 13602 6180
rect 13630 6128 13636 6180
rect 13688 6168 13694 6180
rect 14185 6171 14243 6177
rect 14185 6168 14197 6171
rect 13688 6140 14197 6168
rect 13688 6128 13694 6140
rect 14185 6137 14197 6140
rect 14231 6137 14243 6171
rect 14185 6131 14243 6137
rect 2133 6103 2191 6109
rect 2133 6069 2145 6103
rect 2179 6100 2191 6103
rect 2314 6100 2320 6112
rect 2179 6072 2320 6100
rect 2179 6069 2191 6072
rect 2133 6063 2191 6069
rect 2314 6060 2320 6072
rect 2372 6060 2378 6112
rect 2590 6100 2596 6112
rect 2551 6072 2596 6100
rect 2590 6060 2596 6072
rect 2648 6060 2654 6112
rect 2958 6100 2964 6112
rect 2919 6072 2964 6100
rect 2958 6060 2964 6072
rect 3016 6060 3022 6112
rect 3050 6060 3056 6112
rect 3108 6100 3114 6112
rect 3108 6072 3153 6100
rect 3108 6060 3114 6072
rect 3602 6060 3608 6112
rect 3660 6060 3666 6112
rect 3694 6060 3700 6112
rect 3752 6100 3758 6112
rect 5718 6100 5724 6112
rect 3752 6072 5724 6100
rect 3752 6060 3758 6072
rect 5718 6060 5724 6072
rect 5776 6100 5782 6112
rect 7466 6100 7472 6112
rect 5776 6072 7472 6100
rect 5776 6060 5782 6072
rect 7466 6060 7472 6072
rect 7524 6060 7530 6112
rect 7558 6060 7564 6112
rect 7616 6100 7622 6112
rect 7929 6103 7987 6109
rect 7929 6100 7941 6103
rect 7616 6072 7941 6100
rect 7616 6060 7622 6072
rect 7929 6069 7941 6072
rect 7975 6069 7987 6103
rect 7929 6063 7987 6069
rect 8018 6060 8024 6112
rect 8076 6100 8082 6112
rect 10686 6100 10692 6112
rect 8076 6072 10692 6100
rect 8076 6060 8082 6072
rect 10686 6060 10692 6072
rect 10744 6060 10750 6112
rect 10870 6060 10876 6112
rect 10928 6060 10934 6112
rect 11698 6100 11704 6112
rect 11659 6072 11704 6100
rect 11698 6060 11704 6072
rect 11756 6060 11762 6112
rect 12069 6103 12127 6109
rect 12069 6069 12081 6103
rect 12115 6100 12127 6103
rect 12342 6100 12348 6112
rect 12115 6072 12348 6100
rect 12115 6069 12127 6072
rect 12069 6063 12127 6069
rect 12342 6060 12348 6072
rect 12400 6060 12406 6112
rect 12434 6060 12440 6112
rect 12492 6100 12498 6112
rect 12529 6103 12587 6109
rect 12529 6100 12541 6103
rect 12492 6072 12541 6100
rect 12492 6060 12498 6072
rect 12529 6069 12541 6072
rect 12575 6069 12587 6103
rect 12529 6063 12587 6069
rect 12802 6060 12808 6112
rect 12860 6100 12866 6112
rect 12989 6103 13047 6109
rect 12989 6100 13001 6103
rect 12860 6072 13001 6100
rect 12860 6060 12866 6072
rect 12989 6069 13001 6072
rect 13035 6069 13047 6103
rect 13354 6100 13360 6112
rect 13315 6072 13360 6100
rect 12989 6063 13047 6069
rect 13354 6060 13360 6072
rect 13412 6060 13418 6112
rect 13814 6100 13820 6112
rect 13775 6072 13820 6100
rect 13814 6060 13820 6072
rect 13872 6060 13878 6112
rect 1104 6010 16008 6032
rect 1104 5958 5979 6010
rect 6031 5958 6043 6010
rect 6095 5958 6107 6010
rect 6159 5958 6171 6010
rect 6223 5958 10976 6010
rect 11028 5958 11040 6010
rect 11092 5958 11104 6010
rect 11156 5958 11168 6010
rect 11220 5958 16008 6010
rect 1104 5936 16008 5958
rect 2869 5899 2927 5905
rect 2869 5865 2881 5899
rect 2915 5896 2927 5899
rect 3050 5896 3056 5908
rect 2915 5868 3056 5896
rect 2915 5865 2927 5868
rect 2869 5859 2927 5865
rect 3050 5856 3056 5868
rect 3108 5856 3114 5908
rect 3237 5899 3295 5905
rect 3237 5865 3249 5899
rect 3283 5896 3295 5899
rect 4065 5899 4123 5905
rect 3283 5868 4016 5896
rect 3283 5865 3295 5868
rect 3237 5859 3295 5865
rect 1489 5831 1547 5837
rect 1489 5797 1501 5831
rect 1535 5828 1547 5831
rect 3510 5828 3516 5840
rect 1535 5800 3516 5828
rect 1535 5797 1547 5800
rect 1489 5791 1547 5797
rect 3510 5788 3516 5800
rect 3568 5788 3574 5840
rect 2041 5763 2099 5769
rect 2041 5729 2053 5763
rect 2087 5729 2099 5763
rect 2041 5723 2099 5729
rect 1670 5556 1676 5568
rect 1631 5528 1676 5556
rect 1670 5516 1676 5528
rect 1728 5516 1734 5568
rect 1854 5556 1860 5568
rect 1815 5528 1860 5556
rect 1854 5516 1860 5528
rect 1912 5516 1918 5568
rect 2056 5556 2084 5723
rect 2222 5720 2228 5772
rect 2280 5760 2286 5772
rect 2501 5763 2559 5769
rect 2501 5760 2513 5763
rect 2280 5732 2513 5760
rect 2280 5720 2286 5732
rect 2501 5729 2513 5732
rect 2547 5729 2559 5763
rect 2501 5723 2559 5729
rect 3329 5763 3387 5769
rect 3329 5729 3341 5763
rect 3375 5760 3387 5763
rect 3694 5760 3700 5772
rect 3375 5732 3700 5760
rect 3375 5729 3387 5732
rect 3329 5723 3387 5729
rect 3694 5720 3700 5732
rect 3752 5720 3758 5772
rect 3878 5760 3884 5772
rect 3839 5732 3884 5760
rect 3878 5720 3884 5732
rect 3936 5720 3942 5772
rect 3988 5760 4016 5868
rect 4065 5865 4077 5899
rect 4111 5896 4123 5899
rect 4430 5896 4436 5908
rect 4111 5868 4436 5896
rect 4111 5865 4123 5868
rect 4065 5859 4123 5865
rect 4430 5856 4436 5868
rect 4488 5896 4494 5908
rect 5169 5899 5227 5905
rect 4488 5868 5120 5896
rect 4488 5856 4494 5868
rect 4706 5788 4712 5840
rect 4764 5828 4770 5840
rect 4801 5831 4859 5837
rect 4801 5828 4813 5831
rect 4764 5800 4813 5828
rect 4764 5788 4770 5800
rect 4801 5797 4813 5800
rect 4847 5797 4859 5831
rect 5092 5828 5120 5868
rect 5169 5865 5181 5899
rect 5215 5896 5227 5899
rect 8386 5896 8392 5908
rect 5215 5868 8392 5896
rect 5215 5865 5227 5868
rect 5169 5859 5227 5865
rect 8386 5856 8392 5868
rect 8444 5856 8450 5908
rect 8478 5856 8484 5908
rect 8536 5896 8542 5908
rect 8665 5899 8723 5905
rect 8665 5896 8677 5899
rect 8536 5868 8677 5896
rect 8536 5856 8542 5868
rect 8665 5865 8677 5868
rect 8711 5865 8723 5899
rect 8665 5859 8723 5865
rect 8754 5856 8760 5908
rect 8812 5896 8818 5908
rect 8812 5868 9413 5896
rect 8812 5856 8818 5868
rect 6454 5828 6460 5840
rect 5092 5800 5212 5828
rect 4801 5791 4859 5797
rect 4062 5760 4068 5772
rect 3988 5732 4068 5760
rect 4062 5720 4068 5732
rect 4120 5720 4126 5772
rect 2317 5695 2375 5701
rect 2317 5661 2329 5695
rect 2363 5661 2375 5695
rect 2317 5655 2375 5661
rect 2332 5624 2360 5655
rect 2406 5652 2412 5704
rect 2464 5692 2470 5704
rect 3145 5695 3203 5701
rect 2464 5664 2509 5692
rect 2464 5652 2470 5664
rect 3145 5661 3157 5695
rect 3191 5692 3203 5695
rect 3602 5692 3608 5704
rect 3191 5664 3608 5692
rect 3191 5661 3203 5664
rect 3145 5655 3203 5661
rect 3602 5652 3608 5664
rect 3660 5652 3666 5704
rect 4338 5692 4344 5704
rect 4299 5664 4344 5692
rect 4338 5652 4344 5664
rect 4396 5652 4402 5704
rect 4614 5692 4620 5704
rect 4575 5664 4620 5692
rect 4614 5652 4620 5664
rect 4672 5652 4678 5704
rect 4709 5695 4767 5701
rect 4709 5661 4721 5695
rect 4755 5661 4767 5695
rect 5184 5692 5212 5800
rect 5276 5800 6460 5828
rect 5276 5769 5304 5800
rect 6454 5788 6460 5800
rect 6512 5788 6518 5840
rect 8202 5788 8208 5840
rect 8260 5828 8266 5840
rect 9214 5828 9220 5840
rect 8260 5800 9220 5828
rect 8260 5788 8266 5800
rect 9214 5788 9220 5800
rect 9272 5788 9278 5840
rect 9385 5837 9413 5868
rect 9766 5856 9772 5908
rect 9824 5896 9830 5908
rect 10505 5899 10563 5905
rect 9824 5868 10364 5896
rect 9824 5856 9830 5868
rect 9370 5831 9428 5837
rect 9370 5797 9382 5831
rect 9416 5797 9428 5831
rect 9370 5791 9428 5797
rect 9490 5788 9496 5840
rect 9548 5828 9554 5840
rect 9548 5800 10272 5828
rect 9548 5788 9554 5800
rect 5261 5763 5319 5769
rect 5261 5729 5273 5763
rect 5307 5729 5319 5763
rect 5261 5723 5319 5729
rect 5350 5720 5356 5772
rect 5408 5720 5414 5772
rect 5534 5769 5540 5772
rect 5528 5760 5540 5769
rect 5495 5732 5540 5760
rect 5528 5723 5540 5732
rect 5534 5720 5540 5723
rect 5592 5720 5598 5772
rect 5810 5720 5816 5772
rect 5868 5760 5874 5772
rect 7006 5760 7012 5772
rect 5868 5732 7012 5760
rect 5868 5720 5874 5732
rect 7006 5720 7012 5732
rect 7064 5720 7070 5772
rect 7834 5720 7840 5772
rect 7892 5769 7898 5772
rect 7892 5760 7904 5769
rect 8570 5760 8576 5772
rect 7892 5732 8432 5760
rect 8531 5732 8576 5760
rect 7892 5723 7904 5732
rect 7892 5720 7898 5723
rect 5368 5692 5396 5720
rect 5184 5664 5396 5692
rect 8113 5695 8171 5701
rect 4709 5655 4767 5661
rect 8113 5661 8125 5695
rect 8159 5692 8171 5695
rect 8202 5692 8208 5704
rect 8159 5664 8208 5692
rect 8159 5661 8171 5664
rect 8113 5655 8171 5661
rect 3326 5624 3332 5636
rect 2332 5596 3332 5624
rect 3326 5584 3332 5596
rect 3384 5584 3390 5636
rect 3510 5584 3516 5636
rect 3568 5584 3574 5636
rect 3697 5627 3755 5633
rect 3697 5593 3709 5627
rect 3743 5624 3755 5627
rect 4062 5624 4068 5636
rect 3743 5596 4068 5624
rect 3743 5593 3755 5596
rect 3697 5587 3755 5593
rect 4062 5584 4068 5596
rect 4120 5584 4126 5636
rect 4724 5624 4752 5655
rect 8202 5652 8208 5664
rect 8260 5652 8266 5704
rect 8404 5692 8432 5732
rect 8570 5720 8576 5732
rect 8628 5720 8634 5772
rect 9122 5760 9128 5772
rect 9083 5732 9128 5760
rect 9122 5720 9128 5732
rect 9180 5720 9186 5772
rect 9766 5760 9772 5772
rect 9232 5732 9772 5760
rect 8757 5695 8815 5701
rect 8757 5692 8769 5695
rect 8404 5664 8769 5692
rect 8757 5661 8769 5664
rect 8803 5661 8815 5695
rect 8757 5655 8815 5661
rect 4540 5596 4752 5624
rect 3050 5556 3056 5568
rect 2056 5528 3056 5556
rect 3050 5516 3056 5528
rect 3108 5516 3114 5568
rect 3528 5556 3556 5584
rect 4430 5556 4436 5568
rect 3528 5528 4436 5556
rect 4430 5516 4436 5528
rect 4488 5556 4494 5568
rect 4540 5556 4568 5596
rect 6362 5584 6368 5636
rect 6420 5624 6426 5636
rect 6733 5627 6791 5633
rect 6733 5624 6745 5627
rect 6420 5596 6745 5624
rect 6420 5584 6426 5596
rect 6733 5593 6745 5596
rect 6779 5593 6791 5627
rect 6733 5587 6791 5593
rect 4488 5528 4568 5556
rect 4488 5516 4494 5528
rect 4614 5516 4620 5568
rect 4672 5556 4678 5568
rect 6638 5556 6644 5568
rect 4672 5528 6644 5556
rect 4672 5516 4678 5528
rect 6638 5516 6644 5528
rect 6696 5516 6702 5568
rect 6914 5516 6920 5568
rect 6972 5556 6978 5568
rect 8205 5559 8263 5565
rect 8205 5556 8217 5559
rect 6972 5528 8217 5556
rect 6972 5516 6978 5528
rect 8205 5525 8217 5528
rect 8251 5525 8263 5559
rect 8772 5556 8800 5655
rect 8846 5652 8852 5704
rect 8904 5692 8910 5704
rect 9232 5692 9260 5732
rect 9766 5720 9772 5732
rect 9824 5720 9830 5772
rect 8904 5664 9260 5692
rect 8904 5652 8910 5664
rect 10244 5624 10272 5800
rect 10336 5760 10364 5868
rect 10505 5865 10517 5899
rect 10551 5896 10563 5899
rect 10686 5896 10692 5908
rect 10551 5868 10692 5896
rect 10551 5865 10563 5868
rect 10505 5859 10563 5865
rect 10686 5856 10692 5868
rect 10744 5856 10750 5908
rect 11882 5896 11888 5908
rect 11843 5868 11888 5896
rect 11882 5856 11888 5868
rect 11940 5896 11946 5908
rect 12434 5896 12440 5908
rect 11940 5868 12440 5896
rect 11940 5856 11946 5868
rect 12434 5856 12440 5868
rect 12492 5856 12498 5908
rect 12618 5896 12624 5908
rect 12579 5868 12624 5896
rect 12618 5856 12624 5868
rect 12676 5856 12682 5908
rect 13357 5899 13415 5905
rect 13357 5865 13369 5899
rect 13403 5896 13415 5899
rect 14090 5896 14096 5908
rect 13403 5868 14096 5896
rect 13403 5865 13415 5868
rect 13357 5859 13415 5865
rect 14090 5856 14096 5868
rect 14148 5856 14154 5908
rect 10870 5788 10876 5840
rect 10928 5828 10934 5840
rect 10965 5831 11023 5837
rect 10965 5828 10977 5831
rect 10928 5800 10977 5828
rect 10928 5788 10934 5800
rect 10965 5797 10977 5800
rect 11011 5797 11023 5831
rect 10965 5791 11023 5797
rect 11057 5831 11115 5837
rect 11057 5797 11069 5831
rect 11103 5828 11115 5831
rect 12710 5828 12716 5840
rect 11103 5800 12572 5828
rect 12671 5800 12716 5828
rect 11103 5797 11115 5800
rect 11057 5791 11115 5797
rect 11793 5763 11851 5769
rect 11793 5760 11805 5763
rect 10336 5732 11805 5760
rect 11793 5729 11805 5732
rect 11839 5760 11851 5763
rect 11882 5760 11888 5772
rect 11839 5732 11888 5760
rect 11839 5729 11851 5732
rect 11793 5723 11851 5729
rect 11882 5720 11888 5732
rect 11940 5720 11946 5772
rect 12434 5720 12440 5772
rect 12492 5720 12498 5772
rect 12544 5760 12572 5800
rect 12710 5788 12716 5800
rect 12768 5788 12774 5840
rect 12802 5788 12808 5840
rect 12860 5828 12866 5840
rect 12986 5828 12992 5840
rect 12860 5800 12992 5828
rect 12860 5788 12866 5800
rect 12986 5788 12992 5800
rect 13044 5828 13050 5840
rect 13081 5831 13139 5837
rect 13081 5828 13093 5831
rect 13044 5800 13093 5828
rect 13044 5788 13050 5800
rect 13081 5797 13093 5800
rect 13127 5797 13139 5831
rect 13538 5828 13544 5840
rect 13451 5800 13544 5828
rect 13081 5791 13139 5797
rect 13538 5788 13544 5800
rect 13596 5828 13602 5840
rect 13725 5831 13783 5837
rect 13725 5828 13737 5831
rect 13596 5800 13737 5828
rect 13596 5788 13602 5800
rect 13725 5797 13737 5800
rect 13771 5828 13783 5831
rect 13909 5831 13967 5837
rect 13909 5828 13921 5831
rect 13771 5800 13921 5828
rect 13771 5797 13783 5800
rect 13725 5791 13783 5797
rect 13909 5797 13921 5800
rect 13955 5828 13967 5831
rect 15194 5828 15200 5840
rect 13955 5800 15200 5828
rect 13955 5797 13967 5800
rect 13909 5791 13967 5797
rect 15194 5788 15200 5800
rect 15252 5788 15258 5840
rect 12820 5760 12848 5788
rect 12544 5732 12848 5760
rect 10502 5652 10508 5704
rect 10560 5692 10566 5704
rect 10870 5692 10876 5704
rect 10560 5664 10876 5692
rect 10560 5652 10566 5664
rect 10870 5652 10876 5664
rect 10928 5652 10934 5704
rect 11241 5695 11299 5701
rect 11241 5661 11253 5695
rect 11287 5692 11299 5695
rect 11514 5692 11520 5704
rect 11287 5664 11520 5692
rect 11287 5661 11299 5664
rect 11241 5655 11299 5661
rect 11514 5652 11520 5664
rect 11572 5692 11578 5704
rect 11977 5695 12035 5701
rect 11977 5692 11989 5695
rect 11572 5664 11989 5692
rect 11572 5652 11578 5664
rect 11977 5661 11989 5664
rect 12023 5661 12035 5695
rect 12452 5692 12480 5720
rect 12710 5692 12716 5704
rect 12452 5664 12716 5692
rect 11977 5655 12035 5661
rect 12710 5652 12716 5664
rect 12768 5652 12774 5704
rect 12805 5695 12863 5701
rect 12805 5661 12817 5695
rect 12851 5661 12863 5695
rect 12805 5655 12863 5661
rect 10597 5627 10655 5633
rect 10597 5624 10609 5627
rect 10244 5596 10609 5624
rect 10597 5593 10609 5596
rect 10643 5593 10655 5627
rect 11425 5627 11483 5633
rect 11425 5624 11437 5627
rect 10597 5587 10655 5593
rect 10704 5596 11437 5624
rect 9398 5556 9404 5568
rect 8772 5528 9404 5556
rect 8205 5519 8263 5525
rect 9398 5516 9404 5528
rect 9456 5516 9462 5568
rect 9858 5516 9864 5568
rect 9916 5556 9922 5568
rect 10704 5556 10732 5596
rect 11425 5593 11437 5596
rect 11471 5593 11483 5627
rect 11425 5587 11483 5593
rect 11698 5584 11704 5636
rect 11756 5624 11762 5636
rect 12253 5627 12311 5633
rect 12253 5624 12265 5627
rect 11756 5596 12265 5624
rect 11756 5584 11762 5596
rect 12253 5593 12265 5596
rect 12299 5593 12311 5627
rect 12253 5587 12311 5593
rect 12434 5584 12440 5636
rect 12492 5624 12498 5636
rect 12820 5624 12848 5655
rect 12492 5596 12848 5624
rect 12492 5584 12498 5596
rect 9916 5528 10732 5556
rect 9916 5516 9922 5528
rect 11054 5516 11060 5568
rect 11112 5556 11118 5568
rect 13354 5556 13360 5568
rect 11112 5528 13360 5556
rect 11112 5516 11118 5528
rect 13354 5516 13360 5528
rect 13412 5516 13418 5568
rect 13998 5556 14004 5568
rect 13959 5528 14004 5556
rect 13998 5516 14004 5528
rect 14056 5516 14062 5568
rect 1104 5466 16008 5488
rect 1104 5414 3480 5466
rect 3532 5414 3544 5466
rect 3596 5414 3608 5466
rect 3660 5414 3672 5466
rect 3724 5414 8478 5466
rect 8530 5414 8542 5466
rect 8594 5414 8606 5466
rect 8658 5414 8670 5466
rect 8722 5414 13475 5466
rect 13527 5414 13539 5466
rect 13591 5414 13603 5466
rect 13655 5414 13667 5466
rect 13719 5414 16008 5466
rect 1104 5392 16008 5414
rect 1486 5352 1492 5364
rect 1447 5324 1492 5352
rect 1486 5312 1492 5324
rect 1544 5312 1550 5364
rect 3329 5355 3387 5361
rect 3329 5321 3341 5355
rect 3375 5352 3387 5355
rect 4798 5352 4804 5364
rect 3375 5324 4804 5352
rect 3375 5321 3387 5324
rect 3329 5315 3387 5321
rect 4798 5312 4804 5324
rect 4856 5312 4862 5364
rect 5166 5312 5172 5364
rect 5224 5352 5230 5364
rect 9490 5352 9496 5364
rect 5224 5324 9496 5352
rect 5224 5312 5230 5324
rect 9490 5312 9496 5324
rect 9548 5312 9554 5364
rect 10042 5312 10048 5364
rect 10100 5352 10106 5364
rect 10229 5355 10287 5361
rect 10229 5352 10241 5355
rect 10100 5324 10241 5352
rect 10100 5312 10106 5324
rect 10229 5321 10241 5324
rect 10275 5321 10287 5355
rect 10229 5315 10287 5321
rect 10410 5312 10416 5364
rect 10468 5352 10474 5364
rect 11330 5352 11336 5364
rect 10468 5324 11336 5352
rect 10468 5312 10474 5324
rect 11330 5312 11336 5324
rect 11388 5312 11394 5364
rect 11422 5312 11428 5364
rect 11480 5352 11486 5364
rect 12250 5352 12256 5364
rect 11480 5324 12256 5352
rect 11480 5312 11486 5324
rect 12250 5312 12256 5324
rect 12308 5312 12314 5364
rect 12710 5312 12716 5364
rect 12768 5352 12774 5364
rect 12897 5355 12955 5361
rect 12897 5352 12909 5355
rect 12768 5324 12909 5352
rect 12768 5312 12774 5324
rect 12897 5321 12909 5324
rect 12943 5321 12955 5355
rect 12897 5315 12955 5321
rect 13078 5312 13084 5364
rect 13136 5352 13142 5364
rect 13265 5355 13323 5361
rect 13265 5352 13277 5355
rect 13136 5324 13277 5352
rect 13136 5312 13142 5324
rect 13265 5321 13277 5324
rect 13311 5321 13323 5355
rect 13265 5315 13323 5321
rect 2130 5284 2136 5296
rect 1964 5256 2136 5284
rect 1964 5225 1992 5256
rect 2130 5244 2136 5256
rect 2188 5244 2194 5296
rect 3421 5287 3479 5293
rect 3421 5284 3433 5287
rect 2792 5256 3433 5284
rect 1949 5219 2007 5225
rect 1949 5185 1961 5219
rect 1995 5185 2007 5219
rect 1949 5179 2007 5185
rect 2041 5219 2099 5225
rect 2041 5185 2053 5219
rect 2087 5216 2099 5219
rect 2590 5216 2596 5228
rect 2087 5188 2596 5216
rect 2087 5185 2099 5188
rect 2041 5179 2099 5185
rect 2590 5176 2596 5188
rect 2648 5176 2654 5228
rect 2792 5225 2820 5256
rect 3421 5253 3433 5256
rect 3467 5284 3479 5287
rect 3786 5284 3792 5296
rect 3467 5256 3792 5284
rect 3467 5253 3479 5256
rect 3421 5247 3479 5253
rect 3786 5244 3792 5256
rect 3844 5244 3850 5296
rect 7466 5244 7472 5296
rect 7524 5284 7530 5296
rect 7929 5287 7987 5293
rect 7929 5284 7941 5287
rect 7524 5256 7941 5284
rect 7524 5244 7530 5256
rect 7929 5253 7941 5256
rect 7975 5253 7987 5287
rect 7929 5247 7987 5253
rect 9398 5244 9404 5296
rect 9456 5284 9462 5296
rect 12802 5284 12808 5296
rect 9456 5256 9996 5284
rect 9456 5244 9462 5256
rect 2777 5219 2835 5225
rect 2777 5185 2789 5219
rect 2823 5185 2835 5219
rect 2777 5179 2835 5185
rect 4801 5219 4859 5225
rect 4801 5185 4813 5219
rect 4847 5216 4859 5219
rect 5074 5216 5080 5228
rect 4847 5188 5080 5216
rect 4847 5185 4859 5188
rect 4801 5179 4859 5185
rect 5074 5176 5080 5188
rect 5132 5176 5138 5228
rect 6196 5188 6601 5216
rect 1581 5151 1639 5157
rect 1581 5117 1593 5151
rect 1627 5148 1639 5151
rect 1854 5148 1860 5160
rect 1627 5120 1860 5148
rect 1627 5117 1639 5120
rect 1581 5111 1639 5117
rect 1854 5108 1860 5120
rect 1912 5108 1918 5160
rect 2498 5108 2504 5160
rect 2556 5148 2562 5160
rect 2961 5151 3019 5157
rect 2961 5148 2973 5151
rect 2556 5120 2973 5148
rect 2556 5108 2562 5120
rect 2961 5117 2973 5120
rect 3007 5117 3019 5151
rect 2961 5111 3019 5117
rect 4154 5108 4160 5160
rect 4212 5148 4218 5160
rect 6196 5148 6224 5188
rect 4212 5120 6224 5148
rect 6273 5151 6331 5157
rect 4212 5108 4218 5120
rect 6273 5117 6285 5151
rect 6319 5148 6331 5151
rect 6454 5148 6460 5160
rect 6319 5120 6460 5148
rect 6319 5117 6331 5120
rect 6273 5111 6331 5117
rect 6454 5108 6460 5120
rect 6512 5108 6518 5160
rect 6573 5148 6601 5188
rect 9490 5176 9496 5228
rect 9548 5216 9554 5228
rect 9968 5225 9996 5256
rect 10888 5256 12808 5284
rect 9861 5219 9919 5225
rect 9861 5216 9873 5219
rect 9548 5188 9873 5216
rect 9548 5176 9554 5188
rect 9861 5185 9873 5188
rect 9907 5185 9919 5219
rect 9861 5179 9919 5185
rect 9953 5219 10011 5225
rect 9953 5185 9965 5219
rect 9999 5216 10011 5219
rect 10781 5219 10839 5225
rect 10781 5216 10793 5219
rect 9999 5188 10793 5216
rect 9999 5185 10011 5188
rect 9953 5179 10011 5185
rect 10781 5185 10793 5188
rect 10827 5185 10839 5219
rect 10781 5179 10839 5185
rect 8754 5148 8760 5160
rect 6573 5120 8760 5148
rect 8754 5108 8760 5120
rect 8812 5108 8818 5160
rect 9030 5108 9036 5160
rect 9088 5157 9094 5160
rect 9088 5148 9100 5157
rect 9088 5120 9133 5148
rect 9088 5111 9100 5120
rect 9088 5108 9094 5111
rect 9214 5108 9220 5160
rect 9272 5148 9278 5160
rect 9309 5151 9367 5157
rect 9309 5148 9321 5151
rect 9272 5120 9321 5148
rect 9272 5108 9278 5120
rect 9309 5117 9321 5120
rect 9355 5117 9367 5151
rect 9309 5111 9367 5117
rect 9398 5108 9404 5160
rect 9456 5148 9462 5160
rect 9769 5151 9827 5157
rect 9769 5148 9781 5151
rect 9456 5120 9781 5148
rect 9456 5108 9462 5120
rect 9769 5117 9781 5120
rect 9815 5148 9827 5151
rect 10502 5148 10508 5160
rect 9815 5120 10508 5148
rect 9815 5117 9827 5120
rect 9769 5111 9827 5117
rect 10502 5108 10508 5120
rect 10560 5108 10566 5160
rect 2133 5083 2191 5089
rect 2133 5049 2145 5083
rect 2179 5080 2191 5083
rect 3510 5080 3516 5092
rect 2179 5052 3516 5080
rect 2179 5049 2191 5052
rect 2133 5043 2191 5049
rect 3510 5040 3516 5052
rect 3568 5040 3574 5092
rect 3602 5040 3608 5092
rect 3660 5080 3666 5092
rect 4556 5083 4614 5089
rect 4556 5080 4568 5083
rect 3660 5052 4568 5080
rect 3660 5040 3666 5052
rect 4556 5049 4568 5052
rect 4602 5080 4614 5083
rect 4798 5080 4804 5092
rect 4602 5052 4804 5080
rect 4602 5049 4614 5052
rect 4556 5043 4614 5049
rect 4798 5040 4804 5052
rect 4856 5040 4862 5092
rect 5258 5040 5264 5092
rect 5316 5080 5322 5092
rect 5626 5080 5632 5092
rect 5316 5052 5632 5080
rect 5316 5040 5322 5052
rect 5626 5040 5632 5052
rect 5684 5040 5690 5092
rect 6028 5083 6086 5089
rect 6028 5049 6040 5083
rect 6074 5080 6086 5083
rect 6546 5080 6552 5092
rect 6074 5052 6552 5080
rect 6074 5049 6086 5052
rect 6028 5043 6086 5049
rect 6546 5040 6552 5052
rect 6604 5040 6610 5092
rect 6638 5040 6644 5092
rect 6696 5089 6702 5092
rect 6696 5083 6760 5089
rect 6696 5049 6714 5083
rect 6748 5049 6760 5083
rect 6696 5043 6760 5049
rect 6901 5052 9444 5080
rect 6696 5040 6702 5043
rect 2314 4972 2320 5024
rect 2372 5012 2378 5024
rect 2501 5015 2559 5021
rect 2501 5012 2513 5015
rect 2372 4984 2513 5012
rect 2372 4972 2378 4984
rect 2501 4981 2513 4984
rect 2547 4981 2559 5015
rect 2501 4975 2559 4981
rect 2869 5015 2927 5021
rect 2869 4981 2881 5015
rect 2915 5012 2927 5015
rect 3142 5012 3148 5024
rect 2915 4984 3148 5012
rect 2915 4981 2927 4984
rect 2869 4975 2927 4981
rect 3142 4972 3148 4984
rect 3200 4972 3206 5024
rect 4890 5012 4896 5024
rect 4851 4984 4896 5012
rect 4890 4972 4896 4984
rect 4948 5012 4954 5024
rect 5534 5012 5540 5024
rect 4948 4984 5540 5012
rect 4948 4972 4954 4984
rect 5534 4972 5540 4984
rect 5592 4972 5598 5024
rect 5718 4972 5724 5024
rect 5776 5012 5782 5024
rect 6901 5012 6929 5052
rect 5776 4984 6929 5012
rect 5776 4972 5782 4984
rect 7006 4972 7012 5024
rect 7064 5012 7070 5024
rect 7282 5012 7288 5024
rect 7064 4984 7288 5012
rect 7064 4972 7070 4984
rect 7282 4972 7288 4984
rect 7340 4972 7346 5024
rect 7834 5012 7840 5024
rect 7795 4984 7840 5012
rect 7834 4972 7840 4984
rect 7892 4972 7898 5024
rect 8202 4972 8208 5024
rect 8260 5012 8266 5024
rect 9122 5012 9128 5024
rect 8260 4984 9128 5012
rect 8260 4972 8266 4984
rect 9122 4972 9128 4984
rect 9180 4972 9186 5024
rect 9416 5021 9444 5052
rect 10410 5040 10416 5092
rect 10468 5080 10474 5092
rect 10594 5080 10600 5092
rect 10468 5052 10600 5080
rect 10468 5040 10474 5052
rect 10594 5040 10600 5052
rect 10652 5040 10658 5092
rect 10689 5083 10747 5089
rect 10689 5049 10701 5083
rect 10735 5080 10747 5083
rect 10778 5080 10784 5092
rect 10735 5052 10784 5080
rect 10735 5049 10747 5052
rect 10689 5043 10747 5049
rect 10778 5040 10784 5052
rect 10836 5040 10842 5092
rect 9401 5015 9459 5021
rect 9401 4981 9413 5015
rect 9447 4981 9459 5015
rect 9401 4975 9459 4981
rect 9582 4972 9588 5024
rect 9640 5012 9646 5024
rect 10888 5012 10916 5256
rect 12802 5244 12808 5256
rect 12860 5244 12866 5296
rect 13280 5284 13308 5315
rect 13446 5284 13452 5296
rect 13280 5256 13452 5284
rect 13446 5244 13452 5256
rect 13504 5244 13510 5296
rect 13538 5244 13544 5296
rect 13596 5284 13602 5296
rect 14458 5284 14464 5296
rect 13596 5256 14464 5284
rect 13596 5244 13602 5256
rect 14458 5244 14464 5256
rect 14516 5244 14522 5296
rect 11514 5216 11520 5228
rect 11475 5188 11520 5216
rect 11514 5176 11520 5188
rect 11572 5176 11578 5228
rect 11790 5176 11796 5228
rect 11848 5216 11854 5228
rect 12253 5219 12311 5225
rect 12253 5216 12265 5219
rect 11848 5188 12265 5216
rect 11848 5176 11854 5188
rect 12253 5185 12265 5188
rect 12299 5185 12311 5219
rect 12253 5179 12311 5185
rect 12710 5176 12716 5228
rect 12768 5216 12774 5228
rect 14826 5216 14832 5228
rect 12768 5188 14832 5216
rect 12768 5176 12774 5188
rect 14826 5176 14832 5188
rect 14884 5176 14890 5228
rect 10962 5108 10968 5160
rect 11020 5148 11026 5160
rect 12069 5151 12127 5157
rect 12069 5148 12081 5151
rect 11020 5120 12081 5148
rect 11020 5108 11026 5120
rect 12069 5117 12081 5120
rect 12115 5117 12127 5151
rect 12069 5111 12127 5117
rect 12161 5151 12219 5157
rect 12161 5117 12173 5151
rect 12207 5148 12219 5151
rect 12434 5148 12440 5160
rect 12207 5120 12440 5148
rect 12207 5117 12219 5120
rect 12161 5111 12219 5117
rect 12434 5108 12440 5120
rect 12492 5108 12498 5160
rect 14090 5148 14096 5160
rect 12544 5120 14096 5148
rect 11054 5080 11060 5092
rect 11015 5052 11060 5080
rect 11054 5040 11060 5052
rect 11112 5040 11118 5092
rect 11241 5083 11299 5089
rect 11241 5049 11253 5083
rect 11287 5080 11299 5083
rect 12544 5080 12572 5120
rect 14090 5108 14096 5120
rect 14148 5108 14154 5160
rect 11287 5052 12572 5080
rect 12621 5083 12679 5089
rect 11287 5049 11299 5052
rect 11241 5043 11299 5049
rect 12621 5049 12633 5083
rect 12667 5080 12679 5083
rect 12986 5080 12992 5092
rect 12667 5052 12992 5080
rect 12667 5049 12679 5052
rect 12621 5043 12679 5049
rect 12986 5040 12992 5052
rect 13044 5040 13050 5092
rect 9640 4984 10916 5012
rect 9640 4972 9646 4984
rect 11514 4972 11520 5024
rect 11572 5012 11578 5024
rect 11701 5015 11759 5021
rect 11701 5012 11713 5015
rect 11572 4984 11713 5012
rect 11572 4972 11578 4984
rect 11701 4981 11713 4984
rect 11747 4981 11759 5015
rect 11701 4975 11759 4981
rect 11790 4972 11796 5024
rect 11848 5012 11854 5024
rect 12713 5015 12771 5021
rect 12713 5012 12725 5015
rect 11848 4984 12725 5012
rect 11848 4972 11854 4984
rect 12713 4981 12725 4984
rect 12759 4981 12771 5015
rect 13078 5012 13084 5024
rect 13039 4984 13084 5012
rect 12713 4975 12771 4981
rect 13078 4972 13084 4984
rect 13136 4972 13142 5024
rect 13630 5012 13636 5024
rect 13591 4984 13636 5012
rect 13630 4972 13636 4984
rect 13688 5012 13694 5024
rect 13998 5012 14004 5024
rect 13688 4984 14004 5012
rect 13688 4972 13694 4984
rect 13998 4972 14004 4984
rect 14056 4972 14062 5024
rect 1104 4922 16008 4944
rect 1104 4870 5979 4922
rect 6031 4870 6043 4922
rect 6095 4870 6107 4922
rect 6159 4870 6171 4922
rect 6223 4870 10976 4922
rect 11028 4870 11040 4922
rect 11092 4870 11104 4922
rect 11156 4870 11168 4922
rect 11220 4870 16008 4922
rect 1104 4848 16008 4870
rect 2133 4811 2191 4817
rect 2133 4808 2145 4811
rect 1596 4780 2145 4808
rect 1596 4749 1624 4780
rect 2133 4777 2145 4780
rect 2179 4777 2191 4811
rect 2961 4811 3019 4817
rect 2961 4808 2973 4811
rect 2133 4771 2191 4777
rect 2746 4780 2973 4808
rect 1581 4743 1639 4749
rect 1581 4709 1593 4743
rect 1627 4709 1639 4743
rect 1581 4703 1639 4709
rect 1670 4632 1676 4684
rect 1728 4672 1734 4684
rect 1765 4675 1823 4681
rect 1765 4672 1777 4675
rect 1728 4644 1777 4672
rect 1728 4632 1734 4644
rect 1765 4641 1777 4644
rect 1811 4641 1823 4675
rect 2314 4672 2320 4684
rect 2275 4644 2320 4672
rect 1765 4635 1823 4641
rect 2314 4632 2320 4644
rect 2372 4632 2378 4684
rect 2593 4675 2651 4681
rect 2593 4641 2605 4675
rect 2639 4672 2651 4675
rect 2746 4672 2774 4780
rect 2961 4777 2973 4780
rect 3007 4777 3019 4811
rect 2961 4771 3019 4777
rect 3326 4768 3332 4820
rect 3384 4768 3390 4820
rect 4798 4808 4804 4820
rect 4759 4780 4804 4808
rect 4798 4768 4804 4780
rect 4856 4768 4862 4820
rect 4893 4811 4951 4817
rect 4893 4777 4905 4811
rect 4939 4808 4951 4811
rect 8018 4808 8024 4820
rect 4939 4780 8024 4808
rect 4939 4777 4951 4780
rect 4893 4771 4951 4777
rect 8018 4768 8024 4780
rect 8076 4768 8082 4820
rect 9122 4768 9128 4820
rect 9180 4808 9186 4820
rect 9490 4808 9496 4820
rect 9180 4780 9496 4808
rect 9180 4768 9186 4780
rect 9490 4768 9496 4780
rect 9548 4768 9554 4820
rect 9585 4811 9643 4817
rect 9585 4777 9597 4811
rect 9631 4808 9643 4811
rect 9766 4808 9772 4820
rect 9631 4780 9772 4808
rect 9631 4777 9643 4780
rect 9585 4771 9643 4777
rect 9766 4768 9772 4780
rect 9824 4768 9830 4820
rect 9858 4768 9864 4820
rect 9916 4808 9922 4820
rect 10042 4808 10048 4820
rect 9916 4780 10048 4808
rect 9916 4768 9922 4780
rect 10042 4768 10048 4780
rect 10100 4768 10106 4820
rect 10413 4811 10471 4817
rect 10413 4777 10425 4811
rect 10459 4808 10471 4811
rect 11698 4808 11704 4820
rect 10459 4780 11560 4808
rect 11659 4780 11704 4808
rect 10459 4777 10471 4780
rect 10413 4771 10471 4777
rect 3344 4740 3372 4768
rect 5810 4740 5816 4752
rect 3344 4712 5816 4740
rect 5810 4700 5816 4712
rect 5868 4700 5874 4752
rect 10321 4743 10379 4749
rect 10321 4740 10333 4743
rect 6297 4712 10333 4740
rect 2639 4644 2774 4672
rect 2869 4675 2927 4681
rect 2639 4641 2651 4644
rect 2593 4635 2651 4641
rect 2869 4641 2881 4675
rect 2915 4672 2927 4675
rect 3142 4672 3148 4684
rect 2915 4644 3148 4672
rect 2915 4641 2927 4644
rect 2869 4635 2927 4641
rect 3142 4632 3148 4644
rect 3200 4632 3206 4684
rect 3326 4672 3332 4684
rect 3287 4644 3332 4672
rect 3326 4632 3332 4644
rect 3384 4632 3390 4684
rect 4154 4672 4160 4684
rect 4115 4644 4160 4672
rect 4154 4632 4160 4644
rect 4212 4632 4218 4684
rect 4433 4675 4491 4681
rect 4433 4641 4445 4675
rect 4479 4672 4491 4675
rect 6297 4672 6325 4712
rect 10321 4709 10333 4712
rect 10367 4709 10379 4743
rect 10321 4703 10379 4709
rect 4479 4644 6325 4672
rect 4479 4641 4491 4644
rect 4433 4635 4491 4641
rect 6454 4632 6460 4684
rect 6512 4681 6518 4684
rect 6512 4672 6524 4681
rect 6512 4644 6557 4672
rect 6512 4635 6524 4644
rect 6512 4632 6518 4635
rect 6638 4632 6644 4684
rect 6696 4672 6702 4684
rect 6733 4675 6791 4681
rect 6733 4672 6745 4675
rect 6696 4644 6745 4672
rect 6696 4632 6702 4644
rect 6733 4641 6745 4644
rect 6779 4641 6791 4675
rect 6733 4635 6791 4641
rect 7374 4632 7380 4684
rect 7432 4672 7438 4684
rect 7949 4675 8007 4681
rect 7949 4672 7961 4675
rect 7432 4644 7961 4672
rect 7432 4632 7438 4644
rect 7949 4641 7961 4644
rect 7995 4672 8007 4675
rect 8294 4672 8300 4684
rect 7995 4644 8300 4672
rect 7995 4641 8007 4644
rect 7949 4635 8007 4641
rect 8294 4632 8300 4644
rect 8352 4632 8358 4684
rect 8757 4675 8815 4681
rect 8757 4641 8769 4675
rect 8803 4672 8815 4675
rect 9493 4675 9551 4681
rect 9493 4672 9505 4675
rect 8803 4644 9505 4672
rect 8803 4641 8815 4644
rect 8757 4635 8815 4641
rect 9493 4641 9505 4644
rect 9539 4641 9551 4675
rect 10428 4672 10456 4771
rect 10502 4700 10508 4752
rect 10560 4740 10566 4752
rect 10560 4712 11017 4740
rect 10560 4700 10566 4712
rect 9493 4635 9551 4641
rect 9600 4644 9996 4672
rect 10428 4644 10640 4672
rect 3418 4604 3424 4616
rect 3379 4576 3424 4604
rect 3418 4564 3424 4576
rect 3476 4564 3482 4616
rect 3602 4604 3608 4616
rect 3563 4576 3608 4604
rect 3602 4564 3608 4576
rect 3660 4564 3666 4616
rect 4709 4607 4767 4613
rect 4709 4573 4721 4607
rect 4755 4604 4767 4607
rect 4755 4576 5764 4604
rect 4755 4573 4767 4576
rect 4709 4567 4767 4573
rect 2130 4496 2136 4548
rect 2188 4536 2194 4548
rect 2685 4539 2743 4545
rect 2685 4536 2697 4539
rect 2188 4508 2697 4536
rect 2188 4496 2194 4508
rect 2685 4505 2697 4508
rect 2731 4505 2743 4539
rect 2685 4499 2743 4505
rect 4338 4496 4344 4548
rect 4396 4536 4402 4548
rect 5166 4536 5172 4548
rect 4396 4508 5172 4536
rect 4396 4496 4402 4508
rect 5166 4496 5172 4508
rect 5224 4496 5230 4548
rect 1486 4468 1492 4480
rect 1447 4440 1492 4468
rect 1486 4428 1492 4440
rect 1544 4428 1550 4480
rect 1946 4468 1952 4480
rect 1907 4440 1952 4468
rect 1946 4428 1952 4440
rect 2004 4428 2010 4480
rect 2038 4428 2044 4480
rect 2096 4468 2102 4480
rect 2409 4471 2467 4477
rect 2409 4468 2421 4471
rect 2096 4440 2421 4468
rect 2096 4428 2102 4440
rect 2409 4437 2421 4440
rect 2455 4437 2467 4471
rect 2409 4431 2467 4437
rect 3786 4428 3792 4480
rect 3844 4468 3850 4480
rect 3973 4471 4031 4477
rect 3973 4468 3985 4471
rect 3844 4440 3985 4468
rect 3844 4428 3850 4440
rect 3973 4437 3985 4440
rect 4019 4437 4031 4471
rect 5258 4468 5264 4480
rect 5219 4440 5264 4468
rect 3973 4431 4031 4437
rect 5258 4428 5264 4440
rect 5316 4428 5322 4480
rect 5350 4428 5356 4480
rect 5408 4468 5414 4480
rect 5736 4468 5764 4576
rect 6822 4564 6828 4616
rect 6880 4604 6886 4616
rect 8202 4604 8208 4616
rect 6880 4576 6960 4604
rect 8163 4576 8208 4604
rect 6880 4564 6886 4576
rect 6730 4468 6736 4480
rect 5408 4440 5453 4468
rect 5736 4440 6736 4468
rect 5408 4428 5414 4440
rect 6730 4428 6736 4440
rect 6788 4468 6794 4480
rect 6825 4471 6883 4477
rect 6825 4468 6837 4471
rect 6788 4440 6837 4468
rect 6788 4428 6794 4440
rect 6825 4437 6837 4440
rect 6871 4437 6883 4471
rect 6932 4468 6960 4576
rect 8202 4564 8208 4576
rect 8260 4564 8266 4616
rect 8481 4607 8539 4613
rect 8481 4573 8493 4607
rect 8527 4604 8539 4607
rect 8527 4576 9260 4604
rect 8527 4573 8539 4576
rect 8481 4567 8539 4573
rect 9125 4539 9183 4545
rect 9125 4536 9137 4539
rect 8220 4508 9137 4536
rect 8220 4468 8248 4508
rect 9125 4505 9137 4508
rect 9171 4505 9183 4539
rect 9232 4536 9260 4576
rect 9306 4564 9312 4616
rect 9364 4604 9370 4616
rect 9600 4604 9628 4644
rect 9364 4576 9628 4604
rect 9677 4607 9735 4613
rect 9364 4564 9370 4576
rect 9677 4573 9689 4607
rect 9723 4573 9735 4607
rect 9677 4567 9735 4573
rect 9490 4536 9496 4548
rect 9232 4508 9496 4536
rect 9125 4499 9183 4505
rect 9490 4496 9496 4508
rect 9548 4496 9554 4548
rect 9582 4496 9588 4548
rect 9640 4536 9646 4548
rect 9692 4536 9720 4567
rect 9968 4545 9996 4644
rect 10505 4607 10563 4613
rect 10505 4604 10517 4607
rect 10060 4576 10517 4604
rect 9640 4508 9720 4536
rect 9953 4539 10011 4545
rect 9640 4496 9646 4508
rect 9953 4505 9965 4539
rect 9999 4505 10011 4539
rect 9953 4499 10011 4505
rect 8846 4468 8852 4480
rect 6932 4440 8248 4468
rect 8807 4440 8852 4468
rect 6825 4431 6883 4437
rect 8846 4428 8852 4440
rect 8904 4428 8910 4480
rect 9030 4428 9036 4480
rect 9088 4468 9094 4480
rect 10060 4468 10088 4576
rect 10505 4573 10517 4576
rect 10551 4573 10563 4607
rect 10505 4567 10563 4573
rect 10318 4496 10324 4548
rect 10376 4536 10382 4548
rect 10612 4536 10640 4644
rect 10686 4632 10692 4684
rect 10744 4672 10750 4684
rect 10989 4672 11017 4712
rect 11054 4700 11060 4752
rect 11112 4740 11118 4752
rect 11532 4740 11560 4780
rect 11698 4768 11704 4780
rect 11756 4768 11762 4820
rect 12434 4808 12440 4820
rect 12084 4780 12440 4808
rect 12084 4740 12112 4780
rect 12434 4768 12440 4780
rect 12492 4808 12498 4820
rect 12989 4811 13047 4817
rect 12989 4808 13001 4811
rect 12492 4780 13001 4808
rect 12492 4768 12498 4780
rect 12989 4777 13001 4780
rect 13035 4808 13047 4811
rect 13078 4808 13084 4820
rect 13035 4780 13084 4808
rect 13035 4777 13047 4780
rect 12989 4771 13047 4777
rect 13078 4768 13084 4780
rect 13136 4808 13142 4820
rect 13262 4808 13268 4820
rect 13136 4780 13268 4808
rect 13136 4768 13142 4780
rect 13262 4768 13268 4780
rect 13320 4768 13326 4820
rect 13446 4808 13452 4820
rect 13407 4780 13452 4808
rect 13446 4768 13452 4780
rect 13504 4768 13510 4820
rect 14093 4811 14151 4817
rect 14093 4777 14105 4811
rect 14139 4808 14151 4811
rect 14734 4808 14740 4820
rect 14139 4780 14740 4808
rect 14139 4777 14151 4780
rect 14093 4771 14151 4777
rect 14734 4768 14740 4780
rect 14792 4768 14798 4820
rect 11112 4712 11157 4740
rect 11532 4712 12112 4740
rect 12161 4743 12219 4749
rect 11112 4700 11118 4712
rect 12161 4709 12173 4743
rect 12207 4740 12219 4743
rect 15010 4740 15016 4752
rect 12207 4712 15016 4740
rect 12207 4709 12219 4712
rect 12161 4703 12219 4709
rect 15010 4700 15016 4712
rect 15068 4700 15074 4752
rect 11149 4675 11207 4681
rect 10744 4644 10916 4672
rect 10989 4644 11100 4672
rect 10744 4632 10750 4644
rect 10888 4613 10916 4644
rect 10873 4607 10931 4613
rect 10873 4573 10885 4607
rect 10919 4573 10931 4607
rect 11072 4604 11100 4644
rect 11149 4641 11161 4675
rect 11195 4672 11207 4675
rect 11698 4672 11704 4684
rect 11195 4644 11704 4672
rect 11195 4641 11207 4644
rect 11149 4635 11207 4641
rect 11698 4632 11704 4644
rect 11756 4632 11762 4684
rect 11793 4675 11851 4681
rect 11793 4641 11805 4675
rect 11839 4641 11851 4675
rect 11793 4635 11851 4641
rect 11808 4604 11836 4635
rect 11882 4632 11888 4684
rect 11940 4672 11946 4684
rect 12342 4672 12348 4684
rect 11940 4644 12348 4672
rect 11940 4632 11946 4644
rect 12342 4632 12348 4644
rect 12400 4632 12406 4684
rect 12529 4675 12587 4681
rect 12529 4641 12541 4675
rect 12575 4672 12587 4675
rect 13078 4672 13084 4684
rect 12575 4644 13084 4672
rect 12575 4641 12587 4644
rect 12529 4635 12587 4641
rect 13078 4632 13084 4644
rect 13136 4632 13142 4684
rect 13630 4672 13636 4684
rect 13591 4644 13636 4672
rect 13630 4632 13636 4644
rect 13688 4672 13694 4684
rect 13817 4675 13875 4681
rect 13817 4672 13829 4675
rect 13688 4644 13829 4672
rect 13688 4632 13694 4644
rect 13817 4641 13829 4644
rect 13863 4672 13875 4675
rect 13998 4672 14004 4684
rect 13863 4644 14004 4672
rect 13863 4641 13875 4644
rect 13817 4635 13875 4641
rect 13998 4632 14004 4644
rect 14056 4632 14062 4684
rect 14550 4604 14556 4616
rect 11072 4576 11744 4604
rect 11808 4576 14556 4604
rect 10873 4567 10931 4573
rect 11054 4536 11060 4548
rect 10376 4508 10640 4536
rect 10704 4508 11060 4536
rect 10376 4496 10382 4508
rect 10704 4480 10732 4508
rect 11054 4496 11060 4508
rect 11112 4496 11118 4548
rect 11330 4496 11336 4548
rect 11388 4536 11394 4548
rect 11517 4539 11575 4545
rect 11517 4536 11529 4539
rect 11388 4508 11529 4536
rect 11388 4496 11394 4508
rect 11517 4505 11529 4508
rect 11563 4505 11575 4539
rect 11716 4536 11744 4576
rect 14550 4564 14556 4576
rect 14608 4564 14614 4616
rect 11790 4536 11796 4548
rect 11716 4508 11796 4536
rect 11517 4499 11575 4505
rect 11790 4496 11796 4508
rect 11848 4496 11854 4548
rect 11974 4536 11980 4548
rect 11935 4508 11980 4536
rect 11974 4496 11980 4508
rect 12032 4496 12038 4548
rect 12342 4496 12348 4548
rect 12400 4536 12406 4548
rect 12713 4539 12771 4545
rect 12713 4536 12725 4539
rect 12400 4508 12725 4536
rect 12400 4496 12406 4508
rect 12713 4505 12725 4508
rect 12759 4505 12771 4539
rect 12713 4499 12771 4505
rect 12986 4496 12992 4548
rect 13044 4536 13050 4548
rect 13265 4539 13323 4545
rect 13265 4536 13277 4539
rect 13044 4508 13277 4536
rect 13044 4496 13050 4508
rect 13265 4505 13277 4508
rect 13311 4536 13323 4539
rect 14274 4536 14280 4548
rect 13311 4508 14280 4536
rect 13311 4505 13323 4508
rect 13265 4499 13323 4505
rect 14274 4496 14280 4508
rect 14332 4496 14338 4548
rect 9088 4440 10088 4468
rect 9088 4428 9094 4440
rect 10134 4428 10140 4480
rect 10192 4468 10198 4480
rect 10502 4468 10508 4480
rect 10192 4440 10508 4468
rect 10192 4428 10198 4440
rect 10502 4428 10508 4440
rect 10560 4428 10566 4480
rect 10686 4428 10692 4480
rect 10744 4428 10750 4480
rect 10778 4428 10784 4480
rect 10836 4468 10842 4480
rect 12437 4471 12495 4477
rect 12437 4468 12449 4471
rect 10836 4440 12449 4468
rect 10836 4428 10842 4440
rect 12437 4437 12449 4440
rect 12483 4437 12495 4471
rect 12437 4431 12495 4437
rect 12894 4428 12900 4480
rect 12952 4468 12958 4480
rect 13081 4471 13139 4477
rect 13081 4468 13093 4471
rect 12952 4440 13093 4468
rect 12952 4428 12958 4440
rect 13081 4437 13093 4440
rect 13127 4437 13139 4471
rect 13081 4431 13139 4437
rect 1104 4378 16008 4400
rect 1104 4326 3480 4378
rect 3532 4326 3544 4378
rect 3596 4326 3608 4378
rect 3660 4326 3672 4378
rect 3724 4326 8478 4378
rect 8530 4326 8542 4378
rect 8594 4326 8606 4378
rect 8658 4326 8670 4378
rect 8722 4326 13475 4378
rect 13527 4326 13539 4378
rect 13591 4326 13603 4378
rect 13655 4326 13667 4378
rect 13719 4326 16008 4378
rect 1104 4304 16008 4326
rect 3326 4224 3332 4276
rect 3384 4264 3390 4276
rect 3881 4267 3939 4273
rect 3881 4264 3893 4267
rect 3384 4236 3893 4264
rect 3384 4224 3390 4236
rect 3881 4233 3893 4236
rect 3927 4233 3939 4267
rect 3881 4227 3939 4233
rect 4709 4267 4767 4273
rect 4709 4233 4721 4267
rect 4755 4264 4767 4267
rect 4798 4264 4804 4276
rect 4755 4236 4804 4264
rect 4755 4233 4767 4236
rect 4709 4227 4767 4233
rect 4798 4224 4804 4236
rect 4856 4224 4862 4276
rect 5166 4224 5172 4276
rect 5224 4264 5230 4276
rect 5350 4264 5356 4276
rect 5224 4236 5356 4264
rect 5224 4224 5230 4236
rect 5350 4224 5356 4236
rect 5408 4264 5414 4276
rect 7374 4264 7380 4276
rect 5408 4236 7380 4264
rect 5408 4224 5414 4236
rect 7374 4224 7380 4236
rect 7432 4224 7438 4276
rect 7742 4224 7748 4276
rect 7800 4264 7806 4276
rect 7837 4267 7895 4273
rect 7837 4264 7849 4267
rect 7800 4236 7849 4264
rect 7800 4224 7806 4236
rect 7837 4233 7849 4236
rect 7883 4233 7895 4267
rect 7837 4227 7895 4233
rect 7929 4267 7987 4273
rect 7929 4233 7941 4267
rect 7975 4264 7987 4267
rect 8018 4264 8024 4276
rect 7975 4236 8024 4264
rect 7975 4233 7987 4236
rect 7929 4227 7987 4233
rect 8018 4224 8024 4236
rect 8076 4224 8082 4276
rect 9122 4264 9128 4276
rect 8128 4236 9128 4264
rect 2685 4199 2743 4205
rect 2685 4165 2697 4199
rect 2731 4196 2743 4199
rect 3602 4196 3608 4208
rect 2731 4168 3608 4196
rect 2731 4165 2743 4168
rect 2685 4159 2743 4165
rect 3602 4156 3608 4168
rect 3660 4156 3666 4208
rect 5902 4196 5908 4208
rect 4540 4168 5908 4196
rect 1762 4088 1768 4140
rect 1820 4128 1826 4140
rect 1820 4100 2544 4128
rect 1820 4088 1826 4100
rect 1581 4063 1639 4069
rect 1581 4029 1593 4063
rect 1627 4060 1639 4063
rect 2038 4060 2044 4072
rect 1627 4032 2044 4060
rect 1627 4029 1639 4032
rect 1581 4023 1639 4029
rect 2038 4020 2044 4032
rect 2096 4020 2102 4072
rect 2225 4063 2283 4069
rect 2225 4029 2237 4063
rect 2271 4060 2283 4063
rect 2406 4060 2412 4072
rect 2271 4032 2412 4060
rect 2271 4029 2283 4032
rect 2225 4023 2283 4029
rect 2406 4020 2412 4032
rect 2464 4020 2470 4072
rect 2516 4069 2544 4100
rect 2866 4088 2872 4140
rect 2924 4128 2930 4140
rect 3513 4131 3571 4137
rect 3513 4128 3525 4131
rect 2924 4100 3525 4128
rect 2924 4088 2930 4100
rect 3513 4097 3525 4100
rect 3559 4097 3571 4131
rect 3513 4091 3571 4097
rect 3697 4131 3755 4137
rect 3697 4097 3709 4131
rect 3743 4128 3755 4131
rect 3878 4128 3884 4140
rect 3743 4100 3884 4128
rect 3743 4097 3755 4100
rect 3697 4091 3755 4097
rect 3878 4088 3884 4100
rect 3936 4088 3942 4140
rect 4338 4128 4344 4140
rect 4299 4100 4344 4128
rect 4338 4088 4344 4100
rect 4396 4088 4402 4140
rect 4540 4137 4568 4168
rect 5902 4156 5908 4168
rect 5960 4156 5966 4208
rect 6012 4168 6509 4196
rect 4525 4131 4583 4137
rect 4525 4097 4537 4131
rect 4571 4097 4583 4131
rect 4525 4091 4583 4097
rect 5166 4088 5172 4140
rect 5224 4128 5230 4140
rect 5261 4131 5319 4137
rect 5261 4128 5273 4131
rect 5224 4100 5273 4128
rect 5224 4088 5230 4100
rect 5261 4097 5273 4100
rect 5307 4097 5319 4131
rect 5261 4091 5319 4097
rect 2501 4063 2559 4069
rect 2501 4029 2513 4063
rect 2547 4029 2559 4063
rect 2501 4023 2559 4029
rect 2774 4020 2780 4072
rect 2832 4060 2838 4072
rect 2832 4032 2877 4060
rect 2832 4020 2838 4032
rect 3418 4020 3424 4072
rect 3476 4060 3482 4072
rect 4062 4060 4068 4072
rect 3476 4032 4068 4060
rect 3476 4020 3482 4032
rect 4062 4020 4068 4032
rect 4120 4020 4126 4072
rect 4430 4020 4436 4072
rect 4488 4060 4494 4072
rect 6012 4060 6040 4168
rect 6089 4131 6147 4137
rect 6089 4097 6101 4131
rect 6135 4097 6147 4131
rect 6481 4128 6509 4168
rect 7466 4156 7472 4208
rect 7524 4196 7530 4208
rect 8128 4196 8156 4236
rect 9122 4224 9128 4236
rect 9180 4224 9186 4276
rect 10413 4267 10471 4273
rect 10413 4264 10425 4267
rect 10253 4236 10425 4264
rect 10253 4208 10281 4236
rect 10413 4233 10425 4236
rect 10459 4233 10471 4267
rect 12250 4264 12256 4276
rect 10413 4227 10471 4233
rect 10520 4236 12112 4264
rect 12211 4236 12256 4264
rect 7524 4168 8156 4196
rect 7524 4156 7530 4168
rect 8294 4156 8300 4208
rect 8352 4196 8358 4208
rect 9582 4196 9588 4208
rect 8352 4168 9588 4196
rect 8352 4156 8358 4168
rect 8478 4128 8484 4140
rect 6481 4100 6592 4128
rect 6089 4091 6147 4097
rect 4488 4032 6040 4060
rect 4488 4020 4494 4032
rect 1949 3995 2007 4001
rect 1949 3961 1961 3995
rect 1995 3992 2007 3995
rect 2130 3992 2136 4004
rect 1995 3964 2136 3992
rect 1995 3961 2007 3964
rect 1949 3955 2007 3961
rect 2130 3952 2136 3964
rect 2188 3952 2194 4004
rect 2866 3992 2872 4004
rect 2424 3964 2872 3992
rect 1486 3924 1492 3936
rect 1447 3896 1492 3924
rect 1486 3884 1492 3896
rect 1544 3884 1550 3936
rect 1854 3924 1860 3936
rect 1815 3896 1860 3924
rect 1854 3884 1860 3896
rect 1912 3884 1918 3936
rect 2424 3933 2452 3964
rect 2866 3952 2872 3964
rect 2924 3952 2930 4004
rect 3878 3992 3884 4004
rect 2976 3964 3884 3992
rect 2976 3933 3004 3964
rect 3878 3952 3884 3964
rect 3936 3952 3942 4004
rect 4338 3952 4344 4004
rect 4396 3992 4402 4004
rect 6104 3992 6132 4091
rect 6454 4060 6460 4072
rect 6512 4069 6518 4072
rect 6422 4032 6460 4060
rect 6454 4020 6460 4032
rect 6512 4023 6522 4069
rect 6564 4060 6592 4100
rect 7484 4100 8484 4128
rect 6713 4063 6771 4069
rect 6713 4060 6725 4063
rect 6564 4032 6725 4060
rect 6713 4029 6725 4032
rect 6759 4029 6771 4063
rect 7484 4060 7512 4100
rect 8478 4088 8484 4100
rect 8536 4088 8542 4140
rect 8588 4137 8616 4168
rect 9582 4156 9588 4168
rect 9640 4156 9646 4208
rect 9766 4156 9772 4208
rect 9824 4196 9830 4208
rect 9824 4168 10180 4196
rect 9824 4156 9830 4168
rect 10152 4140 10180 4168
rect 10226 4156 10232 4208
rect 10284 4156 10290 4208
rect 10520 4196 10548 4236
rect 10336 4168 10548 4196
rect 8573 4131 8631 4137
rect 8573 4097 8585 4131
rect 8619 4097 8631 4131
rect 8573 4091 8631 4097
rect 9030 4088 9036 4140
rect 9088 4128 9094 4140
rect 9309 4131 9367 4137
rect 9309 4128 9321 4131
rect 9088 4100 9321 4128
rect 9088 4088 9094 4100
rect 9309 4097 9321 4100
rect 9355 4097 9367 4131
rect 9309 4091 9367 4097
rect 9950 4088 9956 4140
rect 10008 4128 10014 4140
rect 10045 4131 10103 4137
rect 10045 4128 10057 4131
rect 10008 4100 10057 4128
rect 10008 4088 10014 4100
rect 10045 4097 10057 4100
rect 10091 4097 10103 4131
rect 10045 4091 10103 4097
rect 10134 4088 10140 4140
rect 10192 4128 10198 4140
rect 10192 4100 10237 4128
rect 10192 4088 10198 4100
rect 6713 4023 6771 4029
rect 6886 4032 7512 4060
rect 8297 4063 8355 4069
rect 6512 4020 6518 4023
rect 6362 3992 6368 4004
rect 4396 3964 5948 3992
rect 6104 3964 6368 3992
rect 4396 3952 4402 3964
rect 2409 3927 2467 3933
rect 2409 3893 2421 3927
rect 2455 3893 2467 3927
rect 2409 3887 2467 3893
rect 2961 3927 3019 3933
rect 2961 3893 2973 3927
rect 3007 3893 3019 3927
rect 2961 3887 3019 3893
rect 3050 3884 3056 3936
rect 3108 3924 3114 3936
rect 3421 3927 3479 3933
rect 3108 3896 3153 3924
rect 3108 3884 3114 3896
rect 3421 3893 3433 3927
rect 3467 3924 3479 3927
rect 4062 3924 4068 3936
rect 3467 3896 4068 3924
rect 3467 3893 3479 3896
rect 3421 3887 3479 3893
rect 4062 3884 4068 3896
rect 4120 3884 4126 3936
rect 4249 3927 4307 3933
rect 4249 3893 4261 3927
rect 4295 3924 4307 3927
rect 4798 3924 4804 3936
rect 4295 3896 4804 3924
rect 4295 3893 4307 3896
rect 4249 3887 4307 3893
rect 4798 3884 4804 3896
rect 4856 3884 4862 3936
rect 5074 3924 5080 3936
rect 5035 3896 5080 3924
rect 5074 3884 5080 3896
rect 5132 3884 5138 3936
rect 5920 3933 5948 3964
rect 6362 3952 6368 3964
rect 6420 3952 6426 4004
rect 6481 3992 6509 4020
rect 6886 3992 6914 4032
rect 8297 4029 8309 4063
rect 8343 4060 8355 4063
rect 8754 4060 8760 4072
rect 8343 4032 8760 4060
rect 8343 4029 8355 4032
rect 8297 4023 8355 4029
rect 8754 4020 8760 4032
rect 8812 4020 8818 4072
rect 8864 4032 9260 4060
rect 6481 3964 6914 3992
rect 7374 3952 7380 4004
rect 7432 3992 7438 4004
rect 8389 3995 8447 4001
rect 8389 3992 8401 3995
rect 7432 3964 8401 3992
rect 7432 3952 7438 3964
rect 8389 3961 8401 3964
rect 8435 3961 8447 3995
rect 8389 3955 8447 3961
rect 8478 3952 8484 4004
rect 8536 3992 8542 4004
rect 8864 3992 8892 4032
rect 8536 3964 8892 3992
rect 8536 3952 8542 3964
rect 9030 3952 9036 4004
rect 9088 3992 9094 4004
rect 9125 3995 9183 4001
rect 9125 3992 9137 3995
rect 9088 3964 9137 3992
rect 9088 3952 9094 3964
rect 9125 3961 9137 3964
rect 9171 3961 9183 3995
rect 9232 3992 9260 4032
rect 9398 4020 9404 4072
rect 9456 4060 9462 4072
rect 10336 4060 10364 4168
rect 10870 4156 10876 4208
rect 10928 4196 10934 4208
rect 10965 4199 11023 4205
rect 10965 4196 10977 4199
rect 10928 4168 10977 4196
rect 10928 4156 10934 4168
rect 10965 4165 10977 4168
rect 11011 4165 11023 4199
rect 11146 4196 11152 4208
rect 10965 4159 11023 4165
rect 11072 4168 11152 4196
rect 9456 4032 10364 4060
rect 10597 4063 10655 4069
rect 9456 4020 9462 4032
rect 10597 4029 10609 4063
rect 10643 4060 10655 4063
rect 10643 4032 10732 4060
rect 10643 4029 10655 4032
rect 10597 4023 10655 4029
rect 9953 3995 10011 4001
rect 9232 3964 9904 3992
rect 9125 3955 9183 3961
rect 5169 3927 5227 3933
rect 5169 3893 5181 3927
rect 5215 3924 5227 3927
rect 5537 3927 5595 3933
rect 5537 3924 5549 3927
rect 5215 3896 5549 3924
rect 5215 3893 5227 3896
rect 5169 3887 5227 3893
rect 5537 3893 5549 3896
rect 5583 3893 5595 3927
rect 5537 3887 5595 3893
rect 5905 3927 5963 3933
rect 5905 3893 5917 3927
rect 5951 3893 5963 3927
rect 5905 3887 5963 3893
rect 5997 3927 6055 3933
rect 5997 3893 6009 3927
rect 6043 3924 6055 3927
rect 6454 3924 6460 3936
rect 6043 3896 6460 3924
rect 6043 3893 6055 3896
rect 5997 3887 6055 3893
rect 6454 3884 6460 3896
rect 6512 3884 6518 3936
rect 7282 3884 7288 3936
rect 7340 3924 7346 3936
rect 8757 3927 8815 3933
rect 8757 3924 8769 3927
rect 7340 3896 8769 3924
rect 7340 3884 7346 3896
rect 8757 3893 8769 3896
rect 8803 3893 8815 3927
rect 8757 3887 8815 3893
rect 8938 3884 8944 3936
rect 8996 3924 9002 3936
rect 9217 3927 9275 3933
rect 9217 3924 9229 3927
rect 8996 3896 9229 3924
rect 8996 3884 9002 3896
rect 9217 3893 9229 3896
rect 9263 3924 9275 3927
rect 9398 3924 9404 3936
rect 9263 3896 9404 3924
rect 9263 3893 9275 3896
rect 9217 3887 9275 3893
rect 9398 3884 9404 3896
rect 9456 3884 9462 3936
rect 9490 3884 9496 3936
rect 9548 3924 9554 3936
rect 9585 3927 9643 3933
rect 9585 3924 9597 3927
rect 9548 3896 9597 3924
rect 9548 3884 9554 3896
rect 9585 3893 9597 3896
rect 9631 3893 9643 3927
rect 9876 3924 9904 3964
rect 9953 3961 9965 3995
rect 9999 3992 10011 3995
rect 10410 3992 10416 4004
rect 9999 3964 10416 3992
rect 9999 3961 10011 3964
rect 9953 3955 10011 3961
rect 10410 3952 10416 3964
rect 10468 3952 10474 4004
rect 10704 3992 10732 4032
rect 10778 4020 10784 4072
rect 10836 4060 10842 4072
rect 10873 4063 10931 4069
rect 10873 4060 10885 4063
rect 10836 4032 10885 4060
rect 10836 4020 10842 4032
rect 10873 4029 10885 4032
rect 10919 4029 10931 4063
rect 11072 4060 11100 4168
rect 11146 4156 11152 4168
rect 11204 4156 11210 4208
rect 11333 4199 11391 4205
rect 11333 4165 11345 4199
rect 11379 4196 11391 4199
rect 11514 4196 11520 4208
rect 11379 4168 11520 4196
rect 11379 4165 11391 4168
rect 11333 4159 11391 4165
rect 11514 4156 11520 4168
rect 11572 4156 11578 4208
rect 11974 4196 11980 4208
rect 11935 4168 11980 4196
rect 11974 4156 11980 4168
rect 12032 4156 12038 4208
rect 12084 4196 12112 4236
rect 12250 4224 12256 4236
rect 12308 4224 12314 4276
rect 12526 4264 12532 4276
rect 12487 4236 12532 4264
rect 12526 4224 12532 4236
rect 12584 4224 12590 4276
rect 12802 4224 12808 4276
rect 12860 4264 12866 4276
rect 12860 4236 12905 4264
rect 12860 4224 12866 4236
rect 13354 4224 13360 4276
rect 13412 4264 13418 4276
rect 13541 4267 13599 4273
rect 13541 4264 13553 4267
rect 13412 4236 13553 4264
rect 13412 4224 13418 4236
rect 13541 4233 13553 4236
rect 13587 4233 13599 4267
rect 13541 4227 13599 4233
rect 13998 4224 14004 4276
rect 14056 4264 14062 4276
rect 14277 4267 14335 4273
rect 14277 4264 14289 4267
rect 14056 4236 14289 4264
rect 14056 4224 14062 4236
rect 14277 4233 14289 4236
rect 14323 4233 14335 4267
rect 14458 4264 14464 4276
rect 14419 4236 14464 4264
rect 14277 4227 14335 4233
rect 14458 4224 14464 4236
rect 14516 4224 14522 4276
rect 12986 4196 12992 4208
rect 12084 4168 12992 4196
rect 12986 4156 12992 4168
rect 13044 4196 13050 4208
rect 13725 4199 13783 4205
rect 13725 4196 13737 4199
rect 13044 4168 13737 4196
rect 13044 4156 13050 4168
rect 13725 4165 13737 4168
rect 13771 4196 13783 4199
rect 13909 4199 13967 4205
rect 13909 4196 13921 4199
rect 13771 4168 13921 4196
rect 13771 4165 13783 4168
rect 13725 4159 13783 4165
rect 13909 4165 13921 4168
rect 13955 4196 13967 4199
rect 14093 4199 14151 4205
rect 14093 4196 14105 4199
rect 13955 4168 14105 4196
rect 13955 4165 13967 4168
rect 13909 4159 13967 4165
rect 14093 4165 14105 4168
rect 14139 4165 14151 4199
rect 14093 4159 14151 4165
rect 14366 4156 14372 4208
rect 14424 4196 14430 4208
rect 14645 4199 14703 4205
rect 14645 4196 14657 4199
rect 14424 4168 14657 4196
rect 14424 4156 14430 4168
rect 14645 4165 14657 4168
rect 14691 4165 14703 4199
rect 14645 4159 14703 4165
rect 11238 4088 11244 4140
rect 11296 4128 11302 4140
rect 12710 4128 12716 4140
rect 11296 4100 12716 4128
rect 11296 4088 11302 4100
rect 12710 4088 12716 4100
rect 12768 4088 12774 4140
rect 13265 4131 13323 4137
rect 13265 4097 13277 4131
rect 13311 4128 13323 4131
rect 13449 4131 13507 4137
rect 13449 4128 13461 4131
rect 13311 4100 13461 4128
rect 13311 4097 13323 4100
rect 13265 4091 13323 4097
rect 13449 4097 13461 4100
rect 13495 4128 13507 4131
rect 13814 4128 13820 4140
rect 13495 4100 13820 4128
rect 13495 4097 13507 4100
rect 13449 4091 13507 4097
rect 13814 4088 13820 4100
rect 13872 4128 13878 4140
rect 15286 4128 15292 4140
rect 13872 4100 15292 4128
rect 13872 4088 13878 4100
rect 15286 4088 15292 4100
rect 15344 4088 15350 4140
rect 11141 4063 11199 4069
rect 11141 4060 11153 4063
rect 11072 4032 11153 4060
rect 10873 4023 10931 4029
rect 11141 4029 11153 4032
rect 11187 4029 11199 4063
rect 11790 4060 11796 4072
rect 11141 4023 11199 4029
rect 11256 4032 11796 4060
rect 11054 3992 11060 4004
rect 10704 3964 11060 3992
rect 11054 3952 11060 3964
rect 11112 3952 11118 4004
rect 10689 3927 10747 3933
rect 10689 3924 10701 3927
rect 9876 3896 10701 3924
rect 9585 3887 9643 3893
rect 10689 3893 10701 3896
rect 10735 3893 10747 3927
rect 10689 3887 10747 3893
rect 10870 3884 10876 3936
rect 10928 3924 10934 3936
rect 11256 3924 11284 4032
rect 11790 4020 11796 4032
rect 11848 4020 11854 4072
rect 12066 4060 12072 4072
rect 12027 4032 12072 4060
rect 12066 4020 12072 4032
rect 12124 4020 12130 4072
rect 12434 4020 12440 4072
rect 12492 4060 12498 4072
rect 15473 4063 15531 4069
rect 15473 4060 15485 4063
rect 12492 4032 15485 4060
rect 12492 4020 12498 4032
rect 15473 4029 15485 4032
rect 15519 4029 15531 4063
rect 15473 4023 15531 4029
rect 12342 3952 12348 4004
rect 12400 3992 12406 4004
rect 12621 3995 12679 4001
rect 12621 3992 12633 3995
rect 12400 3964 12633 3992
rect 12400 3952 12406 3964
rect 12621 3961 12633 3964
rect 12667 3992 12679 3995
rect 12802 3992 12808 4004
rect 12667 3964 12808 3992
rect 12667 3961 12679 3964
rect 12621 3955 12679 3961
rect 12802 3952 12808 3964
rect 12860 3952 12866 4004
rect 12986 3992 12992 4004
rect 12947 3964 12992 3992
rect 12986 3952 12992 3964
rect 13044 3952 13050 4004
rect 10928 3896 11284 3924
rect 10928 3884 10934 3896
rect 11330 3884 11336 3936
rect 11388 3924 11394 3936
rect 11425 3927 11483 3933
rect 11425 3924 11437 3927
rect 11388 3896 11437 3924
rect 11388 3884 11394 3896
rect 11425 3893 11437 3896
rect 11471 3893 11483 3927
rect 11698 3924 11704 3936
rect 11659 3896 11704 3924
rect 11425 3887 11483 3893
rect 11698 3884 11704 3896
rect 11756 3884 11762 3936
rect 15102 3924 15108 3936
rect 15063 3896 15108 3924
rect 15102 3884 15108 3896
rect 15160 3884 15166 3936
rect 15286 3924 15292 3936
rect 15247 3896 15292 3924
rect 15286 3884 15292 3896
rect 15344 3884 15350 3936
rect 15657 3927 15715 3933
rect 15657 3893 15669 3927
rect 15703 3924 15715 3927
rect 16206 3924 16212 3936
rect 15703 3896 16212 3924
rect 15703 3893 15715 3896
rect 15657 3887 15715 3893
rect 16206 3884 16212 3896
rect 16264 3884 16270 3936
rect 1104 3834 16008 3856
rect 1104 3782 5979 3834
rect 6031 3782 6043 3834
rect 6095 3782 6107 3834
rect 6159 3782 6171 3834
rect 6223 3782 10976 3834
rect 11028 3782 11040 3834
rect 11092 3782 11104 3834
rect 11156 3782 11168 3834
rect 11220 3782 16008 3834
rect 1104 3760 16008 3782
rect 2133 3723 2191 3729
rect 2133 3720 2145 3723
rect 1964 3692 2145 3720
rect 1964 3661 1992 3692
rect 2133 3689 2145 3692
rect 2179 3689 2191 3723
rect 2133 3683 2191 3689
rect 2332 3692 2774 3720
rect 1949 3655 2007 3661
rect 1949 3621 1961 3655
rect 1995 3621 2007 3655
rect 1949 3615 2007 3621
rect 2332 3593 2360 3692
rect 2746 3652 2774 3692
rect 3142 3680 3148 3732
rect 3200 3720 3206 3732
rect 3881 3723 3939 3729
rect 3881 3720 3893 3723
rect 3200 3692 3893 3720
rect 3200 3680 3206 3692
rect 3881 3689 3893 3692
rect 3927 3689 3939 3723
rect 3881 3683 3939 3689
rect 4246 3680 4252 3732
rect 4304 3720 4310 3732
rect 4341 3723 4399 3729
rect 4341 3720 4353 3723
rect 4304 3692 4353 3720
rect 4304 3680 4310 3692
rect 4341 3689 4353 3692
rect 4387 3689 4399 3723
rect 4341 3683 4399 3689
rect 4709 3723 4767 3729
rect 4709 3689 4721 3723
rect 4755 3689 4767 3723
rect 4709 3683 4767 3689
rect 5169 3723 5227 3729
rect 5169 3689 5181 3723
rect 5215 3720 5227 3723
rect 5258 3720 5264 3732
rect 5215 3692 5264 3720
rect 5215 3689 5227 3692
rect 5169 3683 5227 3689
rect 4724 3652 4752 3683
rect 5258 3680 5264 3692
rect 5316 3680 5322 3732
rect 5350 3680 5356 3732
rect 5408 3720 5414 3732
rect 5813 3723 5871 3729
rect 5813 3720 5825 3723
rect 5408 3692 5825 3720
rect 5408 3680 5414 3692
rect 5813 3689 5825 3692
rect 5859 3689 5871 3723
rect 5813 3683 5871 3689
rect 7009 3723 7067 3729
rect 7009 3689 7021 3723
rect 7055 3720 7067 3723
rect 7466 3720 7472 3732
rect 7055 3692 7472 3720
rect 7055 3689 7067 3692
rect 7009 3683 7067 3689
rect 7466 3680 7472 3692
rect 7524 3680 7530 3732
rect 7837 3723 7895 3729
rect 7837 3689 7849 3723
rect 7883 3720 7895 3723
rect 8018 3720 8024 3732
rect 7883 3692 8024 3720
rect 7883 3689 7895 3692
rect 7837 3683 7895 3689
rect 8018 3680 8024 3692
rect 8076 3680 8082 3732
rect 8386 3680 8392 3732
rect 8444 3720 8450 3732
rect 10689 3723 10747 3729
rect 8444 3692 10640 3720
rect 8444 3680 8450 3692
rect 6454 3652 6460 3664
rect 2746 3624 4752 3652
rect 4908 3624 6460 3652
rect 1581 3587 1639 3593
rect 1581 3553 1593 3587
rect 1627 3553 1639 3587
rect 1581 3547 1639 3553
rect 2317 3587 2375 3593
rect 2317 3553 2329 3587
rect 2363 3553 2375 3587
rect 2317 3547 2375 3553
rect 1596 3516 1624 3547
rect 2498 3544 2504 3596
rect 2556 3584 2562 3596
rect 2593 3587 2651 3593
rect 2593 3584 2605 3587
rect 2556 3556 2605 3584
rect 2556 3544 2562 3556
rect 2593 3553 2605 3556
rect 2639 3553 2651 3587
rect 2593 3547 2651 3553
rect 2682 3544 2688 3596
rect 2740 3584 2746 3596
rect 2869 3587 2927 3593
rect 2869 3584 2881 3587
rect 2740 3556 2881 3584
rect 2740 3544 2746 3556
rect 2869 3553 2881 3556
rect 2915 3553 2927 3587
rect 2869 3547 2927 3553
rect 3145 3587 3203 3593
rect 3145 3553 3157 3587
rect 3191 3584 3203 3587
rect 3326 3584 3332 3596
rect 3191 3556 3332 3584
rect 3191 3553 3203 3556
rect 3145 3547 3203 3553
rect 3326 3544 3332 3556
rect 3384 3544 3390 3596
rect 3418 3544 3424 3596
rect 3476 3584 3482 3596
rect 3694 3584 3700 3596
rect 3476 3556 3521 3584
rect 3655 3556 3700 3584
rect 3476 3544 3482 3556
rect 3694 3544 3700 3556
rect 3752 3544 3758 3596
rect 4249 3587 4307 3593
rect 4249 3553 4261 3587
rect 4295 3584 4307 3587
rect 4908 3584 4936 3624
rect 6454 3612 6460 3624
rect 6512 3612 6518 3664
rect 6638 3612 6644 3664
rect 6696 3652 6702 3664
rect 8297 3655 8355 3661
rect 8297 3652 8309 3655
rect 6696 3624 8309 3652
rect 6696 3612 6702 3624
rect 8297 3621 8309 3624
rect 8343 3621 8355 3655
rect 8297 3615 8355 3621
rect 9585 3655 9643 3661
rect 9585 3621 9597 3655
rect 9631 3652 9643 3655
rect 9674 3652 9680 3664
rect 9631 3624 9680 3652
rect 9631 3621 9643 3624
rect 9585 3615 9643 3621
rect 9674 3612 9680 3624
rect 9732 3612 9738 3664
rect 10410 3652 10416 3664
rect 10244 3624 10416 3652
rect 5074 3584 5080 3596
rect 4295 3556 4936 3584
rect 5035 3556 5080 3584
rect 4295 3553 4307 3556
rect 4249 3547 4307 3553
rect 5074 3544 5080 3556
rect 5132 3544 5138 3596
rect 5166 3544 5172 3596
rect 5224 3584 5230 3596
rect 5721 3587 5779 3593
rect 5224 3556 5672 3584
rect 5224 3544 5230 3556
rect 1596 3488 3280 3516
rect 1118 3408 1124 3460
rect 1176 3448 1182 3460
rect 1397 3451 1455 3457
rect 1397 3448 1409 3451
rect 1176 3420 1409 3448
rect 1176 3408 1182 3420
rect 1397 3417 1409 3420
rect 1443 3417 1455 3451
rect 1397 3411 1455 3417
rect 1578 3408 1584 3460
rect 1636 3448 1642 3460
rect 3252 3457 3280 3488
rect 3602 3476 3608 3528
rect 3660 3516 3666 3528
rect 4338 3516 4344 3528
rect 3660 3488 4344 3516
rect 3660 3476 3666 3488
rect 4338 3476 4344 3488
rect 4396 3476 4402 3528
rect 4522 3516 4528 3528
rect 4483 3488 4528 3516
rect 4522 3476 4528 3488
rect 4580 3476 4586 3528
rect 4890 3476 4896 3528
rect 4948 3516 4954 3528
rect 5261 3519 5319 3525
rect 5261 3516 5273 3519
rect 4948 3488 5273 3516
rect 4948 3476 4954 3488
rect 5261 3485 5273 3488
rect 5307 3485 5319 3519
rect 5644 3516 5672 3556
rect 5721 3553 5733 3587
rect 5767 3584 5779 3587
rect 5902 3584 5908 3596
rect 5767 3556 5908 3584
rect 5767 3553 5779 3556
rect 5721 3547 5779 3553
rect 5902 3544 5908 3556
rect 5960 3544 5966 3596
rect 6181 3587 6239 3593
rect 6181 3553 6193 3587
rect 6227 3584 6239 3587
rect 7742 3584 7748 3596
rect 6227 3556 7748 3584
rect 6227 3553 6239 3556
rect 6181 3547 6239 3553
rect 6196 3516 6224 3547
rect 7742 3544 7748 3556
rect 7800 3544 7806 3596
rect 8481 3587 8539 3593
rect 8481 3553 8493 3587
rect 8527 3584 8539 3587
rect 9398 3584 9404 3596
rect 8527 3556 9404 3584
rect 8527 3553 8539 3556
rect 8481 3547 8539 3553
rect 9398 3544 9404 3556
rect 9456 3544 9462 3596
rect 9490 3544 9496 3596
rect 9548 3584 9554 3596
rect 9548 3556 9593 3584
rect 9548 3544 9554 3556
rect 9858 3544 9864 3596
rect 9916 3584 9922 3596
rect 10244 3593 10272 3624
rect 10410 3612 10416 3624
rect 10468 3612 10474 3664
rect 10612 3652 10640 3692
rect 10689 3689 10701 3723
rect 10735 3720 10747 3723
rect 10778 3720 10784 3732
rect 10735 3692 10784 3720
rect 10735 3689 10747 3692
rect 10689 3683 10747 3689
rect 10778 3680 10784 3692
rect 10836 3680 10842 3732
rect 10870 3680 10876 3732
rect 10928 3720 10934 3732
rect 11057 3723 11115 3729
rect 11057 3720 11069 3723
rect 10928 3692 11069 3720
rect 10928 3680 10934 3692
rect 11057 3689 11069 3692
rect 11103 3689 11115 3723
rect 11057 3683 11115 3689
rect 11514 3680 11520 3732
rect 11572 3720 11578 3732
rect 11701 3723 11759 3729
rect 11701 3720 11713 3723
rect 11572 3692 11713 3720
rect 11572 3680 11578 3692
rect 11701 3689 11713 3692
rect 11747 3689 11759 3723
rect 12250 3720 12256 3732
rect 11701 3683 11759 3689
rect 11900 3692 12256 3720
rect 11609 3655 11667 3661
rect 10612 3624 10824 3652
rect 10137 3587 10195 3593
rect 10137 3584 10149 3587
rect 9916 3556 10149 3584
rect 9916 3544 9922 3556
rect 10137 3553 10149 3556
rect 10183 3553 10195 3587
rect 10137 3547 10195 3553
rect 10229 3587 10287 3593
rect 10229 3553 10241 3587
rect 10275 3553 10287 3587
rect 10502 3584 10508 3596
rect 10463 3556 10508 3584
rect 10229 3547 10287 3553
rect 10502 3544 10508 3556
rect 10560 3544 10566 3596
rect 10796 3593 10824 3624
rect 11609 3621 11621 3655
rect 11655 3652 11667 3655
rect 11790 3652 11796 3664
rect 11655 3624 11796 3652
rect 11655 3621 11667 3624
rect 11609 3615 11667 3621
rect 11790 3612 11796 3624
rect 11848 3612 11854 3664
rect 11900 3593 11928 3692
rect 12250 3680 12256 3692
rect 12308 3680 12314 3732
rect 13078 3680 13084 3732
rect 13136 3720 13142 3732
rect 14642 3720 14648 3732
rect 13136 3692 14648 3720
rect 13136 3680 13142 3692
rect 14642 3680 14648 3692
rect 14700 3720 14706 3732
rect 15105 3723 15163 3729
rect 15105 3720 15117 3723
rect 14700 3692 15117 3720
rect 14700 3680 14706 3692
rect 15105 3689 15117 3692
rect 15151 3689 15163 3723
rect 15105 3683 15163 3689
rect 12161 3655 12219 3661
rect 12161 3621 12173 3655
rect 12207 3652 12219 3655
rect 12434 3652 12440 3664
rect 12207 3624 12440 3652
rect 12207 3621 12219 3624
rect 12161 3615 12219 3621
rect 12434 3612 12440 3624
rect 12492 3612 12498 3664
rect 13262 3612 13268 3664
rect 13320 3652 13326 3664
rect 13909 3655 13967 3661
rect 13909 3652 13921 3655
rect 13320 3624 13921 3652
rect 13320 3612 13326 3624
rect 13909 3621 13921 3624
rect 13955 3621 13967 3655
rect 13909 3615 13967 3621
rect 13998 3612 14004 3664
rect 14056 3652 14062 3664
rect 15473 3655 15531 3661
rect 15473 3652 15485 3655
rect 14056 3624 15485 3652
rect 14056 3612 14062 3624
rect 15473 3621 15485 3624
rect 15519 3621 15531 3655
rect 15473 3615 15531 3621
rect 10781 3587 10839 3593
rect 10781 3553 10793 3587
rect 10827 3584 10839 3587
rect 11232 3587 11290 3593
rect 10827 3556 11017 3584
rect 10827 3553 10839 3556
rect 10781 3547 10839 3553
rect 5644 3488 6224 3516
rect 6273 3519 6331 3525
rect 5261 3479 5319 3485
rect 6273 3485 6285 3519
rect 6319 3485 6331 3519
rect 6273 3479 6331 3485
rect 2685 3451 2743 3457
rect 2685 3448 2697 3451
rect 1636 3420 2697 3448
rect 1636 3408 1642 3420
rect 2685 3417 2697 3420
rect 2731 3417 2743 3451
rect 2685 3411 2743 3417
rect 3237 3451 3295 3457
rect 3237 3417 3249 3451
rect 3283 3417 3295 3451
rect 3237 3411 3295 3417
rect 3326 3408 3332 3460
rect 3384 3448 3390 3460
rect 5537 3451 5595 3457
rect 5537 3448 5549 3451
rect 3384 3420 5549 3448
rect 3384 3408 3390 3420
rect 5537 3417 5549 3420
rect 5583 3417 5595 3451
rect 5537 3411 5595 3417
rect 5718 3408 5724 3460
rect 5776 3448 5782 3460
rect 6288 3448 6316 3479
rect 6362 3476 6368 3528
rect 6420 3516 6426 3528
rect 6733 3519 6791 3525
rect 6733 3516 6745 3519
rect 6420 3488 6745 3516
rect 6420 3476 6426 3488
rect 6733 3485 6745 3488
rect 6779 3485 6791 3519
rect 6733 3479 6791 3485
rect 6917 3519 6975 3525
rect 6917 3485 6929 3519
rect 6963 3516 6975 3519
rect 7650 3516 7656 3528
rect 6963 3488 7656 3516
rect 6963 3485 6975 3488
rect 6917 3479 6975 3485
rect 7650 3476 7656 3488
rect 7708 3476 7714 3528
rect 7926 3516 7932 3528
rect 7887 3488 7932 3516
rect 7926 3476 7932 3488
rect 7984 3476 7990 3528
rect 8110 3516 8116 3528
rect 8071 3488 8116 3516
rect 8110 3476 8116 3488
rect 8168 3476 8174 3528
rect 8202 3476 8208 3528
rect 8260 3516 8266 3528
rect 8665 3519 8723 3525
rect 8665 3516 8677 3519
rect 8260 3488 8677 3516
rect 8260 3476 8266 3488
rect 8665 3485 8677 3488
rect 8711 3485 8723 3519
rect 8665 3479 8723 3485
rect 8754 3476 8760 3528
rect 8812 3516 8818 3528
rect 9214 3516 9220 3528
rect 8812 3488 9220 3516
rect 8812 3476 8818 3488
rect 9214 3476 9220 3488
rect 9272 3476 9278 3528
rect 9766 3516 9772 3528
rect 9727 3488 9772 3516
rect 9766 3476 9772 3488
rect 9824 3476 9830 3528
rect 10989 3516 11017 3556
rect 11232 3553 11244 3587
rect 11278 3584 11290 3587
rect 11885 3587 11943 3593
rect 11278 3556 11836 3584
rect 11278 3553 11290 3556
rect 11232 3547 11290 3553
rect 11698 3516 11704 3528
rect 10989 3488 11704 3516
rect 11698 3476 11704 3488
rect 11756 3476 11762 3528
rect 11808 3516 11836 3556
rect 11885 3553 11897 3587
rect 11931 3553 11943 3587
rect 11885 3547 11943 3553
rect 12066 3544 12072 3596
rect 12124 3584 12130 3596
rect 12250 3584 12256 3596
rect 12124 3556 12256 3584
rect 12124 3544 12130 3556
rect 12250 3544 12256 3556
rect 12308 3544 12314 3596
rect 13354 3584 13360 3596
rect 13315 3556 13360 3584
rect 13354 3544 13360 3556
rect 13412 3584 13418 3596
rect 13541 3587 13599 3593
rect 13541 3584 13553 3587
rect 13412 3556 13553 3584
rect 13412 3544 13418 3556
rect 13541 3553 13553 3556
rect 13587 3553 13599 3587
rect 13814 3584 13820 3596
rect 13775 3556 13820 3584
rect 13541 3547 13599 3553
rect 13814 3544 13820 3556
rect 13872 3544 13878 3596
rect 14458 3544 14464 3596
rect 14516 3584 14522 3596
rect 14737 3587 14795 3593
rect 14737 3584 14749 3587
rect 14516 3556 14749 3584
rect 14516 3544 14522 3556
rect 14737 3553 14749 3556
rect 14783 3553 14795 3587
rect 14737 3547 14795 3553
rect 14826 3544 14832 3596
rect 14884 3584 14890 3596
rect 15102 3584 15108 3596
rect 14884 3556 15108 3584
rect 14884 3544 14890 3556
rect 15102 3544 15108 3556
rect 15160 3544 15166 3596
rect 15286 3584 15292 3596
rect 15247 3556 15292 3584
rect 15286 3544 15292 3556
rect 15344 3544 15350 3596
rect 12084 3516 12112 3544
rect 11808 3488 12112 3516
rect 12434 3476 12440 3528
rect 12492 3476 12498 3528
rect 12897 3519 12955 3525
rect 12897 3485 12909 3519
rect 12943 3516 12955 3519
rect 12986 3516 12992 3528
rect 12943 3488 12992 3516
rect 12943 3485 12955 3488
rect 12897 3479 12955 3485
rect 12986 3476 12992 3488
rect 13044 3476 13050 3528
rect 7006 3448 7012 3460
rect 5776 3420 7012 3448
rect 5776 3408 5782 3420
rect 7006 3408 7012 3420
rect 7064 3408 7070 3460
rect 7374 3448 7380 3460
rect 7335 3420 7380 3448
rect 7374 3408 7380 3420
rect 7432 3408 7438 3460
rect 9953 3451 10011 3457
rect 9953 3448 9965 3451
rect 8128 3420 9965 3448
rect 8128 3392 8156 3420
rect 9953 3417 9965 3420
rect 9999 3417 10011 3451
rect 9953 3411 10011 3417
rect 10042 3408 10048 3460
rect 10100 3448 10106 3460
rect 10502 3448 10508 3460
rect 10100 3420 10508 3448
rect 10100 3408 10106 3420
rect 10502 3408 10508 3420
rect 10560 3408 10566 3460
rect 11333 3451 11391 3457
rect 11333 3448 11345 3451
rect 10704 3420 11345 3448
rect 1854 3380 1860 3392
rect 1815 3352 1860 3380
rect 1854 3340 1860 3352
rect 1912 3340 1918 3392
rect 2406 3380 2412 3392
rect 2367 3352 2412 3380
rect 2406 3340 2412 3352
rect 2464 3340 2470 3392
rect 2590 3340 2596 3392
rect 2648 3380 2654 3392
rect 2961 3383 3019 3389
rect 2961 3380 2973 3383
rect 2648 3352 2973 3380
rect 2648 3340 2654 3352
rect 2961 3349 2973 3352
rect 3007 3349 3019 3383
rect 2961 3343 3019 3349
rect 3050 3340 3056 3392
rect 3108 3380 3114 3392
rect 3513 3383 3571 3389
rect 3513 3380 3525 3383
rect 3108 3352 3525 3380
rect 3108 3340 3114 3352
rect 3513 3349 3525 3352
rect 3559 3349 3571 3383
rect 3513 3343 3571 3349
rect 4062 3340 4068 3392
rect 4120 3380 4126 3392
rect 5626 3380 5632 3392
rect 4120 3352 5632 3380
rect 4120 3340 4126 3352
rect 5626 3340 5632 3352
rect 5684 3340 5690 3392
rect 6270 3340 6276 3392
rect 6328 3380 6334 3392
rect 7469 3383 7527 3389
rect 7469 3380 7481 3383
rect 6328 3352 7481 3380
rect 6328 3340 6334 3352
rect 7469 3349 7481 3352
rect 7515 3349 7527 3383
rect 7469 3343 7527 3349
rect 8110 3340 8116 3392
rect 8168 3340 8174 3392
rect 9122 3380 9128 3392
rect 9083 3352 9128 3380
rect 9122 3340 9128 3352
rect 9180 3340 9186 3392
rect 10410 3380 10416 3392
rect 10371 3352 10416 3380
rect 10410 3340 10416 3352
rect 10468 3340 10474 3392
rect 10594 3340 10600 3392
rect 10652 3380 10658 3392
rect 10704 3380 10732 3420
rect 11333 3417 11345 3420
rect 11379 3417 11391 3451
rect 11333 3411 11391 3417
rect 11422 3408 11428 3460
rect 11480 3448 11486 3460
rect 12452 3448 12480 3476
rect 14093 3451 14151 3457
rect 14093 3448 14105 3451
rect 11480 3420 12480 3448
rect 12912 3420 14105 3448
rect 11480 3408 11486 3420
rect 12912 3392 12940 3420
rect 14093 3417 14105 3420
rect 14139 3417 14151 3451
rect 14550 3448 14556 3460
rect 14511 3420 14556 3448
rect 14093 3411 14151 3417
rect 14550 3408 14556 3420
rect 14608 3408 14614 3460
rect 15010 3448 15016 3460
rect 14971 3420 15016 3448
rect 15010 3408 15016 3420
rect 15068 3408 15074 3460
rect 15654 3448 15660 3460
rect 15615 3420 15660 3448
rect 15654 3408 15660 3420
rect 15712 3408 15718 3460
rect 10652 3352 10732 3380
rect 10652 3340 10658 3352
rect 10778 3340 10784 3392
rect 10836 3380 10842 3392
rect 10965 3383 11023 3389
rect 10965 3380 10977 3383
rect 10836 3352 10977 3380
rect 10836 3340 10842 3352
rect 10965 3349 10977 3352
rect 11011 3349 11023 3383
rect 10965 3343 11023 3349
rect 11054 3340 11060 3392
rect 11112 3380 11118 3392
rect 11606 3380 11612 3392
rect 11112 3352 11612 3380
rect 11112 3340 11118 3352
rect 11606 3340 11612 3352
rect 11664 3340 11670 3392
rect 11974 3340 11980 3392
rect 12032 3380 12038 3392
rect 12437 3383 12495 3389
rect 12437 3380 12449 3383
rect 12032 3352 12449 3380
rect 12032 3340 12038 3352
rect 12437 3349 12449 3352
rect 12483 3349 12495 3383
rect 12618 3380 12624 3392
rect 12579 3352 12624 3380
rect 12437 3343 12495 3349
rect 12618 3340 12624 3352
rect 12676 3340 12682 3392
rect 12894 3340 12900 3392
rect 12952 3340 12958 3392
rect 13078 3380 13084 3392
rect 13039 3352 13084 3380
rect 13078 3340 13084 3352
rect 13136 3380 13142 3392
rect 13173 3383 13231 3389
rect 13173 3380 13185 3383
rect 13136 3352 13185 3380
rect 13136 3340 13142 3352
rect 13173 3349 13185 3352
rect 13219 3349 13231 3383
rect 14458 3380 14464 3392
rect 14419 3352 14464 3380
rect 13173 3343 13231 3349
rect 14458 3340 14464 3352
rect 14516 3340 14522 3392
rect 1104 3290 16008 3312
rect 1104 3238 3480 3290
rect 3532 3238 3544 3290
rect 3596 3238 3608 3290
rect 3660 3238 3672 3290
rect 3724 3238 8478 3290
rect 8530 3238 8542 3290
rect 8594 3238 8606 3290
rect 8658 3238 8670 3290
rect 8722 3238 13475 3290
rect 13527 3238 13539 3290
rect 13591 3238 13603 3290
rect 13655 3238 13667 3290
rect 13719 3238 16008 3290
rect 1104 3216 16008 3238
rect 2682 3136 2688 3188
rect 2740 3176 2746 3188
rect 4709 3179 4767 3185
rect 4709 3176 4721 3179
rect 2740 3148 4721 3176
rect 2740 3136 2746 3148
rect 4709 3145 4721 3148
rect 4755 3145 4767 3179
rect 4709 3139 4767 3145
rect 5074 3136 5080 3188
rect 5132 3176 5138 3188
rect 6457 3179 6515 3185
rect 6457 3176 6469 3179
rect 5132 3148 6469 3176
rect 5132 3136 5138 3148
rect 6457 3145 6469 3148
rect 6503 3145 6515 3179
rect 7285 3179 7343 3185
rect 7285 3176 7297 3179
rect 6457 3139 6515 3145
rect 6564 3148 7297 3176
rect 1394 3068 1400 3120
rect 1452 3108 1458 3120
rect 2133 3111 2191 3117
rect 2133 3108 2145 3111
rect 1452 3080 2145 3108
rect 1452 3068 1458 3080
rect 2133 3077 2145 3080
rect 2179 3077 2191 3111
rect 2133 3071 2191 3077
rect 2498 3068 2504 3120
rect 2556 3108 2562 3120
rect 3237 3111 3295 3117
rect 3237 3108 3249 3111
rect 2556 3080 3249 3108
rect 2556 3068 2562 3080
rect 3237 3077 3249 3080
rect 3283 3077 3295 3111
rect 3237 3071 3295 3077
rect 5537 3111 5595 3117
rect 5537 3077 5549 3111
rect 5583 3077 5595 3111
rect 6564 3108 6592 3148
rect 7285 3145 7297 3148
rect 7331 3145 7343 3179
rect 7285 3139 7343 3145
rect 8018 3136 8024 3188
rect 8076 3176 8082 3188
rect 9033 3179 9091 3185
rect 8076 3148 8708 3176
rect 8076 3136 8082 3148
rect 8478 3108 8484 3120
rect 5537 3071 5595 3077
rect 5644 3080 6592 3108
rect 7760 3080 8484 3108
rect 2590 3040 2596 3052
rect 1964 3012 2596 3040
rect 1578 2972 1584 2984
rect 1539 2944 1584 2972
rect 1578 2932 1584 2944
rect 1636 2932 1642 2984
rect 1964 2981 1992 3012
rect 2590 3000 2596 3012
rect 2648 3000 2654 3052
rect 2774 3000 2780 3052
rect 2832 3040 2838 3052
rect 3605 3043 3663 3049
rect 3605 3040 3617 3043
rect 2832 3012 3617 3040
rect 2832 3000 2838 3012
rect 3605 3009 3617 3012
rect 3651 3009 3663 3043
rect 3605 3003 3663 3009
rect 4982 3000 4988 3052
rect 5040 3040 5046 3052
rect 5261 3043 5319 3049
rect 5261 3040 5273 3043
rect 5040 3012 5273 3040
rect 5040 3000 5046 3012
rect 5261 3009 5273 3012
rect 5307 3009 5319 3043
rect 5261 3003 5319 3009
rect 5552 2984 5580 3071
rect 1949 2975 2007 2981
rect 1949 2941 1961 2975
rect 1995 2941 2007 2975
rect 1949 2935 2007 2941
rect 2222 2932 2228 2984
rect 2280 2972 2286 2984
rect 2317 2975 2375 2981
rect 2317 2972 2329 2975
rect 2280 2944 2329 2972
rect 2280 2932 2286 2944
rect 2317 2941 2329 2944
rect 2363 2941 2375 2975
rect 2317 2935 2375 2941
rect 2685 2975 2743 2981
rect 2685 2941 2697 2975
rect 2731 2972 2743 2975
rect 2958 2972 2964 2984
rect 2731 2944 2964 2972
rect 2731 2941 2743 2944
rect 2685 2935 2743 2941
rect 2958 2932 2964 2944
rect 3016 2932 3022 2984
rect 3142 2932 3148 2984
rect 3200 2972 3206 2984
rect 3973 2975 4031 2981
rect 3973 2972 3985 2975
rect 3200 2944 3985 2972
rect 3200 2932 3206 2944
rect 3973 2941 3985 2944
rect 4019 2941 4031 2975
rect 3973 2935 4031 2941
rect 4157 2975 4215 2981
rect 4157 2941 4169 2975
rect 4203 2972 4215 2975
rect 4338 2972 4344 2984
rect 4203 2944 4344 2972
rect 4203 2941 4215 2944
rect 4157 2935 4215 2941
rect 4338 2932 4344 2944
rect 4396 2932 4402 2984
rect 4433 2975 4491 2981
rect 4433 2941 4445 2975
rect 4479 2972 4491 2975
rect 4522 2972 4528 2984
rect 4479 2944 4528 2972
rect 4479 2941 4491 2944
rect 4433 2935 4491 2941
rect 4522 2932 4528 2944
rect 4580 2932 4586 2984
rect 4798 2932 4804 2984
rect 4856 2972 4862 2984
rect 4856 2944 5488 2972
rect 4856 2932 4862 2944
rect 382 2864 388 2916
rect 440 2904 446 2916
rect 1397 2907 1455 2913
rect 1397 2904 1409 2907
rect 440 2876 1409 2904
rect 440 2864 446 2876
rect 1397 2873 1409 2876
rect 1443 2873 1455 2907
rect 1397 2867 1455 2873
rect 1762 2864 1768 2916
rect 1820 2904 1826 2916
rect 1820 2876 1992 2904
rect 1820 2864 1826 2876
rect 750 2796 756 2848
rect 808 2836 814 2848
rect 1857 2839 1915 2845
rect 1857 2836 1869 2839
rect 808 2808 1869 2836
rect 808 2796 814 2808
rect 1857 2805 1869 2808
rect 1903 2805 1915 2839
rect 1964 2836 1992 2876
rect 2130 2864 2136 2916
rect 2188 2904 2194 2916
rect 2869 2907 2927 2913
rect 2869 2904 2881 2907
rect 2188 2876 2881 2904
rect 2188 2864 2194 2876
rect 2869 2873 2881 2876
rect 2915 2873 2927 2907
rect 2869 2867 2927 2873
rect 3053 2907 3111 2913
rect 3053 2873 3065 2907
rect 3099 2904 3111 2907
rect 3326 2904 3332 2916
rect 3099 2876 3332 2904
rect 3099 2873 3111 2876
rect 3053 2867 3111 2873
rect 3326 2864 3332 2876
rect 3384 2864 3390 2916
rect 3421 2907 3479 2913
rect 3421 2873 3433 2907
rect 3467 2904 3479 2907
rect 3694 2904 3700 2916
rect 3467 2876 3700 2904
rect 3467 2873 3479 2876
rect 3421 2867 3479 2873
rect 3694 2864 3700 2876
rect 3752 2864 3758 2916
rect 3789 2907 3847 2913
rect 3789 2873 3801 2907
rect 3835 2904 3847 2907
rect 3878 2904 3884 2916
rect 3835 2876 3884 2904
rect 3835 2873 3847 2876
rect 3789 2867 3847 2873
rect 3878 2864 3884 2876
rect 3936 2864 3942 2916
rect 4617 2907 4675 2913
rect 4617 2873 4629 2907
rect 4663 2904 4675 2907
rect 4890 2904 4896 2916
rect 4663 2876 4896 2904
rect 4663 2873 4675 2876
rect 4617 2867 4675 2873
rect 4890 2864 4896 2876
rect 4948 2864 4954 2916
rect 5074 2904 5080 2916
rect 5035 2876 5080 2904
rect 5074 2864 5080 2876
rect 5132 2864 5138 2916
rect 5166 2864 5172 2916
rect 5224 2904 5230 2916
rect 5460 2904 5488 2944
rect 5534 2932 5540 2984
rect 5592 2932 5598 2984
rect 5644 2904 5672 3080
rect 6178 3040 6184 3052
rect 6139 3012 6184 3040
rect 6178 3000 6184 3012
rect 6236 3000 6242 3052
rect 6270 3000 6276 3052
rect 6328 3040 6334 3052
rect 7760 3049 7788 3080
rect 8478 3068 8484 3080
rect 8536 3068 8542 3120
rect 6917 3043 6975 3049
rect 6917 3040 6929 3043
rect 6328 3012 6929 3040
rect 6328 3000 6334 3012
rect 6917 3009 6929 3012
rect 6963 3009 6975 3043
rect 6917 3003 6975 3009
rect 7009 3043 7067 3049
rect 7009 3009 7021 3043
rect 7055 3009 7067 3043
rect 7009 3003 7067 3009
rect 7745 3043 7803 3049
rect 7745 3009 7757 3043
rect 7791 3009 7803 3043
rect 7745 3003 7803 3009
rect 5810 2932 5816 2984
rect 5868 2972 5874 2984
rect 5905 2975 5963 2981
rect 5905 2972 5917 2975
rect 5868 2944 5917 2972
rect 5868 2932 5874 2944
rect 5905 2941 5917 2944
rect 5951 2941 5963 2975
rect 6822 2972 6828 2984
rect 6783 2944 6828 2972
rect 5905 2935 5963 2941
rect 6822 2932 6828 2944
rect 6880 2932 6886 2984
rect 6362 2904 6368 2916
rect 5224 2876 5269 2904
rect 5460 2876 5672 2904
rect 5920 2876 6368 2904
rect 5224 2864 5230 2876
rect 2593 2839 2651 2845
rect 2593 2836 2605 2839
rect 1964 2808 2605 2836
rect 1857 2799 1915 2805
rect 2593 2805 2605 2808
rect 2639 2805 2651 2839
rect 2593 2799 2651 2805
rect 4062 2796 4068 2848
rect 4120 2836 4126 2848
rect 5920 2836 5948 2876
rect 6362 2864 6368 2876
rect 6420 2864 6426 2916
rect 6730 2864 6736 2916
rect 6788 2904 6794 2916
rect 7024 2904 7052 3003
rect 7834 3000 7840 3052
rect 7892 3040 7898 3052
rect 7892 3012 7937 3040
rect 7892 3000 7898 3012
rect 8018 3000 8024 3052
rect 8076 3040 8082 3052
rect 8680 3049 8708 3148
rect 9033 3145 9045 3179
rect 9079 3176 9091 3179
rect 9306 3176 9312 3188
rect 9079 3148 9312 3176
rect 9079 3145 9091 3148
rect 9033 3139 9091 3145
rect 9306 3136 9312 3148
rect 9364 3136 9370 3188
rect 9398 3136 9404 3188
rect 9456 3176 9462 3188
rect 10781 3179 10839 3185
rect 10781 3176 10793 3179
rect 9456 3148 10793 3176
rect 9456 3136 9462 3148
rect 10781 3145 10793 3148
rect 10827 3145 10839 3179
rect 10781 3139 10839 3145
rect 10888 3148 11184 3176
rect 8754 3068 8760 3120
rect 8812 3108 8818 3120
rect 9674 3108 9680 3120
rect 8812 3080 9680 3108
rect 8812 3068 8818 3080
rect 9646 3068 9680 3080
rect 9732 3068 9738 3120
rect 10888 3108 10916 3148
rect 11054 3108 11060 3120
rect 10529 3080 10916 3108
rect 10980 3080 11060 3108
rect 8665 3043 8723 3049
rect 8076 3012 8524 3040
rect 8076 3000 8082 3012
rect 7653 2975 7711 2981
rect 7653 2941 7665 2975
rect 7699 2972 7711 2975
rect 8202 2972 8208 2984
rect 7699 2944 8208 2972
rect 7699 2941 7711 2944
rect 7653 2935 7711 2941
rect 8202 2932 8208 2944
rect 8260 2932 8266 2984
rect 8496 2981 8524 3012
rect 8665 3009 8677 3043
rect 8711 3009 8723 3043
rect 8938 3040 8944 3052
rect 8665 3003 8723 3009
rect 8864 3012 8944 3040
rect 8481 2975 8539 2981
rect 8481 2941 8493 2975
rect 8527 2972 8539 2975
rect 8864 2972 8892 3012
rect 8938 3000 8944 3012
rect 8996 3000 9002 3052
rect 9030 3000 9036 3052
rect 9088 3040 9094 3052
rect 9309 3043 9367 3049
rect 9309 3040 9321 3043
rect 9088 3012 9321 3040
rect 9088 3000 9094 3012
rect 9309 3009 9321 3012
rect 9355 3009 9367 3043
rect 9646 3040 9674 3068
rect 10529 3040 10557 3080
rect 10980 3040 11008 3080
rect 11054 3068 11060 3080
rect 11112 3068 11118 3120
rect 9646 3012 10557 3040
rect 10888 3012 11008 3040
rect 11156 3040 11184 3148
rect 11440 3148 11744 3176
rect 11333 3111 11391 3117
rect 11333 3077 11345 3111
rect 11379 3108 11391 3111
rect 11440 3108 11468 3148
rect 11379 3080 11468 3108
rect 11379 3077 11391 3080
rect 11333 3071 11391 3077
rect 11606 3040 11612 3052
rect 11156 3012 11612 3040
rect 9309 3003 9367 3009
rect 9125 2975 9183 2981
rect 9125 2972 9137 2975
rect 8527 2944 8892 2972
rect 8956 2944 9137 2972
rect 8527 2941 8539 2944
rect 8481 2935 8539 2941
rect 8956 2916 8984 2944
rect 9125 2941 9137 2944
rect 9171 2972 9183 2975
rect 9766 2972 9772 2984
rect 9171 2944 9772 2972
rect 9171 2941 9183 2944
rect 9125 2935 9183 2941
rect 9766 2932 9772 2944
rect 9824 2932 9830 2984
rect 9858 2932 9864 2984
rect 9916 2972 9922 2984
rect 10152 2981 10180 3012
rect 10137 2975 10195 2981
rect 9916 2944 9961 2972
rect 9916 2932 9922 2944
rect 10137 2941 10149 2975
rect 10183 2941 10195 2975
rect 10137 2935 10195 2941
rect 10226 2932 10232 2984
rect 10284 2972 10290 2984
rect 10405 2975 10463 2981
rect 10405 2972 10417 2975
rect 10284 2944 10417 2972
rect 10284 2932 10290 2944
rect 10405 2941 10417 2944
rect 10451 2941 10463 2975
rect 10405 2935 10463 2941
rect 10511 2932 10517 2984
rect 10569 2972 10575 2984
rect 10569 2944 10613 2972
rect 10569 2932 10575 2944
rect 6788 2876 7052 2904
rect 6788 2864 6794 2876
rect 7282 2864 7288 2916
rect 7340 2864 7346 2916
rect 7374 2864 7380 2916
rect 7432 2904 7438 2916
rect 8846 2904 8852 2916
rect 7432 2876 8852 2904
rect 7432 2864 7438 2876
rect 8846 2864 8852 2876
rect 8904 2864 8910 2916
rect 8938 2864 8944 2916
rect 8996 2864 9002 2916
rect 9493 2907 9551 2913
rect 9493 2873 9505 2907
rect 9539 2904 9551 2907
rect 10888 2904 10916 3012
rect 11606 3000 11612 3012
rect 11664 3000 11670 3052
rect 11716 3040 11744 3148
rect 11790 3136 11796 3188
rect 11848 3136 11854 3188
rect 11885 3179 11943 3185
rect 11885 3145 11897 3179
rect 11931 3176 11943 3179
rect 11974 3176 11980 3188
rect 11931 3148 11980 3176
rect 11931 3145 11943 3148
rect 11885 3139 11943 3145
rect 11974 3136 11980 3148
rect 12032 3136 12038 3188
rect 12069 3179 12127 3185
rect 12069 3145 12081 3179
rect 12115 3176 12127 3179
rect 12342 3176 12348 3188
rect 12115 3148 12348 3176
rect 12115 3145 12127 3148
rect 12069 3139 12127 3145
rect 12342 3136 12348 3148
rect 12400 3136 12406 3188
rect 12437 3179 12495 3185
rect 12437 3145 12449 3179
rect 12483 3176 12495 3179
rect 12710 3176 12716 3188
rect 12483 3148 12716 3176
rect 12483 3145 12495 3148
rect 12437 3139 12495 3145
rect 12710 3136 12716 3148
rect 12768 3136 12774 3188
rect 14090 3176 14096 3188
rect 14051 3148 14096 3176
rect 14090 3136 14096 3148
rect 14148 3136 14154 3188
rect 11808 3108 11836 3136
rect 13814 3108 13820 3120
rect 11808 3080 13820 3108
rect 13814 3068 13820 3080
rect 13872 3068 13878 3120
rect 11790 3040 11796 3052
rect 11716 3012 11796 3040
rect 11790 3000 11796 3012
rect 11848 3000 11854 3052
rect 12342 3000 12348 3052
rect 12400 3040 12406 3052
rect 12713 3043 12771 3049
rect 12713 3040 12725 3043
rect 12400 3012 12725 3040
rect 12400 3000 12406 3012
rect 12713 3009 12725 3012
rect 12759 3009 12771 3043
rect 14550 3040 14556 3052
rect 12713 3003 12771 3009
rect 14384 3012 14556 3040
rect 10965 2975 11023 2981
rect 10965 2941 10977 2975
rect 11011 2972 11023 2975
rect 11146 2972 11152 2984
rect 11011 2944 11152 2972
rect 11011 2941 11023 2944
rect 10965 2935 11023 2941
rect 11146 2932 11152 2944
rect 11204 2932 11210 2984
rect 11241 2975 11299 2981
rect 11241 2941 11253 2975
rect 11287 2972 11299 2975
rect 11347 2972 11353 2984
rect 11287 2944 11353 2972
rect 11287 2941 11299 2944
rect 11241 2935 11299 2941
rect 11347 2932 11353 2944
rect 11405 2932 11411 2984
rect 11517 2975 11575 2981
rect 11517 2941 11529 2975
rect 11563 2941 11575 2975
rect 11698 2972 11704 2984
rect 11659 2944 11704 2972
rect 11517 2935 11575 2941
rect 11532 2904 11560 2935
rect 11698 2932 11704 2944
rect 11756 2932 11762 2984
rect 12066 2932 12072 2984
rect 12124 2972 12130 2984
rect 12253 2975 12311 2981
rect 12253 2972 12265 2975
rect 12124 2944 12265 2972
rect 12124 2932 12130 2944
rect 12253 2941 12265 2944
rect 12299 2941 12311 2975
rect 12253 2935 12311 2941
rect 11606 2904 11612 2916
rect 9539 2876 10916 2904
rect 11072 2876 11468 2904
rect 11532 2876 11612 2904
rect 9539 2873 9551 2876
rect 9493 2867 9551 2873
rect 4120 2808 5948 2836
rect 5997 2839 6055 2845
rect 4120 2796 4126 2808
rect 5997 2805 6009 2839
rect 6043 2836 6055 2839
rect 6914 2836 6920 2848
rect 6043 2808 6920 2836
rect 6043 2805 6055 2808
rect 5997 2799 6055 2805
rect 6914 2796 6920 2808
rect 6972 2796 6978 2848
rect 7300 2836 7328 2864
rect 8113 2839 8171 2845
rect 8113 2836 8125 2839
rect 7300 2808 8125 2836
rect 8113 2805 8125 2808
rect 8159 2805 8171 2839
rect 8113 2799 8171 2805
rect 8573 2839 8631 2845
rect 8573 2805 8585 2839
rect 8619 2836 8631 2839
rect 8662 2836 8668 2848
rect 8619 2808 8668 2836
rect 8619 2805 8631 2808
rect 8573 2799 8631 2805
rect 8662 2796 8668 2808
rect 8720 2796 8726 2848
rect 9030 2796 9036 2848
rect 9088 2836 9094 2848
rect 9508 2836 9536 2867
rect 9674 2836 9680 2848
rect 9088 2808 9536 2836
rect 9635 2808 9680 2836
rect 9088 2796 9094 2808
rect 9674 2796 9680 2808
rect 9732 2796 9738 2848
rect 9950 2836 9956 2848
rect 9911 2808 9956 2836
rect 9950 2796 9956 2808
rect 10008 2796 10014 2848
rect 10226 2836 10232 2848
rect 10187 2808 10232 2836
rect 10226 2796 10232 2808
rect 10284 2796 10290 2848
rect 10689 2839 10747 2845
rect 10689 2805 10701 2839
rect 10735 2836 10747 2839
rect 10870 2836 10876 2848
rect 10735 2808 10876 2836
rect 10735 2805 10747 2808
rect 10689 2799 10747 2805
rect 10870 2796 10876 2808
rect 10928 2796 10934 2848
rect 11072 2845 11100 2876
rect 11057 2839 11115 2845
rect 11057 2805 11069 2839
rect 11103 2805 11115 2839
rect 11440 2836 11468 2876
rect 11606 2864 11612 2876
rect 11664 2904 11670 2916
rect 12268 2904 12296 2935
rect 12434 2932 12440 2984
rect 12492 2972 12498 2984
rect 12621 2975 12679 2981
rect 12621 2972 12633 2975
rect 12492 2944 12633 2972
rect 12492 2932 12498 2944
rect 12621 2941 12633 2944
rect 12667 2972 12679 2975
rect 13081 2975 13139 2981
rect 13081 2972 13093 2975
rect 12667 2944 13093 2972
rect 12667 2941 12679 2944
rect 12621 2935 12679 2941
rect 13081 2941 13093 2944
rect 13127 2941 13139 2975
rect 13081 2935 13139 2941
rect 13170 2932 13176 2984
rect 13228 2972 13234 2984
rect 14384 2981 14412 3012
rect 14550 3000 14556 3012
rect 14608 3000 14614 3052
rect 15197 3043 15255 3049
rect 15197 3040 15209 3043
rect 14752 3012 15209 3040
rect 13541 2975 13599 2981
rect 13541 2972 13553 2975
rect 13228 2944 13553 2972
rect 13228 2932 13234 2944
rect 13541 2941 13553 2944
rect 13587 2941 13599 2975
rect 13541 2935 13599 2941
rect 14268 2975 14326 2981
rect 14268 2941 14280 2975
rect 14314 2941 14326 2975
rect 14268 2935 14326 2941
rect 14377 2975 14435 2981
rect 14377 2941 14389 2975
rect 14423 2941 14435 2975
rect 14642 2972 14648 2984
rect 14603 2944 14648 2972
rect 14377 2935 14435 2941
rect 12897 2907 12955 2913
rect 12897 2904 12909 2907
rect 11664 2876 12112 2904
rect 12268 2876 12909 2904
rect 11664 2864 11670 2876
rect 11974 2836 11980 2848
rect 11440 2808 11980 2836
rect 11057 2799 11115 2805
rect 11974 2796 11980 2808
rect 12032 2796 12038 2848
rect 12084 2836 12112 2876
rect 12897 2873 12909 2876
rect 12943 2873 12955 2907
rect 12897 2867 12955 2873
rect 13446 2864 13452 2916
rect 13504 2904 13510 2916
rect 13725 2907 13783 2913
rect 13725 2904 13737 2907
rect 13504 2876 13737 2904
rect 13504 2864 13510 2876
rect 13725 2873 13737 2876
rect 13771 2873 13783 2907
rect 13725 2867 13783 2873
rect 14182 2864 14188 2916
rect 14240 2904 14246 2916
rect 14292 2904 14320 2935
rect 14642 2932 14648 2944
rect 14700 2932 14706 2984
rect 14752 2904 14780 3012
rect 15197 3009 15209 3012
rect 15243 3009 15255 3043
rect 15197 3003 15255 3009
rect 15010 2932 15016 2984
rect 15068 2972 15074 2984
rect 15105 2975 15163 2981
rect 15105 2972 15117 2975
rect 15068 2944 15117 2972
rect 15068 2932 15074 2944
rect 15105 2941 15117 2944
rect 15151 2941 15163 2975
rect 15105 2935 15163 2941
rect 15473 2907 15531 2913
rect 15473 2904 15485 2907
rect 14240 2876 14780 2904
rect 14844 2876 15485 2904
rect 14240 2864 14246 2876
rect 12618 2836 12624 2848
rect 12084 2808 12624 2836
rect 12618 2796 12624 2808
rect 12676 2796 12682 2848
rect 12802 2796 12808 2848
rect 12860 2836 12866 2848
rect 13265 2839 13323 2845
rect 13265 2836 13277 2839
rect 12860 2808 13277 2836
rect 12860 2796 12866 2808
rect 13265 2805 13277 2808
rect 13311 2805 13323 2839
rect 13265 2799 13323 2805
rect 13814 2796 13820 2848
rect 13872 2836 13878 2848
rect 13909 2839 13967 2845
rect 13909 2836 13921 2839
rect 13872 2808 13921 2836
rect 13872 2796 13878 2808
rect 13909 2805 13921 2808
rect 13955 2805 13967 2839
rect 14550 2836 14556 2848
rect 14511 2808 14556 2836
rect 13909 2799 13967 2805
rect 14550 2796 14556 2808
rect 14608 2796 14614 2848
rect 14844 2845 14872 2876
rect 15473 2873 15485 2876
rect 15519 2873 15531 2907
rect 15473 2867 15531 2873
rect 15657 2907 15715 2913
rect 15657 2873 15669 2907
rect 15703 2904 15715 2907
rect 16942 2904 16948 2916
rect 15703 2876 16948 2904
rect 15703 2873 15715 2876
rect 15657 2867 15715 2873
rect 16942 2864 16948 2876
rect 17000 2864 17006 2916
rect 14829 2839 14887 2845
rect 14829 2805 14841 2839
rect 14875 2805 14887 2839
rect 14829 2799 14887 2805
rect 14918 2796 14924 2848
rect 14976 2836 14982 2848
rect 14976 2808 15021 2836
rect 14976 2796 14982 2808
rect 1104 2746 16008 2768
rect 1104 2694 5979 2746
rect 6031 2694 6043 2746
rect 6095 2694 6107 2746
rect 6159 2694 6171 2746
rect 6223 2694 10976 2746
rect 11028 2694 11040 2746
rect 11092 2694 11104 2746
rect 11156 2694 11168 2746
rect 11220 2694 16008 2746
rect 1104 2672 16008 2694
rect 2406 2632 2412 2644
rect 1596 2604 2412 2632
rect 1596 2573 1624 2604
rect 2406 2592 2412 2604
rect 2464 2592 2470 2644
rect 5353 2635 5411 2641
rect 5353 2632 5365 2635
rect 2746 2604 5365 2632
rect 2746 2576 2774 2604
rect 5353 2601 5365 2604
rect 5399 2601 5411 2635
rect 5626 2632 5632 2644
rect 5587 2604 5632 2632
rect 5353 2595 5411 2601
rect 5626 2592 5632 2604
rect 5684 2592 5690 2644
rect 6454 2592 6460 2644
rect 6512 2632 6518 2644
rect 6549 2635 6607 2641
rect 6549 2632 6561 2635
rect 6512 2604 6561 2632
rect 6512 2592 6518 2604
rect 6549 2601 6561 2604
rect 6595 2601 6607 2635
rect 6549 2595 6607 2601
rect 7009 2635 7067 2641
rect 7009 2601 7021 2635
rect 7055 2632 7067 2635
rect 7098 2632 7104 2644
rect 7055 2604 7104 2632
rect 7055 2601 7067 2604
rect 7009 2595 7067 2601
rect 7098 2592 7104 2604
rect 7156 2592 7162 2644
rect 7377 2635 7435 2641
rect 7377 2601 7389 2635
rect 7423 2601 7435 2635
rect 7377 2595 7435 2601
rect 1581 2567 1639 2573
rect 1581 2533 1593 2567
rect 1627 2533 1639 2567
rect 1581 2527 1639 2533
rect 1946 2524 1952 2576
rect 2004 2564 2010 2576
rect 2004 2536 2176 2564
rect 2004 2524 2010 2536
rect 2038 2496 2044 2508
rect 1999 2468 2044 2496
rect 2038 2456 2044 2468
rect 2096 2456 2102 2508
rect 2148 2496 2176 2536
rect 2682 2524 2688 2576
rect 2740 2536 2774 2576
rect 2740 2524 2746 2536
rect 2866 2524 2872 2576
rect 2924 2564 2930 2576
rect 4433 2567 4491 2573
rect 4433 2564 4445 2567
rect 2924 2536 4445 2564
rect 2924 2524 2930 2536
rect 4433 2533 4445 2536
rect 4479 2533 4491 2567
rect 4433 2527 4491 2533
rect 4614 2524 4620 2576
rect 4672 2564 4678 2576
rect 7392 2564 7420 2595
rect 8662 2592 8668 2644
rect 8720 2632 8726 2644
rect 9490 2632 9496 2644
rect 8720 2604 9496 2632
rect 8720 2592 8726 2604
rect 9490 2592 9496 2604
rect 9548 2592 9554 2644
rect 9582 2592 9588 2644
rect 9640 2632 9646 2644
rect 9677 2635 9735 2641
rect 9677 2632 9689 2635
rect 9640 2604 9689 2632
rect 9640 2592 9646 2604
rect 9677 2601 9689 2604
rect 9723 2601 9735 2635
rect 9677 2595 9735 2601
rect 9953 2635 10011 2641
rect 9953 2601 9965 2635
rect 9999 2632 10011 2635
rect 10318 2632 10324 2644
rect 9999 2604 10324 2632
rect 9999 2601 10011 2604
rect 9953 2595 10011 2601
rect 10318 2592 10324 2604
rect 10376 2592 10382 2644
rect 10410 2592 10416 2644
rect 10468 2632 10474 2644
rect 11514 2632 11520 2644
rect 10468 2604 11017 2632
rect 11475 2604 11520 2632
rect 10468 2592 10474 2604
rect 7742 2564 7748 2576
rect 4672 2536 7420 2564
rect 7703 2536 7748 2564
rect 4672 2524 4678 2536
rect 7742 2524 7748 2536
rect 7800 2524 7806 2576
rect 7837 2567 7895 2573
rect 7837 2533 7849 2567
rect 7883 2564 7895 2567
rect 9122 2564 9128 2576
rect 7883 2536 9128 2564
rect 7883 2533 7895 2536
rect 7837 2527 7895 2533
rect 9122 2524 9128 2536
rect 9180 2524 9186 2576
rect 9214 2524 9220 2576
rect 9272 2564 9278 2576
rect 9272 2536 10456 2564
rect 9272 2524 9278 2536
rect 10428 2508 10456 2536
rect 10870 2524 10876 2576
rect 10928 2524 10934 2576
rect 10989 2564 11017 2604
rect 11514 2592 11520 2604
rect 11572 2592 11578 2644
rect 11790 2592 11796 2644
rect 11848 2632 11854 2644
rect 11974 2632 11980 2644
rect 11848 2604 11980 2632
rect 11848 2592 11854 2604
rect 11974 2592 11980 2604
rect 12032 2592 12038 2644
rect 12526 2592 12532 2644
rect 12584 2632 12590 2644
rect 12897 2635 12955 2641
rect 12897 2632 12909 2635
rect 12584 2604 12909 2632
rect 12584 2592 12590 2604
rect 12897 2601 12909 2604
rect 12943 2601 12955 2635
rect 12897 2595 12955 2601
rect 13265 2635 13323 2641
rect 13265 2601 13277 2635
rect 13311 2632 13323 2635
rect 14090 2632 14096 2644
rect 13311 2604 14096 2632
rect 13311 2601 13323 2604
rect 13265 2595 13323 2601
rect 14090 2592 14096 2604
rect 14148 2592 14154 2644
rect 14369 2635 14427 2641
rect 14369 2601 14381 2635
rect 14415 2632 14427 2635
rect 14415 2604 15516 2632
rect 14415 2601 14427 2604
rect 14369 2595 14427 2601
rect 11054 2564 11060 2576
rect 10989 2536 11060 2564
rect 11054 2524 11060 2536
rect 11112 2524 11118 2576
rect 11146 2524 11152 2576
rect 11204 2564 11210 2576
rect 11333 2567 11391 2573
rect 11333 2564 11345 2567
rect 11204 2536 11345 2564
rect 11204 2524 11210 2536
rect 11333 2533 11345 2536
rect 11379 2533 11391 2567
rect 12437 2567 12495 2573
rect 12437 2564 12449 2567
rect 11333 2527 11391 2533
rect 11440 2536 12449 2564
rect 2573 2499 2631 2505
rect 2573 2496 2585 2499
rect 2148 2468 2585 2496
rect 2573 2465 2585 2468
rect 2619 2465 2631 2499
rect 2573 2459 2631 2465
rect 3786 2456 3792 2508
rect 3844 2496 3850 2508
rect 3881 2499 3939 2505
rect 3881 2496 3893 2499
rect 3844 2468 3893 2496
rect 3844 2456 3850 2468
rect 3881 2465 3893 2468
rect 3927 2465 3939 2499
rect 3881 2459 3939 2465
rect 4065 2499 4123 2505
rect 4065 2465 4077 2499
rect 4111 2496 4123 2499
rect 4246 2496 4252 2508
rect 4111 2468 4252 2496
rect 4111 2465 4123 2468
rect 4065 2459 4123 2465
rect 4246 2456 4252 2468
rect 4304 2456 4310 2508
rect 4798 2496 4804 2508
rect 4759 2468 4804 2496
rect 4798 2456 4804 2468
rect 4856 2456 4862 2508
rect 5166 2496 5172 2508
rect 5127 2468 5172 2496
rect 5166 2456 5172 2468
rect 5224 2456 5230 2508
rect 5537 2499 5595 2505
rect 5537 2465 5549 2499
rect 5583 2496 5595 2499
rect 5994 2496 6000 2508
rect 5583 2468 5856 2496
rect 5955 2468 6000 2496
rect 5583 2465 5595 2468
rect 5537 2459 5595 2465
rect 2314 2428 2320 2440
rect 2275 2400 2320 2428
rect 2314 2388 2320 2400
rect 2372 2388 2378 2440
rect 4890 2428 4896 2440
rect 3620 2400 4896 2428
rect 106 2320 112 2372
rect 164 2360 170 2372
rect 1397 2363 1455 2369
rect 1397 2360 1409 2363
rect 164 2332 1409 2360
rect 164 2320 170 2332
rect 1397 2329 1409 2332
rect 1443 2329 1455 2363
rect 1397 2323 1455 2329
rect 1857 2363 1915 2369
rect 1857 2329 1869 2363
rect 1903 2360 1915 2363
rect 2222 2360 2228 2372
rect 1903 2332 2228 2360
rect 1903 2329 1915 2332
rect 1857 2323 1915 2329
rect 2222 2320 2228 2332
rect 2280 2320 2286 2372
rect 2133 2295 2191 2301
rect 2133 2261 2145 2295
rect 2179 2292 2191 2295
rect 3620 2292 3648 2400
rect 4890 2388 4896 2400
rect 4948 2388 4954 2440
rect 3970 2320 3976 2372
rect 4028 2360 4034 2372
rect 4249 2363 4307 2369
rect 4249 2360 4261 2363
rect 4028 2332 4261 2360
rect 4028 2320 4034 2332
rect 4249 2329 4261 2332
rect 4295 2329 4307 2363
rect 4249 2323 4307 2329
rect 4522 2320 4528 2372
rect 4580 2360 4586 2372
rect 4985 2363 5043 2369
rect 4985 2360 4997 2363
rect 4580 2332 4997 2360
rect 4580 2320 4586 2332
rect 4985 2329 4997 2332
rect 5031 2329 5043 2363
rect 5828 2360 5856 2468
rect 5994 2456 6000 2468
rect 6052 2456 6058 2508
rect 6914 2456 6920 2508
rect 6972 2496 6978 2508
rect 6972 2468 7017 2496
rect 6972 2456 6978 2468
rect 7558 2456 7564 2508
rect 7616 2456 7622 2508
rect 8018 2456 8024 2508
rect 8076 2496 8082 2508
rect 8481 2499 8539 2505
rect 8481 2496 8493 2499
rect 8076 2468 8493 2496
rect 8076 2456 8082 2468
rect 8481 2465 8493 2468
rect 8527 2465 8539 2499
rect 8846 2496 8852 2508
rect 8807 2468 8852 2496
rect 8481 2459 8539 2465
rect 6086 2428 6092 2440
rect 6047 2400 6092 2428
rect 6086 2388 6092 2400
rect 6144 2388 6150 2440
rect 6270 2428 6276 2440
rect 6231 2400 6276 2428
rect 6270 2388 6276 2400
rect 6328 2388 6334 2440
rect 7190 2428 7196 2440
rect 7151 2400 7196 2428
rect 7190 2388 7196 2400
rect 7248 2388 7254 2440
rect 7576 2428 7604 2456
rect 7929 2431 7987 2437
rect 7929 2428 7941 2431
rect 7576 2400 7941 2428
rect 7929 2397 7941 2400
rect 7975 2397 7987 2431
rect 7929 2391 7987 2397
rect 7466 2360 7472 2372
rect 5828 2332 7472 2360
rect 4985 2323 5043 2329
rect 7466 2320 7472 2332
rect 7524 2320 7530 2372
rect 8110 2320 8116 2372
rect 8168 2360 8174 2372
rect 8496 2360 8524 2459
rect 8846 2456 8852 2468
rect 8904 2456 8910 2508
rect 9398 2456 9404 2508
rect 9456 2496 9462 2508
rect 9493 2499 9551 2505
rect 9493 2496 9505 2499
rect 9456 2468 9505 2496
rect 9456 2456 9462 2468
rect 9493 2465 9505 2468
rect 9539 2465 9551 2499
rect 9858 2496 9864 2508
rect 9771 2468 9864 2496
rect 9493 2459 9551 2465
rect 9858 2456 9864 2468
rect 9916 2496 9922 2508
rect 9953 2499 10011 2505
rect 9953 2496 9965 2499
rect 9916 2468 9965 2496
rect 9916 2456 9922 2468
rect 9953 2465 9965 2468
rect 9999 2465 10011 2499
rect 9953 2459 10011 2465
rect 10229 2499 10287 2505
rect 10229 2465 10241 2499
rect 10275 2496 10287 2499
rect 10318 2496 10324 2508
rect 10275 2468 10324 2496
rect 10275 2465 10287 2468
rect 10229 2459 10287 2465
rect 10318 2456 10324 2468
rect 10376 2456 10382 2508
rect 10410 2456 10416 2508
rect 10468 2456 10474 2508
rect 10594 2496 10600 2508
rect 10555 2468 10600 2496
rect 10594 2456 10600 2468
rect 10652 2456 10658 2508
rect 10888 2496 10916 2524
rect 10965 2499 11023 2505
rect 10965 2496 10977 2499
rect 10888 2468 10977 2496
rect 10965 2465 10977 2468
rect 11011 2465 11023 2499
rect 10965 2459 11023 2465
rect 11238 2456 11244 2508
rect 11296 2496 11302 2508
rect 11440 2496 11468 2536
rect 12437 2533 12449 2536
rect 12483 2533 12495 2567
rect 12437 2527 12495 2533
rect 14737 2567 14795 2573
rect 14737 2533 14749 2567
rect 14783 2564 14795 2567
rect 14918 2564 14924 2576
rect 14783 2536 14924 2564
rect 14783 2533 14795 2536
rect 14737 2527 14795 2533
rect 14918 2524 14924 2536
rect 14976 2524 14982 2576
rect 15488 2573 15516 2604
rect 15473 2567 15531 2573
rect 15473 2533 15485 2567
rect 15519 2533 15531 2567
rect 15473 2527 15531 2533
rect 11296 2468 11468 2496
rect 11296 2456 11302 2468
rect 11514 2456 11520 2508
rect 11572 2496 11578 2508
rect 11701 2499 11759 2505
rect 11701 2496 11713 2499
rect 11572 2468 11713 2496
rect 11572 2456 11578 2468
rect 11701 2465 11713 2468
rect 11747 2465 11759 2499
rect 11701 2459 11759 2465
rect 10502 2388 10508 2440
rect 10560 2428 10566 2440
rect 11716 2428 11744 2459
rect 11790 2456 11796 2508
rect 11848 2496 11854 2508
rect 12069 2499 12127 2505
rect 12069 2496 12081 2499
rect 11848 2468 12081 2496
rect 11848 2456 11854 2468
rect 12069 2465 12081 2468
rect 12115 2496 12127 2499
rect 12342 2496 12348 2508
rect 12115 2468 12348 2496
rect 12115 2465 12127 2468
rect 12069 2459 12127 2465
rect 12342 2456 12348 2468
rect 12400 2456 12406 2508
rect 12802 2456 12808 2508
rect 12860 2496 12866 2508
rect 12989 2499 13047 2505
rect 12989 2496 13001 2499
rect 12860 2468 13001 2496
rect 12860 2456 12866 2468
rect 12989 2465 13001 2468
rect 13035 2465 13047 2499
rect 12989 2459 13047 2465
rect 13170 2456 13176 2508
rect 13228 2496 13234 2508
rect 13357 2499 13415 2505
rect 13357 2496 13369 2499
rect 13228 2468 13369 2496
rect 13228 2456 13234 2468
rect 13357 2465 13369 2468
rect 13403 2465 13415 2499
rect 13357 2459 13415 2465
rect 13446 2456 13452 2508
rect 13504 2496 13510 2508
rect 13725 2499 13783 2505
rect 13725 2496 13737 2499
rect 13504 2468 13737 2496
rect 13504 2456 13510 2468
rect 13725 2465 13737 2468
rect 13771 2465 13783 2499
rect 13725 2459 13783 2465
rect 13814 2456 13820 2508
rect 13872 2496 13878 2508
rect 13909 2499 13967 2505
rect 13909 2496 13921 2499
rect 13872 2468 13921 2496
rect 13872 2456 13878 2468
rect 13909 2465 13921 2468
rect 13955 2465 13967 2499
rect 13909 2459 13967 2465
rect 13998 2456 14004 2508
rect 14056 2496 14062 2508
rect 14185 2499 14243 2505
rect 14185 2496 14197 2499
rect 14056 2468 14197 2496
rect 14056 2456 14062 2468
rect 14185 2465 14197 2468
rect 14231 2465 14243 2499
rect 14185 2459 14243 2465
rect 14550 2456 14556 2508
rect 14608 2496 14614 2508
rect 15105 2499 15163 2505
rect 15105 2496 15117 2499
rect 14608 2468 15117 2496
rect 14608 2456 14614 2468
rect 15105 2465 15117 2468
rect 15151 2465 15163 2499
rect 15105 2459 15163 2465
rect 12621 2431 12679 2437
rect 12621 2428 12633 2431
rect 10560 2400 10916 2428
rect 11716 2400 12633 2428
rect 10560 2388 10566 2400
rect 8941 2363 8999 2369
rect 8941 2360 8953 2363
rect 8168 2332 8432 2360
rect 8496 2332 8953 2360
rect 8168 2320 8174 2332
rect 2179 2264 3648 2292
rect 3697 2295 3755 2301
rect 2179 2261 2191 2264
rect 2133 2255 2191 2261
rect 3697 2261 3709 2295
rect 3743 2292 3755 2295
rect 4062 2292 4068 2304
rect 3743 2264 4068 2292
rect 3743 2261 3755 2264
rect 3697 2255 3755 2261
rect 4062 2252 4068 2264
rect 4120 2252 4126 2304
rect 4154 2252 4160 2304
rect 4212 2292 4218 2304
rect 4709 2295 4767 2301
rect 4709 2292 4721 2295
rect 4212 2264 4721 2292
rect 4212 2252 4218 2264
rect 4709 2261 4721 2264
rect 4755 2261 4767 2295
rect 4709 2255 4767 2261
rect 6546 2252 6552 2304
rect 6604 2292 6610 2304
rect 8297 2295 8355 2301
rect 8297 2292 8309 2295
rect 6604 2264 8309 2292
rect 6604 2252 6610 2264
rect 8297 2261 8309 2264
rect 8343 2261 8355 2295
rect 8404 2292 8432 2332
rect 8941 2329 8953 2332
rect 8987 2329 8999 2363
rect 8941 2323 8999 2329
rect 9122 2320 9128 2372
rect 9180 2360 9186 2372
rect 10781 2363 10839 2369
rect 10781 2360 10793 2363
rect 9180 2332 10793 2360
rect 9180 2320 9186 2332
rect 10781 2329 10793 2332
rect 10827 2329 10839 2363
rect 10888 2360 10916 2400
rect 12621 2397 12633 2400
rect 12667 2397 12679 2431
rect 12621 2391 12679 2397
rect 14921 2431 14979 2437
rect 14921 2397 14933 2431
rect 14967 2428 14979 2431
rect 16574 2428 16580 2440
rect 14967 2400 16580 2428
rect 14967 2397 14979 2400
rect 14921 2391 14979 2397
rect 16574 2388 16580 2400
rect 16632 2388 16638 2440
rect 11885 2363 11943 2369
rect 11885 2360 11897 2363
rect 10888 2332 11897 2360
rect 10781 2323 10839 2329
rect 11885 2329 11897 2332
rect 11931 2329 11943 2363
rect 11885 2323 11943 2329
rect 11974 2320 11980 2372
rect 12032 2360 12038 2372
rect 13541 2363 13599 2369
rect 13541 2360 13553 2363
rect 12032 2332 13553 2360
rect 12032 2320 12038 2332
rect 13541 2329 13553 2332
rect 13587 2329 13599 2363
rect 13541 2323 13599 2329
rect 14093 2363 14151 2369
rect 14093 2329 14105 2363
rect 14139 2360 14151 2363
rect 15102 2360 15108 2372
rect 14139 2332 15108 2360
rect 14139 2329 14151 2332
rect 14093 2323 14151 2329
rect 15102 2320 15108 2332
rect 15160 2320 15166 2372
rect 15289 2363 15347 2369
rect 15289 2329 15301 2363
rect 15335 2360 15347 2363
rect 15930 2360 15936 2372
rect 15335 2332 15936 2360
rect 15335 2329 15347 2332
rect 15289 2323 15347 2329
rect 15930 2320 15936 2332
rect 15988 2320 15994 2372
rect 8665 2295 8723 2301
rect 8665 2292 8677 2295
rect 8404 2264 8677 2292
rect 8297 2255 8355 2261
rect 8665 2261 8677 2264
rect 8711 2261 8723 2295
rect 8665 2255 8723 2261
rect 9309 2295 9367 2301
rect 9309 2261 9321 2295
rect 9355 2292 9367 2295
rect 9490 2292 9496 2304
rect 9355 2264 9496 2292
rect 9355 2261 9367 2264
rect 9309 2255 9367 2261
rect 9490 2252 9496 2264
rect 9548 2252 9554 2304
rect 10134 2292 10140 2304
rect 10095 2264 10140 2292
rect 10134 2252 10140 2264
rect 10192 2252 10198 2304
rect 10410 2252 10416 2304
rect 10468 2292 10474 2304
rect 10505 2295 10563 2301
rect 10505 2292 10517 2295
rect 10468 2264 10517 2292
rect 10468 2252 10474 2264
rect 10505 2261 10517 2264
rect 10551 2292 10563 2295
rect 10962 2292 10968 2304
rect 10551 2264 10968 2292
rect 10551 2261 10563 2264
rect 10505 2255 10563 2261
rect 10962 2252 10968 2264
rect 11020 2252 11026 2304
rect 11238 2292 11244 2304
rect 11199 2264 11244 2292
rect 11238 2252 11244 2264
rect 11296 2252 11302 2304
rect 12342 2292 12348 2304
rect 12303 2264 12348 2292
rect 12342 2252 12348 2264
rect 12400 2252 12406 2304
rect 15562 2292 15568 2304
rect 15523 2264 15568 2292
rect 15562 2252 15568 2264
rect 15620 2252 15626 2304
rect 1104 2202 16008 2224
rect 1104 2150 3480 2202
rect 3532 2150 3544 2202
rect 3596 2150 3608 2202
rect 3660 2150 3672 2202
rect 3724 2150 8478 2202
rect 8530 2150 8542 2202
rect 8594 2150 8606 2202
rect 8658 2150 8670 2202
rect 8722 2150 13475 2202
rect 13527 2150 13539 2202
rect 13591 2150 13603 2202
rect 13655 2150 13667 2202
rect 13719 2150 16008 2202
rect 1104 2128 16008 2150
rect 5902 2048 5908 2100
rect 5960 2088 5966 2100
rect 11238 2088 11244 2100
rect 5960 2060 11244 2088
rect 5960 2048 5966 2060
rect 11238 2048 11244 2060
rect 11296 2048 11302 2100
rect 6270 1980 6276 2032
rect 6328 2020 6334 2032
rect 12342 2020 12348 2032
rect 6328 1992 12348 2020
rect 6328 1980 6334 1992
rect 12342 1980 12348 1992
rect 12400 1980 12406 2032
rect 2038 1912 2044 1964
rect 2096 1952 2102 1964
rect 2096 1924 2774 1952
rect 2096 1912 2102 1924
rect 2746 1476 2774 1924
rect 6822 1912 6828 1964
rect 6880 1952 6886 1964
rect 8202 1952 8208 1964
rect 6880 1924 8208 1952
rect 6880 1912 6886 1924
rect 8202 1912 8208 1924
rect 8260 1912 8266 1964
rect 10134 1912 10140 1964
rect 10192 1952 10198 1964
rect 12158 1952 12164 1964
rect 10192 1924 12164 1952
rect 10192 1912 10198 1924
rect 12158 1912 12164 1924
rect 12216 1912 12222 1964
rect 7650 1844 7656 1896
rect 7708 1884 7714 1896
rect 9398 1884 9404 1896
rect 7708 1856 9404 1884
rect 7708 1844 7714 1856
rect 9398 1844 9404 1856
rect 9456 1844 9462 1896
rect 10318 1844 10324 1896
rect 10376 1884 10382 1896
rect 12986 1884 12992 1896
rect 10376 1856 12992 1884
rect 10376 1844 10382 1856
rect 12986 1844 12992 1856
rect 13044 1844 13050 1896
rect 5166 1776 5172 1828
rect 5224 1816 5230 1828
rect 9950 1816 9956 1828
rect 5224 1788 9956 1816
rect 5224 1776 5230 1788
rect 9950 1776 9956 1788
rect 10008 1776 10014 1828
rect 10778 1776 10784 1828
rect 10836 1816 10842 1828
rect 12894 1816 12900 1828
rect 10836 1788 12900 1816
rect 10836 1776 10842 1788
rect 12894 1776 12900 1788
rect 12952 1776 12958 1828
rect 4246 1708 4252 1760
rect 4304 1748 4310 1760
rect 9766 1748 9772 1760
rect 4304 1720 9772 1748
rect 4304 1708 4310 1720
rect 9766 1708 9772 1720
rect 9824 1708 9830 1760
rect 10686 1708 10692 1760
rect 10744 1748 10750 1760
rect 11514 1748 11520 1760
rect 10744 1720 11520 1748
rect 10744 1708 10750 1720
rect 11514 1708 11520 1720
rect 11572 1708 11578 1760
rect 4798 1640 4804 1692
rect 4856 1680 4862 1692
rect 10042 1680 10048 1692
rect 4856 1652 10048 1680
rect 4856 1640 4862 1652
rect 10042 1640 10048 1652
rect 10100 1640 10106 1692
rect 5994 1572 6000 1624
rect 6052 1612 6058 1624
rect 11422 1612 11428 1624
rect 6052 1584 11428 1612
rect 6052 1572 6058 1584
rect 11422 1572 11428 1584
rect 11480 1572 11486 1624
rect 6914 1504 6920 1556
rect 6972 1544 6978 1556
rect 7926 1544 7932 1556
rect 6972 1516 7932 1544
rect 6972 1504 6978 1516
rect 7926 1504 7932 1516
rect 7984 1504 7990 1556
rect 8018 1504 8024 1556
rect 8076 1544 8082 1556
rect 9858 1544 9864 1556
rect 8076 1516 9864 1544
rect 8076 1504 8082 1516
rect 9858 1504 9864 1516
rect 9916 1504 9922 1556
rect 2746 1448 9260 1476
rect 5534 1368 5540 1420
rect 5592 1408 5598 1420
rect 9122 1408 9128 1420
rect 5592 1380 9128 1408
rect 5592 1368 5598 1380
rect 9122 1368 9128 1380
rect 9180 1368 9186 1420
rect 9232 1408 9260 1448
rect 9674 1436 9680 1488
rect 9732 1476 9738 1488
rect 12250 1476 12256 1488
rect 9732 1448 12256 1476
rect 9732 1436 9738 1448
rect 12250 1436 12256 1448
rect 12308 1436 12314 1488
rect 10226 1408 10232 1420
rect 9232 1380 10232 1408
rect 10226 1368 10232 1380
rect 10284 1368 10290 1420
<< via1 >>
rect 8392 17620 8444 17672
rect 8852 17620 8904 17672
rect 3480 17382 3532 17434
rect 3544 17382 3596 17434
rect 3608 17382 3660 17434
rect 3672 17382 3724 17434
rect 8478 17382 8530 17434
rect 8542 17382 8594 17434
rect 8606 17382 8658 17434
rect 8670 17382 8722 17434
rect 13475 17382 13527 17434
rect 13539 17382 13591 17434
rect 13603 17382 13655 17434
rect 13667 17382 13719 17434
rect 2780 17280 2832 17332
rect 2044 17255 2096 17264
rect 2044 17221 2053 17255
rect 2053 17221 2087 17255
rect 2087 17221 2096 17255
rect 2044 17212 2096 17221
rect 2412 17212 2464 17264
rect 3148 17280 3200 17332
rect 4160 17280 4212 17332
rect 2780 17144 2832 17196
rect 2872 17144 2924 17196
rect 1400 17119 1452 17128
rect 1400 17085 1409 17119
rect 1409 17085 1443 17119
rect 1443 17085 1452 17119
rect 1400 17076 1452 17085
rect 2136 17076 2188 17128
rect 2412 17076 2464 17128
rect 3792 17212 3844 17264
rect 4344 17212 4396 17264
rect 6184 17212 6236 17264
rect 6920 17212 6972 17264
rect 7656 17212 7708 17264
rect 8300 17212 8352 17264
rect 9496 17280 9548 17332
rect 13820 17280 13872 17332
rect 14648 17280 14700 17332
rect 8944 17212 8996 17264
rect 2228 17051 2280 17060
rect 2228 17017 2237 17051
rect 2237 17017 2271 17051
rect 2271 17017 2280 17051
rect 2228 17008 2280 17017
rect 2964 17051 3016 17060
rect 2964 17017 2973 17051
rect 2973 17017 3007 17051
rect 3007 17017 3016 17051
rect 2964 17008 3016 17017
rect 4160 17144 4212 17196
rect 4620 17144 4672 17196
rect 9036 17144 9088 17196
rect 3792 17076 3844 17128
rect 6552 17076 6604 17128
rect 7288 17076 7340 17128
rect 8484 17076 8536 17128
rect 9128 17076 9180 17128
rect 9864 17076 9916 17128
rect 10232 17076 10284 17128
rect 10600 17076 10652 17128
rect 10692 17076 10744 17128
rect 11060 17076 11112 17128
rect 11336 17076 11388 17128
rect 11428 17076 11480 17128
rect 12900 17144 12952 17196
rect 14740 17144 14792 17196
rect 11796 17076 11848 17128
rect 13084 17076 13136 17128
rect 13820 17076 13872 17128
rect 14096 17076 14148 17128
rect 4252 17008 4304 17060
rect 4436 17051 4488 17060
rect 4436 17017 4445 17051
rect 4445 17017 4479 17051
rect 4479 17017 4488 17051
rect 4436 17008 4488 17017
rect 4804 17051 4856 17060
rect 4804 17017 4813 17051
rect 4813 17017 4847 17051
rect 4847 17017 4856 17051
rect 4804 17008 4856 17017
rect 5172 17051 5224 17060
rect 5172 17017 5181 17051
rect 5181 17017 5215 17051
rect 5215 17017 5224 17051
rect 5172 17008 5224 17017
rect 5540 17051 5592 17060
rect 5540 17017 5549 17051
rect 5549 17017 5583 17051
rect 5583 17017 5592 17051
rect 5540 17008 5592 17017
rect 5816 17051 5868 17060
rect 5816 17017 5825 17051
rect 5825 17017 5859 17051
rect 5859 17017 5868 17051
rect 5816 17008 5868 17017
rect 6644 17008 6696 17060
rect 7104 17051 7156 17060
rect 2872 16940 2924 16992
rect 3240 16940 3292 16992
rect 7104 17017 7113 17051
rect 7113 17017 7147 17051
rect 7147 17017 7156 17051
rect 7104 17008 7156 17017
rect 7288 16940 7340 16992
rect 8300 17008 8352 17060
rect 8760 17051 8812 17060
rect 8760 17017 8769 17051
rect 8769 17017 8803 17051
rect 8803 17017 8812 17051
rect 8760 17008 8812 17017
rect 8944 17051 8996 17060
rect 8944 17017 8953 17051
rect 8953 17017 8987 17051
rect 8987 17017 8996 17051
rect 8944 17008 8996 17017
rect 9404 17051 9456 17060
rect 9404 17017 9413 17051
rect 9413 17017 9447 17051
rect 9447 17017 9456 17051
rect 9404 17008 9456 17017
rect 12808 17008 12860 17060
rect 14372 17076 14424 17128
rect 8852 16940 8904 16992
rect 9312 16940 9364 16992
rect 10232 16940 10284 16992
rect 10508 16940 10560 16992
rect 10784 16940 10836 16992
rect 11888 16940 11940 16992
rect 12072 16983 12124 16992
rect 12072 16949 12081 16983
rect 12081 16949 12115 16983
rect 12115 16949 12124 16983
rect 12072 16940 12124 16949
rect 12624 16983 12676 16992
rect 12624 16949 12633 16983
rect 12633 16949 12667 16983
rect 12667 16949 12676 16983
rect 12624 16940 12676 16949
rect 14096 16940 14148 16992
rect 14832 17008 14884 17060
rect 15292 17051 15344 17060
rect 15292 17017 15301 17051
rect 15301 17017 15335 17051
rect 15335 17017 15344 17051
rect 15292 17008 15344 17017
rect 16580 16940 16632 16992
rect 5979 16838 6031 16890
rect 6043 16838 6095 16890
rect 6107 16838 6159 16890
rect 6171 16838 6223 16890
rect 10976 16838 11028 16890
rect 11040 16838 11092 16890
rect 11104 16838 11156 16890
rect 11168 16838 11220 16890
rect 572 16736 624 16788
rect 2228 16736 2280 16788
rect 3240 16736 3292 16788
rect 5816 16736 5868 16788
rect 6644 16736 6696 16788
rect 9680 16736 9732 16788
rect 9864 16736 9916 16788
rect 10600 16779 10652 16788
rect 10600 16745 10609 16779
rect 10609 16745 10643 16779
rect 10643 16745 10652 16779
rect 10600 16736 10652 16745
rect 10692 16736 10744 16788
rect 11336 16779 11388 16788
rect 11336 16745 11345 16779
rect 11345 16745 11379 16779
rect 11379 16745 11388 16779
rect 11336 16736 11388 16745
rect 11796 16779 11848 16788
rect 11796 16745 11805 16779
rect 11805 16745 11839 16779
rect 11839 16745 11848 16779
rect 11796 16736 11848 16745
rect 204 16668 256 16720
rect 1308 16600 1360 16652
rect 2412 16600 2464 16652
rect 4988 16711 5040 16720
rect 1676 16532 1728 16584
rect 2872 16600 2924 16652
rect 2044 16464 2096 16516
rect 4988 16677 4997 16711
rect 4997 16677 5031 16711
rect 5031 16677 5040 16711
rect 4988 16668 5040 16677
rect 5356 16711 5408 16720
rect 5356 16677 5365 16711
rect 5365 16677 5399 16711
rect 5399 16677 5408 16711
rect 5356 16668 5408 16677
rect 5724 16711 5776 16720
rect 5724 16677 5733 16711
rect 5733 16677 5767 16711
rect 5767 16677 5776 16711
rect 5724 16668 5776 16677
rect 9956 16668 10008 16720
rect 12164 16668 12216 16720
rect 14004 16736 14056 16788
rect 16212 16736 16264 16788
rect 13360 16668 13412 16720
rect 14556 16711 14608 16720
rect 14556 16677 14565 16711
rect 14565 16677 14599 16711
rect 14599 16677 14608 16711
rect 14556 16668 14608 16677
rect 15200 16668 15252 16720
rect 5816 16600 5868 16652
rect 7012 16600 7064 16652
rect 8484 16600 8536 16652
rect 9036 16600 9088 16652
rect 12532 16600 12584 16652
rect 6460 16532 6512 16584
rect 3884 16464 3936 16516
rect 4528 16464 4580 16516
rect 9772 16532 9824 16584
rect 12808 16600 12860 16652
rect 14372 16600 14424 16652
rect 15476 16600 15528 16652
rect 15660 16643 15712 16652
rect 15660 16609 15669 16643
rect 15669 16609 15703 16643
rect 15703 16609 15712 16643
rect 15660 16600 15712 16609
rect 6920 16464 6972 16516
rect 12164 16507 12216 16516
rect 3792 16396 3844 16448
rect 5080 16396 5132 16448
rect 6736 16439 6788 16448
rect 6736 16405 6745 16439
rect 6745 16405 6779 16439
rect 6779 16405 6788 16439
rect 6736 16396 6788 16405
rect 7196 16396 7248 16448
rect 9772 16396 9824 16448
rect 12164 16473 12173 16507
rect 12173 16473 12207 16507
rect 12207 16473 12216 16507
rect 12164 16464 12216 16473
rect 13268 16507 13320 16516
rect 12808 16396 12860 16448
rect 13268 16473 13277 16507
rect 13277 16473 13311 16507
rect 13311 16473 13320 16507
rect 13268 16464 13320 16473
rect 13912 16464 13964 16516
rect 15108 16507 15160 16516
rect 15108 16473 15117 16507
rect 15117 16473 15151 16507
rect 15151 16473 15160 16507
rect 15108 16464 15160 16473
rect 13176 16396 13228 16448
rect 14464 16439 14516 16448
rect 14464 16405 14473 16439
rect 14473 16405 14507 16439
rect 14507 16405 14516 16439
rect 14464 16396 14516 16405
rect 3480 16294 3532 16346
rect 3544 16294 3596 16346
rect 3608 16294 3660 16346
rect 3672 16294 3724 16346
rect 8478 16294 8530 16346
rect 8542 16294 8594 16346
rect 8606 16294 8658 16346
rect 8670 16294 8722 16346
rect 13475 16294 13527 16346
rect 13539 16294 13591 16346
rect 13603 16294 13655 16346
rect 13667 16294 13719 16346
rect 1492 16235 1544 16244
rect 1492 16201 1501 16235
rect 1501 16201 1535 16235
rect 1535 16201 1544 16235
rect 1492 16192 1544 16201
rect 4804 16192 4856 16244
rect 5816 16192 5868 16244
rect 7012 16235 7064 16244
rect 7012 16201 7021 16235
rect 7021 16201 7055 16235
rect 7055 16201 7064 16235
rect 7012 16192 7064 16201
rect 7288 16235 7340 16244
rect 7288 16201 7297 16235
rect 7297 16201 7331 16235
rect 7331 16201 7340 16235
rect 7288 16192 7340 16201
rect 8944 16192 8996 16244
rect 13360 16192 13412 16244
rect 14556 16235 14608 16244
rect 14556 16201 14565 16235
rect 14565 16201 14599 16235
rect 14599 16201 14608 16235
rect 14556 16192 14608 16201
rect 14740 16235 14792 16244
rect 14740 16201 14749 16235
rect 14749 16201 14783 16235
rect 14783 16201 14792 16235
rect 14740 16192 14792 16201
rect 14924 16235 14976 16244
rect 14924 16201 14933 16235
rect 14933 16201 14967 16235
rect 14967 16201 14976 16235
rect 14924 16192 14976 16201
rect 940 16124 992 16176
rect 6460 16167 6512 16176
rect 6460 16133 6469 16167
rect 6469 16133 6503 16167
rect 6503 16133 6512 16167
rect 6460 16124 6512 16133
rect 12900 16124 12952 16176
rect 1952 16031 2004 16040
rect 1952 15997 1961 16031
rect 1961 15997 1995 16031
rect 1995 15997 2004 16031
rect 1952 15988 2004 15997
rect 2136 15988 2188 16040
rect 3884 15920 3936 15972
rect 2044 15852 2096 15904
rect 2412 15852 2464 15904
rect 2872 15852 2924 15904
rect 4712 15895 4764 15904
rect 4712 15861 4721 15895
rect 4721 15861 4755 15895
rect 4755 15861 4764 15895
rect 4712 15852 4764 15861
rect 6460 15988 6512 16040
rect 6736 15988 6788 16040
rect 6920 16031 6972 16040
rect 6920 15997 6929 16031
rect 6929 15997 6963 16031
rect 6963 15997 6972 16031
rect 6920 15988 6972 15997
rect 9220 16056 9272 16108
rect 7288 15852 7340 15904
rect 7564 15895 7616 15904
rect 7564 15861 7573 15895
rect 7573 15861 7607 15895
rect 7607 15861 7616 15895
rect 7564 15852 7616 15861
rect 9588 15988 9640 16040
rect 11520 15988 11572 16040
rect 15844 15988 15896 16040
rect 8208 15963 8260 15972
rect 8208 15929 8217 15963
rect 8217 15929 8251 15963
rect 8251 15929 8260 15963
rect 8208 15920 8260 15929
rect 9312 15920 9364 15972
rect 13820 15920 13872 15972
rect 16948 15920 17000 15972
rect 7748 15895 7800 15904
rect 7748 15861 7757 15895
rect 7757 15861 7791 15895
rect 7791 15861 7800 15895
rect 7748 15852 7800 15861
rect 7932 15852 7984 15904
rect 9496 15852 9548 15904
rect 10508 15852 10560 15904
rect 15384 15852 15436 15904
rect 5979 15750 6031 15802
rect 6043 15750 6095 15802
rect 6107 15750 6159 15802
rect 6171 15750 6223 15802
rect 10976 15750 11028 15802
rect 11040 15750 11092 15802
rect 11104 15750 11156 15802
rect 11168 15750 11220 15802
rect 2964 15648 3016 15700
rect 4160 15691 4212 15700
rect 4160 15657 4169 15691
rect 4169 15657 4203 15691
rect 4203 15657 4212 15691
rect 4160 15648 4212 15657
rect 4436 15648 4488 15700
rect 5172 15648 5224 15700
rect 5540 15691 5592 15700
rect 5540 15657 5549 15691
rect 5549 15657 5583 15691
rect 5583 15657 5592 15691
rect 5540 15648 5592 15657
rect 6736 15691 6788 15700
rect 6736 15657 6745 15691
rect 6745 15657 6779 15691
rect 6779 15657 6788 15691
rect 6736 15648 6788 15657
rect 7104 15648 7156 15700
rect 8300 15648 8352 15700
rect 9128 15691 9180 15700
rect 9128 15657 9137 15691
rect 9137 15657 9171 15691
rect 9171 15657 9180 15691
rect 9128 15648 9180 15657
rect 9404 15691 9456 15700
rect 9404 15657 9413 15691
rect 9413 15657 9447 15691
rect 9447 15657 9456 15691
rect 9404 15648 9456 15657
rect 9680 15691 9732 15700
rect 9680 15657 9689 15691
rect 9689 15657 9723 15691
rect 9723 15657 9732 15691
rect 9680 15648 9732 15657
rect 9956 15691 10008 15700
rect 9956 15657 9965 15691
rect 9965 15657 9999 15691
rect 9999 15657 10008 15691
rect 9956 15648 10008 15657
rect 15844 15648 15896 15700
rect 1400 15580 1452 15632
rect 4528 15580 4580 15632
rect 2780 15512 2832 15564
rect 4344 15555 4396 15564
rect 4344 15521 4353 15555
rect 4353 15521 4387 15555
rect 4387 15521 4396 15555
rect 4344 15512 4396 15521
rect 4712 15512 4764 15564
rect 7196 15580 7248 15632
rect 7932 15580 7984 15632
rect 6000 15512 6052 15564
rect 6184 15512 6236 15564
rect 7472 15512 7524 15564
rect 1400 15419 1452 15428
rect 1400 15385 1409 15419
rect 1409 15385 1443 15419
rect 1443 15385 1452 15419
rect 1400 15376 1452 15385
rect 4252 15376 4304 15428
rect 5908 15444 5960 15496
rect 7012 15487 7064 15496
rect 6092 15376 6144 15428
rect 7012 15453 7021 15487
rect 7021 15453 7055 15487
rect 7055 15453 7064 15487
rect 7012 15444 7064 15453
rect 6736 15376 6788 15428
rect 5816 15351 5868 15360
rect 5816 15317 5825 15351
rect 5825 15317 5859 15351
rect 5859 15317 5868 15351
rect 5816 15308 5868 15317
rect 6368 15351 6420 15360
rect 6368 15317 6377 15351
rect 6377 15317 6411 15351
rect 6411 15317 6420 15351
rect 6368 15308 6420 15317
rect 6920 15308 6972 15360
rect 7748 15512 7800 15564
rect 8208 15555 8260 15564
rect 8208 15521 8217 15555
rect 8217 15521 8251 15555
rect 8251 15521 8260 15555
rect 8208 15512 8260 15521
rect 8300 15512 8352 15564
rect 8668 15512 8720 15564
rect 11428 15580 11480 15632
rect 15200 15580 15252 15632
rect 9864 15555 9916 15564
rect 7656 15444 7708 15496
rect 8024 15444 8076 15496
rect 8852 15444 8904 15496
rect 9220 15444 9272 15496
rect 9496 15444 9548 15496
rect 9864 15521 9873 15555
rect 9873 15521 9907 15555
rect 9907 15521 9916 15555
rect 9864 15512 9916 15521
rect 10140 15555 10192 15564
rect 10140 15521 10149 15555
rect 10149 15521 10183 15555
rect 10183 15521 10192 15555
rect 10140 15512 10192 15521
rect 15384 15512 15436 15564
rect 11796 15444 11848 15496
rect 15476 15444 15528 15496
rect 12808 15376 12860 15428
rect 9864 15308 9916 15360
rect 10692 15308 10744 15360
rect 3480 15206 3532 15258
rect 3544 15206 3596 15258
rect 3608 15206 3660 15258
rect 3672 15206 3724 15258
rect 8478 15206 8530 15258
rect 8542 15206 8594 15258
rect 8606 15206 8658 15258
rect 8670 15206 8722 15258
rect 13475 15206 13527 15258
rect 13539 15206 13591 15258
rect 13603 15206 13655 15258
rect 13667 15206 13719 15258
rect 3332 15104 3384 15156
rect 7196 15104 7248 15156
rect 9036 15104 9088 15156
rect 9128 15104 9180 15156
rect 9864 15104 9916 15156
rect 5080 14968 5132 15020
rect 7656 15036 7708 15088
rect 6828 14968 6880 15020
rect 4344 14900 4396 14952
rect 5908 14943 5960 14952
rect 5908 14909 5917 14943
rect 5917 14909 5951 14943
rect 5951 14909 5960 14943
rect 5908 14900 5960 14909
rect 6368 14900 6420 14952
rect 2688 14764 2740 14816
rect 6552 14832 6604 14884
rect 4988 14764 5040 14816
rect 5264 14764 5316 14816
rect 5724 14764 5776 14816
rect 7472 14832 7524 14884
rect 10048 15036 10100 15088
rect 8024 14968 8076 15020
rect 8668 15011 8720 15020
rect 8668 14977 8677 15011
rect 8677 14977 8711 15011
rect 8711 14977 8720 15011
rect 8668 14968 8720 14977
rect 8760 14968 8812 15020
rect 12256 14900 12308 14952
rect 8392 14832 8444 14884
rect 7104 14764 7156 14816
rect 7748 14764 7800 14816
rect 9128 14764 9180 14816
rect 14372 14832 14424 14884
rect 14096 14764 14148 14816
rect 14556 14764 14608 14816
rect 5979 14662 6031 14714
rect 6043 14662 6095 14714
rect 6107 14662 6159 14714
rect 6171 14662 6223 14714
rect 10976 14662 11028 14714
rect 11040 14662 11092 14714
rect 11104 14662 11156 14714
rect 11168 14662 11220 14714
rect 4620 14603 4672 14612
rect 4620 14569 4629 14603
rect 4629 14569 4663 14603
rect 4663 14569 4672 14603
rect 4620 14560 4672 14569
rect 4988 14603 5040 14612
rect 4988 14569 4997 14603
rect 4997 14569 5031 14603
rect 5031 14569 5040 14603
rect 4988 14560 5040 14569
rect 2504 14424 2556 14476
rect 4068 14424 4120 14476
rect 6552 14424 6604 14476
rect 7656 14492 7708 14544
rect 7932 14492 7984 14544
rect 8392 14492 8444 14544
rect 9864 14560 9916 14612
rect 3792 14356 3844 14408
rect 5540 14399 5592 14408
rect 5540 14365 5549 14399
rect 5549 14365 5583 14399
rect 5583 14365 5592 14399
rect 5540 14356 5592 14365
rect 1400 14331 1452 14340
rect 1400 14297 1409 14331
rect 1409 14297 1443 14331
rect 1443 14297 1452 14331
rect 1400 14288 1452 14297
rect 4620 14288 4672 14340
rect 7656 14356 7708 14408
rect 6276 14288 6328 14340
rect 4528 14220 4580 14272
rect 5908 14263 5960 14272
rect 5908 14229 5917 14263
rect 5917 14229 5951 14263
rect 5951 14229 5960 14263
rect 5908 14220 5960 14229
rect 7380 14263 7432 14272
rect 7380 14229 7389 14263
rect 7389 14229 7423 14263
rect 7423 14229 7432 14263
rect 7380 14220 7432 14229
rect 7840 14288 7892 14340
rect 8024 14356 8076 14408
rect 8116 14288 8168 14340
rect 8944 14492 8996 14544
rect 9312 14492 9364 14544
rect 10508 14492 10560 14544
rect 8668 14356 8720 14408
rect 9956 14356 10008 14408
rect 9404 14331 9456 14340
rect 9404 14297 9413 14331
rect 9413 14297 9447 14331
rect 9447 14297 9456 14331
rect 9404 14288 9456 14297
rect 9680 14288 9732 14340
rect 10232 14288 10284 14340
rect 10876 14288 10928 14340
rect 8208 14220 8260 14272
rect 9036 14220 9088 14272
rect 9312 14220 9364 14272
rect 10048 14220 10100 14272
rect 10508 14220 10560 14272
rect 3480 14118 3532 14170
rect 3544 14118 3596 14170
rect 3608 14118 3660 14170
rect 3672 14118 3724 14170
rect 8478 14118 8530 14170
rect 8542 14118 8594 14170
rect 8606 14118 8658 14170
rect 8670 14118 8722 14170
rect 13475 14118 13527 14170
rect 13539 14118 13591 14170
rect 13603 14118 13655 14170
rect 13667 14118 13719 14170
rect 2504 14059 2556 14068
rect 2504 14025 2513 14059
rect 2513 14025 2547 14059
rect 2547 14025 2556 14059
rect 2504 14016 2556 14025
rect 2780 14059 2832 14068
rect 2780 14025 2789 14059
rect 2789 14025 2823 14059
rect 2823 14025 2832 14059
rect 2780 14016 2832 14025
rect 5540 14016 5592 14068
rect 9496 14016 9548 14068
rect 11336 14016 11388 14068
rect 3516 13880 3568 13932
rect 4528 13923 4580 13932
rect 4528 13889 4537 13923
rect 4537 13889 4571 13923
rect 4571 13889 4580 13923
rect 4528 13880 4580 13889
rect 4712 13923 4764 13932
rect 4712 13889 4721 13923
rect 4721 13889 4755 13923
rect 4755 13889 4764 13923
rect 4712 13880 4764 13889
rect 6276 13948 6328 14000
rect 7932 13991 7984 14000
rect 7932 13957 7941 13991
rect 7941 13957 7975 13991
rect 7975 13957 7984 13991
rect 7932 13948 7984 13957
rect 8208 13948 8260 14000
rect 14188 13948 14240 14000
rect 2964 13855 3016 13864
rect 2964 13821 2973 13855
rect 2973 13821 3007 13855
rect 3007 13821 3016 13855
rect 2964 13812 3016 13821
rect 4896 13855 4948 13864
rect 4896 13821 4905 13855
rect 4905 13821 4939 13855
rect 4939 13821 4948 13855
rect 4896 13812 4948 13821
rect 5908 13812 5960 13864
rect 2780 13744 2832 13796
rect 6276 13812 6328 13864
rect 6736 13812 6788 13864
rect 8116 13880 8168 13932
rect 9036 13880 9088 13932
rect 7104 13812 7156 13864
rect 7840 13855 7892 13864
rect 7840 13821 7849 13855
rect 7849 13821 7883 13855
rect 7883 13821 7892 13855
rect 7840 13812 7892 13821
rect 8392 13812 8444 13864
rect 12348 13880 12400 13932
rect 8208 13744 8260 13796
rect 2504 13676 2556 13728
rect 5632 13676 5684 13728
rect 7564 13676 7616 13728
rect 8484 13676 8536 13728
rect 8668 13744 8720 13796
rect 14280 13812 14332 13864
rect 14464 13812 14516 13864
rect 11704 13744 11756 13796
rect 8944 13676 8996 13728
rect 9128 13719 9180 13728
rect 9128 13685 9137 13719
rect 9137 13685 9171 13719
rect 9171 13685 9180 13719
rect 9128 13676 9180 13685
rect 9312 13676 9364 13728
rect 9680 13676 9732 13728
rect 10416 13719 10468 13728
rect 10416 13685 10425 13719
rect 10425 13685 10459 13719
rect 10459 13685 10468 13719
rect 10416 13676 10468 13685
rect 10508 13676 10560 13728
rect 14464 13676 14516 13728
rect 14832 13676 14884 13728
rect 5979 13574 6031 13626
rect 6043 13574 6095 13626
rect 6107 13574 6159 13626
rect 6171 13574 6223 13626
rect 10976 13574 11028 13626
rect 11040 13574 11092 13626
rect 11104 13574 11156 13626
rect 11168 13574 11220 13626
rect 3424 13515 3476 13524
rect 3424 13481 3433 13515
rect 3433 13481 3467 13515
rect 3467 13481 3476 13515
rect 3424 13472 3476 13481
rect 3884 13515 3936 13524
rect 3884 13481 3893 13515
rect 3893 13481 3927 13515
rect 3927 13481 3936 13515
rect 3884 13472 3936 13481
rect 4896 13472 4948 13524
rect 1400 13379 1452 13388
rect 1400 13345 1409 13379
rect 1409 13345 1443 13379
rect 1443 13345 1452 13379
rect 1400 13336 1452 13345
rect 2596 13336 2648 13388
rect 6828 13404 6880 13456
rect 7196 13447 7248 13456
rect 7196 13413 7230 13447
rect 7230 13413 7248 13447
rect 7196 13404 7248 13413
rect 8024 13404 8076 13456
rect 8392 13472 8444 13524
rect 8668 13472 8720 13524
rect 9036 13472 9088 13524
rect 9864 13472 9916 13524
rect 10232 13472 10284 13524
rect 10784 13472 10836 13524
rect 11612 13472 11664 13524
rect 8944 13404 8996 13456
rect 9404 13404 9456 13456
rect 9588 13404 9640 13456
rect 3056 13268 3108 13320
rect 3516 13311 3568 13320
rect 3516 13277 3525 13311
rect 3525 13277 3559 13311
rect 3559 13277 3568 13311
rect 3516 13268 3568 13277
rect 2136 13132 2188 13184
rect 4620 13336 4672 13388
rect 4252 13268 4304 13320
rect 5816 13268 5868 13320
rect 4160 13200 4212 13252
rect 4988 13132 5040 13184
rect 5448 13175 5500 13184
rect 5448 13141 5457 13175
rect 5457 13141 5491 13175
rect 5491 13141 5500 13175
rect 5448 13132 5500 13141
rect 7656 13132 7708 13184
rect 7840 13132 7892 13184
rect 8852 13336 8904 13388
rect 9772 13336 9824 13388
rect 11060 13404 11112 13456
rect 11336 13336 11388 13388
rect 8852 13200 8904 13252
rect 9128 13243 9180 13252
rect 9128 13209 9137 13243
rect 9137 13209 9171 13243
rect 9171 13209 9180 13243
rect 9128 13200 9180 13209
rect 9404 13268 9456 13320
rect 9864 13200 9916 13252
rect 12348 13268 12400 13320
rect 10508 13200 10560 13252
rect 11612 13200 11664 13252
rect 10048 13132 10100 13184
rect 11152 13175 11204 13184
rect 11152 13141 11161 13175
rect 11161 13141 11195 13175
rect 11195 13141 11204 13175
rect 11152 13132 11204 13141
rect 11244 13132 11296 13184
rect 11428 13132 11480 13184
rect 3480 13030 3532 13082
rect 3544 13030 3596 13082
rect 3608 13030 3660 13082
rect 3672 13030 3724 13082
rect 8478 13030 8530 13082
rect 8542 13030 8594 13082
rect 8606 13030 8658 13082
rect 8670 13030 8722 13082
rect 13475 13030 13527 13082
rect 13539 13030 13591 13082
rect 13603 13030 13655 13082
rect 13667 13030 13719 13082
rect 2596 12971 2648 12980
rect 2596 12937 2605 12971
rect 2605 12937 2639 12971
rect 2639 12937 2648 12971
rect 2596 12928 2648 12937
rect 2964 12860 3016 12912
rect 5632 12928 5684 12980
rect 7196 12928 7248 12980
rect 8116 12928 8168 12980
rect 9680 12928 9732 12980
rect 10048 12928 10100 12980
rect 11428 12971 11480 12980
rect 11428 12937 11437 12971
rect 11437 12937 11471 12971
rect 11471 12937 11480 12971
rect 11428 12928 11480 12937
rect 9128 12860 9180 12912
rect 10600 12860 10652 12912
rect 2136 12767 2188 12776
rect 2136 12733 2145 12767
rect 2145 12733 2179 12767
rect 2179 12733 2188 12767
rect 2136 12724 2188 12733
rect 2780 12724 2832 12776
rect 9036 12792 9088 12844
rect 14464 12860 14516 12912
rect 10876 12835 10928 12844
rect 10876 12801 10885 12835
rect 10885 12801 10919 12835
rect 10919 12801 10928 12835
rect 10876 12792 10928 12801
rect 11612 12792 11664 12844
rect 12440 12792 12492 12844
rect 3516 12656 3568 12708
rect 3608 12656 3660 12708
rect 4068 12656 4120 12708
rect 4528 12699 4580 12708
rect 4528 12665 4546 12699
rect 4546 12665 4580 12699
rect 4528 12656 4580 12665
rect 4896 12767 4948 12776
rect 4896 12733 4905 12767
rect 4905 12733 4939 12767
rect 4939 12733 4948 12767
rect 4896 12724 4948 12733
rect 6460 12767 6512 12776
rect 6460 12733 6469 12767
rect 6469 12733 6503 12767
rect 6503 12733 6512 12767
rect 6460 12724 6512 12733
rect 7656 12724 7708 12776
rect 7840 12724 7892 12776
rect 9680 12724 9732 12776
rect 9772 12767 9824 12776
rect 9772 12733 9781 12767
rect 9781 12733 9815 12767
rect 9815 12733 9824 12767
rect 9772 12724 9824 12733
rect 10416 12724 10468 12776
rect 12164 12724 12216 12776
rect 12256 12724 12308 12776
rect 14096 12724 14148 12776
rect 5448 12656 5500 12708
rect 5816 12656 5868 12708
rect 8024 12656 8076 12708
rect 8760 12656 8812 12708
rect 8944 12656 8996 12708
rect 9864 12699 9916 12708
rect 2044 12631 2096 12640
rect 2044 12597 2053 12631
rect 2053 12597 2087 12631
rect 2087 12597 2096 12631
rect 2044 12588 2096 12597
rect 4712 12588 4764 12640
rect 4988 12588 5040 12640
rect 9312 12588 9364 12640
rect 9864 12665 9873 12699
rect 9873 12665 9907 12699
rect 9907 12665 9916 12699
rect 9864 12656 9916 12665
rect 10600 12631 10652 12640
rect 10600 12597 10609 12631
rect 10609 12597 10643 12631
rect 10643 12597 10652 12631
rect 10600 12588 10652 12597
rect 10784 12588 10836 12640
rect 11244 12656 11296 12708
rect 11520 12656 11572 12708
rect 11980 12656 12032 12708
rect 12256 12588 12308 12640
rect 5979 12486 6031 12538
rect 6043 12486 6095 12538
rect 6107 12486 6159 12538
rect 6171 12486 6223 12538
rect 10976 12486 11028 12538
rect 11040 12486 11092 12538
rect 11104 12486 11156 12538
rect 11168 12486 11220 12538
rect 1400 12359 1452 12368
rect 1400 12325 1409 12359
rect 1409 12325 1443 12359
rect 1443 12325 1452 12359
rect 1400 12316 1452 12325
rect 3608 12384 3660 12436
rect 3884 12384 3936 12436
rect 4068 12427 4120 12436
rect 4068 12393 4077 12427
rect 4077 12393 4111 12427
rect 4111 12393 4120 12427
rect 4068 12384 4120 12393
rect 4436 12384 4488 12436
rect 5264 12384 5316 12436
rect 5816 12384 5868 12436
rect 4160 12316 4212 12368
rect 5908 12316 5960 12368
rect 3148 12248 3200 12300
rect 2320 12223 2372 12232
rect 2320 12189 2329 12223
rect 2329 12189 2363 12223
rect 2363 12189 2372 12223
rect 2320 12180 2372 12189
rect 2412 12223 2464 12232
rect 2412 12189 2421 12223
rect 2421 12189 2455 12223
rect 2455 12189 2464 12223
rect 2412 12180 2464 12189
rect 3240 12223 3292 12232
rect 2596 12112 2648 12164
rect 3240 12189 3249 12223
rect 3249 12189 3283 12223
rect 3283 12189 3292 12223
rect 3240 12180 3292 12189
rect 4344 12180 4396 12232
rect 3148 12112 3200 12164
rect 6736 12384 6788 12436
rect 6828 12384 6880 12436
rect 7748 12384 7800 12436
rect 10692 12384 10744 12436
rect 11428 12384 11480 12436
rect 11796 12427 11848 12436
rect 11796 12393 11805 12427
rect 11805 12393 11839 12427
rect 11839 12393 11848 12427
rect 11796 12384 11848 12393
rect 12256 12427 12308 12436
rect 12256 12393 12265 12427
rect 12265 12393 12299 12427
rect 12299 12393 12308 12427
rect 12256 12384 12308 12393
rect 12716 12427 12768 12436
rect 12716 12393 12725 12427
rect 12725 12393 12759 12427
rect 12759 12393 12768 12427
rect 12716 12384 12768 12393
rect 12992 12384 13044 12436
rect 13268 12384 13320 12436
rect 4528 12180 4580 12232
rect 5908 12180 5960 12232
rect 7196 12291 7248 12300
rect 7196 12257 7214 12291
rect 7214 12257 7248 12291
rect 7196 12248 7248 12257
rect 7656 12248 7708 12300
rect 8852 12248 8904 12300
rect 9312 12316 9364 12368
rect 9956 12248 10008 12300
rect 7932 12044 7984 12096
rect 10968 12180 11020 12232
rect 11796 12180 11848 12232
rect 12348 12180 12400 12232
rect 9312 12044 9364 12096
rect 9496 12044 9548 12096
rect 11244 12044 11296 12096
rect 11428 12087 11480 12096
rect 11428 12053 11437 12087
rect 11437 12053 11471 12087
rect 11471 12053 11480 12087
rect 11428 12044 11480 12053
rect 11796 12044 11848 12096
rect 12072 12044 12124 12096
rect 13360 12044 13412 12096
rect 14004 12044 14056 12096
rect 14648 12044 14700 12096
rect 3480 11942 3532 11994
rect 3544 11942 3596 11994
rect 3608 11942 3660 11994
rect 3672 11942 3724 11994
rect 8478 11942 8530 11994
rect 8542 11942 8594 11994
rect 8606 11942 8658 11994
rect 8670 11942 8722 11994
rect 13475 11942 13527 11994
rect 13539 11942 13591 11994
rect 13603 11942 13655 11994
rect 13667 11942 13719 11994
rect 2044 11840 2096 11892
rect 3792 11840 3844 11892
rect 3976 11883 4028 11892
rect 3976 11849 3985 11883
rect 3985 11849 4019 11883
rect 4019 11849 4028 11883
rect 3976 11840 4028 11849
rect 7932 11883 7984 11892
rect 7932 11849 7941 11883
rect 7941 11849 7975 11883
rect 7975 11849 7984 11883
rect 7932 11840 7984 11849
rect 11336 11840 11388 11892
rect 11704 11883 11756 11892
rect 11704 11849 11713 11883
rect 11713 11849 11747 11883
rect 11747 11849 11756 11883
rect 11704 11840 11756 11849
rect 12532 11883 12584 11892
rect 12532 11849 12541 11883
rect 12541 11849 12575 11883
rect 12575 11849 12584 11883
rect 12532 11840 12584 11849
rect 13360 11883 13412 11892
rect 13360 11849 13369 11883
rect 13369 11849 13403 11883
rect 13403 11849 13412 11883
rect 13360 11840 13412 11849
rect 3056 11747 3108 11756
rect 3056 11713 3065 11747
rect 3065 11713 3099 11747
rect 3099 11713 3108 11747
rect 3056 11704 3108 11713
rect 3148 11704 3200 11756
rect 4344 11704 4396 11756
rect 4804 11772 4856 11824
rect 4620 11747 4672 11756
rect 4620 11713 4629 11747
rect 4629 11713 4663 11747
rect 4663 11713 4672 11747
rect 6460 11747 6512 11756
rect 4620 11704 4672 11713
rect 4528 11636 4580 11688
rect 4896 11679 4948 11688
rect 4896 11645 4905 11679
rect 4905 11645 4939 11679
rect 4939 11645 4948 11679
rect 4896 11636 4948 11645
rect 6460 11713 6469 11747
rect 6469 11713 6503 11747
rect 6503 11713 6512 11747
rect 6460 11704 6512 11713
rect 9312 11747 9364 11756
rect 9312 11713 9321 11747
rect 9321 11713 9355 11747
rect 9355 11713 9364 11747
rect 9312 11704 9364 11713
rect 9680 11704 9732 11756
rect 5448 11636 5500 11688
rect 8300 11636 8352 11688
rect 9036 11679 9088 11688
rect 10232 11772 10284 11824
rect 9036 11645 9054 11679
rect 9054 11645 9088 11679
rect 9036 11636 9088 11645
rect 1952 11611 2004 11620
rect 1952 11577 1961 11611
rect 1961 11577 1995 11611
rect 1995 11577 2004 11611
rect 1952 11568 2004 11577
rect 2228 11500 2280 11552
rect 3332 11568 3384 11620
rect 4344 11568 4396 11620
rect 5816 11568 5868 11620
rect 3608 11543 3660 11552
rect 3608 11509 3617 11543
rect 3617 11509 3651 11543
rect 3651 11509 3660 11543
rect 3608 11500 3660 11509
rect 4068 11543 4120 11552
rect 4068 11509 4077 11543
rect 4077 11509 4111 11543
rect 4111 11509 4120 11543
rect 4068 11500 4120 11509
rect 4528 11543 4580 11552
rect 4528 11509 4537 11543
rect 4537 11509 4571 11543
rect 4571 11509 4580 11543
rect 4528 11500 4580 11509
rect 4804 11500 4856 11552
rect 10600 11704 10652 11756
rect 11980 11772 12032 11824
rect 12440 11772 12492 11824
rect 12992 11772 13044 11824
rect 11244 11704 11296 11756
rect 11612 11704 11664 11756
rect 12716 11704 12768 11756
rect 14004 11704 14056 11756
rect 11060 11679 11112 11688
rect 11060 11645 11069 11679
rect 11069 11645 11103 11679
rect 11103 11645 11112 11679
rect 11060 11636 11112 11645
rect 11428 11636 11480 11688
rect 7840 11543 7892 11552
rect 7840 11509 7849 11543
rect 7849 11509 7883 11543
rect 7883 11509 7892 11543
rect 7840 11500 7892 11509
rect 8392 11500 8444 11552
rect 8852 11500 8904 11552
rect 9404 11543 9456 11552
rect 9404 11509 9413 11543
rect 9413 11509 9447 11543
rect 9447 11509 9456 11543
rect 9404 11500 9456 11509
rect 9496 11500 9548 11552
rect 10232 11543 10284 11552
rect 10232 11509 10241 11543
rect 10241 11509 10275 11543
rect 10275 11509 10284 11543
rect 10232 11500 10284 11509
rect 10692 11543 10744 11552
rect 10692 11509 10701 11543
rect 10701 11509 10735 11543
rect 10735 11509 10744 11543
rect 10692 11500 10744 11509
rect 10876 11500 10928 11552
rect 14740 11636 14792 11688
rect 12624 11568 12676 11620
rect 13176 11568 13228 11620
rect 14648 11568 14700 11620
rect 11704 11500 11756 11552
rect 13084 11500 13136 11552
rect 14464 11500 14516 11552
rect 5979 11398 6031 11450
rect 6043 11398 6095 11450
rect 6107 11398 6159 11450
rect 6171 11398 6223 11450
rect 10976 11398 11028 11450
rect 11040 11398 11092 11450
rect 11104 11398 11156 11450
rect 11168 11398 11220 11450
rect 1492 11339 1544 11348
rect 1492 11305 1501 11339
rect 1501 11305 1535 11339
rect 1535 11305 1544 11339
rect 1492 11296 1544 11305
rect 4068 11296 4120 11348
rect 4160 11296 4212 11348
rect 9496 11296 9548 11348
rect 10784 11296 10836 11348
rect 11520 11296 11572 11348
rect 11980 11296 12032 11348
rect 14372 11339 14424 11348
rect 14372 11305 14381 11339
rect 14381 11305 14415 11339
rect 14415 11305 14424 11339
rect 14372 11296 14424 11305
rect 14740 11339 14792 11348
rect 14740 11305 14749 11339
rect 14749 11305 14783 11339
rect 14783 11305 14792 11339
rect 14740 11296 14792 11305
rect 15292 11339 15344 11348
rect 15292 11305 15301 11339
rect 15301 11305 15335 11339
rect 15335 11305 15344 11339
rect 15292 11296 15344 11305
rect 3608 11228 3660 11280
rect 2504 11203 2556 11212
rect 2504 11169 2513 11203
rect 2513 11169 2547 11203
rect 2547 11169 2556 11203
rect 2504 11160 2556 11169
rect 3332 11203 3384 11212
rect 3332 11169 3341 11203
rect 3341 11169 3375 11203
rect 3375 11169 3384 11203
rect 3332 11160 3384 11169
rect 2596 11135 2648 11144
rect 2596 11101 2605 11135
rect 2605 11101 2639 11135
rect 2639 11101 2648 11135
rect 2596 11092 2648 11101
rect 4804 11160 4856 11212
rect 5264 11160 5316 11212
rect 2136 10999 2188 11008
rect 2136 10965 2145 10999
rect 2145 10965 2179 10999
rect 2179 10965 2188 10999
rect 2136 10956 2188 10965
rect 5540 11092 5592 11144
rect 3792 11024 3844 11076
rect 6460 11228 6512 11280
rect 6276 11160 6328 11212
rect 7840 11228 7892 11280
rect 8208 11228 8260 11280
rect 9956 11228 10008 11280
rect 10692 11228 10744 11280
rect 10876 11228 10928 11280
rect 10968 11228 11020 11280
rect 4436 10956 4488 11008
rect 4620 10956 4672 11008
rect 7196 11024 7248 11076
rect 7932 10956 7984 11008
rect 9588 11160 9640 11212
rect 11060 11160 11112 11212
rect 11980 11203 12032 11212
rect 11980 11169 11989 11203
rect 11989 11169 12023 11203
rect 12023 11169 12032 11203
rect 11980 11160 12032 11169
rect 9772 11135 9824 11144
rect 9772 11101 9781 11135
rect 9781 11101 9815 11135
rect 9815 11101 9824 11135
rect 9772 11092 9824 11101
rect 10600 11135 10652 11144
rect 10600 11101 10609 11135
rect 10609 11101 10643 11135
rect 10643 11101 10652 11135
rect 10600 11092 10652 11101
rect 10876 11092 10928 11144
rect 11520 11092 11572 11144
rect 11888 11135 11940 11144
rect 11888 11101 11897 11135
rect 11897 11101 11931 11135
rect 11931 11101 11940 11135
rect 11888 11092 11940 11101
rect 12256 11228 12308 11280
rect 12532 11228 12584 11280
rect 12992 11228 13044 11280
rect 13176 11228 13228 11280
rect 12716 11092 12768 11144
rect 14740 11160 14792 11212
rect 13268 11092 13320 11144
rect 10324 11024 10376 11076
rect 12164 11024 12216 11076
rect 12440 11067 12492 11076
rect 12440 11033 12449 11067
rect 12449 11033 12483 11067
rect 12483 11033 12492 11067
rect 12440 11024 12492 11033
rect 9496 10956 9548 11008
rect 9588 10956 9640 11008
rect 9772 10956 9824 11008
rect 9956 10999 10008 11008
rect 9956 10965 9965 10999
rect 9965 10965 9999 10999
rect 9999 10965 10008 10999
rect 9956 10956 10008 10965
rect 10784 10999 10836 11008
rect 10784 10965 10793 10999
rect 10793 10965 10827 10999
rect 10827 10965 10836 10999
rect 10784 10956 10836 10965
rect 11612 10956 11664 11008
rect 13360 10956 13412 11008
rect 14004 11024 14056 11076
rect 14556 11024 14608 11076
rect 15108 10956 15160 11008
rect 3480 10854 3532 10906
rect 3544 10854 3596 10906
rect 3608 10854 3660 10906
rect 3672 10854 3724 10906
rect 8478 10854 8530 10906
rect 8542 10854 8594 10906
rect 8606 10854 8658 10906
rect 8670 10854 8722 10906
rect 13475 10854 13527 10906
rect 13539 10854 13591 10906
rect 13603 10854 13655 10906
rect 13667 10854 13719 10906
rect 2596 10752 2648 10804
rect 3332 10795 3384 10804
rect 3332 10761 3341 10795
rect 3341 10761 3375 10795
rect 3375 10761 3384 10795
rect 3332 10752 3384 10761
rect 2688 10616 2740 10668
rect 9496 10752 9548 10804
rect 10692 10752 10744 10804
rect 11060 10795 11112 10804
rect 11060 10761 11069 10795
rect 11069 10761 11103 10795
rect 11103 10761 11112 10795
rect 11060 10752 11112 10761
rect 11428 10795 11480 10804
rect 11428 10761 11437 10795
rect 11437 10761 11471 10795
rect 11471 10761 11480 10795
rect 11428 10752 11480 10761
rect 12072 10752 12124 10804
rect 12624 10752 12676 10804
rect 12808 10752 12860 10804
rect 13084 10752 13136 10804
rect 14188 10795 14240 10804
rect 14188 10761 14197 10795
rect 14197 10761 14231 10795
rect 14231 10761 14240 10795
rect 14188 10752 14240 10761
rect 9312 10727 9364 10736
rect 4896 10659 4948 10668
rect 4896 10625 4905 10659
rect 4905 10625 4939 10659
rect 4939 10625 4948 10659
rect 4896 10616 4948 10625
rect 5908 10616 5960 10668
rect 9312 10693 9321 10727
rect 9321 10693 9355 10727
rect 9355 10693 9364 10727
rect 9312 10684 9364 10693
rect 1860 10480 1912 10532
rect 3240 10480 3292 10532
rect 3424 10591 3476 10600
rect 3424 10557 3433 10591
rect 3433 10557 3467 10591
rect 3467 10557 3476 10591
rect 3424 10548 3476 10557
rect 4620 10548 4672 10600
rect 4804 10548 4856 10600
rect 3792 10480 3844 10532
rect 3976 10480 4028 10532
rect 4436 10480 4488 10532
rect 5540 10548 5592 10600
rect 7932 10591 7984 10600
rect 7932 10557 7941 10591
rect 7941 10557 7975 10591
rect 7975 10557 7984 10591
rect 7932 10548 7984 10557
rect 9128 10616 9180 10668
rect 9772 10684 9824 10736
rect 10600 10684 10652 10736
rect 9680 10616 9732 10668
rect 5908 10480 5960 10532
rect 6552 10480 6604 10532
rect 8024 10480 8076 10532
rect 8668 10548 8720 10600
rect 9588 10548 9640 10600
rect 10232 10616 10284 10668
rect 10876 10659 10928 10668
rect 10876 10625 10885 10659
rect 10885 10625 10919 10659
rect 10919 10625 10928 10659
rect 10876 10616 10928 10625
rect 10416 10548 10468 10600
rect 11244 10727 11296 10736
rect 11244 10693 11253 10727
rect 11253 10693 11287 10727
rect 11287 10693 11296 10727
rect 11244 10684 11296 10693
rect 11612 10616 11664 10668
rect 12900 10684 12952 10736
rect 13912 10684 13964 10736
rect 12624 10616 12676 10668
rect 14740 10659 14792 10668
rect 14740 10625 14749 10659
rect 14749 10625 14783 10659
rect 14783 10625 14792 10659
rect 14740 10616 14792 10625
rect 14004 10548 14056 10600
rect 14096 10548 14148 10600
rect 1492 10455 1544 10464
rect 1492 10421 1501 10455
rect 1501 10421 1535 10455
rect 1535 10421 1544 10455
rect 1492 10412 1544 10421
rect 2044 10455 2096 10464
rect 2044 10421 2053 10455
rect 2053 10421 2087 10455
rect 2087 10421 2096 10455
rect 2044 10412 2096 10421
rect 4160 10412 4212 10464
rect 4988 10412 5040 10464
rect 6276 10412 6328 10464
rect 8668 10412 8720 10464
rect 8852 10412 8904 10464
rect 10324 10412 10376 10464
rect 12256 10480 12308 10532
rect 13268 10480 13320 10532
rect 13360 10480 13412 10532
rect 12440 10455 12492 10464
rect 12440 10421 12449 10455
rect 12449 10421 12483 10455
rect 12483 10421 12492 10455
rect 12440 10412 12492 10421
rect 12808 10412 12860 10464
rect 13728 10412 13780 10464
rect 14096 10455 14148 10464
rect 14096 10421 14105 10455
rect 14105 10421 14139 10455
rect 14139 10421 14148 10455
rect 14096 10412 14148 10421
rect 14556 10412 14608 10464
rect 5979 10310 6031 10362
rect 6043 10310 6095 10362
rect 6107 10310 6159 10362
rect 6171 10310 6223 10362
rect 10976 10310 11028 10362
rect 11040 10310 11092 10362
rect 11104 10310 11156 10362
rect 11168 10310 11220 10362
rect 1860 10251 1912 10260
rect 1860 10217 1869 10251
rect 1869 10217 1903 10251
rect 1903 10217 1912 10251
rect 1860 10208 1912 10217
rect 2044 10208 2096 10260
rect 2412 10072 2464 10124
rect 2688 10072 2740 10124
rect 2596 10047 2648 10056
rect 2596 10013 2605 10047
rect 2605 10013 2639 10047
rect 2639 10013 2648 10047
rect 2596 10004 2648 10013
rect 4528 10208 4580 10260
rect 4620 10208 4672 10260
rect 5264 10208 5316 10260
rect 5632 10208 5684 10260
rect 4436 10140 4488 10192
rect 6460 10140 6512 10192
rect 3148 10072 3200 10124
rect 3700 10072 3752 10124
rect 3884 10072 3936 10124
rect 4528 10072 4580 10124
rect 5080 10072 5132 10124
rect 5816 10072 5868 10124
rect 8300 10208 8352 10260
rect 9404 10208 9456 10260
rect 9956 10208 10008 10260
rect 10232 10208 10284 10260
rect 8944 10140 8996 10192
rect 9036 10140 9088 10192
rect 2872 10004 2924 10056
rect 3056 10004 3108 10056
rect 4160 10004 4212 10056
rect 5172 10047 5224 10056
rect 1584 9936 1636 9988
rect 1768 9911 1820 9920
rect 1768 9877 1777 9911
rect 1777 9877 1811 9911
rect 1811 9877 1820 9911
rect 1768 9868 1820 9877
rect 2872 9868 2924 9920
rect 4712 9936 4764 9988
rect 4528 9868 4580 9920
rect 5172 10013 5181 10047
rect 5181 10013 5215 10047
rect 5215 10013 5224 10047
rect 5172 10004 5224 10013
rect 8668 10047 8720 10056
rect 6276 9868 6328 9920
rect 6552 9911 6604 9920
rect 6552 9877 6561 9911
rect 6561 9877 6595 9911
rect 6595 9877 6604 9911
rect 6552 9868 6604 9877
rect 8668 10013 8677 10047
rect 8677 10013 8711 10047
rect 8711 10013 8720 10047
rect 8668 10004 8720 10013
rect 8852 10072 8904 10124
rect 9128 10004 9180 10056
rect 10416 10072 10468 10124
rect 10140 10004 10192 10056
rect 10784 10140 10836 10192
rect 11060 10072 11112 10124
rect 12256 10208 12308 10260
rect 12072 10183 12124 10192
rect 12072 10149 12081 10183
rect 12081 10149 12115 10183
rect 12115 10149 12124 10183
rect 12072 10140 12124 10149
rect 11980 10072 12032 10124
rect 12348 10072 12400 10124
rect 12532 10208 12584 10260
rect 13268 10251 13320 10260
rect 13268 10217 13277 10251
rect 13277 10217 13311 10251
rect 13311 10217 13320 10251
rect 13268 10208 13320 10217
rect 13820 10208 13872 10260
rect 14096 10208 14148 10260
rect 12440 10004 12492 10056
rect 8024 9979 8076 9988
rect 8024 9945 8033 9979
rect 8033 9945 8067 9979
rect 8067 9945 8076 9979
rect 8024 9936 8076 9945
rect 7932 9868 7984 9920
rect 9036 9868 9088 9920
rect 9312 9868 9364 9920
rect 9680 9868 9732 9920
rect 10048 9868 10100 9920
rect 10508 9936 10560 9988
rect 11244 9936 11296 9988
rect 12716 9936 12768 9988
rect 10600 9868 10652 9920
rect 11060 9868 11112 9920
rect 11152 9868 11204 9920
rect 13268 10072 13320 10124
rect 14280 10140 14332 10192
rect 13912 10072 13964 10124
rect 14188 10072 14240 10124
rect 15476 10115 15528 10124
rect 15476 10081 15485 10115
rect 15485 10081 15519 10115
rect 15519 10081 15528 10115
rect 15476 10072 15528 10081
rect 13452 10004 13504 10056
rect 14832 10004 14884 10056
rect 14372 9979 14424 9988
rect 14372 9945 14381 9979
rect 14381 9945 14415 9979
rect 14415 9945 14424 9979
rect 14372 9936 14424 9945
rect 15660 9979 15712 9988
rect 15660 9945 15669 9979
rect 15669 9945 15703 9979
rect 15703 9945 15712 9979
rect 15660 9936 15712 9945
rect 14004 9868 14056 9920
rect 3480 9766 3532 9818
rect 3544 9766 3596 9818
rect 3608 9766 3660 9818
rect 3672 9766 3724 9818
rect 8478 9766 8530 9818
rect 8542 9766 8594 9818
rect 8606 9766 8658 9818
rect 8670 9766 8722 9818
rect 13475 9766 13527 9818
rect 13539 9766 13591 9818
rect 13603 9766 13655 9818
rect 13667 9766 13719 9818
rect 2228 9596 2280 9648
rect 2780 9596 2832 9648
rect 3240 9664 3292 9716
rect 11244 9664 11296 9716
rect 11612 9664 11664 9716
rect 11704 9707 11756 9716
rect 11704 9673 11713 9707
rect 11713 9673 11747 9707
rect 11747 9673 11756 9707
rect 11704 9664 11756 9673
rect 11980 9664 12032 9716
rect 12900 9664 12952 9716
rect 3332 9596 3384 9648
rect 2320 9528 2372 9580
rect 2872 9528 2924 9580
rect 3240 9571 3292 9580
rect 3240 9537 3249 9571
rect 3249 9537 3283 9571
rect 3283 9537 3292 9571
rect 3240 9528 3292 9537
rect 4620 9596 4672 9648
rect 6276 9639 6328 9648
rect 6276 9605 6285 9639
rect 6285 9605 6319 9639
rect 6319 9605 6328 9639
rect 6276 9596 6328 9605
rect 6460 9639 6512 9648
rect 6460 9605 6469 9639
rect 6469 9605 6503 9639
rect 6503 9605 6512 9639
rect 6460 9596 6512 9605
rect 1400 9503 1452 9512
rect 1400 9469 1409 9503
rect 1409 9469 1443 9503
rect 1443 9469 1452 9503
rect 1400 9460 1452 9469
rect 4436 9528 4488 9580
rect 4896 9503 4948 9512
rect 4896 9469 4905 9503
rect 4905 9469 4939 9503
rect 4939 9469 4948 9503
rect 4896 9460 4948 9469
rect 6552 9528 6604 9580
rect 7656 9596 7708 9648
rect 9404 9596 9456 9648
rect 10508 9596 10560 9648
rect 12164 9571 12216 9580
rect 1860 9392 1912 9444
rect 2964 9367 3016 9376
rect 2964 9333 2973 9367
rect 2973 9333 3007 9367
rect 3007 9333 3016 9367
rect 2964 9324 3016 9333
rect 3056 9367 3108 9376
rect 3056 9333 3065 9367
rect 3065 9333 3099 9367
rect 3099 9333 3108 9367
rect 4252 9392 4304 9444
rect 3056 9324 3108 9333
rect 4804 9324 4856 9376
rect 5448 9324 5500 9376
rect 5540 9324 5592 9376
rect 6828 9367 6880 9376
rect 6828 9333 6837 9367
rect 6837 9333 6871 9367
rect 6871 9333 6880 9367
rect 6828 9324 6880 9333
rect 7472 9324 7524 9376
rect 7840 9460 7892 9512
rect 9128 9460 9180 9512
rect 9036 9392 9088 9444
rect 9312 9392 9364 9444
rect 11152 9460 11204 9512
rect 11336 9503 11388 9512
rect 11336 9469 11345 9503
rect 11345 9469 11379 9503
rect 11379 9469 11388 9503
rect 11336 9460 11388 9469
rect 9588 9392 9640 9444
rect 9772 9392 9824 9444
rect 10968 9392 11020 9444
rect 12164 9537 12173 9571
rect 12173 9537 12207 9571
rect 12207 9537 12216 9571
rect 12164 9528 12216 9537
rect 12348 9571 12400 9580
rect 12348 9537 12357 9571
rect 12357 9537 12391 9571
rect 12391 9537 12400 9571
rect 12348 9528 12400 9537
rect 12256 9460 12308 9512
rect 12532 9528 12584 9580
rect 12716 9528 12768 9580
rect 15476 9664 15528 9716
rect 14280 9571 14332 9580
rect 14280 9537 14289 9571
rect 14289 9537 14323 9571
rect 14323 9537 14332 9571
rect 14280 9528 14332 9537
rect 12808 9503 12860 9512
rect 12808 9469 12817 9503
rect 12817 9469 12851 9503
rect 12851 9469 12860 9503
rect 12808 9460 12860 9469
rect 15108 9460 15160 9512
rect 11888 9324 11940 9376
rect 12900 9367 12952 9376
rect 12900 9333 12909 9367
rect 12909 9333 12943 9367
rect 12943 9333 12952 9367
rect 15476 9435 15528 9444
rect 15476 9401 15485 9435
rect 15485 9401 15519 9435
rect 15519 9401 15528 9435
rect 15476 9392 15528 9401
rect 12900 9324 12952 9333
rect 13728 9367 13780 9376
rect 13728 9333 13737 9367
rect 13737 9333 13771 9367
rect 13771 9333 13780 9367
rect 13728 9324 13780 9333
rect 14464 9367 14516 9376
rect 14464 9333 14473 9367
rect 14473 9333 14507 9367
rect 14507 9333 14516 9367
rect 14464 9324 14516 9333
rect 14740 9324 14792 9376
rect 15108 9324 15160 9376
rect 5979 9222 6031 9274
rect 6043 9222 6095 9274
rect 6107 9222 6159 9274
rect 6171 9222 6223 9274
rect 10976 9222 11028 9274
rect 11040 9222 11092 9274
rect 11104 9222 11156 9274
rect 11168 9222 11220 9274
rect 1492 9163 1544 9172
rect 1492 9129 1501 9163
rect 1501 9129 1535 9163
rect 1535 9129 1544 9163
rect 1492 9120 1544 9129
rect 1860 9163 1912 9172
rect 1860 9129 1869 9163
rect 1869 9129 1903 9163
rect 1903 9129 1912 9163
rect 1860 9120 1912 9129
rect 3056 9120 3108 9172
rect 3608 9120 3660 9172
rect 3976 9163 4028 9172
rect 3976 9129 3985 9163
rect 3985 9129 4019 9163
rect 4019 9129 4028 9163
rect 3976 9120 4028 9129
rect 2964 9052 3016 9104
rect 4988 9052 5040 9104
rect 6276 9052 6328 9104
rect 7932 9052 7984 9104
rect 1584 9027 1636 9036
rect 1584 8993 1593 9027
rect 1593 8993 1627 9027
rect 1627 8993 1636 9027
rect 1584 8984 1636 8993
rect 2136 8984 2188 9036
rect 2412 9027 2464 9036
rect 2412 8993 2421 9027
rect 2421 8993 2455 9027
rect 2455 8993 2464 9027
rect 2412 8984 2464 8993
rect 2504 9027 2556 9036
rect 2504 8993 2513 9027
rect 2513 8993 2547 9027
rect 2547 8993 2556 9027
rect 2504 8984 2556 8993
rect 4068 8984 4120 9036
rect 4344 8984 4396 9036
rect 1860 8780 1912 8832
rect 2136 8780 2188 8832
rect 3240 8848 3292 8900
rect 4160 8916 4212 8968
rect 5356 8959 5408 8968
rect 5356 8925 5365 8959
rect 5365 8925 5399 8959
rect 5399 8925 5408 8959
rect 5356 8916 5408 8925
rect 4344 8848 4396 8900
rect 8208 8984 8260 9036
rect 9772 9120 9824 9172
rect 10784 9120 10836 9172
rect 11336 9163 11388 9172
rect 9312 9052 9364 9104
rect 9496 9052 9548 9104
rect 11060 9052 11112 9104
rect 4160 8780 4212 8832
rect 5172 8780 5224 8832
rect 6920 8823 6972 8832
rect 6920 8789 6929 8823
rect 6929 8789 6963 8823
rect 6963 8789 6972 8823
rect 6920 8780 6972 8789
rect 7932 8780 7984 8832
rect 9036 8916 9088 8968
rect 9128 8959 9180 8968
rect 9128 8925 9137 8959
rect 9137 8925 9171 8959
rect 9171 8925 9180 8959
rect 9128 8916 9180 8925
rect 10508 8984 10560 9036
rect 10968 9027 11020 9036
rect 10600 8916 10652 8968
rect 10968 8993 10977 9027
rect 10977 8993 11011 9027
rect 11011 8993 11020 9027
rect 10968 8984 11020 8993
rect 11336 9129 11345 9163
rect 11345 9129 11379 9163
rect 11379 9129 11388 9163
rect 11336 9120 11388 9129
rect 11244 9052 11296 9104
rect 11980 9120 12032 9172
rect 12624 9120 12676 9172
rect 12808 9120 12860 9172
rect 13452 9120 13504 9172
rect 13912 9120 13964 9172
rect 14740 9163 14792 9172
rect 14740 9129 14749 9163
rect 14749 9129 14783 9163
rect 14783 9129 14792 9163
rect 14740 9120 14792 9129
rect 11336 8916 11388 8968
rect 11520 8959 11572 8968
rect 11520 8925 11529 8959
rect 11529 8925 11563 8959
rect 11563 8925 11572 8959
rect 11520 8916 11572 8925
rect 11704 8984 11756 9036
rect 11888 8984 11940 9036
rect 12348 8916 12400 8968
rect 12716 8959 12768 8968
rect 12716 8925 12725 8959
rect 12725 8925 12759 8959
rect 12759 8925 12768 8959
rect 12900 8959 12952 8968
rect 12716 8916 12768 8925
rect 12900 8925 12909 8959
rect 12909 8925 12943 8959
rect 12943 8925 12952 8959
rect 12900 8916 12952 8925
rect 13360 8916 13412 8968
rect 13820 8916 13872 8968
rect 12992 8848 13044 8900
rect 13452 8848 13504 8900
rect 14832 8959 14884 8968
rect 14832 8925 14841 8959
rect 14841 8925 14875 8959
rect 14875 8925 14884 8959
rect 14832 8916 14884 8925
rect 15200 8984 15252 9036
rect 14372 8848 14424 8900
rect 8852 8780 8904 8832
rect 9496 8780 9548 8832
rect 12532 8780 12584 8832
rect 13360 8780 13412 8832
rect 14096 8823 14148 8832
rect 14096 8789 14105 8823
rect 14105 8789 14139 8823
rect 14139 8789 14148 8823
rect 14096 8780 14148 8789
rect 3480 8678 3532 8730
rect 3544 8678 3596 8730
rect 3608 8678 3660 8730
rect 3672 8678 3724 8730
rect 8478 8678 8530 8730
rect 8542 8678 8594 8730
rect 8606 8678 8658 8730
rect 8670 8678 8722 8730
rect 13475 8678 13527 8730
rect 13539 8678 13591 8730
rect 13603 8678 13655 8730
rect 13667 8678 13719 8730
rect 1860 8576 1912 8628
rect 2228 8576 2280 8628
rect 3332 8508 3384 8560
rect 3240 8483 3292 8492
rect 3240 8449 3249 8483
rect 3249 8449 3283 8483
rect 3283 8449 3292 8483
rect 3240 8440 3292 8449
rect 2136 8415 2188 8424
rect 2136 8381 2145 8415
rect 2145 8381 2179 8415
rect 2179 8381 2188 8415
rect 2136 8372 2188 8381
rect 2320 8372 2372 8424
rect 4896 8415 4948 8424
rect 4896 8381 4905 8415
rect 4905 8381 4939 8415
rect 4939 8381 4948 8415
rect 6552 8508 6604 8560
rect 8392 8551 8444 8560
rect 8392 8517 8401 8551
rect 8401 8517 8435 8551
rect 8435 8517 8444 8551
rect 8392 8508 8444 8517
rect 10508 8576 10560 8628
rect 10600 8576 10652 8628
rect 11336 8619 11388 8628
rect 11336 8585 11345 8619
rect 11345 8585 11379 8619
rect 11379 8585 11388 8619
rect 11336 8576 11388 8585
rect 12164 8576 12216 8628
rect 12348 8576 12400 8628
rect 13912 8576 13964 8628
rect 14832 8576 14884 8628
rect 12532 8551 12584 8560
rect 12532 8517 12541 8551
rect 12541 8517 12575 8551
rect 12575 8517 12584 8551
rect 12532 8508 12584 8517
rect 13360 8551 13412 8560
rect 13360 8517 13369 8551
rect 13369 8517 13403 8551
rect 13403 8517 13412 8551
rect 13360 8508 13412 8517
rect 13544 8508 13596 8560
rect 8760 8440 8812 8492
rect 9772 8483 9824 8492
rect 9772 8449 9781 8483
rect 9781 8449 9815 8483
rect 9815 8449 9824 8483
rect 9772 8440 9824 8449
rect 11244 8483 11296 8492
rect 11244 8449 11253 8483
rect 11253 8449 11287 8483
rect 11287 8449 11296 8483
rect 11244 8440 11296 8449
rect 4896 8372 4948 8381
rect 1400 8347 1452 8356
rect 1400 8313 1409 8347
rect 1409 8313 1443 8347
rect 1443 8313 1452 8347
rect 1400 8304 1452 8313
rect 3516 8304 3568 8356
rect 9680 8372 9732 8424
rect 12440 8440 12492 8492
rect 12900 8440 12952 8492
rect 13636 8440 13688 8492
rect 13820 8440 13872 8492
rect 14280 8483 14332 8492
rect 14280 8449 14289 8483
rect 14289 8449 14323 8483
rect 14323 8449 14332 8483
rect 14280 8440 14332 8449
rect 15200 8483 15252 8492
rect 15200 8449 15209 8483
rect 15209 8449 15243 8483
rect 15243 8449 15252 8483
rect 15200 8440 15252 8449
rect 2044 8236 2096 8288
rect 2964 8279 3016 8288
rect 2964 8245 2973 8279
rect 2973 8245 3007 8279
rect 3007 8245 3016 8279
rect 2964 8236 3016 8245
rect 3056 8279 3108 8288
rect 3056 8245 3065 8279
rect 3065 8245 3099 8279
rect 3099 8245 3108 8279
rect 3056 8236 3108 8245
rect 3332 8236 3384 8288
rect 5172 8347 5224 8356
rect 5172 8313 5206 8347
rect 5206 8313 5224 8347
rect 5172 8304 5224 8313
rect 5448 8304 5500 8356
rect 9312 8304 9364 8356
rect 10416 8304 10468 8356
rect 10876 8304 10928 8356
rect 11152 8304 11204 8356
rect 11980 8372 12032 8424
rect 12164 8372 12216 8424
rect 11704 8304 11756 8356
rect 12532 8372 12584 8424
rect 12624 8372 12676 8424
rect 13544 8372 13596 8424
rect 14004 8372 14056 8424
rect 3700 8236 3752 8288
rect 4528 8236 4580 8288
rect 6644 8236 6696 8288
rect 8116 8236 8168 8288
rect 8668 8236 8720 8288
rect 11980 8236 12032 8288
rect 13452 8304 13504 8356
rect 14096 8304 14148 8356
rect 14280 8304 14332 8356
rect 12348 8236 12400 8288
rect 13268 8236 13320 8288
rect 13728 8236 13780 8288
rect 14832 8236 14884 8288
rect 5979 8134 6031 8186
rect 6043 8134 6095 8186
rect 6107 8134 6159 8186
rect 6171 8134 6223 8186
rect 10976 8134 11028 8186
rect 11040 8134 11092 8186
rect 11104 8134 11156 8186
rect 11168 8134 11220 8186
rect 1492 8075 1544 8084
rect 1492 8041 1501 8075
rect 1501 8041 1535 8075
rect 1535 8041 1544 8075
rect 1492 8032 1544 8041
rect 1860 8032 1912 8084
rect 2688 8032 2740 8084
rect 3056 8032 3108 8084
rect 3240 8075 3292 8084
rect 3240 8041 3249 8075
rect 3249 8041 3283 8075
rect 3283 8041 3292 8075
rect 3240 8032 3292 8041
rect 3516 8032 3568 8084
rect 1584 7964 1636 8016
rect 2044 7939 2096 7948
rect 2044 7905 2053 7939
rect 2053 7905 2087 7939
rect 2087 7905 2096 7939
rect 2044 7896 2096 7905
rect 2412 7939 2464 7948
rect 2412 7905 2421 7939
rect 2421 7905 2455 7939
rect 2455 7905 2464 7939
rect 2412 7896 2464 7905
rect 2780 7964 2832 8016
rect 2964 7896 3016 7948
rect 3608 7896 3660 7948
rect 3976 7964 4028 8016
rect 5080 8032 5132 8084
rect 5172 8032 5224 8084
rect 8300 8032 8352 8084
rect 8852 8032 8904 8084
rect 2688 7828 2740 7880
rect 3056 7871 3108 7880
rect 3056 7837 3065 7871
rect 3065 7837 3099 7871
rect 3099 7837 3108 7871
rect 3056 7828 3108 7837
rect 6920 7964 6972 8016
rect 5724 7896 5776 7948
rect 7840 7896 7892 7948
rect 8392 7964 8444 8016
rect 8668 7939 8720 7948
rect 8668 7905 8686 7939
rect 8686 7905 8720 7939
rect 8668 7896 8720 7905
rect 4528 7828 4580 7880
rect 3608 7760 3660 7812
rect 4344 7760 4396 7812
rect 1768 7692 1820 7744
rect 3884 7692 3936 7744
rect 4068 7692 4120 7744
rect 5816 7828 5868 7880
rect 5632 7760 5684 7812
rect 7932 7828 7984 7880
rect 9404 8032 9456 8084
rect 10600 8032 10652 8084
rect 11796 8075 11848 8084
rect 9036 7964 9088 8016
rect 10968 8007 11020 8016
rect 10968 7973 10977 8007
rect 10977 7973 11011 8007
rect 11011 7973 11020 8007
rect 10968 7964 11020 7973
rect 11796 8041 11805 8075
rect 11805 8041 11839 8075
rect 11839 8041 11848 8075
rect 11796 8032 11848 8041
rect 12256 8032 12308 8084
rect 12348 8032 12400 8084
rect 13728 7964 13780 8016
rect 15016 7964 15068 8016
rect 12532 7896 12584 7948
rect 10508 7871 10560 7880
rect 10508 7837 10517 7871
rect 10517 7837 10551 7871
rect 10551 7837 10560 7871
rect 10508 7828 10560 7837
rect 10784 7828 10836 7880
rect 4896 7692 4948 7744
rect 6000 7735 6052 7744
rect 6000 7701 6009 7735
rect 6009 7701 6043 7735
rect 6043 7701 6052 7735
rect 6000 7692 6052 7701
rect 6460 7692 6512 7744
rect 6828 7692 6880 7744
rect 7196 7692 7248 7744
rect 10876 7760 10928 7812
rect 11152 7871 11204 7880
rect 11152 7837 11161 7871
rect 11161 7837 11195 7871
rect 11195 7837 11204 7871
rect 11980 7871 12032 7880
rect 11152 7828 11204 7837
rect 11980 7837 11989 7871
rect 11989 7837 12023 7871
rect 12023 7837 12032 7871
rect 11980 7828 12032 7837
rect 12440 7828 12492 7880
rect 13084 7896 13136 7948
rect 13176 7896 13228 7948
rect 13820 7896 13872 7948
rect 14188 7896 14240 7948
rect 12900 7871 12952 7880
rect 12256 7803 12308 7812
rect 10600 7735 10652 7744
rect 10600 7701 10609 7735
rect 10609 7701 10643 7735
rect 10643 7701 10652 7735
rect 10600 7692 10652 7701
rect 10784 7692 10836 7744
rect 11244 7692 11296 7744
rect 11428 7735 11480 7744
rect 11428 7701 11437 7735
rect 11437 7701 11471 7735
rect 11471 7701 11480 7735
rect 11428 7692 11480 7701
rect 12256 7769 12265 7803
rect 12265 7769 12299 7803
rect 12299 7769 12308 7803
rect 12256 7760 12308 7769
rect 12900 7837 12909 7871
rect 12909 7837 12943 7871
rect 12943 7837 12952 7871
rect 12900 7828 12952 7837
rect 13636 7871 13688 7880
rect 13636 7837 13645 7871
rect 13645 7837 13679 7871
rect 13679 7837 13688 7871
rect 13636 7828 13688 7837
rect 14096 7760 14148 7812
rect 12348 7692 12400 7744
rect 12532 7692 12584 7744
rect 12992 7692 13044 7744
rect 13084 7735 13136 7744
rect 13084 7701 13093 7735
rect 13093 7701 13127 7735
rect 13127 7701 13136 7735
rect 13084 7692 13136 7701
rect 14188 7735 14240 7744
rect 14188 7701 14197 7735
rect 14197 7701 14231 7735
rect 14231 7701 14240 7735
rect 14188 7692 14240 7701
rect 14740 7735 14792 7744
rect 14740 7701 14749 7735
rect 14749 7701 14783 7735
rect 14783 7701 14792 7735
rect 14740 7692 14792 7701
rect 14924 7735 14976 7744
rect 14924 7701 14933 7735
rect 14933 7701 14967 7735
rect 14967 7701 14976 7735
rect 14924 7692 14976 7701
rect 3480 7590 3532 7642
rect 3544 7590 3596 7642
rect 3608 7590 3660 7642
rect 3672 7590 3724 7642
rect 8478 7590 8530 7642
rect 8542 7590 8594 7642
rect 8606 7590 8658 7642
rect 8670 7590 8722 7642
rect 13475 7590 13527 7642
rect 13539 7590 13591 7642
rect 13603 7590 13655 7642
rect 13667 7590 13719 7642
rect 3240 7488 3292 7540
rect 3148 7420 3200 7472
rect 1400 7395 1452 7404
rect 1400 7361 1409 7395
rect 1409 7361 1443 7395
rect 1443 7361 1452 7395
rect 1400 7352 1452 7361
rect 2688 7352 2740 7404
rect 2964 7352 3016 7404
rect 10600 7488 10652 7540
rect 10876 7488 10928 7540
rect 1768 7284 1820 7336
rect 4896 7327 4948 7336
rect 4896 7293 4905 7327
rect 4905 7293 4939 7327
rect 4939 7293 4948 7327
rect 4896 7284 4948 7293
rect 1676 7216 1728 7268
rect 2136 7191 2188 7200
rect 2136 7157 2145 7191
rect 2145 7157 2179 7191
rect 2179 7157 2188 7191
rect 2136 7148 2188 7157
rect 2872 7191 2924 7200
rect 2872 7157 2881 7191
rect 2881 7157 2915 7191
rect 2915 7157 2924 7191
rect 2872 7148 2924 7157
rect 3056 7216 3108 7268
rect 5448 7284 5500 7336
rect 6368 7420 6420 7472
rect 10416 7420 10468 7472
rect 9404 7395 9456 7404
rect 9404 7361 9413 7395
rect 9413 7361 9447 7395
rect 9447 7361 9456 7395
rect 9404 7352 9456 7361
rect 10508 7352 10560 7404
rect 10968 7352 11020 7404
rect 6000 7284 6052 7336
rect 7564 7259 7616 7268
rect 4160 7148 4212 7200
rect 4988 7148 5040 7200
rect 5080 7148 5132 7200
rect 5632 7148 5684 7200
rect 5816 7148 5868 7200
rect 7564 7225 7582 7259
rect 7582 7225 7616 7259
rect 7564 7216 7616 7225
rect 7932 7327 7984 7336
rect 7932 7293 7941 7327
rect 7941 7293 7975 7327
rect 7975 7293 7984 7327
rect 7932 7284 7984 7293
rect 10784 7284 10836 7336
rect 10876 7327 10928 7336
rect 10876 7293 10885 7327
rect 10885 7293 10919 7327
rect 10919 7293 10928 7327
rect 12532 7488 12584 7540
rect 12716 7488 12768 7540
rect 14004 7488 14056 7540
rect 14280 7488 14332 7540
rect 14740 7488 14792 7540
rect 11244 7420 11296 7472
rect 12992 7420 13044 7472
rect 13084 7395 13136 7404
rect 10876 7284 10928 7293
rect 11336 7284 11388 7336
rect 11980 7284 12032 7336
rect 13084 7361 13093 7395
rect 13093 7361 13127 7395
rect 13127 7361 13136 7395
rect 13084 7352 13136 7361
rect 12900 7284 12952 7336
rect 14004 7284 14056 7336
rect 14648 7284 14700 7336
rect 9680 7259 9732 7268
rect 9680 7225 9714 7259
rect 9714 7225 9732 7259
rect 9680 7216 9732 7225
rect 10048 7216 10100 7268
rect 12624 7216 12676 7268
rect 14464 7216 14516 7268
rect 9220 7148 9272 7200
rect 9312 7191 9364 7200
rect 9312 7157 9321 7191
rect 9321 7157 9355 7191
rect 9355 7157 9364 7191
rect 9312 7148 9364 7157
rect 10324 7148 10376 7200
rect 11428 7148 11480 7200
rect 11704 7191 11756 7200
rect 11704 7157 11713 7191
rect 11713 7157 11747 7191
rect 11747 7157 11756 7191
rect 11704 7148 11756 7157
rect 12164 7148 12216 7200
rect 12348 7148 12400 7200
rect 12900 7191 12952 7200
rect 12900 7157 12909 7191
rect 12909 7157 12943 7191
rect 12943 7157 12952 7191
rect 12900 7148 12952 7157
rect 12992 7191 13044 7200
rect 12992 7157 13001 7191
rect 13001 7157 13035 7191
rect 13035 7157 13044 7191
rect 13820 7191 13872 7200
rect 12992 7148 13044 7157
rect 13820 7157 13829 7191
rect 13829 7157 13863 7191
rect 13863 7157 13872 7191
rect 13820 7148 13872 7157
rect 14372 7191 14424 7200
rect 14372 7157 14381 7191
rect 14381 7157 14415 7191
rect 14415 7157 14424 7191
rect 14372 7148 14424 7157
rect 5979 7046 6031 7098
rect 6043 7046 6095 7098
rect 6107 7046 6159 7098
rect 6171 7046 6223 7098
rect 10976 7046 11028 7098
rect 11040 7046 11092 7098
rect 11104 7046 11156 7098
rect 11168 7046 11220 7098
rect 1676 6944 1728 6996
rect 1492 6876 1544 6928
rect 2596 6944 2648 6996
rect 2504 6919 2556 6928
rect 2504 6885 2513 6919
rect 2513 6885 2547 6919
rect 2547 6885 2556 6919
rect 2504 6876 2556 6885
rect 2964 6944 3016 6996
rect 1584 6808 1636 6860
rect 2320 6808 2372 6860
rect 4252 6851 4304 6860
rect 4252 6817 4261 6851
rect 4261 6817 4295 6851
rect 4295 6817 4304 6851
rect 4252 6808 4304 6817
rect 2228 6783 2280 6792
rect 2228 6749 2237 6783
rect 2237 6749 2271 6783
rect 2271 6749 2280 6783
rect 2228 6740 2280 6749
rect 2412 6783 2464 6792
rect 2412 6749 2421 6783
rect 2421 6749 2455 6783
rect 2455 6749 2464 6783
rect 2412 6740 2464 6749
rect 3608 6783 3660 6792
rect 1860 6647 1912 6656
rect 1860 6613 1869 6647
rect 1869 6613 1903 6647
rect 1903 6613 1912 6647
rect 1860 6604 1912 6613
rect 2044 6604 2096 6656
rect 2872 6647 2924 6656
rect 2872 6613 2881 6647
rect 2881 6613 2915 6647
rect 2915 6613 2924 6647
rect 2872 6604 2924 6613
rect 3056 6604 3108 6656
rect 3608 6749 3617 6783
rect 3617 6749 3651 6783
rect 3651 6749 3660 6783
rect 3608 6740 3660 6749
rect 4712 6987 4764 6996
rect 4712 6953 4721 6987
rect 4721 6953 4755 6987
rect 4755 6953 4764 6987
rect 4712 6944 4764 6953
rect 4804 6919 4856 6928
rect 4804 6885 4813 6919
rect 4813 6885 4847 6919
rect 4847 6885 4856 6919
rect 4804 6876 4856 6885
rect 8392 6944 8444 6996
rect 8760 6944 8812 6996
rect 11980 6944 12032 6996
rect 12256 6987 12308 6996
rect 12256 6953 12265 6987
rect 12265 6953 12299 6987
rect 12299 6953 12308 6987
rect 12256 6944 12308 6953
rect 12716 6944 12768 6996
rect 13176 6944 13228 6996
rect 14096 6944 14148 6996
rect 5264 6876 5316 6928
rect 6092 6876 6144 6928
rect 6460 6876 6512 6928
rect 7564 6876 7616 6928
rect 5724 6808 5776 6860
rect 7932 6876 7984 6928
rect 7748 6851 7800 6860
rect 8208 6876 8260 6928
rect 7748 6817 7766 6851
rect 7766 6817 7800 6851
rect 7748 6808 7800 6817
rect 5540 6740 5592 6792
rect 8116 6808 8168 6860
rect 8852 6876 8904 6928
rect 9312 6876 9364 6928
rect 10048 6876 10100 6928
rect 11612 6876 11664 6928
rect 11796 6876 11848 6928
rect 12348 6919 12400 6928
rect 9864 6808 9916 6860
rect 10416 6808 10468 6860
rect 10508 6808 10560 6860
rect 11152 6808 11204 6860
rect 11980 6808 12032 6860
rect 12348 6885 12357 6919
rect 12357 6885 12391 6919
rect 12391 6885 12400 6919
rect 12348 6876 12400 6885
rect 14924 6876 14976 6928
rect 12808 6808 12860 6860
rect 8208 6740 8260 6792
rect 3976 6672 4028 6724
rect 4068 6715 4120 6724
rect 4068 6681 4077 6715
rect 4077 6681 4111 6715
rect 4111 6681 4120 6715
rect 4068 6672 4120 6681
rect 4712 6672 4764 6724
rect 4252 6604 4304 6656
rect 4528 6604 4580 6656
rect 6736 6672 6788 6724
rect 8024 6672 8076 6724
rect 8852 6740 8904 6792
rect 9036 6672 9088 6724
rect 9404 6783 9456 6792
rect 9404 6749 9413 6783
rect 9413 6749 9447 6783
rect 9447 6749 9456 6783
rect 9404 6740 9456 6749
rect 11520 6740 11572 6792
rect 11704 6783 11756 6792
rect 11704 6749 11713 6783
rect 11713 6749 11747 6783
rect 11747 6749 11756 6783
rect 11704 6740 11756 6749
rect 11796 6740 11848 6792
rect 12624 6740 12676 6792
rect 13268 6783 13320 6792
rect 13268 6749 13277 6783
rect 13277 6749 13311 6783
rect 13311 6749 13320 6783
rect 13268 6740 13320 6749
rect 9680 6672 9732 6724
rect 12256 6672 12308 6724
rect 7012 6604 7064 6656
rect 7104 6604 7156 6656
rect 8208 6604 8260 6656
rect 10416 6604 10468 6656
rect 10876 6604 10928 6656
rect 11060 6647 11112 6656
rect 11060 6613 11069 6647
rect 11069 6613 11103 6647
rect 11103 6613 11112 6647
rect 11060 6604 11112 6613
rect 11152 6604 11204 6656
rect 14280 6604 14332 6656
rect 14740 6647 14792 6656
rect 14740 6613 14749 6647
rect 14749 6613 14783 6647
rect 14783 6613 14792 6647
rect 14740 6604 14792 6613
rect 3480 6502 3532 6554
rect 3544 6502 3596 6554
rect 3608 6502 3660 6554
rect 3672 6502 3724 6554
rect 8478 6502 8530 6554
rect 8542 6502 8594 6554
rect 8606 6502 8658 6554
rect 8670 6502 8722 6554
rect 13475 6502 13527 6554
rect 13539 6502 13591 6554
rect 13603 6502 13655 6554
rect 13667 6502 13719 6554
rect 1492 6443 1544 6452
rect 1492 6409 1501 6443
rect 1501 6409 1535 6443
rect 1535 6409 1544 6443
rect 1492 6400 1544 6409
rect 2412 6400 2464 6452
rect 3792 6400 3844 6452
rect 4436 6400 4488 6452
rect 5264 6400 5316 6452
rect 5540 6400 5592 6452
rect 8024 6400 8076 6452
rect 8300 6400 8352 6452
rect 10048 6400 10100 6452
rect 10416 6400 10468 6452
rect 11796 6400 11848 6452
rect 2228 6332 2280 6384
rect 3608 6332 3660 6384
rect 5080 6332 5132 6384
rect 9404 6375 9456 6384
rect 9404 6341 9413 6375
rect 9413 6341 9447 6375
rect 9447 6341 9456 6375
rect 9404 6332 9456 6341
rect 10784 6332 10836 6384
rect 10876 6332 10928 6384
rect 11888 6332 11940 6384
rect 1860 6196 1912 6248
rect 2044 6307 2096 6316
rect 2044 6273 2053 6307
rect 2053 6273 2087 6307
rect 2087 6273 2096 6307
rect 2044 6264 2096 6273
rect 2320 6264 2372 6316
rect 2688 6264 2740 6316
rect 3332 6264 3384 6316
rect 4896 6196 4948 6248
rect 5080 6196 5132 6248
rect 6460 6239 6512 6248
rect 6460 6205 6469 6239
rect 6469 6205 6503 6239
rect 6503 6205 6512 6239
rect 6460 6196 6512 6205
rect 11152 6264 11204 6316
rect 12992 6400 13044 6452
rect 12624 6332 12676 6384
rect 12716 6264 12768 6316
rect 13084 6307 13136 6316
rect 13084 6273 13093 6307
rect 13093 6273 13127 6307
rect 13127 6273 13136 6307
rect 13084 6264 13136 6273
rect 14372 6307 14424 6316
rect 14372 6273 14381 6307
rect 14381 6273 14415 6307
rect 14415 6273 14424 6307
rect 14372 6264 14424 6273
rect 8760 6196 8812 6248
rect 9220 6196 9272 6248
rect 5448 6128 5500 6180
rect 5816 6128 5868 6180
rect 6368 6128 6420 6180
rect 6552 6128 6604 6180
rect 7012 6128 7064 6180
rect 8300 6128 8352 6180
rect 8852 6128 8904 6180
rect 9680 6128 9732 6180
rect 10232 6128 10284 6180
rect 10324 6128 10376 6180
rect 12624 6196 12676 6248
rect 12992 6196 13044 6248
rect 10968 6128 11020 6180
rect 11428 6171 11480 6180
rect 11428 6137 11437 6171
rect 11437 6137 11471 6171
rect 11471 6137 11480 6171
rect 11428 6128 11480 6137
rect 11980 6128 12032 6180
rect 13544 6128 13596 6180
rect 13636 6128 13688 6180
rect 2320 6060 2372 6112
rect 2596 6103 2648 6112
rect 2596 6069 2605 6103
rect 2605 6069 2639 6103
rect 2639 6069 2648 6103
rect 2596 6060 2648 6069
rect 2964 6103 3016 6112
rect 2964 6069 2973 6103
rect 2973 6069 3007 6103
rect 3007 6069 3016 6103
rect 2964 6060 3016 6069
rect 3056 6103 3108 6112
rect 3056 6069 3065 6103
rect 3065 6069 3099 6103
rect 3099 6069 3108 6103
rect 3056 6060 3108 6069
rect 3608 6060 3660 6112
rect 3700 6060 3752 6112
rect 5724 6060 5776 6112
rect 7472 6060 7524 6112
rect 7564 6060 7616 6112
rect 8024 6060 8076 6112
rect 10692 6060 10744 6112
rect 10876 6060 10928 6112
rect 11704 6103 11756 6112
rect 11704 6069 11713 6103
rect 11713 6069 11747 6103
rect 11747 6069 11756 6103
rect 11704 6060 11756 6069
rect 12348 6060 12400 6112
rect 12440 6060 12492 6112
rect 12808 6060 12860 6112
rect 13360 6103 13412 6112
rect 13360 6069 13369 6103
rect 13369 6069 13403 6103
rect 13403 6069 13412 6103
rect 13360 6060 13412 6069
rect 13820 6103 13872 6112
rect 13820 6069 13829 6103
rect 13829 6069 13863 6103
rect 13863 6069 13872 6103
rect 13820 6060 13872 6069
rect 5979 5958 6031 6010
rect 6043 5958 6095 6010
rect 6107 5958 6159 6010
rect 6171 5958 6223 6010
rect 10976 5958 11028 6010
rect 11040 5958 11092 6010
rect 11104 5958 11156 6010
rect 11168 5958 11220 6010
rect 3056 5856 3108 5908
rect 3516 5788 3568 5840
rect 1676 5559 1728 5568
rect 1676 5525 1685 5559
rect 1685 5525 1719 5559
rect 1719 5525 1728 5559
rect 1676 5516 1728 5525
rect 1860 5559 1912 5568
rect 1860 5525 1869 5559
rect 1869 5525 1903 5559
rect 1903 5525 1912 5559
rect 1860 5516 1912 5525
rect 2228 5720 2280 5772
rect 3700 5720 3752 5772
rect 3884 5763 3936 5772
rect 3884 5729 3893 5763
rect 3893 5729 3927 5763
rect 3927 5729 3936 5763
rect 3884 5720 3936 5729
rect 4436 5856 4488 5908
rect 4712 5788 4764 5840
rect 8392 5856 8444 5908
rect 8484 5856 8536 5908
rect 8760 5856 8812 5908
rect 4068 5720 4120 5772
rect 2412 5695 2464 5704
rect 2412 5661 2421 5695
rect 2421 5661 2455 5695
rect 2455 5661 2464 5695
rect 2412 5652 2464 5661
rect 3608 5652 3660 5704
rect 4344 5695 4396 5704
rect 4344 5661 4353 5695
rect 4353 5661 4387 5695
rect 4387 5661 4396 5695
rect 4344 5652 4396 5661
rect 4620 5695 4672 5704
rect 4620 5661 4629 5695
rect 4629 5661 4663 5695
rect 4663 5661 4672 5695
rect 4620 5652 4672 5661
rect 6460 5788 6512 5840
rect 8208 5788 8260 5840
rect 9220 5788 9272 5840
rect 9772 5856 9824 5908
rect 9496 5788 9548 5840
rect 5356 5720 5408 5772
rect 5540 5763 5592 5772
rect 5540 5729 5574 5763
rect 5574 5729 5592 5763
rect 5540 5720 5592 5729
rect 5816 5720 5868 5772
rect 7012 5720 7064 5772
rect 7840 5763 7892 5772
rect 7840 5729 7858 5763
rect 7858 5729 7892 5763
rect 8576 5763 8628 5772
rect 7840 5720 7892 5729
rect 3332 5584 3384 5636
rect 3516 5584 3568 5636
rect 4068 5584 4120 5636
rect 8208 5652 8260 5704
rect 8576 5729 8585 5763
rect 8585 5729 8619 5763
rect 8619 5729 8628 5763
rect 8576 5720 8628 5729
rect 9128 5763 9180 5772
rect 9128 5729 9137 5763
rect 9137 5729 9171 5763
rect 9171 5729 9180 5763
rect 9128 5720 9180 5729
rect 3056 5516 3108 5568
rect 4436 5516 4488 5568
rect 6368 5584 6420 5636
rect 4620 5516 4672 5568
rect 6644 5559 6696 5568
rect 6644 5525 6653 5559
rect 6653 5525 6687 5559
rect 6687 5525 6696 5559
rect 6644 5516 6696 5525
rect 6920 5516 6972 5568
rect 8852 5652 8904 5704
rect 9772 5720 9824 5772
rect 10692 5856 10744 5908
rect 11888 5899 11940 5908
rect 11888 5865 11897 5899
rect 11897 5865 11931 5899
rect 11931 5865 11940 5899
rect 11888 5856 11940 5865
rect 12440 5856 12492 5908
rect 12624 5899 12676 5908
rect 12624 5865 12633 5899
rect 12633 5865 12667 5899
rect 12667 5865 12676 5899
rect 12624 5856 12676 5865
rect 14096 5856 14148 5908
rect 10876 5788 10928 5840
rect 12716 5831 12768 5840
rect 11888 5720 11940 5772
rect 12440 5720 12492 5772
rect 12716 5797 12725 5831
rect 12725 5797 12759 5831
rect 12759 5797 12768 5831
rect 12716 5788 12768 5797
rect 12808 5788 12860 5840
rect 12992 5788 13044 5840
rect 13544 5831 13596 5840
rect 13544 5797 13553 5831
rect 13553 5797 13587 5831
rect 13587 5797 13596 5831
rect 13544 5788 13596 5797
rect 15200 5788 15252 5840
rect 10508 5652 10560 5704
rect 10876 5652 10928 5704
rect 11520 5652 11572 5704
rect 12716 5652 12768 5704
rect 9404 5516 9456 5568
rect 9864 5516 9916 5568
rect 11704 5584 11756 5636
rect 12440 5584 12492 5636
rect 11060 5516 11112 5568
rect 13360 5516 13412 5568
rect 14004 5559 14056 5568
rect 14004 5525 14013 5559
rect 14013 5525 14047 5559
rect 14047 5525 14056 5559
rect 14004 5516 14056 5525
rect 3480 5414 3532 5466
rect 3544 5414 3596 5466
rect 3608 5414 3660 5466
rect 3672 5414 3724 5466
rect 8478 5414 8530 5466
rect 8542 5414 8594 5466
rect 8606 5414 8658 5466
rect 8670 5414 8722 5466
rect 13475 5414 13527 5466
rect 13539 5414 13591 5466
rect 13603 5414 13655 5466
rect 13667 5414 13719 5466
rect 1492 5355 1544 5364
rect 1492 5321 1501 5355
rect 1501 5321 1535 5355
rect 1535 5321 1544 5355
rect 1492 5312 1544 5321
rect 4804 5312 4856 5364
rect 5172 5312 5224 5364
rect 9496 5312 9548 5364
rect 10048 5312 10100 5364
rect 10416 5312 10468 5364
rect 11336 5312 11388 5364
rect 11428 5312 11480 5364
rect 12256 5312 12308 5364
rect 12716 5312 12768 5364
rect 13084 5312 13136 5364
rect 2136 5244 2188 5296
rect 2596 5176 2648 5228
rect 3792 5244 3844 5296
rect 7472 5244 7524 5296
rect 9404 5244 9456 5296
rect 5080 5176 5132 5228
rect 1860 5108 1912 5160
rect 2504 5108 2556 5160
rect 4160 5108 4212 5160
rect 6460 5151 6512 5160
rect 6460 5117 6469 5151
rect 6469 5117 6503 5151
rect 6503 5117 6512 5151
rect 6460 5108 6512 5117
rect 9496 5176 9548 5228
rect 8760 5108 8812 5160
rect 9036 5151 9088 5160
rect 9036 5117 9054 5151
rect 9054 5117 9088 5151
rect 9036 5108 9088 5117
rect 9220 5108 9272 5160
rect 9404 5108 9456 5160
rect 10508 5108 10560 5160
rect 3516 5040 3568 5092
rect 3608 5040 3660 5092
rect 4804 5040 4856 5092
rect 5264 5040 5316 5092
rect 5632 5040 5684 5092
rect 6552 5040 6604 5092
rect 6644 5040 6696 5092
rect 2320 4972 2372 5024
rect 3148 4972 3200 5024
rect 4896 5015 4948 5024
rect 4896 4981 4905 5015
rect 4905 4981 4939 5015
rect 4939 4981 4948 5015
rect 4896 4972 4948 4981
rect 5540 4972 5592 5024
rect 5724 4972 5776 5024
rect 7012 4972 7064 5024
rect 7288 4972 7340 5024
rect 7840 5015 7892 5024
rect 7840 4981 7849 5015
rect 7849 4981 7883 5015
rect 7883 4981 7892 5015
rect 7840 4972 7892 4981
rect 8208 4972 8260 5024
rect 9128 4972 9180 5024
rect 10416 5040 10468 5092
rect 10600 5083 10652 5092
rect 10600 5049 10609 5083
rect 10609 5049 10643 5083
rect 10643 5049 10652 5083
rect 10600 5040 10652 5049
rect 10784 5040 10836 5092
rect 9588 4972 9640 5024
rect 12808 5244 12860 5296
rect 13452 5244 13504 5296
rect 13544 5287 13596 5296
rect 13544 5253 13553 5287
rect 13553 5253 13587 5287
rect 13587 5253 13596 5287
rect 13544 5244 13596 5253
rect 14464 5244 14516 5296
rect 11520 5219 11572 5228
rect 11520 5185 11529 5219
rect 11529 5185 11563 5219
rect 11563 5185 11572 5219
rect 11520 5176 11572 5185
rect 11796 5176 11848 5228
rect 12716 5176 12768 5228
rect 14832 5176 14884 5228
rect 10968 5108 11020 5160
rect 12440 5108 12492 5160
rect 11060 5083 11112 5092
rect 11060 5049 11069 5083
rect 11069 5049 11103 5083
rect 11103 5049 11112 5083
rect 11060 5040 11112 5049
rect 14096 5108 14148 5160
rect 12992 5040 13044 5092
rect 11520 4972 11572 5024
rect 11796 4972 11848 5024
rect 13084 5015 13136 5024
rect 13084 4981 13093 5015
rect 13093 4981 13127 5015
rect 13127 4981 13136 5015
rect 13084 4972 13136 4981
rect 13636 5015 13688 5024
rect 13636 4981 13645 5015
rect 13645 4981 13679 5015
rect 13679 4981 13688 5015
rect 13636 4972 13688 4981
rect 14004 4972 14056 5024
rect 5979 4870 6031 4922
rect 6043 4870 6095 4922
rect 6107 4870 6159 4922
rect 6171 4870 6223 4922
rect 10976 4870 11028 4922
rect 11040 4870 11092 4922
rect 11104 4870 11156 4922
rect 11168 4870 11220 4922
rect 1676 4632 1728 4684
rect 2320 4675 2372 4684
rect 2320 4641 2329 4675
rect 2329 4641 2363 4675
rect 2363 4641 2372 4675
rect 2320 4632 2372 4641
rect 3332 4768 3384 4820
rect 4804 4811 4856 4820
rect 4804 4777 4813 4811
rect 4813 4777 4847 4811
rect 4847 4777 4856 4811
rect 4804 4768 4856 4777
rect 8024 4768 8076 4820
rect 9128 4768 9180 4820
rect 9496 4768 9548 4820
rect 9772 4768 9824 4820
rect 9864 4768 9916 4820
rect 10048 4768 10100 4820
rect 11704 4811 11756 4820
rect 5816 4700 5868 4752
rect 3148 4632 3200 4684
rect 3332 4675 3384 4684
rect 3332 4641 3341 4675
rect 3341 4641 3375 4675
rect 3375 4641 3384 4675
rect 3332 4632 3384 4641
rect 4160 4675 4212 4684
rect 4160 4641 4169 4675
rect 4169 4641 4203 4675
rect 4203 4641 4212 4675
rect 4160 4632 4212 4641
rect 6460 4675 6512 4684
rect 6460 4641 6478 4675
rect 6478 4641 6512 4675
rect 6460 4632 6512 4641
rect 6644 4632 6696 4684
rect 7380 4632 7432 4684
rect 8300 4632 8352 4684
rect 10508 4700 10560 4752
rect 3424 4607 3476 4616
rect 3424 4573 3433 4607
rect 3433 4573 3467 4607
rect 3467 4573 3476 4607
rect 3424 4564 3476 4573
rect 3608 4607 3660 4616
rect 3608 4573 3617 4607
rect 3617 4573 3651 4607
rect 3651 4573 3660 4607
rect 3608 4564 3660 4573
rect 2136 4496 2188 4548
rect 4344 4496 4396 4548
rect 5172 4496 5224 4548
rect 1492 4471 1544 4480
rect 1492 4437 1501 4471
rect 1501 4437 1535 4471
rect 1535 4437 1544 4471
rect 1492 4428 1544 4437
rect 1952 4471 2004 4480
rect 1952 4437 1961 4471
rect 1961 4437 1995 4471
rect 1995 4437 2004 4471
rect 1952 4428 2004 4437
rect 2044 4428 2096 4480
rect 3792 4428 3844 4480
rect 5264 4471 5316 4480
rect 5264 4437 5273 4471
rect 5273 4437 5307 4471
rect 5307 4437 5316 4471
rect 5264 4428 5316 4437
rect 5356 4471 5408 4480
rect 5356 4437 5365 4471
rect 5365 4437 5399 4471
rect 5399 4437 5408 4471
rect 6828 4564 6880 4616
rect 8208 4607 8260 4616
rect 5356 4428 5408 4437
rect 6736 4428 6788 4480
rect 8208 4573 8217 4607
rect 8217 4573 8251 4607
rect 8251 4573 8260 4607
rect 8208 4564 8260 4573
rect 9312 4564 9364 4616
rect 9496 4496 9548 4548
rect 9588 4496 9640 4548
rect 8852 4471 8904 4480
rect 8852 4437 8861 4471
rect 8861 4437 8895 4471
rect 8895 4437 8904 4471
rect 8852 4428 8904 4437
rect 9036 4428 9088 4480
rect 10324 4496 10376 4548
rect 10692 4632 10744 4684
rect 11060 4743 11112 4752
rect 11060 4709 11069 4743
rect 11069 4709 11103 4743
rect 11103 4709 11112 4743
rect 11704 4777 11713 4811
rect 11713 4777 11747 4811
rect 11747 4777 11756 4811
rect 11704 4768 11756 4777
rect 12440 4768 12492 4820
rect 13084 4768 13136 4820
rect 13268 4768 13320 4820
rect 13452 4811 13504 4820
rect 13452 4777 13461 4811
rect 13461 4777 13495 4811
rect 13495 4777 13504 4811
rect 13452 4768 13504 4777
rect 14740 4768 14792 4820
rect 11060 4700 11112 4709
rect 15016 4700 15068 4752
rect 11704 4632 11756 4684
rect 11888 4632 11940 4684
rect 12348 4632 12400 4684
rect 13084 4632 13136 4684
rect 13636 4675 13688 4684
rect 13636 4641 13645 4675
rect 13645 4641 13679 4675
rect 13679 4641 13688 4675
rect 13636 4632 13688 4641
rect 14004 4632 14056 4684
rect 11060 4496 11112 4548
rect 11336 4496 11388 4548
rect 14556 4564 14608 4616
rect 11796 4496 11848 4548
rect 11980 4539 12032 4548
rect 11980 4505 11989 4539
rect 11989 4505 12023 4539
rect 12023 4505 12032 4539
rect 11980 4496 12032 4505
rect 12348 4496 12400 4548
rect 12992 4496 13044 4548
rect 14280 4496 14332 4548
rect 10140 4428 10192 4480
rect 10508 4428 10560 4480
rect 10692 4428 10744 4480
rect 10784 4428 10836 4480
rect 12900 4428 12952 4480
rect 3480 4326 3532 4378
rect 3544 4326 3596 4378
rect 3608 4326 3660 4378
rect 3672 4326 3724 4378
rect 8478 4326 8530 4378
rect 8542 4326 8594 4378
rect 8606 4326 8658 4378
rect 8670 4326 8722 4378
rect 13475 4326 13527 4378
rect 13539 4326 13591 4378
rect 13603 4326 13655 4378
rect 13667 4326 13719 4378
rect 3332 4224 3384 4276
rect 4804 4224 4856 4276
rect 5172 4224 5224 4276
rect 5356 4224 5408 4276
rect 7380 4224 7432 4276
rect 7748 4224 7800 4276
rect 8024 4224 8076 4276
rect 3608 4156 3660 4208
rect 1768 4088 1820 4140
rect 2044 4020 2096 4072
rect 2412 4020 2464 4072
rect 2872 4088 2924 4140
rect 3884 4088 3936 4140
rect 4344 4131 4396 4140
rect 4344 4097 4353 4131
rect 4353 4097 4387 4131
rect 4387 4097 4396 4131
rect 4344 4088 4396 4097
rect 5908 4156 5960 4208
rect 5172 4088 5224 4140
rect 2780 4063 2832 4072
rect 2780 4029 2789 4063
rect 2789 4029 2823 4063
rect 2823 4029 2832 4063
rect 2780 4020 2832 4029
rect 3424 4020 3476 4072
rect 4068 4020 4120 4072
rect 4436 4020 4488 4072
rect 7472 4156 7524 4208
rect 9128 4224 9180 4276
rect 12256 4267 12308 4276
rect 8300 4156 8352 4208
rect 2136 3952 2188 4004
rect 1492 3927 1544 3936
rect 1492 3893 1501 3927
rect 1501 3893 1535 3927
rect 1535 3893 1544 3927
rect 1492 3884 1544 3893
rect 1860 3927 1912 3936
rect 1860 3893 1869 3927
rect 1869 3893 1903 3927
rect 1903 3893 1912 3927
rect 1860 3884 1912 3893
rect 2872 3952 2924 4004
rect 3884 3952 3936 4004
rect 4344 3952 4396 4004
rect 6460 4063 6512 4072
rect 6460 4029 6476 4063
rect 6476 4029 6510 4063
rect 6510 4029 6512 4063
rect 6460 4020 6512 4029
rect 8484 4088 8536 4140
rect 9588 4156 9640 4208
rect 9772 4156 9824 4208
rect 10232 4156 10284 4208
rect 9036 4088 9088 4140
rect 9956 4088 10008 4140
rect 10140 4131 10192 4140
rect 10140 4097 10149 4131
rect 10149 4097 10183 4131
rect 10183 4097 10192 4131
rect 10140 4088 10192 4097
rect 3056 3927 3108 3936
rect 3056 3893 3065 3927
rect 3065 3893 3099 3927
rect 3099 3893 3108 3927
rect 3056 3884 3108 3893
rect 4068 3884 4120 3936
rect 4804 3884 4856 3936
rect 5080 3927 5132 3936
rect 5080 3893 5089 3927
rect 5089 3893 5123 3927
rect 5123 3893 5132 3927
rect 5080 3884 5132 3893
rect 6368 3952 6420 4004
rect 8760 4020 8812 4072
rect 7380 3952 7432 4004
rect 8484 3952 8536 4004
rect 9036 3952 9088 4004
rect 9404 4020 9456 4072
rect 10876 4156 10928 4208
rect 6460 3884 6512 3936
rect 7288 3884 7340 3936
rect 8944 3884 8996 3936
rect 9404 3884 9456 3936
rect 9496 3884 9548 3936
rect 10416 3952 10468 4004
rect 10784 4020 10836 4072
rect 11152 4156 11204 4208
rect 11520 4156 11572 4208
rect 11980 4199 12032 4208
rect 11980 4165 11989 4199
rect 11989 4165 12023 4199
rect 12023 4165 12032 4199
rect 11980 4156 12032 4165
rect 12256 4233 12265 4267
rect 12265 4233 12299 4267
rect 12299 4233 12308 4267
rect 12256 4224 12308 4233
rect 12532 4267 12584 4276
rect 12532 4233 12541 4267
rect 12541 4233 12575 4267
rect 12575 4233 12584 4267
rect 12532 4224 12584 4233
rect 12808 4267 12860 4276
rect 12808 4233 12817 4267
rect 12817 4233 12851 4267
rect 12851 4233 12860 4267
rect 12808 4224 12860 4233
rect 13360 4224 13412 4276
rect 14004 4224 14056 4276
rect 14464 4267 14516 4276
rect 14464 4233 14473 4267
rect 14473 4233 14507 4267
rect 14507 4233 14516 4267
rect 14464 4224 14516 4233
rect 12992 4156 13044 4208
rect 14372 4156 14424 4208
rect 11244 4088 11296 4140
rect 12716 4088 12768 4140
rect 13820 4088 13872 4140
rect 15292 4088 15344 4140
rect 11060 3952 11112 4004
rect 10876 3884 10928 3936
rect 11796 4020 11848 4072
rect 12072 4063 12124 4072
rect 12072 4029 12081 4063
rect 12081 4029 12115 4063
rect 12115 4029 12124 4063
rect 12072 4020 12124 4029
rect 12440 4020 12492 4072
rect 12348 3952 12400 4004
rect 12808 3952 12860 4004
rect 12992 3995 13044 4004
rect 12992 3961 13001 3995
rect 13001 3961 13035 3995
rect 13035 3961 13044 3995
rect 12992 3952 13044 3961
rect 11336 3884 11388 3936
rect 11704 3927 11756 3936
rect 11704 3893 11713 3927
rect 11713 3893 11747 3927
rect 11747 3893 11756 3927
rect 11704 3884 11756 3893
rect 15108 3927 15160 3936
rect 15108 3893 15117 3927
rect 15117 3893 15151 3927
rect 15151 3893 15160 3927
rect 15108 3884 15160 3893
rect 15292 3927 15344 3936
rect 15292 3893 15301 3927
rect 15301 3893 15335 3927
rect 15335 3893 15344 3927
rect 15292 3884 15344 3893
rect 16212 3884 16264 3936
rect 5979 3782 6031 3834
rect 6043 3782 6095 3834
rect 6107 3782 6159 3834
rect 6171 3782 6223 3834
rect 10976 3782 11028 3834
rect 11040 3782 11092 3834
rect 11104 3782 11156 3834
rect 11168 3782 11220 3834
rect 3148 3680 3200 3732
rect 4252 3680 4304 3732
rect 5264 3680 5316 3732
rect 5356 3680 5408 3732
rect 7472 3680 7524 3732
rect 8024 3680 8076 3732
rect 8392 3680 8444 3732
rect 2504 3544 2556 3596
rect 2688 3544 2740 3596
rect 3332 3544 3384 3596
rect 3424 3587 3476 3596
rect 3424 3553 3433 3587
rect 3433 3553 3467 3587
rect 3467 3553 3476 3587
rect 3700 3587 3752 3596
rect 3424 3544 3476 3553
rect 3700 3553 3709 3587
rect 3709 3553 3743 3587
rect 3743 3553 3752 3587
rect 3700 3544 3752 3553
rect 6460 3612 6512 3664
rect 6644 3612 6696 3664
rect 9680 3612 9732 3664
rect 5080 3587 5132 3596
rect 5080 3553 5089 3587
rect 5089 3553 5123 3587
rect 5123 3553 5132 3587
rect 5080 3544 5132 3553
rect 5172 3544 5224 3596
rect 1124 3408 1176 3460
rect 1584 3408 1636 3460
rect 3608 3476 3660 3528
rect 4344 3476 4396 3528
rect 4528 3519 4580 3528
rect 4528 3485 4537 3519
rect 4537 3485 4571 3519
rect 4571 3485 4580 3519
rect 4528 3476 4580 3485
rect 4896 3476 4948 3528
rect 5908 3544 5960 3596
rect 7748 3544 7800 3596
rect 9404 3544 9456 3596
rect 9496 3587 9548 3596
rect 9496 3553 9505 3587
rect 9505 3553 9539 3587
rect 9539 3553 9548 3587
rect 9496 3544 9548 3553
rect 9864 3544 9916 3596
rect 10416 3612 10468 3664
rect 10784 3680 10836 3732
rect 10876 3680 10928 3732
rect 11520 3680 11572 3732
rect 10508 3587 10560 3596
rect 10508 3553 10517 3587
rect 10517 3553 10551 3587
rect 10551 3553 10560 3587
rect 10508 3544 10560 3553
rect 11796 3612 11848 3664
rect 12256 3680 12308 3732
rect 13084 3680 13136 3732
rect 14648 3680 14700 3732
rect 12440 3612 12492 3664
rect 13268 3612 13320 3664
rect 14004 3612 14056 3664
rect 3332 3408 3384 3460
rect 5724 3408 5776 3460
rect 6368 3519 6420 3528
rect 6368 3485 6377 3519
rect 6377 3485 6411 3519
rect 6411 3485 6420 3519
rect 6368 3476 6420 3485
rect 7656 3476 7708 3528
rect 7932 3519 7984 3528
rect 7932 3485 7941 3519
rect 7941 3485 7975 3519
rect 7975 3485 7984 3519
rect 7932 3476 7984 3485
rect 8116 3519 8168 3528
rect 8116 3485 8125 3519
rect 8125 3485 8159 3519
rect 8159 3485 8168 3519
rect 8116 3476 8168 3485
rect 8208 3476 8260 3528
rect 8760 3476 8812 3528
rect 9220 3476 9272 3528
rect 9772 3519 9824 3528
rect 9772 3485 9781 3519
rect 9781 3485 9815 3519
rect 9815 3485 9824 3519
rect 9772 3476 9824 3485
rect 11704 3476 11756 3528
rect 12072 3544 12124 3596
rect 12256 3544 12308 3596
rect 13360 3587 13412 3596
rect 13360 3553 13369 3587
rect 13369 3553 13403 3587
rect 13403 3553 13412 3587
rect 13360 3544 13412 3553
rect 13820 3587 13872 3596
rect 13820 3553 13829 3587
rect 13829 3553 13863 3587
rect 13863 3553 13872 3587
rect 13820 3544 13872 3553
rect 14464 3544 14516 3596
rect 14832 3587 14884 3596
rect 14832 3553 14841 3587
rect 14841 3553 14875 3587
rect 14875 3553 14884 3587
rect 14832 3544 14884 3553
rect 15108 3544 15160 3596
rect 15292 3587 15344 3596
rect 15292 3553 15301 3587
rect 15301 3553 15335 3587
rect 15335 3553 15344 3587
rect 15292 3544 15344 3553
rect 12440 3476 12492 3528
rect 12992 3476 13044 3528
rect 7012 3408 7064 3460
rect 7380 3451 7432 3460
rect 7380 3417 7389 3451
rect 7389 3417 7423 3451
rect 7423 3417 7432 3451
rect 7380 3408 7432 3417
rect 10048 3408 10100 3460
rect 10508 3408 10560 3460
rect 1860 3383 1912 3392
rect 1860 3349 1869 3383
rect 1869 3349 1903 3383
rect 1903 3349 1912 3383
rect 1860 3340 1912 3349
rect 2412 3383 2464 3392
rect 2412 3349 2421 3383
rect 2421 3349 2455 3383
rect 2455 3349 2464 3383
rect 2412 3340 2464 3349
rect 2596 3340 2648 3392
rect 3056 3340 3108 3392
rect 4068 3340 4120 3392
rect 5632 3340 5684 3392
rect 6276 3340 6328 3392
rect 8116 3340 8168 3392
rect 9128 3383 9180 3392
rect 9128 3349 9137 3383
rect 9137 3349 9171 3383
rect 9171 3349 9180 3383
rect 9128 3340 9180 3349
rect 10416 3383 10468 3392
rect 10416 3349 10425 3383
rect 10425 3349 10459 3383
rect 10459 3349 10468 3383
rect 10416 3340 10468 3349
rect 10600 3340 10652 3392
rect 11428 3408 11480 3460
rect 14556 3451 14608 3460
rect 14556 3417 14565 3451
rect 14565 3417 14599 3451
rect 14599 3417 14608 3451
rect 14556 3408 14608 3417
rect 15016 3451 15068 3460
rect 15016 3417 15025 3451
rect 15025 3417 15059 3451
rect 15059 3417 15068 3451
rect 15016 3408 15068 3417
rect 15660 3451 15712 3460
rect 15660 3417 15669 3451
rect 15669 3417 15703 3451
rect 15703 3417 15712 3451
rect 15660 3408 15712 3417
rect 10784 3340 10836 3392
rect 11060 3340 11112 3392
rect 11612 3340 11664 3392
rect 11980 3340 12032 3392
rect 12624 3383 12676 3392
rect 12624 3349 12633 3383
rect 12633 3349 12667 3383
rect 12667 3349 12676 3383
rect 12624 3340 12676 3349
rect 12900 3340 12952 3392
rect 13084 3383 13136 3392
rect 13084 3349 13093 3383
rect 13093 3349 13127 3383
rect 13127 3349 13136 3383
rect 13084 3340 13136 3349
rect 14464 3383 14516 3392
rect 14464 3349 14473 3383
rect 14473 3349 14507 3383
rect 14507 3349 14516 3383
rect 14464 3340 14516 3349
rect 3480 3238 3532 3290
rect 3544 3238 3596 3290
rect 3608 3238 3660 3290
rect 3672 3238 3724 3290
rect 8478 3238 8530 3290
rect 8542 3238 8594 3290
rect 8606 3238 8658 3290
rect 8670 3238 8722 3290
rect 13475 3238 13527 3290
rect 13539 3238 13591 3290
rect 13603 3238 13655 3290
rect 13667 3238 13719 3290
rect 2688 3136 2740 3188
rect 5080 3136 5132 3188
rect 1400 3068 1452 3120
rect 2504 3068 2556 3120
rect 8024 3136 8076 3188
rect 1584 2975 1636 2984
rect 1584 2941 1593 2975
rect 1593 2941 1627 2975
rect 1627 2941 1636 2975
rect 1584 2932 1636 2941
rect 2596 3000 2648 3052
rect 2780 3000 2832 3052
rect 4988 3000 5040 3052
rect 2228 2932 2280 2984
rect 2964 2932 3016 2984
rect 3148 2932 3200 2984
rect 4344 2932 4396 2984
rect 4528 2932 4580 2984
rect 4804 2932 4856 2984
rect 388 2864 440 2916
rect 1768 2864 1820 2916
rect 756 2796 808 2848
rect 2136 2864 2188 2916
rect 3332 2864 3384 2916
rect 3700 2864 3752 2916
rect 3884 2864 3936 2916
rect 4896 2864 4948 2916
rect 5080 2907 5132 2916
rect 5080 2873 5089 2907
rect 5089 2873 5123 2907
rect 5123 2873 5132 2907
rect 5080 2864 5132 2873
rect 5172 2907 5224 2916
rect 5172 2873 5181 2907
rect 5181 2873 5215 2907
rect 5215 2873 5224 2907
rect 5540 2932 5592 2984
rect 6184 3043 6236 3052
rect 6184 3009 6193 3043
rect 6193 3009 6227 3043
rect 6227 3009 6236 3043
rect 6184 3000 6236 3009
rect 6276 3000 6328 3052
rect 8484 3068 8536 3120
rect 5816 2932 5868 2984
rect 6828 2975 6880 2984
rect 6828 2941 6837 2975
rect 6837 2941 6871 2975
rect 6871 2941 6880 2975
rect 6828 2932 6880 2941
rect 5172 2864 5224 2873
rect 4068 2796 4120 2848
rect 6368 2864 6420 2916
rect 6736 2864 6788 2916
rect 7840 3043 7892 3052
rect 7840 3009 7849 3043
rect 7849 3009 7883 3043
rect 7883 3009 7892 3043
rect 7840 3000 7892 3009
rect 8024 3000 8076 3052
rect 9312 3136 9364 3188
rect 9404 3136 9456 3188
rect 8760 3068 8812 3120
rect 9680 3068 9732 3120
rect 8208 2932 8260 2984
rect 8944 3000 8996 3052
rect 9036 3000 9088 3052
rect 11060 3068 11112 3120
rect 9772 2932 9824 2984
rect 9864 2975 9916 2984
rect 9864 2941 9873 2975
rect 9873 2941 9907 2975
rect 9907 2941 9916 2975
rect 9864 2932 9916 2941
rect 10232 2932 10284 2984
rect 10517 2975 10569 2984
rect 10517 2941 10525 2975
rect 10525 2941 10559 2975
rect 10559 2941 10569 2975
rect 10517 2932 10569 2941
rect 7288 2864 7340 2916
rect 7380 2864 7432 2916
rect 8852 2864 8904 2916
rect 8944 2864 8996 2916
rect 11612 3000 11664 3052
rect 11796 3136 11848 3188
rect 11980 3136 12032 3188
rect 12348 3136 12400 3188
rect 12716 3136 12768 3188
rect 14096 3179 14148 3188
rect 14096 3145 14105 3179
rect 14105 3145 14139 3179
rect 14139 3145 14148 3179
rect 14096 3136 14148 3145
rect 13820 3068 13872 3120
rect 11796 3000 11848 3052
rect 12348 3000 12400 3052
rect 11152 2932 11204 2984
rect 11353 2932 11405 2984
rect 11704 2975 11756 2984
rect 11704 2941 11713 2975
rect 11713 2941 11747 2975
rect 11747 2941 11756 2975
rect 11704 2932 11756 2941
rect 12072 2932 12124 2984
rect 6920 2796 6972 2848
rect 8668 2796 8720 2848
rect 9036 2796 9088 2848
rect 9680 2839 9732 2848
rect 9680 2805 9689 2839
rect 9689 2805 9723 2839
rect 9723 2805 9732 2839
rect 9680 2796 9732 2805
rect 9956 2839 10008 2848
rect 9956 2805 9965 2839
rect 9965 2805 9999 2839
rect 9999 2805 10008 2839
rect 9956 2796 10008 2805
rect 10232 2839 10284 2848
rect 10232 2805 10241 2839
rect 10241 2805 10275 2839
rect 10275 2805 10284 2839
rect 10232 2796 10284 2805
rect 10876 2796 10928 2848
rect 11612 2864 11664 2916
rect 12440 2932 12492 2984
rect 13176 2932 13228 2984
rect 14556 3000 14608 3052
rect 14648 2975 14700 2984
rect 11980 2796 12032 2848
rect 13452 2864 13504 2916
rect 14188 2864 14240 2916
rect 14648 2941 14657 2975
rect 14657 2941 14691 2975
rect 14691 2941 14700 2975
rect 14648 2932 14700 2941
rect 15016 2932 15068 2984
rect 12624 2796 12676 2848
rect 12808 2796 12860 2848
rect 13820 2796 13872 2848
rect 14556 2839 14608 2848
rect 14556 2805 14565 2839
rect 14565 2805 14599 2839
rect 14599 2805 14608 2839
rect 14556 2796 14608 2805
rect 16948 2864 17000 2916
rect 14924 2839 14976 2848
rect 14924 2805 14933 2839
rect 14933 2805 14967 2839
rect 14967 2805 14976 2839
rect 14924 2796 14976 2805
rect 5979 2694 6031 2746
rect 6043 2694 6095 2746
rect 6107 2694 6159 2746
rect 6171 2694 6223 2746
rect 10976 2694 11028 2746
rect 11040 2694 11092 2746
rect 11104 2694 11156 2746
rect 11168 2694 11220 2746
rect 2412 2592 2464 2644
rect 5632 2635 5684 2644
rect 5632 2601 5641 2635
rect 5641 2601 5675 2635
rect 5675 2601 5684 2635
rect 5632 2592 5684 2601
rect 6460 2592 6512 2644
rect 7104 2592 7156 2644
rect 1952 2524 2004 2576
rect 2044 2499 2096 2508
rect 2044 2465 2053 2499
rect 2053 2465 2087 2499
rect 2087 2465 2096 2499
rect 2044 2456 2096 2465
rect 2688 2524 2740 2576
rect 2872 2524 2924 2576
rect 4620 2524 4672 2576
rect 8668 2592 8720 2644
rect 9496 2592 9548 2644
rect 9588 2592 9640 2644
rect 10324 2592 10376 2644
rect 10416 2592 10468 2644
rect 11520 2635 11572 2644
rect 7748 2567 7800 2576
rect 7748 2533 7757 2567
rect 7757 2533 7791 2567
rect 7791 2533 7800 2567
rect 7748 2524 7800 2533
rect 9128 2524 9180 2576
rect 9220 2524 9272 2576
rect 10876 2524 10928 2576
rect 11520 2601 11529 2635
rect 11529 2601 11563 2635
rect 11563 2601 11572 2635
rect 11520 2592 11572 2601
rect 11796 2592 11848 2644
rect 11980 2592 12032 2644
rect 12532 2592 12584 2644
rect 14096 2592 14148 2644
rect 11060 2524 11112 2576
rect 11152 2524 11204 2576
rect 3792 2456 3844 2508
rect 4252 2456 4304 2508
rect 4804 2499 4856 2508
rect 4804 2465 4813 2499
rect 4813 2465 4847 2499
rect 4847 2465 4856 2499
rect 4804 2456 4856 2465
rect 5172 2499 5224 2508
rect 5172 2465 5181 2499
rect 5181 2465 5215 2499
rect 5215 2465 5224 2499
rect 5172 2456 5224 2465
rect 6000 2499 6052 2508
rect 2320 2431 2372 2440
rect 2320 2397 2329 2431
rect 2329 2397 2363 2431
rect 2363 2397 2372 2431
rect 2320 2388 2372 2397
rect 112 2320 164 2372
rect 2228 2320 2280 2372
rect 4896 2388 4948 2440
rect 3976 2320 4028 2372
rect 4528 2320 4580 2372
rect 6000 2465 6009 2499
rect 6009 2465 6043 2499
rect 6043 2465 6052 2499
rect 6000 2456 6052 2465
rect 6920 2499 6972 2508
rect 6920 2465 6929 2499
rect 6929 2465 6963 2499
rect 6963 2465 6972 2499
rect 6920 2456 6972 2465
rect 7564 2456 7616 2508
rect 8024 2456 8076 2508
rect 8852 2499 8904 2508
rect 6092 2431 6144 2440
rect 6092 2397 6101 2431
rect 6101 2397 6135 2431
rect 6135 2397 6144 2431
rect 6092 2388 6144 2397
rect 6276 2431 6328 2440
rect 6276 2397 6285 2431
rect 6285 2397 6319 2431
rect 6319 2397 6328 2431
rect 6276 2388 6328 2397
rect 7196 2431 7248 2440
rect 7196 2397 7205 2431
rect 7205 2397 7239 2431
rect 7239 2397 7248 2431
rect 7196 2388 7248 2397
rect 7472 2320 7524 2372
rect 8116 2320 8168 2372
rect 8852 2465 8861 2499
rect 8861 2465 8895 2499
rect 8895 2465 8904 2499
rect 8852 2456 8904 2465
rect 9404 2456 9456 2508
rect 9864 2499 9916 2508
rect 9864 2465 9873 2499
rect 9873 2465 9907 2499
rect 9907 2465 9916 2499
rect 9864 2456 9916 2465
rect 10324 2456 10376 2508
rect 10416 2456 10468 2508
rect 10600 2499 10652 2508
rect 10600 2465 10609 2499
rect 10609 2465 10643 2499
rect 10643 2465 10652 2499
rect 10600 2456 10652 2465
rect 11244 2456 11296 2508
rect 14924 2524 14976 2576
rect 11520 2456 11572 2508
rect 10508 2388 10560 2440
rect 11796 2456 11848 2508
rect 12348 2456 12400 2508
rect 12808 2456 12860 2508
rect 13176 2456 13228 2508
rect 13452 2456 13504 2508
rect 13820 2456 13872 2508
rect 14004 2456 14056 2508
rect 14556 2456 14608 2508
rect 4068 2252 4120 2304
rect 4160 2252 4212 2304
rect 6552 2252 6604 2304
rect 9128 2320 9180 2372
rect 16580 2388 16632 2440
rect 11980 2320 12032 2372
rect 15108 2320 15160 2372
rect 15936 2320 15988 2372
rect 9496 2252 9548 2304
rect 10140 2295 10192 2304
rect 10140 2261 10149 2295
rect 10149 2261 10183 2295
rect 10183 2261 10192 2295
rect 10140 2252 10192 2261
rect 10416 2252 10468 2304
rect 10968 2252 11020 2304
rect 11244 2295 11296 2304
rect 11244 2261 11253 2295
rect 11253 2261 11287 2295
rect 11287 2261 11296 2295
rect 11244 2252 11296 2261
rect 12348 2295 12400 2304
rect 12348 2261 12357 2295
rect 12357 2261 12391 2295
rect 12391 2261 12400 2295
rect 12348 2252 12400 2261
rect 15568 2295 15620 2304
rect 15568 2261 15577 2295
rect 15577 2261 15611 2295
rect 15611 2261 15620 2295
rect 15568 2252 15620 2261
rect 3480 2150 3532 2202
rect 3544 2150 3596 2202
rect 3608 2150 3660 2202
rect 3672 2150 3724 2202
rect 8478 2150 8530 2202
rect 8542 2150 8594 2202
rect 8606 2150 8658 2202
rect 8670 2150 8722 2202
rect 13475 2150 13527 2202
rect 13539 2150 13591 2202
rect 13603 2150 13655 2202
rect 13667 2150 13719 2202
rect 5908 2048 5960 2100
rect 11244 2048 11296 2100
rect 6276 1980 6328 2032
rect 12348 1980 12400 2032
rect 2044 1912 2096 1964
rect 6828 1912 6880 1964
rect 8208 1912 8260 1964
rect 10140 1912 10192 1964
rect 12164 1912 12216 1964
rect 7656 1844 7708 1896
rect 9404 1844 9456 1896
rect 10324 1844 10376 1896
rect 12992 1844 13044 1896
rect 5172 1776 5224 1828
rect 9956 1776 10008 1828
rect 10784 1776 10836 1828
rect 12900 1776 12952 1828
rect 4252 1708 4304 1760
rect 9772 1708 9824 1760
rect 10692 1708 10744 1760
rect 11520 1708 11572 1760
rect 4804 1640 4856 1692
rect 10048 1640 10100 1692
rect 6000 1572 6052 1624
rect 11428 1572 11480 1624
rect 6920 1504 6972 1556
rect 7932 1504 7984 1556
rect 8024 1504 8076 1556
rect 9864 1504 9916 1556
rect 5540 1368 5592 1420
rect 9128 1368 9180 1420
rect 9680 1436 9732 1488
rect 12256 1436 12308 1488
rect 10232 1368 10284 1420
<< metal2 >>
rect 202 19200 258 20000
rect 570 19200 626 20000
rect 938 19200 994 20000
rect 1306 19200 1362 20000
rect 1398 19408 1454 19417
rect 1398 19343 1454 19352
rect 216 16726 244 19200
rect 584 16794 612 19200
rect 572 16788 624 16794
rect 572 16730 624 16736
rect 204 16720 256 16726
rect 204 16662 256 16668
rect 952 16182 980 19200
rect 1320 16658 1348 19200
rect 1412 17134 1440 19343
rect 1674 19200 1730 20000
rect 2042 19200 2098 20000
rect 2410 19200 2466 20000
rect 2778 19200 2834 20000
rect 3146 19200 3202 20000
rect 3514 19200 3570 20000
rect 3882 19200 3938 20000
rect 4250 19200 4306 20000
rect 4618 19200 4674 20000
rect 4986 19200 5042 20000
rect 5354 19200 5410 20000
rect 5722 19200 5778 20000
rect 6182 19200 6238 20000
rect 6550 19200 6606 20000
rect 6918 19200 6974 20000
rect 7286 19200 7342 20000
rect 7654 19200 7710 20000
rect 8022 19200 8078 20000
rect 8390 19200 8446 20000
rect 8758 19200 8814 20000
rect 9126 19200 9182 20000
rect 9494 19200 9550 20000
rect 9862 19200 9918 20000
rect 10230 19200 10286 20000
rect 10598 19200 10654 20000
rect 10966 19200 11022 20000
rect 11334 19200 11390 20000
rect 11794 19200 11850 20000
rect 12162 19200 12218 20000
rect 12530 19200 12586 20000
rect 12898 19200 12954 20000
rect 13266 19200 13322 20000
rect 13634 19200 13690 20000
rect 14002 19200 14058 20000
rect 14370 19200 14426 20000
rect 14738 19200 14794 20000
rect 15106 19200 15162 20000
rect 15474 19200 15530 20000
rect 15842 19200 15898 20000
rect 16210 19200 16266 20000
rect 16578 19200 16634 20000
rect 16946 19200 17002 20000
rect 1400 17128 1452 17134
rect 1400 17070 1452 17076
rect 1308 16652 1360 16658
rect 1308 16594 1360 16600
rect 940 16176 992 16182
rect 940 16118 992 16124
rect 1412 15638 1440 17070
rect 1688 16590 1716 19200
rect 1950 17368 2006 17377
rect 1950 17303 2006 17312
rect 1676 16584 1728 16590
rect 1676 16526 1728 16532
rect 1490 16416 1546 16425
rect 1490 16351 1546 16360
rect 1504 16250 1532 16351
rect 1492 16244 1544 16250
rect 1492 16186 1544 16192
rect 1964 16046 1992 17303
rect 2056 17270 2084 19200
rect 2424 17270 2452 19200
rect 2792 18578 2820 19200
rect 2792 18550 2912 18578
rect 2778 18456 2834 18465
rect 2778 18391 2834 18400
rect 2792 17338 2820 18391
rect 2780 17332 2832 17338
rect 2780 17274 2832 17280
rect 2044 17264 2096 17270
rect 2044 17206 2096 17212
rect 2412 17264 2464 17270
rect 2412 17206 2464 17212
rect 2884 17202 2912 18550
rect 3160 17338 3188 19200
rect 3528 17626 3556 19200
rect 3528 17598 3832 17626
rect 3454 17436 3750 17456
rect 3510 17434 3534 17436
rect 3590 17434 3614 17436
rect 3670 17434 3694 17436
rect 3532 17382 3534 17434
rect 3596 17382 3608 17434
rect 3670 17382 3672 17434
rect 3510 17380 3534 17382
rect 3590 17380 3614 17382
rect 3670 17380 3694 17382
rect 3454 17360 3750 17380
rect 3148 17332 3200 17338
rect 3148 17274 3200 17280
rect 3804 17270 3832 17598
rect 3896 17320 3924 19200
rect 4160 17332 4212 17338
rect 3896 17292 4160 17320
rect 4160 17274 4212 17280
rect 3792 17264 3844 17270
rect 4264 17252 4292 19200
rect 4344 17264 4396 17270
rect 4264 17224 4344 17252
rect 3792 17206 3844 17212
rect 4344 17206 4396 17212
rect 4632 17202 4660 19200
rect 2780 17196 2832 17202
rect 2780 17138 2832 17144
rect 2872 17196 2924 17202
rect 2872 17138 2924 17144
rect 4160 17196 4212 17202
rect 4160 17138 4212 17144
rect 4620 17196 4672 17202
rect 4620 17138 4672 17144
rect 2136 17128 2188 17134
rect 2136 17070 2188 17076
rect 2412 17128 2464 17134
rect 2412 17070 2464 17076
rect 2044 16516 2096 16522
rect 2044 16458 2096 16464
rect 1952 16040 2004 16046
rect 1952 15982 2004 15988
rect 2056 15910 2084 16458
rect 2148 16046 2176 17070
rect 2228 17060 2280 17066
rect 2228 17002 2280 17008
rect 2240 16794 2268 17002
rect 2228 16788 2280 16794
rect 2228 16730 2280 16736
rect 2424 16658 2452 17070
rect 2792 16980 2820 17138
rect 3792 17128 3844 17134
rect 3792 17070 3844 17076
rect 2964 17060 3016 17066
rect 2964 17002 3016 17008
rect 2872 16992 2924 16998
rect 2792 16952 2872 16980
rect 2872 16934 2924 16940
rect 2412 16652 2464 16658
rect 2412 16594 2464 16600
rect 2872 16652 2924 16658
rect 2872 16594 2924 16600
rect 2136 16040 2188 16046
rect 2136 15982 2188 15988
rect 2884 15910 2912 16594
rect 2044 15904 2096 15910
rect 2044 15846 2096 15852
rect 2412 15904 2464 15910
rect 2412 15846 2464 15852
rect 2872 15904 2924 15910
rect 2872 15846 2924 15852
rect 1400 15632 1452 15638
rect 2424 15586 2452 15846
rect 1400 15574 1452 15580
rect 2332 15558 2452 15586
rect 2780 15564 2832 15570
rect 1398 15464 1454 15473
rect 1398 15399 1400 15408
rect 1452 15399 1454 15408
rect 1400 15370 1452 15376
rect 1398 14376 1454 14385
rect 1398 14311 1400 14320
rect 1452 14311 1454 14320
rect 1400 14282 1452 14288
rect 1398 13424 1454 13433
rect 1398 13359 1400 13368
rect 1452 13359 1454 13368
rect 1400 13330 1452 13336
rect 2136 13184 2188 13190
rect 2136 13126 2188 13132
rect 2148 12782 2176 13126
rect 2136 12776 2188 12782
rect 2136 12718 2188 12724
rect 2044 12640 2096 12646
rect 2044 12582 2096 12588
rect 1398 12472 1454 12481
rect 1398 12407 1454 12416
rect 1412 12374 1440 12407
rect 1400 12368 1452 12374
rect 1400 12310 1452 12316
rect 2056 11898 2084 12582
rect 2332 12434 2360 15558
rect 2780 15506 2832 15512
rect 2688 14816 2740 14822
rect 2688 14758 2740 14764
rect 2504 14476 2556 14482
rect 2504 14418 2556 14424
rect 2516 14074 2544 14418
rect 2504 14068 2556 14074
rect 2504 14010 2556 14016
rect 2504 13728 2556 13734
rect 2504 13670 2556 13676
rect 2410 12608 2466 12617
rect 2410 12543 2466 12552
rect 2148 12406 2360 12434
rect 2044 11892 2096 11898
rect 2044 11834 2096 11840
rect 1950 11656 2006 11665
rect 1950 11591 1952 11600
rect 2004 11591 2006 11600
rect 1952 11562 2004 11568
rect 2148 11506 2176 12406
rect 2424 12356 2452 12543
rect 2516 12424 2544 13670
rect 2596 13388 2648 13394
rect 2596 13330 2648 13336
rect 2608 12986 2636 13330
rect 2596 12980 2648 12986
rect 2596 12922 2648 12928
rect 2516 12396 2636 12424
rect 2332 12328 2452 12356
rect 2332 12238 2360 12328
rect 2320 12232 2372 12238
rect 2320 12174 2372 12180
rect 2412 12232 2464 12238
rect 2412 12174 2464 12180
rect 2424 11801 2452 12174
rect 2608 12170 2636 12396
rect 2596 12164 2648 12170
rect 2596 12106 2648 12112
rect 2410 11792 2466 11801
rect 2410 11727 2466 11736
rect 1964 11478 2176 11506
rect 2228 11552 2280 11558
rect 2700 11506 2728 14758
rect 2792 14074 2820 15506
rect 2780 14068 2832 14074
rect 2780 14010 2832 14016
rect 2780 13796 2832 13802
rect 2780 13738 2832 13744
rect 2792 12782 2820 13738
rect 2780 12776 2832 12782
rect 2780 12718 2832 12724
rect 2884 12434 2912 15846
rect 2976 15706 3004 17002
rect 3240 16992 3292 16998
rect 3240 16934 3292 16940
rect 3252 16794 3280 16934
rect 3240 16788 3292 16794
rect 3240 16730 3292 16736
rect 2964 15700 3016 15706
rect 2964 15642 3016 15648
rect 2964 13864 3016 13870
rect 2964 13806 3016 13812
rect 2976 12918 3004 13806
rect 3146 13424 3202 13433
rect 3146 13359 3202 13368
rect 3056 13320 3108 13326
rect 3056 13262 3108 13268
rect 2964 12912 3016 12918
rect 2964 12854 3016 12860
rect 2228 11494 2280 11500
rect 1490 11384 1546 11393
rect 1490 11319 1492 11328
rect 1544 11319 1546 11328
rect 1492 11290 1544 11296
rect 1860 10532 1912 10538
rect 1860 10474 1912 10480
rect 1492 10464 1544 10470
rect 1490 10432 1492 10441
rect 1544 10432 1546 10441
rect 1490 10367 1546 10376
rect 1872 10266 1900 10474
rect 1860 10260 1912 10266
rect 1860 10202 1912 10208
rect 1584 9988 1636 9994
rect 1584 9930 1636 9936
rect 1400 9512 1452 9518
rect 1398 9480 1400 9489
rect 1452 9480 1454 9489
rect 1398 9415 1454 9424
rect 1490 9344 1546 9353
rect 1490 9279 1546 9288
rect 1504 9178 1532 9279
rect 1492 9172 1544 9178
rect 1492 9114 1544 9120
rect 1398 8392 1454 8401
rect 1398 8327 1400 8336
rect 1452 8327 1454 8336
rect 1400 8298 1452 8304
rect 1504 8090 1532 9114
rect 1596 9042 1624 9930
rect 1768 9920 1820 9926
rect 1768 9862 1820 9868
rect 1584 9036 1636 9042
rect 1584 8978 1636 8984
rect 1492 8084 1544 8090
rect 1780 8072 1808 9862
rect 1860 9444 1912 9450
rect 1860 9386 1912 9392
rect 1872 9178 1900 9386
rect 1860 9172 1912 9178
rect 1860 9114 1912 9120
rect 1860 8832 1912 8838
rect 1860 8774 1912 8780
rect 1872 8634 1900 8774
rect 1860 8628 1912 8634
rect 1860 8570 1912 8576
rect 1860 8084 1912 8090
rect 1780 8044 1860 8072
rect 1492 8026 1544 8032
rect 1860 8026 1912 8032
rect 1398 7440 1454 7449
rect 1398 7375 1400 7384
rect 1452 7375 1454 7384
rect 1400 7346 1452 7352
rect 1504 6934 1532 8026
rect 1584 8016 1636 8022
rect 1584 7958 1636 7964
rect 1492 6928 1544 6934
rect 1492 6870 1544 6876
rect 1596 6866 1624 7958
rect 1768 7744 1820 7750
rect 1768 7686 1820 7692
rect 1780 7342 1808 7686
rect 1768 7336 1820 7342
rect 1768 7278 1820 7284
rect 1676 7268 1728 7274
rect 1676 7210 1728 7216
rect 1688 7002 1716 7210
rect 1872 7188 1900 8026
rect 1780 7160 1900 7188
rect 1676 6996 1728 7002
rect 1676 6938 1728 6944
rect 1584 6860 1636 6866
rect 1584 6802 1636 6808
rect 1490 6488 1546 6497
rect 1490 6423 1492 6432
rect 1544 6423 1546 6432
rect 1492 6394 1544 6400
rect 1676 5568 1728 5574
rect 1676 5510 1728 5516
rect 1490 5400 1546 5409
rect 1490 5335 1492 5344
rect 1544 5335 1546 5344
rect 1492 5306 1544 5312
rect 1688 4690 1716 5510
rect 1676 4684 1728 4690
rect 1676 4626 1728 4632
rect 1492 4480 1544 4486
rect 1490 4448 1492 4457
rect 1544 4448 1546 4457
rect 1490 4383 1546 4392
rect 1492 3936 1544 3942
rect 1492 3878 1544 3884
rect 1124 3460 1176 3466
rect 1124 3402 1176 3408
rect 388 2916 440 2922
rect 388 2858 440 2864
rect 112 2372 164 2378
rect 112 2314 164 2320
rect 124 800 152 2314
rect 400 800 428 2858
rect 756 2848 808 2854
rect 756 2790 808 2796
rect 768 800 796 2790
rect 1136 800 1164 3402
rect 1400 3120 1452 3126
rect 1400 3062 1452 3068
rect 1412 800 1440 3062
rect 1504 2417 1532 3878
rect 1584 3460 1636 3466
rect 1584 3402 1636 3408
rect 1596 2990 1624 3402
rect 1584 2984 1636 2990
rect 1584 2926 1636 2932
rect 1490 2408 1546 2417
rect 1490 2343 1546 2352
rect 110 0 166 800
rect 386 0 442 800
rect 754 0 810 800
rect 1122 0 1178 800
rect 1398 0 1454 800
rect 1688 513 1716 4626
rect 1780 4146 1808 7160
rect 1860 6656 1912 6662
rect 1860 6598 1912 6604
rect 1872 6254 1900 6598
rect 1860 6248 1912 6254
rect 1860 6190 1912 6196
rect 1860 5568 1912 5574
rect 1860 5510 1912 5516
rect 1872 5166 1900 5510
rect 1860 5160 1912 5166
rect 1860 5102 1912 5108
rect 1964 5001 1992 11478
rect 2136 11008 2188 11014
rect 2136 10950 2188 10956
rect 2044 10464 2096 10470
rect 2044 10406 2096 10412
rect 2056 10266 2084 10406
rect 2044 10260 2096 10266
rect 2044 10202 2096 10208
rect 2148 9042 2176 10950
rect 2240 10033 2268 11494
rect 2424 11478 2728 11506
rect 2792 12406 2912 12434
rect 2424 10130 2452 11478
rect 2504 11212 2556 11218
rect 2504 11154 2556 11160
rect 2412 10124 2464 10130
rect 2412 10066 2464 10072
rect 2226 10024 2282 10033
rect 2226 9959 2282 9968
rect 2228 9648 2280 9654
rect 2228 9590 2280 9596
rect 2136 9036 2188 9042
rect 2136 8978 2188 8984
rect 2136 8832 2188 8838
rect 2136 8774 2188 8780
rect 2148 8430 2176 8774
rect 2240 8634 2268 9590
rect 2320 9580 2372 9586
rect 2320 9522 2372 9528
rect 2228 8628 2280 8634
rect 2228 8570 2280 8576
rect 2332 8430 2360 9522
rect 2516 9217 2544 11154
rect 2596 11144 2648 11150
rect 2596 11086 2648 11092
rect 2608 10810 2636 11086
rect 2596 10804 2648 10810
rect 2596 10746 2648 10752
rect 2688 10668 2740 10674
rect 2688 10610 2740 10616
rect 2700 10577 2728 10610
rect 2686 10568 2742 10577
rect 2686 10503 2742 10512
rect 2688 10124 2740 10130
rect 2688 10066 2740 10072
rect 2596 10056 2648 10062
rect 2596 9998 2648 10004
rect 2608 9489 2636 9998
rect 2594 9480 2650 9489
rect 2594 9415 2650 9424
rect 2502 9208 2558 9217
rect 2502 9143 2558 9152
rect 2410 9072 2466 9081
rect 2410 9007 2412 9016
rect 2464 9007 2466 9016
rect 2504 9036 2556 9042
rect 2412 8978 2464 8984
rect 2504 8978 2556 8984
rect 2136 8424 2188 8430
rect 2136 8366 2188 8372
rect 2320 8424 2372 8430
rect 2320 8366 2372 8372
rect 2044 8288 2096 8294
rect 2516 8265 2544 8978
rect 2700 8945 2728 10066
rect 2792 10044 2820 12406
rect 2870 12336 2926 12345
rect 2870 12271 2926 12280
rect 2884 10146 2912 12271
rect 3068 11762 3096 13262
rect 3160 12306 3188 13359
rect 3252 12345 3280 16730
rect 3804 16454 3832 17070
rect 3884 16516 3936 16522
rect 3884 16458 3936 16464
rect 3792 16448 3844 16454
rect 3896 16425 3924 16458
rect 3792 16390 3844 16396
rect 3882 16416 3938 16425
rect 3454 16348 3750 16368
rect 3882 16351 3938 16360
rect 3510 16346 3534 16348
rect 3590 16346 3614 16348
rect 3670 16346 3694 16348
rect 3532 16294 3534 16346
rect 3596 16294 3608 16346
rect 3670 16294 3672 16346
rect 3510 16292 3534 16294
rect 3590 16292 3614 16294
rect 3670 16292 3694 16294
rect 3454 16272 3750 16292
rect 3884 15972 3936 15978
rect 3884 15914 3936 15920
rect 3454 15260 3750 15280
rect 3510 15258 3534 15260
rect 3590 15258 3614 15260
rect 3670 15258 3694 15260
rect 3532 15206 3534 15258
rect 3596 15206 3608 15258
rect 3670 15206 3672 15258
rect 3510 15204 3534 15206
rect 3590 15204 3614 15206
rect 3670 15204 3694 15206
rect 3454 15184 3750 15204
rect 3332 15156 3384 15162
rect 3332 15098 3384 15104
rect 3238 12336 3294 12345
rect 3148 12300 3200 12306
rect 3238 12271 3294 12280
rect 3148 12242 3200 12248
rect 3240 12232 3292 12238
rect 3238 12200 3240 12209
rect 3292 12200 3294 12209
rect 3148 12164 3200 12170
rect 3238 12135 3294 12144
rect 3148 12106 3200 12112
rect 3160 11762 3188 12106
rect 3056 11756 3108 11762
rect 3056 11698 3108 11704
rect 3148 11756 3200 11762
rect 3148 11698 3200 11704
rect 3344 11626 3372 15098
rect 3792 14408 3844 14414
rect 3792 14350 3844 14356
rect 3454 14172 3750 14192
rect 3510 14170 3534 14172
rect 3590 14170 3614 14172
rect 3670 14170 3694 14172
rect 3532 14118 3534 14170
rect 3596 14118 3608 14170
rect 3670 14118 3672 14170
rect 3510 14116 3534 14118
rect 3590 14116 3614 14118
rect 3670 14116 3694 14118
rect 3454 14096 3750 14116
rect 3516 13932 3568 13938
rect 3516 13874 3568 13880
rect 3422 13832 3478 13841
rect 3422 13767 3478 13776
rect 3436 13530 3464 13767
rect 3424 13524 3476 13530
rect 3424 13466 3476 13472
rect 3528 13326 3556 13874
rect 3516 13320 3568 13326
rect 3516 13262 3568 13268
rect 3454 13084 3750 13104
rect 3510 13082 3534 13084
rect 3590 13082 3614 13084
rect 3670 13082 3694 13084
rect 3532 13030 3534 13082
rect 3596 13030 3608 13082
rect 3670 13030 3672 13082
rect 3510 13028 3534 13030
rect 3590 13028 3614 13030
rect 3670 13028 3694 13030
rect 3454 13008 3750 13028
rect 3514 12880 3570 12889
rect 3514 12815 3570 12824
rect 3528 12714 3556 12815
rect 3516 12708 3568 12714
rect 3516 12650 3568 12656
rect 3608 12708 3660 12714
rect 3608 12650 3660 12656
rect 3620 12442 3648 12650
rect 3608 12436 3660 12442
rect 3608 12378 3660 12384
rect 3454 11996 3750 12016
rect 3510 11994 3534 11996
rect 3590 11994 3614 11996
rect 3670 11994 3694 11996
rect 3532 11942 3534 11994
rect 3596 11942 3608 11994
rect 3670 11942 3672 11994
rect 3510 11940 3534 11942
rect 3590 11940 3614 11942
rect 3670 11940 3694 11942
rect 3454 11920 3750 11940
rect 3804 11898 3832 14350
rect 3896 13530 3924 15914
rect 4172 15706 4200 17138
rect 4252 17060 4304 17066
rect 4252 17002 4304 17008
rect 4436 17060 4488 17066
rect 4436 17002 4488 17008
rect 4804 17060 4856 17066
rect 4804 17002 4856 17008
rect 4160 15700 4212 15706
rect 4160 15642 4212 15648
rect 4264 15434 4292 17002
rect 4448 15706 4476 17002
rect 4528 16516 4580 16522
rect 4528 16458 4580 16464
rect 4436 15700 4488 15706
rect 4436 15642 4488 15648
rect 4540 15638 4568 16458
rect 4816 16250 4844 17002
rect 5000 16726 5028 19200
rect 5172 17060 5224 17066
rect 5172 17002 5224 17008
rect 4988 16720 5040 16726
rect 4988 16662 5040 16668
rect 5080 16448 5132 16454
rect 5080 16390 5132 16396
rect 4804 16244 4856 16250
rect 4804 16186 4856 16192
rect 4712 15904 4764 15910
rect 4712 15846 4764 15852
rect 4528 15632 4580 15638
rect 4528 15574 4580 15580
rect 4724 15570 4752 15846
rect 5092 15586 5120 16390
rect 5184 15706 5212 17002
rect 5368 16726 5396 19200
rect 5540 17060 5592 17066
rect 5540 17002 5592 17008
rect 5356 16720 5408 16726
rect 5356 16662 5408 16668
rect 5552 15706 5580 17002
rect 5736 16726 5764 19200
rect 6196 17270 6224 19200
rect 6184 17264 6236 17270
rect 6184 17206 6236 17212
rect 6564 17134 6592 19200
rect 6932 17270 6960 19200
rect 6920 17264 6972 17270
rect 6920 17206 6972 17212
rect 7300 17134 7328 19200
rect 7668 17270 7696 19200
rect 7656 17264 7708 17270
rect 8036 17252 8064 19200
rect 8404 17678 8432 19200
rect 8772 17762 8800 19200
rect 8772 17734 8984 17762
rect 8392 17672 8444 17678
rect 8392 17614 8444 17620
rect 8852 17672 8904 17678
rect 8852 17614 8904 17620
rect 8452 17436 8748 17456
rect 8508 17434 8532 17436
rect 8588 17434 8612 17436
rect 8668 17434 8692 17436
rect 8530 17382 8532 17434
rect 8594 17382 8606 17434
rect 8668 17382 8670 17434
rect 8508 17380 8532 17382
rect 8588 17380 8612 17382
rect 8668 17380 8692 17382
rect 8452 17360 8748 17380
rect 8300 17264 8352 17270
rect 8036 17224 8300 17252
rect 7656 17206 7708 17212
rect 8300 17206 8352 17212
rect 6552 17128 6604 17134
rect 6552 17070 6604 17076
rect 7288 17128 7340 17134
rect 7288 17070 7340 17076
rect 8484 17128 8536 17134
rect 8864 17082 8892 17614
rect 8956 17270 8984 17734
rect 8944 17264 8996 17270
rect 9140 17218 9168 19200
rect 9508 17338 9536 19200
rect 9496 17332 9548 17338
rect 9496 17274 9548 17280
rect 8944 17206 8996 17212
rect 9048 17202 9168 17218
rect 9036 17196 9168 17202
rect 9088 17190 9168 17196
rect 9036 17138 9088 17144
rect 9876 17134 9904 19200
rect 10244 17134 10272 19200
rect 10612 17626 10640 19200
rect 10612 17598 10732 17626
rect 10704 17134 10732 17598
rect 8484 17070 8536 17076
rect 5816 17060 5868 17066
rect 5816 17002 5868 17008
rect 6644 17060 6696 17066
rect 6644 17002 6696 17008
rect 7104 17060 7156 17066
rect 7104 17002 7156 17008
rect 8300 17060 8352 17066
rect 8300 17002 8352 17008
rect 5828 16794 5856 17002
rect 5953 16892 6249 16912
rect 6009 16890 6033 16892
rect 6089 16890 6113 16892
rect 6169 16890 6193 16892
rect 6031 16838 6033 16890
rect 6095 16838 6107 16890
rect 6169 16838 6171 16890
rect 6009 16836 6033 16838
rect 6089 16836 6113 16838
rect 6169 16836 6193 16838
rect 5953 16816 6249 16836
rect 6656 16794 6684 17002
rect 5816 16788 5868 16794
rect 5816 16730 5868 16736
rect 6644 16788 6696 16794
rect 6644 16730 6696 16736
rect 5724 16720 5776 16726
rect 5724 16662 5776 16668
rect 5816 16652 5868 16658
rect 5816 16594 5868 16600
rect 7012 16652 7064 16658
rect 7012 16594 7064 16600
rect 5828 16250 5856 16594
rect 6460 16584 6512 16590
rect 6460 16526 6512 16532
rect 5816 16244 5868 16250
rect 5816 16186 5868 16192
rect 6472 16182 6500 16526
rect 6920 16516 6972 16522
rect 6920 16458 6972 16464
rect 6736 16448 6788 16454
rect 6736 16390 6788 16396
rect 6460 16176 6512 16182
rect 6460 16118 6512 16124
rect 6748 16046 6776 16390
rect 6932 16046 6960 16458
rect 7024 16250 7052 16594
rect 7012 16244 7064 16250
rect 7012 16186 7064 16192
rect 6460 16040 6512 16046
rect 6460 15982 6512 15988
rect 6736 16040 6788 16046
rect 6736 15982 6788 15988
rect 6920 16040 6972 16046
rect 6920 15982 6972 15988
rect 5953 15804 6249 15824
rect 6009 15802 6033 15804
rect 6089 15802 6113 15804
rect 6169 15802 6193 15804
rect 6031 15750 6033 15802
rect 6095 15750 6107 15802
rect 6169 15750 6171 15802
rect 6009 15748 6033 15750
rect 6089 15748 6113 15750
rect 6169 15748 6193 15750
rect 5953 15728 6249 15748
rect 5172 15700 5224 15706
rect 5172 15642 5224 15648
rect 5540 15700 5592 15706
rect 5540 15642 5592 15648
rect 4344 15564 4396 15570
rect 4344 15506 4396 15512
rect 4712 15564 4764 15570
rect 5092 15558 5212 15586
rect 4712 15506 4764 15512
rect 4252 15428 4304 15434
rect 4252 15370 4304 15376
rect 4356 14958 4384 15506
rect 4618 15056 4674 15065
rect 4618 14991 4674 15000
rect 5080 15020 5132 15026
rect 4344 14952 4396 14958
rect 4344 14894 4396 14900
rect 4632 14618 4660 14991
rect 5080 14962 5132 14968
rect 4988 14816 5040 14822
rect 4988 14758 5040 14764
rect 5000 14618 5028 14758
rect 4620 14612 4672 14618
rect 4620 14554 4672 14560
rect 4988 14612 5040 14618
rect 4988 14554 5040 14560
rect 4068 14476 4120 14482
rect 4068 14418 4120 14424
rect 3884 13524 3936 13530
rect 3884 13466 3936 13472
rect 4080 13274 4108 14418
rect 4620 14340 4672 14346
rect 4620 14282 4672 14288
rect 4528 14272 4580 14278
rect 4528 14214 4580 14220
rect 4540 13938 4568 14214
rect 4528 13932 4580 13938
rect 4528 13874 4580 13880
rect 4632 13818 4660 14282
rect 4712 13932 4764 13938
rect 4712 13874 4764 13880
rect 4540 13790 4660 13818
rect 3988 13246 4108 13274
rect 4252 13320 4304 13326
rect 4252 13262 4304 13268
rect 4160 13252 4212 13258
rect 3884 12436 3936 12442
rect 3988 12424 4016 13246
rect 4160 13194 4212 13200
rect 4066 13152 4122 13161
rect 4066 13087 4122 13096
rect 4080 12714 4108 13087
rect 4068 12708 4120 12714
rect 4068 12650 4120 12656
rect 3936 12396 4016 12424
rect 4068 12436 4120 12442
rect 3884 12378 3936 12384
rect 4068 12378 4120 12384
rect 4080 12345 4108 12378
rect 4172 12374 4200 13194
rect 4160 12368 4212 12374
rect 4066 12336 4122 12345
rect 3896 12294 4066 12322
rect 3792 11892 3844 11898
rect 3792 11834 3844 11840
rect 3332 11620 3384 11626
rect 3332 11562 3384 11568
rect 3608 11552 3660 11558
rect 3608 11494 3660 11500
rect 3620 11286 3648 11494
rect 3608 11280 3660 11286
rect 3608 11222 3660 11228
rect 3332 11212 3384 11218
rect 3332 11154 3384 11160
rect 3344 10810 3372 11154
rect 3804 11082 3832 11834
rect 3792 11076 3844 11082
rect 3792 11018 3844 11024
rect 3454 10908 3750 10928
rect 3510 10906 3534 10908
rect 3590 10906 3614 10908
rect 3670 10906 3694 10908
rect 3532 10854 3534 10906
rect 3596 10854 3608 10906
rect 3670 10854 3672 10906
rect 3510 10852 3534 10854
rect 3590 10852 3614 10854
rect 3670 10852 3694 10854
rect 3454 10832 3750 10852
rect 3332 10804 3384 10810
rect 3332 10746 3384 10752
rect 3424 10600 3476 10606
rect 3344 10560 3424 10588
rect 3240 10532 3292 10538
rect 3240 10474 3292 10480
rect 2884 10118 3004 10146
rect 2872 10056 2924 10062
rect 2792 10016 2872 10044
rect 2872 9998 2924 10004
rect 2872 9920 2924 9926
rect 2872 9862 2924 9868
rect 2780 9648 2832 9654
rect 2780 9590 2832 9596
rect 2686 8936 2742 8945
rect 2686 8871 2742 8880
rect 2686 8392 2742 8401
rect 2686 8327 2742 8336
rect 2044 8230 2096 8236
rect 2502 8256 2558 8265
rect 2056 7954 2084 8230
rect 2502 8191 2558 8200
rect 2700 8090 2728 8327
rect 2688 8084 2740 8090
rect 2688 8026 2740 8032
rect 2792 8022 2820 9590
rect 2884 9586 2912 9862
rect 2872 9580 2924 9586
rect 2872 9522 2924 9528
rect 2976 9466 3004 10118
rect 3148 10124 3200 10130
rect 3148 10066 3200 10072
rect 3056 10056 3108 10062
rect 3056 9998 3108 10004
rect 3068 9625 3096 9998
rect 3054 9616 3110 9625
rect 3054 9551 3110 9560
rect 2884 9438 3004 9466
rect 2780 8016 2832 8022
rect 2410 7984 2466 7993
rect 2044 7948 2096 7954
rect 2780 7958 2832 7964
rect 2410 7919 2412 7928
rect 2044 7890 2096 7896
rect 2464 7919 2466 7928
rect 2412 7890 2464 7896
rect 2688 7880 2740 7886
rect 2884 7868 2912 9438
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 3056 9376 3108 9382
rect 3056 9318 3108 9324
rect 2976 9110 3004 9318
rect 3068 9178 3096 9318
rect 3056 9172 3108 9178
rect 3056 9114 3108 9120
rect 2964 9104 3016 9110
rect 2964 9046 3016 9052
rect 2964 8288 3016 8294
rect 2962 8256 2964 8265
rect 3056 8288 3108 8294
rect 3016 8256 3018 8265
rect 3056 8230 3108 8236
rect 2962 8191 3018 8200
rect 3068 8090 3096 8230
rect 3056 8084 3108 8090
rect 3056 8026 3108 8032
rect 2962 7984 3018 7993
rect 2962 7919 2964 7928
rect 3016 7919 3018 7928
rect 2964 7890 3016 7896
rect 2688 7822 2740 7828
rect 2792 7840 2912 7868
rect 3056 7880 3108 7886
rect 2700 7410 2728 7822
rect 2688 7404 2740 7410
rect 2688 7346 2740 7352
rect 2136 7200 2188 7206
rect 2136 7142 2188 7148
rect 2044 6656 2096 6662
rect 2044 6598 2096 6604
rect 2056 6322 2084 6598
rect 2044 6316 2096 6322
rect 2044 6258 2096 6264
rect 2148 6089 2176 7142
rect 2596 6996 2648 7002
rect 2596 6938 2648 6944
rect 2504 6928 2556 6934
rect 2502 6896 2504 6905
rect 2556 6896 2558 6905
rect 2320 6860 2372 6866
rect 2502 6831 2558 6840
rect 2320 6802 2372 6808
rect 2228 6792 2280 6798
rect 2228 6734 2280 6740
rect 2240 6390 2268 6734
rect 2228 6384 2280 6390
rect 2228 6326 2280 6332
rect 2332 6322 2360 6802
rect 2412 6792 2464 6798
rect 2412 6734 2464 6740
rect 2424 6458 2452 6734
rect 2412 6452 2464 6458
rect 2412 6394 2464 6400
rect 2320 6316 2372 6322
rect 2320 6258 2372 6264
rect 2226 6216 2282 6225
rect 2608 6202 2636 6938
rect 2688 6316 2740 6322
rect 2688 6258 2740 6264
rect 2226 6151 2282 6160
rect 2516 6174 2636 6202
rect 2134 6080 2190 6089
rect 2134 6015 2190 6024
rect 2134 5944 2190 5953
rect 2134 5879 2190 5888
rect 2148 5302 2176 5879
rect 2240 5778 2268 6151
rect 2320 6112 2372 6118
rect 2320 6054 2372 6060
rect 2228 5772 2280 5778
rect 2228 5714 2280 5720
rect 2136 5296 2188 5302
rect 2136 5238 2188 5244
rect 2332 5114 2360 6054
rect 2410 5808 2466 5817
rect 2410 5743 2466 5752
rect 2424 5710 2452 5743
rect 2412 5704 2464 5710
rect 2412 5646 2464 5652
rect 2516 5166 2544 6174
rect 2596 6112 2648 6118
rect 2596 6054 2648 6060
rect 2608 5234 2636 6054
rect 2596 5228 2648 5234
rect 2596 5170 2648 5176
rect 2240 5086 2360 5114
rect 2504 5160 2556 5166
rect 2504 5102 2556 5108
rect 1950 4992 2006 5001
rect 1950 4927 2006 4936
rect 2136 4548 2188 4554
rect 2136 4490 2188 4496
rect 1952 4480 2004 4486
rect 1952 4422 2004 4428
rect 2044 4480 2096 4486
rect 2044 4422 2096 4428
rect 1768 4140 1820 4146
rect 1768 4082 1820 4088
rect 1860 3936 1912 3942
rect 1860 3878 1912 3884
rect 1872 3505 1900 3878
rect 1858 3496 1914 3505
rect 1858 3431 1914 3440
rect 1860 3392 1912 3398
rect 1860 3334 1912 3340
rect 1768 2916 1820 2922
rect 1768 2858 1820 2864
rect 1780 800 1808 2858
rect 1872 1465 1900 3334
rect 1964 2582 1992 4422
rect 2056 4078 2084 4422
rect 2044 4072 2096 4078
rect 2044 4014 2096 4020
rect 2148 4010 2176 4490
rect 2136 4004 2188 4010
rect 2136 3946 2188 3952
rect 2240 3097 2268 5086
rect 2320 5024 2372 5030
rect 2320 4966 2372 4972
rect 2332 4690 2360 4966
rect 2320 4684 2372 4690
rect 2320 4626 2372 4632
rect 2412 4072 2464 4078
rect 2410 4040 2412 4049
rect 2464 4040 2466 4049
rect 2410 3975 2466 3984
rect 2516 3913 2544 5102
rect 2700 4978 2728 6258
rect 2608 4950 2728 4978
rect 2502 3904 2558 3913
rect 2502 3839 2558 3848
rect 2516 3602 2544 3839
rect 2504 3596 2556 3602
rect 2332 3556 2504 3584
rect 2226 3088 2282 3097
rect 2226 3023 2282 3032
rect 2228 2984 2280 2990
rect 2228 2926 2280 2932
rect 2136 2916 2188 2922
rect 2136 2858 2188 2864
rect 1952 2576 2004 2582
rect 1952 2518 2004 2524
rect 2044 2508 2096 2514
rect 2044 2450 2096 2456
rect 2056 1970 2084 2450
rect 2044 1964 2096 1970
rect 2044 1906 2096 1912
rect 1858 1456 1914 1465
rect 1858 1391 1914 1400
rect 2148 800 2176 2858
rect 2240 2689 2268 2926
rect 2226 2680 2282 2689
rect 2226 2615 2282 2624
rect 2332 2530 2360 3556
rect 2504 3538 2556 3544
rect 2608 3482 2636 4950
rect 2686 4856 2742 4865
rect 2686 4791 2742 4800
rect 2700 3602 2728 4791
rect 2792 4729 2820 7840
rect 3160 7857 3188 10066
rect 3252 9722 3280 10474
rect 3240 9716 3292 9722
rect 3240 9658 3292 9664
rect 3344 9654 3372 10560
rect 3424 10542 3476 10548
rect 3804 10538 3832 11018
rect 3792 10532 3844 10538
rect 3792 10474 3844 10480
rect 3896 10130 3924 12294
rect 4160 12310 4212 12316
rect 4066 12271 4122 12280
rect 4264 12220 4292 13262
rect 4540 12714 4568 13790
rect 4620 13388 4672 13394
rect 4620 13330 4672 13336
rect 4528 12708 4580 12714
rect 4528 12650 4580 12656
rect 4540 12617 4568 12650
rect 4526 12608 4582 12617
rect 4526 12543 4582 12552
rect 4436 12436 4488 12442
rect 4436 12378 4488 12384
rect 3988 12192 4292 12220
rect 4344 12232 4396 12238
rect 3988 11898 4016 12192
rect 4344 12174 4396 12180
rect 4356 12050 4384 12174
rect 4172 12022 4384 12050
rect 3976 11892 4028 11898
rect 3976 11834 4028 11840
rect 4068 11552 4120 11558
rect 4068 11494 4120 11500
rect 4172 11506 4200 12022
rect 4342 11928 4398 11937
rect 4342 11863 4398 11872
rect 4356 11762 4384 11863
rect 4344 11756 4396 11762
rect 4344 11698 4396 11704
rect 4344 11620 4396 11626
rect 4448 11608 4476 12378
rect 4528 12232 4580 12238
rect 4528 12174 4580 12180
rect 4540 11694 4568 12174
rect 4632 11880 4660 13330
rect 4724 13297 4752 13874
rect 4896 13864 4948 13870
rect 4896 13806 4948 13812
rect 4908 13530 4936 13806
rect 4896 13524 4948 13530
rect 4896 13466 4948 13472
rect 4710 13288 4766 13297
rect 4710 13223 4766 13232
rect 4724 12646 4752 13223
rect 4908 12782 4936 13466
rect 4988 13184 5040 13190
rect 4988 13126 5040 13132
rect 4896 12776 4948 12782
rect 4802 12744 4858 12753
rect 4896 12718 4948 12724
rect 4802 12679 4858 12688
rect 4712 12640 4764 12646
rect 4712 12582 4764 12588
rect 4632 11852 4752 11880
rect 4620 11756 4672 11762
rect 4620 11698 4672 11704
rect 4528 11688 4580 11694
rect 4528 11630 4580 11636
rect 4396 11580 4476 11608
rect 4344 11562 4396 11568
rect 4528 11552 4580 11558
rect 4080 11354 4108 11494
rect 4172 11478 4292 11506
rect 4528 11494 4580 11500
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 4160 11348 4212 11354
rect 4160 11290 4212 11296
rect 3976 10532 4028 10538
rect 3976 10474 4028 10480
rect 3700 10124 3752 10130
rect 3700 10066 3752 10072
rect 3884 10124 3936 10130
rect 3884 10066 3936 10072
rect 3712 9908 3740 10066
rect 3712 9880 3924 9908
rect 3454 9820 3750 9840
rect 3510 9818 3534 9820
rect 3590 9818 3614 9820
rect 3670 9818 3694 9820
rect 3532 9766 3534 9818
rect 3596 9766 3608 9818
rect 3670 9766 3672 9818
rect 3510 9764 3534 9766
rect 3590 9764 3614 9766
rect 3670 9764 3694 9766
rect 3454 9744 3750 9764
rect 3332 9648 3384 9654
rect 3238 9616 3294 9625
rect 3332 9590 3384 9596
rect 3238 9551 3240 9560
rect 3292 9551 3294 9560
rect 3240 9522 3292 9528
rect 3608 9172 3660 9178
rect 3608 9114 3660 9120
rect 3240 8900 3292 8906
rect 3240 8842 3292 8848
rect 3252 8498 3280 8842
rect 3620 8820 3648 9114
rect 3620 8792 3832 8820
rect 3454 8732 3750 8752
rect 3510 8730 3534 8732
rect 3590 8730 3614 8732
rect 3670 8730 3694 8732
rect 3532 8678 3534 8730
rect 3596 8678 3608 8730
rect 3670 8678 3672 8730
rect 3510 8676 3534 8678
rect 3590 8676 3614 8678
rect 3670 8676 3694 8678
rect 3454 8656 3750 8676
rect 3332 8560 3384 8566
rect 3332 8502 3384 8508
rect 3240 8492 3292 8498
rect 3240 8434 3292 8440
rect 3344 8294 3372 8502
rect 3516 8356 3568 8362
rect 3516 8298 3568 8304
rect 3332 8288 3384 8294
rect 3332 8230 3384 8236
rect 3528 8090 3556 8298
rect 3700 8288 3752 8294
rect 3700 8230 3752 8236
rect 3240 8084 3292 8090
rect 3240 8026 3292 8032
rect 3516 8084 3568 8090
rect 3516 8026 3568 8032
rect 3056 7822 3108 7828
rect 3146 7848 3202 7857
rect 2964 7404 3016 7410
rect 2964 7346 3016 7352
rect 2872 7200 2924 7206
rect 2872 7142 2924 7148
rect 2884 6769 2912 7142
rect 2976 7002 3004 7346
rect 3068 7274 3096 7822
rect 3146 7783 3202 7792
rect 3252 7546 3280 8026
rect 3712 7993 3740 8230
rect 3698 7984 3754 7993
rect 3608 7948 3660 7954
rect 3698 7919 3754 7928
rect 3608 7890 3660 7896
rect 3620 7818 3648 7890
rect 3608 7812 3660 7818
rect 3608 7754 3660 7760
rect 3454 7644 3750 7664
rect 3510 7642 3534 7644
rect 3590 7642 3614 7644
rect 3670 7642 3694 7644
rect 3532 7590 3534 7642
rect 3596 7590 3608 7642
rect 3670 7590 3672 7642
rect 3510 7588 3534 7590
rect 3590 7588 3614 7590
rect 3670 7588 3694 7590
rect 3454 7568 3750 7588
rect 3240 7540 3292 7546
rect 3240 7482 3292 7488
rect 3148 7472 3200 7478
rect 3148 7414 3200 7420
rect 3056 7268 3108 7274
rect 3056 7210 3108 7216
rect 2964 6996 3016 7002
rect 2964 6938 3016 6944
rect 2870 6760 2926 6769
rect 2870 6695 2926 6704
rect 2872 6656 2924 6662
rect 2872 6598 2924 6604
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 2778 4720 2834 4729
rect 2778 4655 2834 4664
rect 2884 4146 2912 6598
rect 3068 6236 3096 6598
rect 3160 6304 3188 7414
rect 3804 7313 3832 8792
rect 3896 8537 3924 9880
rect 3988 9178 4016 10474
rect 4172 10470 4200 11290
rect 4160 10464 4212 10470
rect 4160 10406 4212 10412
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 4172 9761 4200 9998
rect 4158 9752 4214 9761
rect 4158 9687 4214 9696
rect 4264 9450 4292 11478
rect 4436 11008 4488 11014
rect 4436 10950 4488 10956
rect 4342 10568 4398 10577
rect 4448 10538 4476 10950
rect 4342 10503 4398 10512
rect 4436 10532 4488 10538
rect 4252 9444 4304 9450
rect 4252 9386 4304 9392
rect 3976 9172 4028 9178
rect 3976 9114 4028 9120
rect 4068 9036 4120 9042
rect 4068 8978 4120 8984
rect 3882 8528 3938 8537
rect 3882 8463 3938 8472
rect 3976 8016 4028 8022
rect 3882 7984 3938 7993
rect 3976 7958 4028 7964
rect 3882 7919 3938 7928
rect 3896 7750 3924 7919
rect 3884 7744 3936 7750
rect 3884 7686 3936 7692
rect 3790 7304 3846 7313
rect 3790 7239 3846 7248
rect 3606 7168 3662 7177
rect 3606 7103 3662 7112
rect 3330 7032 3386 7041
rect 3330 6967 3386 6976
rect 3344 6322 3372 6967
rect 3620 6798 3648 7103
rect 3882 6896 3938 6905
rect 3882 6831 3938 6840
rect 3608 6792 3660 6798
rect 3608 6734 3660 6740
rect 3454 6556 3750 6576
rect 3510 6554 3534 6556
rect 3590 6554 3614 6556
rect 3670 6554 3694 6556
rect 3532 6502 3534 6554
rect 3596 6502 3608 6554
rect 3670 6502 3672 6554
rect 3510 6500 3534 6502
rect 3590 6500 3614 6502
rect 3670 6500 3694 6502
rect 3454 6480 3750 6500
rect 3896 6497 3924 6831
rect 3988 6730 4016 7958
rect 4080 7857 4108 8978
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 4172 8838 4200 8910
rect 4160 8832 4212 8838
rect 4160 8774 4212 8780
rect 4066 7848 4122 7857
rect 4066 7783 4122 7792
rect 4068 7744 4120 7750
rect 4068 7686 4120 7692
rect 4158 7712 4214 7721
rect 4080 6984 4108 7686
rect 4158 7647 4214 7656
rect 4172 7206 4200 7647
rect 4160 7200 4212 7206
rect 4160 7142 4212 7148
rect 4080 6956 4200 6984
rect 4066 6896 4122 6905
rect 4066 6831 4122 6840
rect 4080 6730 4108 6831
rect 3976 6724 4028 6730
rect 3976 6666 4028 6672
rect 4068 6724 4120 6730
rect 4068 6666 4120 6672
rect 3882 6488 3938 6497
rect 3792 6452 3844 6458
rect 3882 6423 3938 6432
rect 3792 6394 3844 6400
rect 3608 6384 3660 6390
rect 3608 6326 3660 6332
rect 3332 6316 3384 6322
rect 3160 6276 3280 6304
rect 3068 6208 3188 6236
rect 2964 6112 3016 6118
rect 2964 6054 3016 6060
rect 3056 6112 3108 6118
rect 3056 6054 3108 6060
rect 2976 4185 3004 6054
rect 3068 5914 3096 6054
rect 3056 5908 3108 5914
rect 3056 5850 3108 5856
rect 3056 5568 3108 5574
rect 3056 5510 3108 5516
rect 2962 4176 3018 4185
rect 2872 4140 2924 4146
rect 2962 4111 3018 4120
rect 2872 4082 2924 4088
rect 2780 4072 2832 4078
rect 2780 4014 2832 4020
rect 2688 3596 2740 3602
rect 2688 3538 2740 3544
rect 2792 3505 2820 4014
rect 2872 4004 2924 4010
rect 2872 3946 2924 3952
rect 2778 3496 2834 3505
rect 2608 3454 2728 3482
rect 2412 3392 2464 3398
rect 2412 3334 2464 3340
rect 2596 3392 2648 3398
rect 2596 3334 2648 3340
rect 2424 2650 2452 3334
rect 2504 3120 2556 3126
rect 2504 3062 2556 3068
rect 2412 2644 2464 2650
rect 2412 2586 2464 2592
rect 2240 2502 2360 2530
rect 2240 2378 2268 2502
rect 2320 2440 2372 2446
rect 2318 2408 2320 2417
rect 2372 2408 2374 2417
rect 2228 2372 2280 2378
rect 2318 2343 2374 2352
rect 2228 2314 2280 2320
rect 2516 800 2544 3062
rect 2608 3058 2636 3334
rect 2700 3194 2728 3454
rect 2778 3431 2834 3440
rect 2688 3188 2740 3194
rect 2688 3130 2740 3136
rect 2596 3052 2648 3058
rect 2596 2994 2648 3000
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 2686 2680 2742 2689
rect 2686 2615 2742 2624
rect 2700 2582 2728 2615
rect 2688 2576 2740 2582
rect 2688 2518 2740 2524
rect 2792 800 2820 2994
rect 2884 2582 2912 3946
rect 3068 3942 3096 5510
rect 3160 5030 3188 6208
rect 3148 5024 3200 5030
rect 3146 4992 3148 5001
rect 3200 4992 3202 5001
rect 3146 4927 3202 4936
rect 3148 4684 3200 4690
rect 3148 4626 3200 4632
rect 3056 3936 3108 3942
rect 3056 3878 3108 3884
rect 3160 3738 3188 4626
rect 3148 3732 3200 3738
rect 3148 3674 3200 3680
rect 3056 3392 3108 3398
rect 3056 3334 3108 3340
rect 2964 2984 3016 2990
rect 3068 2972 3096 3334
rect 3016 2944 3096 2972
rect 3148 2984 3200 2990
rect 2964 2926 3016 2932
rect 3252 2961 3280 6276
rect 3332 6258 3384 6264
rect 3620 6118 3648 6326
rect 3608 6112 3660 6118
rect 3608 6054 3660 6060
rect 3700 6112 3752 6118
rect 3700 6054 3752 6060
rect 3712 5930 3740 6054
rect 3620 5902 3740 5930
rect 3516 5840 3568 5846
rect 3516 5782 3568 5788
rect 3528 5642 3556 5782
rect 3620 5710 3648 5902
rect 3700 5772 3752 5778
rect 3700 5714 3752 5720
rect 3608 5704 3660 5710
rect 3608 5646 3660 5652
rect 3332 5636 3384 5642
rect 3332 5578 3384 5584
rect 3516 5636 3568 5642
rect 3516 5578 3568 5584
rect 3344 4826 3372 5578
rect 3712 5556 3740 5714
rect 3804 5624 3832 6394
rect 4080 6372 4108 6666
rect 4172 6633 4200 6956
rect 4264 6866 4292 9386
rect 4356 9042 4384 10503
rect 4436 10474 4488 10480
rect 4540 10266 4568 11494
rect 4632 11014 4660 11698
rect 4620 11008 4672 11014
rect 4620 10950 4672 10956
rect 4632 10606 4660 10950
rect 4620 10600 4672 10606
rect 4620 10542 4672 10548
rect 4528 10260 4580 10266
rect 4528 10202 4580 10208
rect 4620 10260 4672 10266
rect 4620 10202 4672 10208
rect 4436 10192 4488 10198
rect 4436 10134 4488 10140
rect 4526 10160 4582 10169
rect 4448 9586 4476 10134
rect 4526 10095 4528 10104
rect 4580 10095 4582 10104
rect 4528 10066 4580 10072
rect 4540 9926 4568 10066
rect 4528 9920 4580 9926
rect 4528 9862 4580 9868
rect 4436 9580 4488 9586
rect 4436 9522 4488 9528
rect 4344 9036 4396 9042
rect 4344 8978 4396 8984
rect 4344 8900 4396 8906
rect 4344 8842 4396 8848
rect 4356 8673 4384 8842
rect 4342 8664 4398 8673
rect 4342 8599 4398 8608
rect 4540 8294 4568 9862
rect 4632 9654 4660 10202
rect 4724 9994 4752 11852
rect 4816 11830 4844 12679
rect 4804 11824 4856 11830
rect 4804 11766 4856 11772
rect 4908 11694 4936 12718
rect 5000 12646 5028 13126
rect 4988 12640 5040 12646
rect 4988 12582 5040 12588
rect 4896 11688 4948 11694
rect 4896 11630 4948 11636
rect 4804 11552 4856 11558
rect 4804 11494 4856 11500
rect 4816 11218 4844 11494
rect 4804 11212 4856 11218
rect 4804 11154 4856 11160
rect 4908 10674 4936 11630
rect 4896 10668 4948 10674
rect 4896 10610 4948 10616
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 4712 9988 4764 9994
rect 4712 9930 4764 9936
rect 4620 9648 4672 9654
rect 4620 9590 4672 9596
rect 4816 9382 4844 10542
rect 4988 10464 5040 10470
rect 5092 10452 5120 14962
rect 5184 11121 5212 15558
rect 6000 15564 6052 15570
rect 6184 15564 6236 15570
rect 6000 15506 6052 15512
rect 6104 15524 6184 15552
rect 5908 15496 5960 15502
rect 5908 15438 5960 15444
rect 5816 15360 5868 15366
rect 5816 15302 5868 15308
rect 5264 14816 5316 14822
rect 5264 14758 5316 14764
rect 5724 14816 5776 14822
rect 5724 14758 5776 14764
rect 5276 12442 5304 14758
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5552 14074 5580 14350
rect 5540 14068 5592 14074
rect 5540 14010 5592 14016
rect 5632 13728 5684 13734
rect 5632 13670 5684 13676
rect 5448 13184 5500 13190
rect 5448 13126 5500 13132
rect 5460 12714 5488 13126
rect 5644 12986 5672 13670
rect 5632 12980 5684 12986
rect 5632 12922 5684 12928
rect 5448 12708 5500 12714
rect 5448 12650 5500 12656
rect 5264 12436 5316 12442
rect 5264 12378 5316 12384
rect 5446 11928 5502 11937
rect 5446 11863 5502 11872
rect 5460 11694 5488 11863
rect 5448 11688 5500 11694
rect 5448 11630 5500 11636
rect 5262 11248 5318 11257
rect 5262 11183 5264 11192
rect 5316 11183 5318 11192
rect 5264 11154 5316 11160
rect 5170 11112 5226 11121
rect 5170 11047 5226 11056
rect 5040 10424 5120 10452
rect 4988 10406 5040 10412
rect 5092 10130 5120 10424
rect 5276 10266 5304 11154
rect 5540 11144 5592 11150
rect 5540 11086 5592 11092
rect 5552 10606 5580 11086
rect 5540 10600 5592 10606
rect 5540 10542 5592 10548
rect 5264 10260 5316 10266
rect 5264 10202 5316 10208
rect 5080 10124 5132 10130
rect 5080 10066 5132 10072
rect 5172 10056 5224 10062
rect 5552 10044 5580 10542
rect 5644 10266 5672 12922
rect 5736 12889 5764 14758
rect 5828 13977 5856 15302
rect 5920 14958 5948 15438
rect 6012 15194 6040 15506
rect 6104 15434 6132 15524
rect 6184 15506 6236 15512
rect 6092 15428 6144 15434
rect 6092 15370 6144 15376
rect 6368 15360 6420 15366
rect 6368 15302 6420 15308
rect 6012 15166 6316 15194
rect 5908 14952 5960 14958
rect 5908 14894 5960 14900
rect 5953 14716 6249 14736
rect 6009 14714 6033 14716
rect 6089 14714 6113 14716
rect 6169 14714 6193 14716
rect 6031 14662 6033 14714
rect 6095 14662 6107 14714
rect 6169 14662 6171 14714
rect 6009 14660 6033 14662
rect 6089 14660 6113 14662
rect 6169 14660 6193 14662
rect 5953 14640 6249 14660
rect 6288 14464 6316 15166
rect 6380 14958 6408 15302
rect 6368 14952 6420 14958
rect 6368 14894 6420 14900
rect 6288 14436 6408 14464
rect 6276 14340 6328 14346
rect 6276 14282 6328 14288
rect 5908 14272 5960 14278
rect 5908 14214 5960 14220
rect 5814 13968 5870 13977
rect 5814 13903 5870 13912
rect 5920 13870 5948 14214
rect 6288 14006 6316 14282
rect 6276 14000 6328 14006
rect 6276 13942 6328 13948
rect 5908 13864 5960 13870
rect 5908 13806 5960 13812
rect 6276 13864 6328 13870
rect 6276 13806 6328 13812
rect 5953 13628 6249 13648
rect 6009 13626 6033 13628
rect 6089 13626 6113 13628
rect 6169 13626 6193 13628
rect 6031 13574 6033 13626
rect 6095 13574 6107 13626
rect 6169 13574 6171 13626
rect 6009 13572 6033 13574
rect 6089 13572 6113 13574
rect 6169 13572 6193 13574
rect 5953 13552 6249 13572
rect 5816 13320 5868 13326
rect 5816 13262 5868 13268
rect 5722 12880 5778 12889
rect 5722 12815 5778 12824
rect 5828 12714 5856 13262
rect 5816 12708 5868 12714
rect 5816 12650 5868 12656
rect 5828 12442 5856 12650
rect 5953 12540 6249 12560
rect 6009 12538 6033 12540
rect 6089 12538 6113 12540
rect 6169 12538 6193 12540
rect 6031 12486 6033 12538
rect 6095 12486 6107 12538
rect 6169 12486 6171 12538
rect 6009 12484 6033 12486
rect 6089 12484 6113 12486
rect 6169 12484 6193 12486
rect 5953 12464 6249 12484
rect 5816 12436 5868 12442
rect 5816 12378 5868 12384
rect 5908 12368 5960 12374
rect 5908 12310 5960 12316
rect 5920 12238 5948 12310
rect 5908 12232 5960 12238
rect 5908 12174 5960 12180
rect 5816 11620 5868 11626
rect 5816 11562 5868 11568
rect 5632 10260 5684 10266
rect 5632 10202 5684 10208
rect 5828 10130 5856 11562
rect 5953 11452 6249 11472
rect 6009 11450 6033 11452
rect 6089 11450 6113 11452
rect 6169 11450 6193 11452
rect 6031 11398 6033 11450
rect 6095 11398 6107 11450
rect 6169 11398 6171 11450
rect 6009 11396 6033 11398
rect 6089 11396 6113 11398
rect 6169 11396 6193 11398
rect 5953 11376 6249 11396
rect 6288 11370 6316 13806
rect 6380 12617 6408 14436
rect 6472 14362 6500 15982
rect 6734 15736 6790 15745
rect 7116 15706 7144 17002
rect 7288 16992 7340 16998
rect 7288 16934 7340 16940
rect 7196 16448 7248 16454
rect 7196 16390 7248 16396
rect 6734 15671 6736 15680
rect 6788 15671 6790 15680
rect 7104 15700 7156 15706
rect 6736 15642 6788 15648
rect 7104 15642 7156 15648
rect 7208 15638 7236 16390
rect 7300 16250 7328 16934
rect 7288 16244 7340 16250
rect 7288 16186 7340 16192
rect 8208 15972 8260 15978
rect 8208 15914 8260 15920
rect 7288 15904 7340 15910
rect 7288 15846 7340 15852
rect 7564 15904 7616 15910
rect 7564 15846 7616 15852
rect 7748 15904 7800 15910
rect 7748 15846 7800 15852
rect 7932 15904 7984 15910
rect 7932 15846 7984 15852
rect 7196 15632 7248 15638
rect 7196 15574 7248 15580
rect 7012 15496 7064 15502
rect 7012 15438 7064 15444
rect 6736 15428 6788 15434
rect 6736 15370 6788 15376
rect 6552 14884 6604 14890
rect 6552 14826 6604 14832
rect 6564 14482 6592 14826
rect 6552 14476 6604 14482
rect 6552 14418 6604 14424
rect 6748 14385 6776 15370
rect 6920 15360 6972 15366
rect 6920 15302 6972 15308
rect 6828 15020 6880 15026
rect 6828 14962 6880 14968
rect 6734 14376 6790 14385
rect 6472 14334 6684 14362
rect 6460 12776 6512 12782
rect 6460 12718 6512 12724
rect 6366 12608 6422 12617
rect 6366 12543 6422 12552
rect 6472 11762 6500 12718
rect 6460 11756 6512 11762
rect 6460 11698 6512 11704
rect 6288 11342 6408 11370
rect 6276 11212 6328 11218
rect 6276 11154 6328 11160
rect 5908 10668 5960 10674
rect 5908 10610 5960 10616
rect 5920 10538 5948 10610
rect 5908 10532 5960 10538
rect 5908 10474 5960 10480
rect 6288 10470 6316 11154
rect 6276 10464 6328 10470
rect 6276 10406 6328 10412
rect 5953 10364 6249 10384
rect 6009 10362 6033 10364
rect 6089 10362 6113 10364
rect 6169 10362 6193 10364
rect 6031 10310 6033 10362
rect 6095 10310 6107 10362
rect 6169 10310 6171 10362
rect 6009 10308 6033 10310
rect 6089 10308 6113 10310
rect 6169 10308 6193 10310
rect 5953 10288 6249 10308
rect 5816 10124 5868 10130
rect 5816 10066 5868 10072
rect 5224 10016 5580 10044
rect 5172 9998 5224 10004
rect 5184 9674 5212 9998
rect 4908 9646 5212 9674
rect 4908 9518 4936 9646
rect 4896 9512 4948 9518
rect 4896 9454 4948 9460
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 4988 9104 5040 9110
rect 4988 9046 5040 9052
rect 4896 8424 4948 8430
rect 4896 8366 4948 8372
rect 4528 8288 4580 8294
rect 4528 8230 4580 8236
rect 4540 7993 4568 8230
rect 4526 7984 4582 7993
rect 4526 7919 4582 7928
rect 4710 7984 4766 7993
rect 4710 7919 4766 7928
rect 4528 7880 4580 7886
rect 4448 7840 4528 7868
rect 4344 7812 4396 7818
rect 4344 7754 4396 7760
rect 4252 6860 4304 6866
rect 4252 6802 4304 6808
rect 4252 6656 4304 6662
rect 4158 6624 4214 6633
rect 4252 6598 4304 6604
rect 4158 6559 4214 6568
rect 3896 6344 4108 6372
rect 3896 5778 3924 6344
rect 4264 5930 4292 6598
rect 4356 6066 4384 7754
rect 4448 6458 4476 7840
rect 4528 7822 4580 7828
rect 4724 7002 4752 7919
rect 4908 7750 4936 8366
rect 4896 7744 4948 7750
rect 4896 7686 4948 7692
rect 4908 7342 4936 7686
rect 4896 7336 4948 7342
rect 4896 7278 4948 7284
rect 4712 6996 4764 7002
rect 4712 6938 4764 6944
rect 4804 6928 4856 6934
rect 4804 6870 4856 6876
rect 4712 6724 4764 6730
rect 4712 6666 4764 6672
rect 4528 6656 4580 6662
rect 4528 6598 4580 6604
rect 4436 6452 4488 6458
rect 4436 6394 4488 6400
rect 4356 6038 4476 6066
rect 4080 5902 4292 5930
rect 4448 5914 4476 6038
rect 4436 5908 4488 5914
rect 4080 5778 4108 5902
rect 4436 5850 4488 5856
rect 3884 5772 3936 5778
rect 3884 5714 3936 5720
rect 4068 5772 4120 5778
rect 4068 5714 4120 5720
rect 4344 5704 4396 5710
rect 4342 5672 4344 5681
rect 4396 5672 4398 5681
rect 4068 5636 4120 5642
rect 3804 5596 4016 5624
rect 3712 5545 3924 5556
rect 3712 5536 3938 5545
rect 3712 5528 3882 5536
rect 3454 5468 3750 5488
rect 3882 5471 3938 5480
rect 3510 5466 3534 5468
rect 3590 5466 3614 5468
rect 3670 5466 3694 5468
rect 3532 5414 3534 5466
rect 3596 5414 3608 5466
rect 3670 5414 3672 5466
rect 3510 5412 3534 5414
rect 3590 5412 3614 5414
rect 3670 5412 3694 5414
rect 3454 5392 3750 5412
rect 3882 5400 3938 5409
rect 3882 5335 3938 5344
rect 3792 5296 3844 5302
rect 3896 5284 3924 5335
rect 3844 5256 3924 5284
rect 3792 5238 3844 5244
rect 3988 5216 4016 5596
rect 4342 5607 4398 5616
rect 4068 5578 4120 5584
rect 4080 5250 4108 5578
rect 4436 5568 4488 5574
rect 4436 5510 4488 5516
rect 4080 5222 4292 5250
rect 3896 5188 4016 5216
rect 3516 5092 3568 5098
rect 3516 5034 3568 5040
rect 3608 5092 3660 5098
rect 3608 5034 3660 5040
rect 3528 5001 3556 5034
rect 3514 4992 3570 5001
rect 3514 4927 3570 4936
rect 3332 4820 3384 4826
rect 3332 4762 3384 4768
rect 3332 4684 3384 4690
rect 3332 4626 3384 4632
rect 3344 4282 3372 4626
rect 3620 4622 3648 5034
rect 3424 4616 3476 4622
rect 3422 4584 3424 4593
rect 3608 4616 3660 4622
rect 3476 4584 3478 4593
rect 3608 4558 3660 4564
rect 3422 4519 3478 4528
rect 3792 4480 3844 4486
rect 3792 4422 3844 4428
rect 3454 4380 3750 4400
rect 3510 4378 3534 4380
rect 3590 4378 3614 4380
rect 3670 4378 3694 4380
rect 3532 4326 3534 4378
rect 3596 4326 3608 4378
rect 3670 4326 3672 4378
rect 3510 4324 3534 4326
rect 3590 4324 3614 4326
rect 3670 4324 3694 4326
rect 3454 4304 3750 4324
rect 3332 4276 3384 4282
rect 3332 4218 3384 4224
rect 3608 4208 3660 4214
rect 3608 4150 3660 4156
rect 3424 4072 3476 4078
rect 3424 4014 3476 4020
rect 3330 3768 3386 3777
rect 3330 3703 3386 3712
rect 3344 3602 3372 3703
rect 3436 3602 3464 4014
rect 3332 3596 3384 3602
rect 3332 3538 3384 3544
rect 3424 3596 3476 3602
rect 3424 3538 3476 3544
rect 3620 3534 3648 4150
rect 3698 3632 3754 3641
rect 3698 3567 3700 3576
rect 3752 3567 3754 3576
rect 3700 3538 3752 3544
rect 3608 3528 3660 3534
rect 3608 3470 3660 3476
rect 3332 3460 3384 3466
rect 3332 3402 3384 3408
rect 3148 2926 3200 2932
rect 3238 2952 3294 2961
rect 2872 2576 2924 2582
rect 2872 2518 2924 2524
rect 3160 800 3188 2926
rect 3344 2922 3372 3402
rect 3454 3292 3750 3312
rect 3510 3290 3534 3292
rect 3590 3290 3614 3292
rect 3670 3290 3694 3292
rect 3532 3238 3534 3290
rect 3596 3238 3608 3290
rect 3670 3238 3672 3290
rect 3510 3236 3534 3238
rect 3590 3236 3614 3238
rect 3670 3236 3694 3238
rect 3454 3216 3750 3236
rect 3804 2938 3832 4422
rect 3896 4146 3924 5188
rect 4160 5160 4212 5166
rect 4160 5102 4212 5108
rect 4172 4690 4200 5102
rect 4160 4684 4212 4690
rect 4160 4626 4212 4632
rect 4066 4584 4122 4593
rect 4066 4519 4122 4528
rect 3884 4140 3936 4146
rect 3884 4082 3936 4088
rect 4080 4078 4108 4519
rect 4068 4072 4120 4078
rect 4068 4014 4120 4020
rect 3884 4004 3936 4010
rect 3884 3946 3936 3952
rect 3712 2922 3832 2938
rect 3896 2922 3924 3946
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 4080 3398 4108 3878
rect 4264 3738 4292 5222
rect 4344 4548 4396 4554
rect 4344 4490 4396 4496
rect 4356 4146 4384 4490
rect 4448 4321 4476 5510
rect 4434 4312 4490 4321
rect 4434 4247 4490 4256
rect 4344 4140 4396 4146
rect 4344 4082 4396 4088
rect 4436 4072 4488 4078
rect 4540 4060 4568 6598
rect 4724 5846 4752 6666
rect 4712 5840 4764 5846
rect 4712 5782 4764 5788
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 4632 5574 4660 5646
rect 4620 5568 4672 5574
rect 4620 5510 4672 5516
rect 4618 4992 4674 5001
rect 4618 4927 4674 4936
rect 4488 4032 4568 4060
rect 4436 4014 4488 4020
rect 4344 4004 4396 4010
rect 4344 3946 4396 3952
rect 4356 3913 4384 3946
rect 4342 3904 4398 3913
rect 4342 3839 4398 3848
rect 4252 3732 4304 3738
rect 4252 3674 4304 3680
rect 4540 3534 4568 4032
rect 4344 3528 4396 3534
rect 4344 3470 4396 3476
rect 4528 3528 4580 3534
rect 4528 3470 4580 3476
rect 4068 3392 4120 3398
rect 4068 3334 4120 3340
rect 4356 2990 4384 3470
rect 4526 3224 4582 3233
rect 4526 3159 4582 3168
rect 4540 2990 4568 3159
rect 4344 2984 4396 2990
rect 4344 2926 4396 2932
rect 4528 2984 4580 2990
rect 4528 2926 4580 2932
rect 3238 2887 3294 2896
rect 3332 2916 3384 2922
rect 3332 2858 3384 2864
rect 3700 2916 3832 2922
rect 3752 2910 3832 2916
rect 3884 2916 3936 2922
rect 3700 2858 3752 2864
rect 3884 2858 3936 2864
rect 4068 2848 4120 2854
rect 4068 2790 4120 2796
rect 3792 2508 3844 2514
rect 3792 2450 3844 2456
rect 3454 2204 3750 2224
rect 3510 2202 3534 2204
rect 3590 2202 3614 2204
rect 3670 2202 3694 2204
rect 3532 2150 3534 2202
rect 3596 2150 3608 2202
rect 3670 2150 3672 2202
rect 3510 2148 3534 2150
rect 3590 2148 3614 2150
rect 3670 2148 3694 2150
rect 3454 2128 3750 2148
rect 3804 1170 3832 2450
rect 3976 2372 4028 2378
rect 3976 2314 4028 2320
rect 3988 1170 4016 2314
rect 4080 2310 4108 2790
rect 4632 2582 4660 4927
rect 4724 4865 4752 5782
rect 4816 5370 4844 6870
rect 4908 6254 4936 7278
rect 5000 7206 5028 9046
rect 5368 8974 5396 10016
rect 6288 9926 6316 10406
rect 6380 10169 6408 11342
rect 6472 11286 6500 11698
rect 6460 11280 6512 11286
rect 6460 11222 6512 11228
rect 6552 10532 6604 10538
rect 6552 10474 6604 10480
rect 6460 10192 6512 10198
rect 6366 10160 6422 10169
rect 6460 10134 6512 10140
rect 6366 10095 6422 10104
rect 6276 9920 6328 9926
rect 6276 9862 6328 9868
rect 6472 9654 6500 10134
rect 6564 9926 6592 10474
rect 6552 9920 6604 9926
rect 6552 9862 6604 9868
rect 6276 9648 6328 9654
rect 5630 9616 5686 9625
rect 6276 9590 6328 9596
rect 6460 9648 6512 9654
rect 6460 9590 6512 9596
rect 5630 9551 5686 9560
rect 5448 9376 5500 9382
rect 5540 9376 5592 9382
rect 5448 9318 5500 9324
rect 5538 9344 5540 9353
rect 5592 9344 5594 9353
rect 5356 8968 5408 8974
rect 5356 8910 5408 8916
rect 5172 8832 5224 8838
rect 5078 8800 5134 8809
rect 5172 8774 5224 8780
rect 5078 8735 5134 8744
rect 5092 8090 5120 8735
rect 5184 8362 5212 8774
rect 5460 8362 5488 9318
rect 5538 9279 5594 9288
rect 5644 9081 5672 9551
rect 5953 9276 6249 9296
rect 6009 9274 6033 9276
rect 6089 9274 6113 9276
rect 6169 9274 6193 9276
rect 6031 9222 6033 9274
rect 6095 9222 6107 9274
rect 6169 9222 6171 9274
rect 6009 9220 6033 9222
rect 6089 9220 6113 9222
rect 6169 9220 6193 9222
rect 5953 9200 6249 9220
rect 6288 9110 6316 9590
rect 6564 9586 6592 9862
rect 6552 9580 6604 9586
rect 6552 9522 6604 9528
rect 6276 9104 6328 9110
rect 5630 9072 5686 9081
rect 6276 9046 6328 9052
rect 5630 9007 5686 9016
rect 6550 8664 6606 8673
rect 6550 8599 6606 8608
rect 6564 8566 6592 8599
rect 6552 8560 6604 8566
rect 6552 8502 6604 8508
rect 5172 8356 5224 8362
rect 5172 8298 5224 8304
rect 5448 8356 5500 8362
rect 5448 8298 5500 8304
rect 5184 8090 5212 8298
rect 6656 8294 6684 14334
rect 6734 14311 6790 14320
rect 6748 13870 6776 14311
rect 6736 13864 6788 13870
rect 6736 13806 6788 13812
rect 6840 13462 6868 14962
rect 6828 13456 6880 13462
rect 6828 13398 6880 13404
rect 6840 12442 6868 13398
rect 6932 12753 6960 15302
rect 7024 12889 7052 15438
rect 7196 15156 7248 15162
rect 7196 15098 7248 15104
rect 7104 14816 7156 14822
rect 7104 14758 7156 14764
rect 7116 13870 7144 14758
rect 7104 13864 7156 13870
rect 7208 13841 7236 15098
rect 7104 13806 7156 13812
rect 7194 13832 7250 13841
rect 7194 13767 7250 13776
rect 7196 13456 7248 13462
rect 7196 13398 7248 13404
rect 7208 12986 7236 13398
rect 7196 12980 7248 12986
rect 7196 12922 7248 12928
rect 7010 12880 7066 12889
rect 7010 12815 7066 12824
rect 6918 12744 6974 12753
rect 6918 12679 6974 12688
rect 6736 12436 6788 12442
rect 6736 12378 6788 12384
rect 6828 12436 6880 12442
rect 6828 12378 6880 12384
rect 6748 11529 6776 12378
rect 7196 12300 7248 12306
rect 7196 12242 7248 12248
rect 6734 11520 6790 11529
rect 6734 11455 6790 11464
rect 7208 11082 7236 12242
rect 7196 11076 7248 11082
rect 7196 11018 7248 11024
rect 7208 10305 7236 11018
rect 7194 10296 7250 10305
rect 7194 10231 7250 10240
rect 6826 10160 6882 10169
rect 6826 10095 6882 10104
rect 6840 9382 6868 10095
rect 7194 9752 7250 9761
rect 7194 9687 7250 9696
rect 6828 9376 6880 9382
rect 6828 9318 6880 9324
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6644 8288 6696 8294
rect 5814 8256 5870 8265
rect 6644 8230 6696 8236
rect 5814 8191 5870 8200
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 5172 8084 5224 8090
rect 5172 8026 5224 8032
rect 5170 7984 5226 7993
rect 5170 7919 5226 7928
rect 5724 7948 5776 7954
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 5080 7200 5132 7206
rect 5080 7142 5132 7148
rect 4896 6248 4948 6254
rect 4896 6190 4948 6196
rect 4804 5364 4856 5370
rect 4804 5306 4856 5312
rect 4804 5092 4856 5098
rect 4804 5034 4856 5040
rect 4816 5001 4844 5034
rect 4896 5024 4948 5030
rect 4802 4992 4858 5001
rect 4896 4966 4948 4972
rect 4802 4927 4858 4936
rect 4710 4856 4766 4865
rect 4710 4791 4766 4800
rect 4804 4820 4856 4826
rect 4804 4762 4856 4768
rect 4710 4312 4766 4321
rect 4816 4282 4844 4762
rect 4710 4247 4766 4256
rect 4804 4276 4856 4282
rect 4620 2576 4672 2582
rect 4620 2518 4672 2524
rect 4252 2508 4304 2514
rect 4252 2450 4304 2456
rect 4068 2304 4120 2310
rect 4068 2246 4120 2252
rect 4160 2304 4212 2310
rect 4160 2246 4212 2252
rect 3528 1142 3832 1170
rect 3896 1142 4016 1170
rect 3528 800 3556 1142
rect 3896 800 3924 1142
rect 4172 800 4200 2246
rect 4264 1766 4292 2450
rect 4724 2417 4752 4247
rect 4804 4218 4856 4224
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 4816 2990 4844 3878
rect 4908 3534 4936 4966
rect 4896 3528 4948 3534
rect 4896 3470 4948 3476
rect 5000 3058 5028 7142
rect 5092 6390 5120 7142
rect 5080 6384 5132 6390
rect 5080 6326 5132 6332
rect 5080 6248 5132 6254
rect 5080 6190 5132 6196
rect 5092 5234 5120 6190
rect 5184 5556 5212 7919
rect 5724 7890 5776 7896
rect 5632 7812 5684 7818
rect 5632 7754 5684 7760
rect 5448 7336 5500 7342
rect 5448 7278 5500 7284
rect 5262 7032 5318 7041
rect 5262 6967 5318 6976
rect 5276 6934 5304 6967
rect 5264 6928 5316 6934
rect 5264 6870 5316 6876
rect 5264 6452 5316 6458
rect 5264 6394 5316 6400
rect 5276 5624 5304 6394
rect 5460 6186 5488 7278
rect 5644 7206 5672 7754
rect 5632 7200 5684 7206
rect 5736 7177 5764 7890
rect 5828 7886 5856 8191
rect 5953 8188 6249 8208
rect 6009 8186 6033 8188
rect 6089 8186 6113 8188
rect 6169 8186 6193 8188
rect 6031 8134 6033 8186
rect 6095 8134 6107 8186
rect 6169 8134 6171 8186
rect 6009 8132 6033 8134
rect 6089 8132 6113 8134
rect 6169 8132 6193 8134
rect 5953 8112 6249 8132
rect 6932 8022 6960 8774
rect 6920 8016 6972 8022
rect 6920 7958 6972 7964
rect 5816 7880 5868 7886
rect 5816 7822 5868 7828
rect 7208 7750 7236 9687
rect 7300 9024 7328 15846
rect 7472 15564 7524 15570
rect 7576 15552 7604 15846
rect 7760 15570 7788 15846
rect 7944 15638 7972 15846
rect 8220 15745 8248 15914
rect 8206 15736 8262 15745
rect 8312 15706 8340 17002
rect 8496 16658 8524 17070
rect 8772 17066 8892 17082
rect 9128 17128 9180 17134
rect 9128 17070 9180 17076
rect 9864 17128 9916 17134
rect 9864 17070 9916 17076
rect 10232 17128 10284 17134
rect 10232 17070 10284 17076
rect 10600 17128 10652 17134
rect 10600 17070 10652 17076
rect 10692 17128 10744 17134
rect 10980 17116 11008 19200
rect 11348 17320 11376 19200
rect 11348 17292 11468 17320
rect 11440 17134 11468 17292
rect 11808 17134 11836 19200
rect 11060 17128 11112 17134
rect 10980 17088 11060 17116
rect 10692 17070 10744 17076
rect 11060 17070 11112 17076
rect 11336 17128 11388 17134
rect 11336 17070 11388 17076
rect 11428 17128 11480 17134
rect 11428 17070 11480 17076
rect 11796 17128 11848 17134
rect 11796 17070 11848 17076
rect 8760 17060 8892 17066
rect 8812 17054 8892 17060
rect 8944 17060 8996 17066
rect 8760 17002 8812 17008
rect 8944 17002 8996 17008
rect 8852 16992 8904 16998
rect 8852 16934 8904 16940
rect 8484 16652 8536 16658
rect 8484 16594 8536 16600
rect 8452 16348 8748 16368
rect 8508 16346 8532 16348
rect 8588 16346 8612 16348
rect 8668 16346 8692 16348
rect 8530 16294 8532 16346
rect 8594 16294 8606 16346
rect 8668 16294 8670 16346
rect 8508 16292 8532 16294
rect 8588 16292 8612 16294
rect 8668 16292 8692 16294
rect 8452 16272 8748 16292
rect 8206 15671 8262 15680
rect 8300 15700 8352 15706
rect 8300 15642 8352 15648
rect 7932 15632 7984 15638
rect 7932 15574 7984 15580
rect 7524 15524 7604 15552
rect 7472 15506 7524 15512
rect 7472 14884 7524 14890
rect 7472 14826 7524 14832
rect 7380 14272 7432 14278
rect 7380 14214 7432 14220
rect 7392 13161 7420 14214
rect 7484 13569 7512 14826
rect 7576 13734 7604 15524
rect 7748 15564 7800 15570
rect 7748 15506 7800 15512
rect 7656 15496 7708 15502
rect 7656 15438 7708 15444
rect 7668 15094 7696 15438
rect 7656 15088 7708 15094
rect 7656 15030 7708 15036
rect 7668 14550 7696 15030
rect 7748 14816 7800 14822
rect 7748 14758 7800 14764
rect 7656 14544 7708 14550
rect 7656 14486 7708 14492
rect 7656 14408 7708 14414
rect 7656 14350 7708 14356
rect 7564 13728 7616 13734
rect 7564 13670 7616 13676
rect 7470 13560 7526 13569
rect 7470 13495 7526 13504
rect 7378 13152 7434 13161
rect 7378 13087 7434 13096
rect 7472 9376 7524 9382
rect 7576 9364 7604 13670
rect 7668 13190 7696 14350
rect 7656 13184 7708 13190
rect 7656 13126 7708 13132
rect 7656 12776 7708 12782
rect 7656 12718 7708 12724
rect 7668 12306 7696 12718
rect 7760 12442 7788 14758
rect 7944 14550 7972 15574
rect 8208 15564 8260 15570
rect 8208 15506 8260 15512
rect 8300 15564 8352 15570
rect 8300 15506 8352 15512
rect 8668 15564 8720 15570
rect 8668 15506 8720 15512
rect 8024 15496 8076 15502
rect 8220 15473 8248 15506
rect 8024 15438 8076 15444
rect 8206 15464 8262 15473
rect 8036 15026 8064 15438
rect 8206 15399 8262 15408
rect 8024 15020 8076 15026
rect 8024 14962 8076 14968
rect 7932 14544 7984 14550
rect 7932 14486 7984 14492
rect 8024 14408 8076 14414
rect 7838 14376 7894 14385
rect 8024 14350 8076 14356
rect 7838 14311 7840 14320
rect 7892 14311 7894 14320
rect 7840 14282 7892 14288
rect 7932 14000 7984 14006
rect 7932 13942 7984 13948
rect 7840 13864 7892 13870
rect 7840 13806 7892 13812
rect 7852 13190 7880 13806
rect 7840 13184 7892 13190
rect 7840 13126 7892 13132
rect 7852 12782 7880 13126
rect 7840 12776 7892 12782
rect 7840 12718 7892 12724
rect 7748 12436 7800 12442
rect 7748 12378 7800 12384
rect 7656 12300 7708 12306
rect 7656 12242 7708 12248
rect 7944 12209 7972 13942
rect 8036 13462 8064 14350
rect 8116 14340 8168 14346
rect 8116 14282 8168 14288
rect 8128 13938 8156 14282
rect 8208 14272 8260 14278
rect 8208 14214 8260 14220
rect 8220 14006 8248 14214
rect 8208 14000 8260 14006
rect 8208 13942 8260 13948
rect 8116 13932 8168 13938
rect 8116 13874 8168 13880
rect 8024 13456 8076 13462
rect 8024 13398 8076 13404
rect 8022 13288 8078 13297
rect 8022 13223 8078 13232
rect 8036 12714 8064 13223
rect 8128 12986 8156 13874
rect 8208 13796 8260 13802
rect 8208 13738 8260 13744
rect 8220 13705 8248 13738
rect 8206 13696 8262 13705
rect 8206 13631 8262 13640
rect 8116 12980 8168 12986
rect 8116 12922 8168 12928
rect 8024 12708 8076 12714
rect 8024 12650 8076 12656
rect 7930 12200 7986 12209
rect 7930 12135 7986 12144
rect 7932 12096 7984 12102
rect 7932 12038 7984 12044
rect 7944 11898 7972 12038
rect 7932 11892 7984 11898
rect 7932 11834 7984 11840
rect 8312 11778 8340 15506
rect 8680 15348 8708 15506
rect 8864 15502 8892 16934
rect 8956 16250 8984 17002
rect 9036 16652 9088 16658
rect 9036 16594 9088 16600
rect 8944 16244 8996 16250
rect 8944 16186 8996 16192
rect 8852 15496 8904 15502
rect 8852 15438 8904 15444
rect 8680 15320 8892 15348
rect 8452 15260 8748 15280
rect 8508 15258 8532 15260
rect 8588 15258 8612 15260
rect 8668 15258 8692 15260
rect 8530 15206 8532 15258
rect 8594 15206 8606 15258
rect 8668 15206 8670 15258
rect 8508 15204 8532 15206
rect 8588 15204 8612 15206
rect 8668 15204 8692 15206
rect 8452 15184 8748 15204
rect 8758 15056 8814 15065
rect 8668 15020 8720 15026
rect 8758 14991 8760 15000
rect 8668 14962 8720 14968
rect 8812 14991 8814 15000
rect 8760 14962 8812 14968
rect 8392 14884 8444 14890
rect 8392 14826 8444 14832
rect 8404 14550 8432 14826
rect 8392 14544 8444 14550
rect 8392 14486 8444 14492
rect 8680 14414 8708 14962
rect 8668 14408 8720 14414
rect 8668 14350 8720 14356
rect 8452 14172 8748 14192
rect 8508 14170 8532 14172
rect 8588 14170 8612 14172
rect 8668 14170 8692 14172
rect 8530 14118 8532 14170
rect 8594 14118 8606 14170
rect 8668 14118 8670 14170
rect 8508 14116 8532 14118
rect 8588 14116 8612 14118
rect 8668 14116 8692 14118
rect 8452 14096 8748 14116
rect 8392 13864 8444 13870
rect 8392 13806 8444 13812
rect 8482 13832 8538 13841
rect 8404 13530 8432 13806
rect 8482 13767 8538 13776
rect 8668 13796 8720 13802
rect 8496 13734 8524 13767
rect 8668 13738 8720 13744
rect 8484 13728 8536 13734
rect 8484 13670 8536 13676
rect 8680 13530 8708 13738
rect 8392 13524 8444 13530
rect 8392 13466 8444 13472
rect 8668 13524 8720 13530
rect 8668 13466 8720 13472
rect 8864 13394 8892 15320
rect 9048 15162 9076 16594
rect 9140 15706 9168 17070
rect 9404 17060 9456 17066
rect 9404 17002 9456 17008
rect 9312 16992 9364 16998
rect 9312 16934 9364 16940
rect 9220 16108 9272 16114
rect 9220 16050 9272 16056
rect 9128 15700 9180 15706
rect 9128 15642 9180 15648
rect 9232 15502 9260 16050
rect 9324 15978 9352 16934
rect 9312 15972 9364 15978
rect 9312 15914 9364 15920
rect 9220 15496 9272 15502
rect 9220 15438 9272 15444
rect 9036 15156 9088 15162
rect 9036 15098 9088 15104
rect 9128 15156 9180 15162
rect 9128 15098 9180 15104
rect 9140 14822 9168 15098
rect 9128 14816 9180 14822
rect 9128 14758 9180 14764
rect 9324 14550 9352 15914
rect 9416 15706 9444 17002
rect 9876 16794 9904 17070
rect 10232 16992 10284 16998
rect 10232 16934 10284 16940
rect 10508 16992 10560 16998
rect 10508 16934 10560 16940
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 9864 16788 9916 16794
rect 9864 16730 9916 16736
rect 9588 16040 9640 16046
rect 9588 15982 9640 15988
rect 9496 15904 9548 15910
rect 9494 15872 9496 15881
rect 9548 15872 9550 15881
rect 9494 15807 9550 15816
rect 9404 15700 9456 15706
rect 9404 15642 9456 15648
rect 9496 15496 9548 15502
rect 9496 15438 9548 15444
rect 8944 14544 8996 14550
rect 8944 14486 8996 14492
rect 9312 14544 9364 14550
rect 9312 14486 9364 14492
rect 8956 13734 8984 14486
rect 9404 14340 9456 14346
rect 9404 14282 9456 14288
rect 9036 14272 9088 14278
rect 9036 14214 9088 14220
rect 9312 14272 9364 14278
rect 9312 14214 9364 14220
rect 9057 14090 9085 14214
rect 9048 14062 9085 14090
rect 9048 13938 9076 14062
rect 9126 13968 9182 13977
rect 9036 13932 9088 13938
rect 9126 13903 9182 13912
rect 9036 13874 9088 13880
rect 9140 13734 9168 13903
rect 9324 13841 9352 14214
rect 9310 13832 9366 13841
rect 9310 13767 9366 13776
rect 8944 13728 8996 13734
rect 9128 13728 9180 13734
rect 8944 13670 8996 13676
rect 9034 13696 9090 13705
rect 9128 13670 9180 13676
rect 9312 13728 9364 13734
rect 9312 13670 9364 13676
rect 9034 13631 9090 13640
rect 9048 13530 9076 13631
rect 9126 13560 9182 13569
rect 9036 13524 9088 13530
rect 9126 13495 9182 13504
rect 9036 13466 9088 13472
rect 8944 13456 8996 13462
rect 8944 13398 8996 13404
rect 8852 13388 8904 13394
rect 8852 13330 8904 13336
rect 8852 13252 8904 13258
rect 8852 13194 8904 13200
rect 8452 13084 8748 13104
rect 8508 13082 8532 13084
rect 8588 13082 8612 13084
rect 8668 13082 8692 13084
rect 8530 13030 8532 13082
rect 8594 13030 8606 13082
rect 8668 13030 8670 13082
rect 8508 13028 8532 13030
rect 8588 13028 8612 13030
rect 8668 13028 8692 13030
rect 8452 13008 8748 13028
rect 8760 12708 8812 12714
rect 8760 12650 8812 12656
rect 8772 12481 8800 12650
rect 8758 12472 8814 12481
rect 8758 12407 8814 12416
rect 8864 12306 8892 13194
rect 8956 12714 8984 13398
rect 9140 13258 9168 13495
rect 9324 13297 9352 13670
rect 9416 13462 9444 14282
rect 9508 14074 9536 15438
rect 9496 14068 9548 14074
rect 9496 14010 9548 14016
rect 9600 13954 9628 15982
rect 9692 15706 9720 16730
rect 9956 16720 10008 16726
rect 9956 16662 10008 16668
rect 9772 16584 9824 16590
rect 9770 16552 9772 16561
rect 9824 16552 9826 16561
rect 9770 16487 9826 16496
rect 9772 16448 9824 16454
rect 9772 16390 9824 16396
rect 9680 15700 9732 15706
rect 9680 15642 9732 15648
rect 9784 15065 9812 16390
rect 9968 15706 9996 16662
rect 9956 15700 10008 15706
rect 9956 15642 10008 15648
rect 9864 15564 9916 15570
rect 9864 15506 9916 15512
rect 10140 15564 10192 15570
rect 10140 15506 10192 15512
rect 9876 15366 9904 15506
rect 9864 15360 9916 15366
rect 9864 15302 9916 15308
rect 9876 15162 9904 15302
rect 9864 15156 9916 15162
rect 9864 15098 9916 15104
rect 10048 15088 10100 15094
rect 9770 15056 9826 15065
rect 10048 15030 10100 15036
rect 9770 14991 9826 15000
rect 9864 14612 9916 14618
rect 9864 14554 9916 14560
rect 9678 14376 9734 14385
rect 9678 14311 9680 14320
rect 9732 14311 9734 14320
rect 9680 14282 9732 14288
rect 9678 13968 9734 13977
rect 9600 13926 9678 13954
rect 9678 13903 9734 13912
rect 9494 13832 9550 13841
rect 9494 13767 9550 13776
rect 9404 13456 9456 13462
rect 9404 13398 9456 13404
rect 9404 13320 9456 13326
rect 9310 13288 9366 13297
rect 9128 13252 9180 13258
rect 9404 13262 9456 13268
rect 9310 13223 9366 13232
rect 9128 13194 9180 13200
rect 9128 12912 9180 12918
rect 9126 12880 9128 12889
rect 9180 12880 9182 12889
rect 9416 12866 9444 13262
rect 9036 12844 9088 12850
rect 9182 12838 9260 12866
rect 9126 12815 9182 12824
rect 9036 12786 9088 12792
rect 8944 12708 8996 12714
rect 8944 12650 8996 12656
rect 8942 12608 8998 12617
rect 8942 12543 8998 12552
rect 8852 12300 8904 12306
rect 8852 12242 8904 12248
rect 8452 11996 8748 12016
rect 8508 11994 8532 11996
rect 8588 11994 8612 11996
rect 8668 11994 8692 11996
rect 8530 11942 8532 11994
rect 8594 11942 8606 11994
rect 8668 11942 8670 11994
rect 8508 11940 8532 11942
rect 8588 11940 8612 11942
rect 8668 11940 8692 11942
rect 8452 11920 8748 11940
rect 8312 11750 8432 11778
rect 8300 11688 8352 11694
rect 8300 11630 8352 11636
rect 7840 11552 7892 11558
rect 7840 11494 7892 11500
rect 7852 11286 7880 11494
rect 7840 11280 7892 11286
rect 8208 11280 8260 11286
rect 7840 11222 7892 11228
rect 7944 11240 8208 11268
rect 7944 11098 7972 11240
rect 8208 11222 8260 11228
rect 7668 11070 7972 11098
rect 8114 11112 8170 11121
rect 7668 9654 7696 11070
rect 8114 11047 8170 11056
rect 7932 11008 7984 11014
rect 7932 10950 7984 10956
rect 7944 10606 7972 10950
rect 7932 10600 7984 10606
rect 7932 10542 7984 10548
rect 7746 10432 7802 10441
rect 7746 10367 7802 10376
rect 7656 9648 7708 9654
rect 7656 9590 7708 9596
rect 7524 9336 7604 9364
rect 7472 9318 7524 9324
rect 7300 8996 7420 9024
rect 7286 8936 7342 8945
rect 7286 8871 7342 8880
rect 7300 8401 7328 8871
rect 7392 8650 7420 8996
rect 7484 8809 7512 9318
rect 7760 8922 7788 10367
rect 7944 9926 7972 10542
rect 8024 10532 8076 10538
rect 8024 10474 8076 10480
rect 8036 9994 8064 10474
rect 8024 9988 8076 9994
rect 8024 9930 8076 9936
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 7840 9512 7892 9518
rect 7944 9500 7972 9862
rect 7892 9472 7972 9500
rect 8128 9489 8156 11047
rect 8312 10266 8340 11630
rect 8404 11558 8432 11750
rect 8392 11552 8444 11558
rect 8392 11494 8444 11500
rect 8852 11552 8904 11558
rect 8852 11494 8904 11500
rect 8452 10908 8748 10928
rect 8508 10906 8532 10908
rect 8588 10906 8612 10908
rect 8668 10906 8692 10908
rect 8530 10854 8532 10906
rect 8594 10854 8606 10906
rect 8668 10854 8670 10906
rect 8508 10852 8532 10854
rect 8588 10852 8612 10854
rect 8668 10852 8692 10854
rect 8452 10832 8748 10852
rect 8668 10600 8720 10606
rect 8668 10542 8720 10548
rect 8680 10470 8708 10542
rect 8864 10470 8892 11494
rect 8668 10464 8720 10470
rect 8852 10464 8904 10470
rect 8668 10406 8720 10412
rect 8850 10432 8852 10441
rect 8904 10432 8906 10441
rect 8300 10260 8352 10266
rect 8300 10202 8352 10208
rect 8680 10062 8708 10406
rect 8850 10367 8906 10376
rect 8850 10296 8906 10305
rect 8850 10231 8906 10240
rect 8864 10130 8892 10231
rect 8956 10198 8984 12543
rect 9048 11694 9076 12786
rect 9126 12608 9182 12617
rect 9126 12543 9182 12552
rect 9036 11688 9088 11694
rect 9036 11630 9088 11636
rect 9034 11520 9090 11529
rect 9034 11455 9090 11464
rect 9048 10198 9076 11455
rect 9140 11132 9168 12543
rect 9232 12356 9260 12838
rect 9324 12838 9444 12866
rect 9324 12646 9352 12838
rect 9312 12640 9364 12646
rect 9312 12582 9364 12588
rect 9312 12368 9364 12374
rect 9232 12328 9312 12356
rect 9312 12310 9364 12316
rect 9508 12102 9536 13767
rect 9680 13728 9732 13734
rect 9678 13696 9680 13705
rect 9732 13696 9734 13705
rect 9678 13631 9734 13640
rect 9876 13530 9904 14554
rect 9956 14408 10008 14414
rect 9956 14350 10008 14356
rect 9864 13524 9916 13530
rect 9864 13466 9916 13472
rect 9588 13456 9640 13462
rect 9588 13398 9640 13404
rect 9312 12096 9364 12102
rect 9312 12038 9364 12044
rect 9496 12096 9548 12102
rect 9496 12038 9548 12044
rect 9324 11762 9352 12038
rect 9312 11756 9364 11762
rect 9312 11698 9364 11704
rect 9508 11558 9536 12038
rect 9404 11552 9456 11558
rect 9404 11494 9456 11500
rect 9496 11552 9548 11558
rect 9496 11494 9548 11500
rect 9140 11104 9260 11132
rect 9128 10668 9180 10674
rect 9128 10610 9180 10616
rect 8944 10192 8996 10198
rect 8944 10134 8996 10140
rect 9036 10192 9088 10198
rect 9036 10134 9088 10140
rect 8852 10124 8904 10130
rect 8852 10066 8904 10072
rect 8668 10056 8720 10062
rect 8668 9998 8720 10004
rect 8452 9820 8748 9840
rect 8508 9818 8532 9820
rect 8588 9818 8612 9820
rect 8668 9818 8692 9820
rect 8530 9766 8532 9818
rect 8594 9766 8606 9818
rect 8668 9766 8670 9818
rect 8508 9764 8532 9766
rect 8588 9764 8612 9766
rect 8668 9764 8692 9766
rect 8452 9744 8748 9764
rect 8114 9480 8170 9489
rect 7840 9454 7892 9460
rect 8114 9415 8170 9424
rect 8114 9208 8170 9217
rect 8114 9143 8170 9152
rect 7932 9104 7984 9110
rect 8128 9092 8156 9143
rect 7984 9064 8156 9092
rect 7932 9046 7984 9052
rect 8208 9036 8260 9042
rect 8208 8978 8260 8984
rect 7760 8894 8064 8922
rect 7932 8832 7984 8838
rect 7470 8800 7526 8809
rect 7932 8774 7984 8780
rect 7470 8735 7526 8744
rect 7392 8622 7696 8650
rect 7286 8392 7342 8401
rect 7286 8327 7342 8336
rect 6000 7744 6052 7750
rect 6000 7686 6052 7692
rect 6460 7744 6512 7750
rect 6460 7686 6512 7692
rect 6828 7744 6880 7750
rect 7196 7744 7248 7750
rect 6880 7704 6960 7732
rect 6828 7686 6880 7692
rect 6012 7342 6040 7686
rect 6368 7472 6420 7478
rect 6368 7414 6420 7420
rect 6000 7336 6052 7342
rect 6000 7278 6052 7284
rect 5816 7200 5868 7206
rect 5632 7142 5684 7148
rect 5722 7168 5778 7177
rect 6380 7177 6408 7414
rect 5816 7142 5868 7148
rect 6366 7168 6422 7177
rect 5722 7103 5778 7112
rect 5724 6860 5776 6866
rect 5724 6802 5776 6808
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 5552 6458 5580 6734
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5448 6180 5500 6186
rect 5448 6122 5500 6128
rect 5736 6118 5764 6802
rect 5828 6186 5856 7142
rect 5953 7100 6249 7120
rect 6366 7103 6422 7112
rect 6009 7098 6033 7100
rect 6089 7098 6113 7100
rect 6169 7098 6193 7100
rect 6031 7046 6033 7098
rect 6095 7046 6107 7098
rect 6169 7046 6171 7098
rect 6009 7044 6033 7046
rect 6089 7044 6113 7046
rect 6169 7044 6193 7046
rect 5953 7024 6249 7044
rect 6472 7041 6500 7686
rect 6458 7032 6514 7041
rect 6458 6967 6514 6976
rect 6092 6928 6144 6934
rect 6460 6928 6512 6934
rect 6288 6888 6460 6916
rect 6288 6882 6316 6888
rect 6144 6876 6316 6882
rect 6092 6870 6316 6876
rect 6460 6870 6512 6876
rect 6104 6854 6316 6870
rect 6736 6724 6788 6730
rect 6736 6666 6788 6672
rect 6460 6248 6512 6254
rect 6460 6190 6512 6196
rect 5816 6180 5868 6186
rect 5816 6122 5868 6128
rect 6368 6180 6420 6186
rect 6368 6122 6420 6128
rect 5724 6112 5776 6118
rect 5724 6054 5776 6060
rect 5828 5953 5856 6122
rect 5953 6012 6249 6032
rect 6009 6010 6033 6012
rect 6089 6010 6113 6012
rect 6169 6010 6193 6012
rect 6031 5958 6033 6010
rect 6095 5958 6107 6010
rect 6169 5958 6171 6010
rect 6009 5956 6033 5958
rect 6089 5956 6113 5958
rect 6169 5956 6193 5958
rect 5814 5944 5870 5953
rect 5953 5936 6249 5956
rect 5814 5879 5870 5888
rect 5356 5772 5408 5778
rect 5540 5772 5592 5778
rect 5408 5732 5488 5760
rect 5356 5714 5408 5720
rect 5276 5596 5396 5624
rect 5184 5528 5304 5556
rect 5172 5364 5224 5370
rect 5172 5306 5224 5312
rect 5080 5228 5132 5234
rect 5080 5170 5132 5176
rect 5184 4554 5212 5306
rect 5276 5098 5304 5528
rect 5264 5092 5316 5098
rect 5264 5034 5316 5040
rect 5368 5001 5396 5596
rect 5354 4992 5410 5001
rect 5354 4927 5410 4936
rect 5172 4548 5224 4554
rect 5172 4490 5224 4496
rect 5264 4480 5316 4486
rect 5264 4422 5316 4428
rect 5356 4480 5408 4486
rect 5356 4422 5408 4428
rect 5172 4276 5224 4282
rect 5172 4218 5224 4224
rect 5184 4146 5212 4218
rect 5172 4140 5224 4146
rect 5172 4082 5224 4088
rect 5080 3936 5132 3942
rect 5078 3904 5080 3913
rect 5132 3904 5134 3913
rect 5078 3839 5134 3848
rect 5170 3768 5226 3777
rect 5276 3738 5304 4422
rect 5368 4282 5396 4422
rect 5356 4276 5408 4282
rect 5356 4218 5408 4224
rect 5354 3904 5410 3913
rect 5354 3839 5410 3848
rect 5368 3738 5396 3839
rect 5170 3703 5226 3712
rect 5264 3732 5316 3738
rect 5184 3602 5212 3703
rect 5264 3674 5316 3680
rect 5356 3732 5408 3738
rect 5356 3674 5408 3680
rect 5080 3596 5132 3602
rect 5080 3538 5132 3544
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 5092 3194 5120 3538
rect 5460 3369 5488 5732
rect 5540 5714 5592 5720
rect 5816 5772 5868 5778
rect 5816 5714 5868 5720
rect 5552 5030 5580 5714
rect 5828 5658 5856 5714
rect 5644 5630 5856 5658
rect 6380 5642 6408 6122
rect 6472 5846 6500 6190
rect 6552 6180 6604 6186
rect 6552 6122 6604 6128
rect 6460 5840 6512 5846
rect 6460 5782 6512 5788
rect 6368 5636 6420 5642
rect 5644 5545 5672 5630
rect 6288 5596 6368 5624
rect 5630 5536 5686 5545
rect 5630 5471 5686 5480
rect 5814 5536 5870 5545
rect 5814 5471 5870 5480
rect 5632 5092 5684 5098
rect 5632 5034 5684 5040
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5538 4448 5594 4457
rect 5538 4383 5594 4392
rect 5170 3360 5226 3369
rect 5170 3295 5226 3304
rect 5446 3360 5502 3369
rect 5446 3295 5502 3304
rect 5080 3188 5132 3194
rect 5080 3130 5132 3136
rect 4988 3052 5040 3058
rect 4988 2994 5040 3000
rect 4804 2984 4856 2990
rect 4804 2926 4856 2932
rect 5078 2952 5134 2961
rect 4896 2916 4948 2922
rect 5184 2922 5212 3295
rect 5552 2990 5580 4383
rect 5644 3482 5672 5034
rect 5724 5024 5776 5030
rect 5724 4966 5776 4972
rect 5736 3584 5764 4966
rect 5828 4758 5856 5471
rect 5953 4924 6249 4944
rect 6009 4922 6033 4924
rect 6089 4922 6113 4924
rect 6169 4922 6193 4924
rect 6031 4870 6033 4922
rect 6095 4870 6107 4922
rect 6169 4870 6171 4922
rect 6009 4868 6033 4870
rect 6089 4868 6113 4870
rect 6169 4868 6193 4870
rect 5953 4848 6249 4868
rect 5816 4752 5868 4758
rect 5816 4694 5868 4700
rect 5814 4448 5870 4457
rect 5814 4383 5870 4392
rect 5828 3720 5856 4383
rect 5908 4208 5960 4214
rect 6288 4196 6316 5596
rect 6368 5578 6420 5584
rect 6472 5166 6500 5782
rect 6564 5409 6592 6122
rect 6644 5568 6696 5574
rect 6748 5545 6776 6666
rect 6932 6089 6960 7704
rect 7196 7686 7248 7692
rect 7564 7268 7616 7274
rect 7564 7210 7616 7216
rect 7576 6934 7604 7210
rect 7564 6928 7616 6934
rect 7564 6870 7616 6876
rect 7012 6656 7064 6662
rect 7012 6598 7064 6604
rect 7104 6656 7156 6662
rect 7104 6598 7156 6604
rect 7024 6186 7052 6598
rect 7012 6180 7064 6186
rect 7012 6122 7064 6128
rect 6918 6080 6974 6089
rect 6918 6015 6974 6024
rect 7012 5772 7064 5778
rect 7012 5714 7064 5720
rect 6920 5568 6972 5574
rect 6644 5510 6696 5516
rect 6734 5536 6790 5545
rect 6550 5400 6606 5409
rect 6550 5335 6606 5344
rect 6460 5160 6512 5166
rect 6460 5102 6512 5108
rect 6472 4842 6500 5102
rect 6656 5098 6684 5510
rect 6920 5510 6972 5516
rect 6734 5471 6790 5480
rect 6552 5092 6604 5098
rect 6552 5034 6604 5040
rect 6644 5092 6696 5098
rect 6644 5034 6696 5040
rect 6564 4978 6592 5034
rect 6564 4950 6776 4978
rect 6472 4814 6592 4842
rect 6460 4684 6512 4690
rect 5960 4168 6316 4196
rect 5908 4150 5960 4156
rect 5953 3836 6249 3856
rect 6009 3834 6033 3836
rect 6089 3834 6113 3836
rect 6169 3834 6193 3836
rect 6031 3782 6033 3834
rect 6095 3782 6107 3834
rect 6169 3782 6171 3834
rect 6009 3780 6033 3782
rect 6089 3780 6113 3782
rect 6169 3780 6193 3782
rect 5953 3760 6249 3780
rect 6288 3720 6316 4168
rect 6380 4644 6460 4672
rect 6380 4010 6408 4644
rect 6564 4672 6592 4814
rect 6644 4684 6696 4690
rect 6564 4644 6644 4672
rect 6460 4626 6512 4632
rect 6644 4626 6696 4632
rect 6458 4312 6514 4321
rect 6656 4298 6684 4626
rect 6748 4486 6776 4950
rect 6828 4616 6880 4622
rect 6828 4558 6880 4564
rect 6736 4480 6788 4486
rect 6736 4422 6788 4428
rect 6514 4270 6684 4298
rect 6458 4247 6514 4256
rect 6472 4078 6500 4247
rect 6460 4072 6512 4078
rect 6460 4014 6512 4020
rect 6368 4004 6420 4010
rect 6368 3946 6420 3952
rect 5828 3692 5948 3720
rect 5920 3602 5948 3692
rect 6196 3692 6316 3720
rect 5908 3596 5960 3602
rect 5736 3556 5856 3584
rect 5644 3466 5764 3482
rect 5644 3460 5776 3466
rect 5644 3454 5724 3460
rect 5724 3402 5776 3408
rect 5632 3392 5684 3398
rect 5632 3334 5684 3340
rect 5540 2984 5592 2990
rect 5540 2926 5592 2932
rect 5078 2887 5080 2896
rect 4896 2858 4948 2864
rect 5132 2887 5134 2896
rect 5172 2916 5224 2922
rect 5080 2858 5132 2864
rect 5172 2858 5224 2864
rect 4908 2774 4936 2858
rect 4908 2746 5304 2774
rect 4804 2508 4856 2514
rect 4804 2450 4856 2456
rect 5172 2508 5224 2514
rect 5172 2450 5224 2456
rect 4710 2408 4766 2417
rect 4528 2372 4580 2378
rect 4710 2343 4766 2352
rect 4528 2314 4580 2320
rect 4252 1760 4304 1766
rect 4252 1702 4304 1708
rect 4540 800 4568 2314
rect 4816 1698 4844 2450
rect 4896 2440 4948 2446
rect 4896 2382 4948 2388
rect 4804 1692 4856 1698
rect 4804 1634 4856 1640
rect 4908 800 4936 2382
rect 5184 1834 5212 2450
rect 5172 1828 5224 1834
rect 5172 1770 5224 1776
rect 5276 800 5304 2746
rect 5644 2650 5672 3334
rect 5828 2990 5856 3556
rect 5908 3538 5960 3544
rect 6196 3058 6224 3692
rect 6380 3534 6408 3946
rect 6460 3936 6512 3942
rect 6458 3904 6460 3913
rect 6512 3904 6514 3913
rect 6458 3839 6514 3848
rect 6550 3768 6606 3777
rect 6550 3703 6606 3712
rect 6460 3664 6512 3670
rect 6460 3606 6512 3612
rect 6368 3528 6420 3534
rect 6368 3470 6420 3476
rect 6276 3392 6328 3398
rect 6276 3334 6328 3340
rect 6288 3058 6316 3334
rect 6184 3052 6236 3058
rect 6184 2994 6236 3000
rect 6276 3052 6328 3058
rect 6276 2994 6328 3000
rect 5816 2984 5868 2990
rect 5816 2926 5868 2932
rect 6274 2952 6330 2961
rect 6380 2922 6408 3470
rect 6274 2887 6330 2896
rect 6368 2916 6420 2922
rect 5953 2748 6249 2768
rect 6009 2746 6033 2748
rect 6089 2746 6113 2748
rect 6169 2746 6193 2748
rect 6031 2694 6033 2746
rect 6095 2694 6107 2746
rect 6169 2694 6171 2746
rect 6009 2692 6033 2694
rect 6089 2692 6113 2694
rect 6169 2692 6193 2694
rect 5953 2672 6249 2692
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 5908 2100 5960 2106
rect 5908 2042 5960 2048
rect 5540 1420 5592 1426
rect 5540 1362 5592 1368
rect 5552 800 5580 1362
rect 5920 800 5948 2042
rect 6012 1630 6040 2450
rect 6288 2446 6316 2887
rect 6368 2858 6420 2864
rect 6472 2650 6500 3606
rect 6564 3369 6592 3703
rect 6644 3664 6696 3670
rect 6644 3606 6696 3612
rect 6550 3360 6606 3369
rect 6550 3295 6606 3304
rect 6550 2816 6606 2825
rect 6550 2751 6606 2760
rect 6460 2644 6512 2650
rect 6460 2586 6512 2592
rect 6564 2553 6592 2751
rect 6550 2544 6606 2553
rect 6550 2479 6606 2488
rect 6092 2440 6144 2446
rect 6090 2408 6092 2417
rect 6276 2440 6328 2446
rect 6144 2408 6146 2417
rect 6276 2382 6328 2388
rect 6090 2343 6146 2352
rect 6564 2310 6592 2479
rect 6552 2304 6604 2310
rect 6552 2246 6604 2252
rect 6276 2032 6328 2038
rect 6276 1974 6328 1980
rect 6000 1624 6052 1630
rect 6000 1566 6052 1572
rect 6288 800 6316 1974
rect 6656 800 6684 3606
rect 6748 2922 6776 4422
rect 6840 2990 6868 4558
rect 6828 2984 6880 2990
rect 6828 2926 6880 2932
rect 6736 2916 6788 2922
rect 6736 2858 6788 2864
rect 6932 2854 6960 5510
rect 7024 5030 7052 5714
rect 7012 5024 7064 5030
rect 7012 4966 7064 4972
rect 7012 3460 7064 3466
rect 7012 3402 7064 3408
rect 6920 2848 6972 2854
rect 7024 2825 7052 3402
rect 6920 2790 6972 2796
rect 7010 2816 7066 2825
rect 7010 2751 7066 2760
rect 7116 2650 7144 6598
rect 7378 6488 7434 6497
rect 7378 6423 7434 6432
rect 7392 5953 7420 6423
rect 7576 6118 7604 6870
rect 7472 6112 7524 6118
rect 7472 6054 7524 6060
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 7378 5944 7434 5953
rect 7378 5879 7434 5888
rect 7484 5302 7512 6054
rect 7472 5296 7524 5302
rect 7208 5256 7472 5284
rect 7104 2644 7156 2650
rect 7104 2586 7156 2592
rect 6920 2508 6972 2514
rect 6840 2468 6920 2496
rect 6840 1970 6868 2468
rect 6920 2450 6972 2456
rect 7208 2446 7236 5256
rect 7472 5238 7524 5244
rect 7288 5024 7340 5030
rect 7288 4966 7340 4972
rect 7300 3942 7328 4966
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 7392 4282 7420 4626
rect 7380 4276 7432 4282
rect 7380 4218 7432 4224
rect 7472 4208 7524 4214
rect 7472 4150 7524 4156
rect 7380 4004 7432 4010
rect 7380 3946 7432 3952
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 7392 3466 7420 3946
rect 7484 3738 7512 4150
rect 7472 3732 7524 3738
rect 7472 3674 7524 3680
rect 7380 3460 7432 3466
rect 7380 3402 7432 3408
rect 7286 3088 7342 3097
rect 7286 3023 7342 3032
rect 7300 2922 7328 3023
rect 7288 2916 7340 2922
rect 7288 2858 7340 2864
rect 7380 2916 7432 2922
rect 7380 2858 7432 2864
rect 7392 2774 7420 2858
rect 7300 2746 7420 2774
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 6828 1964 6880 1970
rect 6828 1906 6880 1912
rect 6920 1556 6972 1562
rect 6920 1498 6972 1504
rect 6932 800 6960 1498
rect 7300 800 7328 2746
rect 7484 2378 7512 3674
rect 7576 2514 7604 6054
rect 7668 3534 7696 8622
rect 7840 7948 7892 7954
rect 7840 7890 7892 7896
rect 7748 6860 7800 6866
rect 7748 6802 7800 6808
rect 7760 4282 7788 6802
rect 7852 5896 7880 7890
rect 7944 7886 7972 8774
rect 7932 7880 7984 7886
rect 7932 7822 7984 7828
rect 7944 7342 7972 7822
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 7944 6934 7972 7278
rect 8036 7256 8064 8894
rect 8116 8288 8168 8294
rect 8116 8230 8168 8236
rect 8128 8129 8156 8230
rect 8114 8120 8170 8129
rect 8114 8055 8170 8064
rect 8220 8004 8248 8978
rect 8852 8832 8904 8838
rect 8298 8800 8354 8809
rect 8852 8774 8904 8780
rect 8298 8735 8354 8744
rect 8312 8090 8340 8735
rect 8452 8732 8748 8752
rect 8508 8730 8532 8732
rect 8588 8730 8612 8732
rect 8668 8730 8692 8732
rect 8530 8678 8532 8730
rect 8594 8678 8606 8730
rect 8668 8678 8670 8730
rect 8508 8676 8532 8678
rect 8588 8676 8612 8678
rect 8668 8676 8692 8678
rect 8452 8656 8748 8676
rect 8392 8560 8444 8566
rect 8392 8502 8444 8508
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 8404 8022 8432 8502
rect 8760 8492 8812 8498
rect 8864 8480 8892 8774
rect 8812 8452 8892 8480
rect 8760 8434 8812 8440
rect 8668 8288 8720 8294
rect 8668 8230 8720 8236
rect 8128 7976 8248 8004
rect 8392 8016 8444 8022
rect 8128 7460 8156 7976
rect 8392 7958 8444 7964
rect 8680 7954 8708 8230
rect 8852 8084 8904 8090
rect 8852 8026 8904 8032
rect 8668 7948 8720 7954
rect 8668 7890 8720 7896
rect 8864 7721 8892 8026
rect 8850 7712 8906 7721
rect 8452 7644 8748 7664
rect 8850 7647 8906 7656
rect 8508 7642 8532 7644
rect 8588 7642 8612 7644
rect 8668 7642 8692 7644
rect 8530 7590 8532 7642
rect 8594 7590 8606 7642
rect 8668 7590 8670 7642
rect 8508 7588 8532 7590
rect 8588 7588 8612 7590
rect 8668 7588 8692 7590
rect 8206 7576 8262 7585
rect 8452 7568 8748 7588
rect 8850 7576 8906 7585
rect 8262 7520 8850 7528
rect 8206 7511 8906 7520
rect 8220 7500 8892 7511
rect 8128 7432 8800 7460
rect 8036 7228 8248 7256
rect 8114 7168 8170 7177
rect 8114 7103 8170 7112
rect 7932 6928 7984 6934
rect 7932 6870 7984 6876
rect 8128 6866 8156 7103
rect 8220 6934 8248 7228
rect 8772 7002 8800 7432
rect 8392 6996 8444 7002
rect 8760 6996 8812 7002
rect 8444 6956 8708 6984
rect 8392 6938 8444 6944
rect 8208 6928 8260 6934
rect 8680 6882 8708 6956
rect 8760 6938 8812 6944
rect 8852 6928 8904 6934
rect 8208 6870 8260 6876
rect 8116 6860 8168 6866
rect 8116 6802 8168 6808
rect 8312 6854 8616 6882
rect 8680 6876 8852 6882
rect 8680 6870 8904 6876
rect 8680 6854 8892 6870
rect 8024 6724 8076 6730
rect 8024 6666 8076 6672
rect 8036 6458 8064 6666
rect 8024 6452 8076 6458
rect 8024 6394 8076 6400
rect 8024 6112 8076 6118
rect 7944 6072 8024 6100
rect 7944 5896 7972 6072
rect 8024 6054 8076 6060
rect 7852 5868 7972 5896
rect 7840 5772 7892 5778
rect 7840 5714 7892 5720
rect 7852 5030 7880 5714
rect 7840 5024 7892 5030
rect 7840 4966 7892 4972
rect 7748 4276 7800 4282
rect 7748 4218 7800 4224
rect 7748 3596 7800 3602
rect 7748 3538 7800 3544
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 7668 2689 7696 3470
rect 7760 2938 7788 3538
rect 7852 3058 7880 4966
rect 7944 3618 7972 5868
rect 8024 4820 8076 4826
rect 8024 4762 8076 4768
rect 8036 4282 8064 4762
rect 8128 4457 8156 6802
rect 8208 6792 8260 6798
rect 8312 6780 8340 6854
rect 8260 6752 8340 6780
rect 8588 6780 8616 6854
rect 8852 6792 8904 6798
rect 8588 6752 8852 6780
rect 8208 6734 8260 6740
rect 8852 6734 8904 6740
rect 8208 6656 8260 6662
rect 8312 6633 8892 6644
rect 8208 6598 8260 6604
rect 8298 6624 8906 6633
rect 8220 6361 8248 6598
rect 8354 6616 8850 6624
rect 8298 6559 8354 6568
rect 8452 6556 8748 6576
rect 8850 6559 8906 6568
rect 8508 6554 8532 6556
rect 8588 6554 8612 6556
rect 8668 6554 8692 6556
rect 8530 6502 8532 6554
rect 8594 6502 8606 6554
rect 8668 6502 8670 6554
rect 8508 6500 8532 6502
rect 8588 6500 8612 6502
rect 8668 6500 8692 6502
rect 8452 6480 8748 6500
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 8206 6352 8262 6361
rect 8206 6287 8262 6296
rect 8312 6186 8340 6394
rect 8760 6248 8812 6254
rect 8666 6216 8722 6225
rect 8300 6180 8352 6186
rect 8300 6122 8352 6128
rect 8588 6174 8666 6202
rect 8392 5908 8444 5914
rect 8484 5908 8536 5914
rect 8444 5868 8484 5896
rect 8392 5850 8444 5856
rect 8484 5850 8536 5856
rect 8208 5840 8260 5846
rect 8206 5808 8208 5817
rect 8260 5808 8262 5817
rect 8206 5743 8262 5752
rect 8390 5808 8446 5817
rect 8588 5778 8616 6174
rect 8760 6190 8812 6196
rect 8666 6151 8722 6160
rect 8772 5914 8800 6190
rect 8852 6180 8904 6186
rect 8852 6122 8904 6128
rect 8760 5908 8812 5914
rect 8760 5850 8812 5856
rect 8864 5817 8892 6122
rect 8850 5808 8906 5817
rect 8390 5743 8446 5752
rect 8576 5772 8628 5778
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 8220 5030 8248 5646
rect 8404 5624 8432 5743
rect 8850 5743 8906 5752
rect 8576 5714 8628 5720
rect 8852 5704 8904 5710
rect 8852 5646 8904 5652
rect 8312 5596 8432 5624
rect 8312 5545 8340 5596
rect 8298 5536 8354 5545
rect 8298 5471 8354 5480
rect 8452 5468 8748 5488
rect 8508 5466 8532 5468
rect 8588 5466 8612 5468
rect 8668 5466 8692 5468
rect 8530 5414 8532 5466
rect 8594 5414 8606 5466
rect 8668 5414 8670 5466
rect 8508 5412 8532 5414
rect 8588 5412 8612 5414
rect 8668 5412 8692 5414
rect 8452 5392 8748 5412
rect 8760 5160 8812 5166
rect 8864 5148 8892 5646
rect 8812 5120 8892 5148
rect 8760 5102 8812 5108
rect 8208 5024 8260 5030
rect 8208 4966 8260 4972
rect 8220 4622 8248 4966
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 8114 4448 8170 4457
rect 8114 4383 8170 4392
rect 8024 4276 8076 4282
rect 8024 4218 8076 4224
rect 8312 4214 8340 4626
rect 8852 4480 8904 4486
rect 8852 4422 8904 4428
rect 8452 4380 8748 4400
rect 8508 4378 8532 4380
rect 8588 4378 8612 4380
rect 8668 4378 8692 4380
rect 8530 4326 8532 4378
rect 8594 4326 8606 4378
rect 8668 4326 8670 4378
rect 8508 4324 8532 4326
rect 8588 4324 8612 4326
rect 8668 4324 8692 4326
rect 8452 4304 8748 4324
rect 8300 4208 8352 4214
rect 8128 4168 8300 4196
rect 8022 3904 8078 3913
rect 8022 3839 8078 3848
rect 8036 3738 8064 3839
rect 8024 3732 8076 3738
rect 8024 3674 8076 3680
rect 7944 3590 8064 3618
rect 7932 3528 7984 3534
rect 7932 3470 7984 3476
rect 7944 3097 7972 3470
rect 8036 3194 8064 3590
rect 8128 3534 8156 4168
rect 8300 4150 8352 4156
rect 8484 4140 8536 4146
rect 8484 4082 8536 4088
rect 8496 4010 8524 4082
rect 8760 4072 8812 4078
rect 8760 4014 8812 4020
rect 8484 4004 8536 4010
rect 8484 3946 8536 3952
rect 8392 3732 8444 3738
rect 8312 3692 8392 3720
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8116 3392 8168 3398
rect 8116 3334 8168 3340
rect 8128 3233 8156 3334
rect 8114 3224 8170 3233
rect 8024 3188 8076 3194
rect 8114 3159 8170 3168
rect 8024 3130 8076 3136
rect 7930 3088 7986 3097
rect 7840 3052 7892 3058
rect 7930 3023 7986 3032
rect 8024 3052 8076 3058
rect 7840 2994 7892 3000
rect 8024 2994 8076 3000
rect 8036 2938 8064 2994
rect 8220 2990 8248 3470
rect 8208 2984 8260 2990
rect 7760 2910 8064 2938
rect 8114 2952 8170 2961
rect 8208 2926 8260 2932
rect 8114 2887 8170 2896
rect 7654 2680 7710 2689
rect 7654 2615 7710 2624
rect 7748 2576 7800 2582
rect 7748 2518 7800 2524
rect 7564 2508 7616 2514
rect 7564 2450 7616 2456
rect 7472 2372 7524 2378
rect 7472 2314 7524 2320
rect 7760 2009 7788 2518
rect 8024 2508 8076 2514
rect 7944 2468 8024 2496
rect 7746 2000 7802 2009
rect 7746 1935 7802 1944
rect 7656 1896 7708 1902
rect 7656 1838 7708 1844
rect 7668 800 7696 1838
rect 7944 1562 7972 2468
rect 8024 2450 8076 2456
rect 8128 2378 8156 2887
rect 8206 2544 8262 2553
rect 8206 2479 8262 2488
rect 8116 2372 8168 2378
rect 8116 2314 8168 2320
rect 8128 2281 8156 2314
rect 8114 2272 8170 2281
rect 8114 2207 8170 2216
rect 8220 1970 8248 2479
rect 8208 1964 8260 1970
rect 8208 1906 8260 1912
rect 7932 1556 7984 1562
rect 7932 1498 7984 1504
rect 8024 1556 8076 1562
rect 8024 1498 8076 1504
rect 8036 800 8064 1498
rect 8312 800 8340 3692
rect 8392 3674 8444 3680
rect 8772 3534 8800 4014
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 8452 3292 8748 3312
rect 8508 3290 8532 3292
rect 8588 3290 8612 3292
rect 8668 3290 8692 3292
rect 8530 3238 8532 3290
rect 8594 3238 8606 3290
rect 8668 3238 8670 3290
rect 8508 3236 8532 3238
rect 8588 3236 8612 3238
rect 8668 3236 8692 3238
rect 8452 3216 8748 3236
rect 8484 3120 8536 3126
rect 8760 3120 8812 3126
rect 8536 3080 8760 3108
rect 8484 3062 8536 3068
rect 8760 3062 8812 3068
rect 8864 2922 8892 4422
rect 8956 4026 8984 10134
rect 9140 10062 9168 10610
rect 9128 10056 9180 10062
rect 9128 9998 9180 10004
rect 9036 9920 9088 9926
rect 9036 9862 9088 9868
rect 9048 9450 9076 9862
rect 9140 9761 9168 9998
rect 9126 9752 9182 9761
rect 9126 9687 9182 9696
rect 9128 9512 9180 9518
rect 9128 9454 9180 9460
rect 9036 9444 9088 9450
rect 9036 9386 9088 9392
rect 9140 9353 9168 9454
rect 9126 9344 9182 9353
rect 9126 9279 9182 9288
rect 9140 8974 9168 9279
rect 9036 8968 9088 8974
rect 9036 8910 9088 8916
rect 9128 8968 9180 8974
rect 9128 8910 9180 8916
rect 9048 8022 9076 8910
rect 9232 8673 9260 11104
rect 9312 10736 9364 10742
rect 9310 10704 9312 10713
rect 9364 10704 9366 10713
rect 9310 10639 9366 10648
rect 9324 9926 9352 10639
rect 9416 10266 9444 11494
rect 9496 11348 9548 11354
rect 9496 11290 9548 11296
rect 9508 11121 9536 11290
rect 9600 11218 9628 13398
rect 9772 13388 9824 13394
rect 9772 13330 9824 13336
rect 9784 13297 9812 13330
rect 9770 13288 9826 13297
rect 9770 13223 9826 13232
rect 9864 13252 9916 13258
rect 9864 13194 9916 13200
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 9692 12782 9720 12922
rect 9876 12889 9904 13194
rect 9862 12880 9918 12889
rect 9862 12815 9918 12824
rect 9680 12776 9732 12782
rect 9680 12718 9732 12724
rect 9772 12776 9824 12782
rect 9772 12718 9824 12724
rect 9862 12744 9918 12753
rect 9692 11762 9720 12718
rect 9680 11756 9732 11762
rect 9680 11698 9732 11704
rect 9784 11234 9812 12718
rect 9862 12679 9864 12688
rect 9916 12679 9918 12688
rect 9864 12650 9916 12656
rect 9862 12336 9918 12345
rect 9968 12306 9996 14350
rect 10060 14278 10088 15030
rect 10048 14272 10100 14278
rect 10048 14214 10100 14220
rect 10048 13184 10100 13190
rect 10048 13126 10100 13132
rect 10060 12986 10088 13126
rect 10048 12980 10100 12986
rect 10048 12922 10100 12928
rect 9862 12271 9918 12280
rect 9956 12300 10008 12306
rect 9588 11212 9640 11218
rect 9588 11154 9640 11160
rect 9692 11206 9812 11234
rect 9494 11112 9550 11121
rect 9494 11047 9550 11056
rect 9496 11008 9548 11014
rect 9496 10950 9548 10956
rect 9588 11008 9640 11014
rect 9588 10950 9640 10956
rect 9508 10810 9536 10950
rect 9496 10804 9548 10810
rect 9496 10746 9548 10752
rect 9600 10606 9628 10950
rect 9692 10674 9720 11206
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 9784 11014 9812 11086
rect 9772 11008 9824 11014
rect 9772 10950 9824 10956
rect 9770 10840 9826 10849
rect 9770 10775 9826 10784
rect 9784 10742 9812 10775
rect 9772 10736 9824 10742
rect 9772 10678 9824 10684
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 9588 10600 9640 10606
rect 9588 10542 9640 10548
rect 9404 10260 9456 10266
rect 9404 10202 9456 10208
rect 9402 10160 9458 10169
rect 9402 10095 9458 10104
rect 9312 9920 9364 9926
rect 9312 9862 9364 9868
rect 9416 9654 9444 10095
rect 9692 9926 9720 10610
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9404 9648 9456 9654
rect 9404 9590 9456 9596
rect 9312 9444 9364 9450
rect 9312 9386 9364 9392
rect 9588 9444 9640 9450
rect 9588 9386 9640 9392
rect 9772 9444 9824 9450
rect 9772 9386 9824 9392
rect 9324 9110 9352 9386
rect 9494 9208 9550 9217
rect 9494 9143 9550 9152
rect 9508 9110 9536 9143
rect 9312 9104 9364 9110
rect 9312 9046 9364 9052
rect 9496 9104 9548 9110
rect 9496 9046 9548 9052
rect 9496 8832 9548 8838
rect 9600 8820 9628 9386
rect 9678 9344 9734 9353
rect 9678 9279 9734 9288
rect 9548 8792 9628 8820
rect 9496 8774 9548 8780
rect 9218 8664 9274 8673
rect 9218 8599 9274 8608
rect 9692 8514 9720 9279
rect 9784 9178 9812 9386
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9692 8498 9812 8514
rect 9692 8492 9824 8498
rect 9692 8486 9772 8492
rect 9772 8434 9824 8440
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 9312 8356 9364 8362
rect 9312 8298 9364 8304
rect 9036 8016 9088 8022
rect 9036 7958 9088 7964
rect 9324 7290 9352 8298
rect 9404 8084 9456 8090
rect 9404 8026 9456 8032
rect 9416 7410 9444 8026
rect 9404 7404 9456 7410
rect 9404 7346 9456 7352
rect 9324 7262 9444 7290
rect 9692 7274 9720 8366
rect 9220 7200 9272 7206
rect 9220 7142 9272 7148
rect 9312 7200 9364 7206
rect 9312 7142 9364 7148
rect 9036 6724 9088 6730
rect 9036 6666 9088 6672
rect 9048 5166 9076 6666
rect 9232 6644 9260 7142
rect 9324 6934 9352 7142
rect 9312 6928 9364 6934
rect 9312 6870 9364 6876
rect 9416 6798 9444 7262
rect 9680 7268 9732 7274
rect 9680 7210 9732 7216
rect 9876 6866 9904 12271
rect 9956 12242 10008 12248
rect 10046 12200 10102 12209
rect 10046 12135 10102 12144
rect 9954 11384 10010 11393
rect 9954 11319 10010 11328
rect 9968 11286 9996 11319
rect 9956 11280 10008 11286
rect 9956 11222 10008 11228
rect 9956 11008 10008 11014
rect 9956 10950 10008 10956
rect 9968 10266 9996 10950
rect 9956 10260 10008 10266
rect 9956 10202 10008 10208
rect 10060 10146 10088 12135
rect 9968 10118 10088 10146
rect 10152 10146 10180 15506
rect 10244 14346 10272 16934
rect 10520 15910 10548 16934
rect 10612 16794 10640 17070
rect 10704 16794 10732 17070
rect 10784 16992 10836 16998
rect 10784 16934 10836 16940
rect 10600 16788 10652 16794
rect 10600 16730 10652 16736
rect 10692 16788 10744 16794
rect 10692 16730 10744 16736
rect 10508 15904 10560 15910
rect 10508 15846 10560 15852
rect 10322 15464 10378 15473
rect 10322 15399 10378 15408
rect 10232 14340 10284 14346
rect 10232 14282 10284 14288
rect 10232 13524 10284 13530
rect 10232 13466 10284 13472
rect 10244 11830 10272 13466
rect 10336 12594 10364 15399
rect 10520 14550 10548 15846
rect 10692 15360 10744 15366
rect 10692 15302 10744 15308
rect 10508 14544 10560 14550
rect 10508 14486 10560 14492
rect 10508 14272 10560 14278
rect 10508 14214 10560 14220
rect 10520 13920 10548 14214
rect 10520 13892 10640 13920
rect 10414 13832 10470 13841
rect 10414 13767 10470 13776
rect 10428 13734 10456 13767
rect 10416 13728 10468 13734
rect 10416 13670 10468 13676
rect 10508 13728 10560 13734
rect 10508 13670 10560 13676
rect 10520 13546 10548 13670
rect 10428 13518 10548 13546
rect 10428 12782 10456 13518
rect 10508 13252 10560 13258
rect 10508 13194 10560 13200
rect 10416 12776 10468 12782
rect 10416 12718 10468 12724
rect 10336 12566 10456 12594
rect 10232 11824 10284 11830
rect 10232 11766 10284 11772
rect 10232 11552 10284 11558
rect 10232 11494 10284 11500
rect 10244 10674 10272 11494
rect 10324 11076 10376 11082
rect 10324 11018 10376 11024
rect 10232 10668 10284 10674
rect 10232 10610 10284 10616
rect 10336 10554 10364 11018
rect 10428 10985 10456 12566
rect 10414 10976 10470 10985
rect 10414 10911 10470 10920
rect 10428 10606 10456 10911
rect 10244 10526 10364 10554
rect 10416 10600 10468 10606
rect 10416 10542 10468 10548
rect 10244 10266 10272 10526
rect 10324 10464 10376 10470
rect 10324 10406 10376 10412
rect 10414 10432 10470 10441
rect 10232 10260 10284 10266
rect 10232 10202 10284 10208
rect 10152 10118 10272 10146
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 9404 6792 9456 6798
rect 9404 6734 9456 6740
rect 9770 6760 9826 6769
rect 9680 6724 9732 6730
rect 9770 6695 9826 6704
rect 9680 6666 9732 6672
rect 9232 6616 9444 6644
rect 9416 6390 9444 6616
rect 9494 6624 9550 6633
rect 9692 6610 9720 6666
rect 9550 6582 9720 6610
rect 9494 6559 9550 6568
rect 9404 6384 9456 6390
rect 9404 6326 9456 6332
rect 9220 6248 9272 6254
rect 9140 6208 9220 6236
rect 9140 5778 9168 6208
rect 9784 6225 9812 6695
rect 9220 6190 9272 6196
rect 9770 6216 9826 6225
rect 9680 6180 9732 6186
rect 9770 6151 9826 6160
rect 9680 6122 9732 6128
rect 9220 5840 9272 5846
rect 9496 5840 9548 5846
rect 9272 5800 9496 5828
rect 9220 5782 9272 5788
rect 9496 5782 9548 5788
rect 9128 5772 9180 5778
rect 9128 5714 9180 5720
rect 9036 5160 9088 5166
rect 9036 5102 9088 5108
rect 9140 5148 9168 5714
rect 9404 5568 9456 5574
rect 9404 5510 9456 5516
rect 9416 5302 9444 5510
rect 9494 5400 9550 5409
rect 9494 5335 9496 5344
rect 9548 5335 9550 5344
rect 9496 5306 9548 5312
rect 9404 5296 9456 5302
rect 9310 5264 9366 5273
rect 9404 5238 9456 5244
rect 9494 5264 9550 5273
rect 9310 5199 9366 5208
rect 9494 5199 9496 5208
rect 9220 5160 9272 5166
rect 9140 5120 9220 5148
rect 9048 4486 9076 5102
rect 9140 5030 9168 5120
rect 9220 5102 9272 5108
rect 9128 5024 9180 5030
rect 9128 4966 9180 4972
rect 9324 4865 9352 5199
rect 9548 5199 9550 5208
rect 9496 5170 9548 5176
rect 9404 5160 9456 5166
rect 9404 5102 9456 5108
rect 9310 4856 9366 4865
rect 9128 4820 9180 4826
rect 9310 4791 9366 4800
rect 9128 4762 9180 4768
rect 9140 4593 9168 4762
rect 9312 4616 9364 4622
rect 9126 4584 9182 4593
rect 9312 4558 9364 4564
rect 9126 4519 9182 4528
rect 9036 4480 9088 4486
rect 9324 4457 9352 4558
rect 9036 4422 9088 4428
rect 9310 4448 9366 4457
rect 9048 4146 9076 4422
rect 9310 4383 9366 4392
rect 9126 4312 9182 4321
rect 9126 4247 9128 4256
rect 9180 4247 9182 4256
rect 9128 4218 9180 4224
rect 9416 4154 9444 5102
rect 9508 4826 9536 5170
rect 9588 5024 9640 5030
rect 9588 4966 9640 4972
rect 9496 4820 9548 4826
rect 9496 4762 9548 4768
rect 9600 4706 9628 4966
rect 9508 4678 9628 4706
rect 9508 4554 9536 4678
rect 9496 4548 9548 4554
rect 9496 4490 9548 4496
rect 9588 4548 9640 4554
rect 9588 4490 9640 4496
rect 9600 4214 9628 4490
rect 9588 4208 9640 4214
rect 9036 4140 9088 4146
rect 9036 4082 9088 4088
rect 9324 4126 9444 4154
rect 9494 4176 9550 4185
rect 8956 4010 9076 4026
rect 8956 4004 9088 4010
rect 8956 3998 9036 4004
rect 9036 3946 9088 3952
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 8956 3058 8984 3878
rect 9048 3058 9076 3946
rect 9220 3528 9272 3534
rect 9220 3470 9272 3476
rect 9128 3392 9180 3398
rect 9128 3334 9180 3340
rect 8944 3052 8996 3058
rect 8944 2994 8996 3000
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 8852 2916 8904 2922
rect 8852 2858 8904 2864
rect 8944 2916 8996 2922
rect 8944 2858 8996 2864
rect 8668 2848 8720 2854
rect 8666 2816 8668 2825
rect 8720 2816 8722 2825
rect 8666 2751 8722 2760
rect 8680 2650 8708 2751
rect 8668 2644 8720 2650
rect 8668 2586 8720 2592
rect 8864 2514 8892 2858
rect 8852 2508 8904 2514
rect 8852 2450 8904 2456
rect 8452 2204 8748 2224
rect 8508 2202 8532 2204
rect 8588 2202 8612 2204
rect 8668 2202 8692 2204
rect 8530 2150 8532 2202
rect 8594 2150 8606 2202
rect 8668 2150 8670 2202
rect 8508 2148 8532 2150
rect 8588 2148 8612 2150
rect 8668 2148 8692 2150
rect 8452 2128 8748 2148
rect 8956 1952 8984 2858
rect 9036 2848 9088 2854
rect 9036 2790 9088 2796
rect 8680 1924 8984 1952
rect 8680 800 8708 1924
rect 9048 800 9076 2790
rect 9140 2582 9168 3334
rect 9232 2582 9260 3470
rect 9324 3194 9352 4126
rect 9588 4150 9640 4156
rect 9494 4111 9550 4120
rect 9404 4072 9456 4078
rect 9404 4014 9456 4020
rect 9416 3942 9444 4014
rect 9508 3942 9536 4111
rect 9692 4026 9720 6122
rect 9772 5908 9824 5914
rect 9772 5850 9824 5856
rect 9784 5778 9812 5850
rect 9772 5772 9824 5778
rect 9772 5714 9824 5720
rect 9968 5658 9996 10118
rect 10140 10056 10192 10062
rect 10140 9998 10192 10004
rect 10048 9920 10100 9926
rect 10048 9862 10100 9868
rect 10060 7274 10088 9862
rect 10152 8809 10180 9998
rect 10138 8800 10194 8809
rect 10138 8735 10194 8744
rect 10048 7268 10100 7274
rect 10048 7210 10100 7216
rect 10060 7177 10088 7210
rect 10046 7168 10102 7177
rect 10046 7103 10102 7112
rect 10048 6928 10100 6934
rect 10048 6870 10100 6876
rect 10060 6633 10088 6870
rect 10046 6624 10102 6633
rect 10046 6559 10102 6568
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 10060 6225 10088 6394
rect 10046 6216 10102 6225
rect 10046 6151 10102 6160
rect 9784 5630 9996 5658
rect 9784 4826 9812 5630
rect 9864 5568 9916 5574
rect 9916 5528 9996 5556
rect 9864 5510 9916 5516
rect 9772 4820 9824 4826
rect 9772 4762 9824 4768
rect 9864 4820 9916 4826
rect 9864 4762 9916 4768
rect 9784 4457 9812 4762
rect 9770 4448 9826 4457
rect 9770 4383 9826 4392
rect 9772 4208 9824 4214
rect 9772 4150 9824 4156
rect 9600 3998 9720 4026
rect 9404 3936 9456 3942
rect 9404 3878 9456 3884
rect 9496 3936 9548 3942
rect 9496 3878 9548 3884
rect 9404 3596 9456 3602
rect 9404 3538 9456 3544
rect 9496 3596 9548 3602
rect 9600 3584 9628 3998
rect 9680 3664 9732 3670
rect 9680 3606 9732 3612
rect 9548 3556 9628 3584
rect 9496 3538 9548 3544
rect 9416 3194 9444 3538
rect 9508 3233 9536 3538
rect 9586 3360 9642 3369
rect 9586 3295 9642 3304
rect 9494 3224 9550 3233
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 9404 3188 9456 3194
rect 9494 3159 9550 3168
rect 9404 3130 9456 3136
rect 9600 2650 9628 3295
rect 9692 3126 9720 3606
rect 9784 3534 9812 4150
rect 9876 3602 9904 4762
rect 9968 4146 9996 5528
rect 10046 5400 10102 5409
rect 10046 5335 10048 5344
rect 10100 5335 10102 5344
rect 10048 5306 10100 5312
rect 10152 5250 10180 8735
rect 10244 8673 10272 10118
rect 10230 8664 10286 8673
rect 10230 8599 10286 8608
rect 10244 6186 10272 8599
rect 10336 8265 10364 10406
rect 10414 10367 10470 10376
rect 10428 10130 10456 10367
rect 10416 10124 10468 10130
rect 10416 10066 10468 10072
rect 10520 9994 10548 13194
rect 10612 12918 10640 13892
rect 10704 13025 10732 15302
rect 10796 13530 10824 16934
rect 10950 16892 11246 16912
rect 11006 16890 11030 16892
rect 11086 16890 11110 16892
rect 11166 16890 11190 16892
rect 11028 16838 11030 16890
rect 11092 16838 11104 16890
rect 11166 16838 11168 16890
rect 11006 16836 11030 16838
rect 11086 16836 11110 16838
rect 11166 16836 11190 16838
rect 10950 16816 11246 16836
rect 11348 16794 11376 17070
rect 11808 16794 11836 17070
rect 11888 16992 11940 16998
rect 12072 16992 12124 16998
rect 11940 16952 12020 16980
rect 11888 16934 11940 16940
rect 11336 16788 11388 16794
rect 11336 16730 11388 16736
rect 11796 16788 11848 16794
rect 11796 16730 11848 16736
rect 11520 16040 11572 16046
rect 11520 15982 11572 15988
rect 10950 15804 11246 15824
rect 11006 15802 11030 15804
rect 11086 15802 11110 15804
rect 11166 15802 11190 15804
rect 11028 15750 11030 15802
rect 11092 15750 11104 15802
rect 11166 15750 11168 15802
rect 11006 15748 11030 15750
rect 11086 15748 11110 15750
rect 11166 15748 11190 15750
rect 10950 15728 11246 15748
rect 11428 15632 11480 15638
rect 11428 15574 11480 15580
rect 10950 14716 11246 14736
rect 11006 14714 11030 14716
rect 11086 14714 11110 14716
rect 11166 14714 11190 14716
rect 11028 14662 11030 14714
rect 11092 14662 11104 14714
rect 11166 14662 11168 14714
rect 11006 14660 11030 14662
rect 11086 14660 11110 14662
rect 11166 14660 11190 14662
rect 10950 14640 11246 14660
rect 10876 14340 10928 14346
rect 10876 14282 10928 14288
rect 10784 13524 10836 13530
rect 10784 13466 10836 13472
rect 10888 13410 10916 14282
rect 11336 14068 11388 14074
rect 11336 14010 11388 14016
rect 10950 13628 11246 13648
rect 11006 13626 11030 13628
rect 11086 13626 11110 13628
rect 11166 13626 11190 13628
rect 11028 13574 11030 13626
rect 11092 13574 11104 13626
rect 11166 13574 11168 13626
rect 11006 13572 11030 13574
rect 11086 13572 11110 13574
rect 11166 13572 11190 13574
rect 10950 13552 11246 13572
rect 11348 13512 11376 14010
rect 11256 13484 11376 13512
rect 10796 13382 10916 13410
rect 11060 13456 11112 13462
rect 11256 13410 11284 13484
rect 11112 13404 11284 13410
rect 11060 13398 11284 13404
rect 11072 13382 11284 13398
rect 11336 13388 11388 13394
rect 10690 13016 10746 13025
rect 10690 12951 10746 12960
rect 10600 12912 10652 12918
rect 10600 12854 10652 12860
rect 10796 12646 10824 13382
rect 11164 13190 11192 13382
rect 11336 13330 11388 13336
rect 11152 13184 11204 13190
rect 11150 13152 11152 13161
rect 11244 13184 11296 13190
rect 11204 13152 11206 13161
rect 11244 13126 11296 13132
rect 11150 13087 11206 13096
rect 10874 12880 10930 12889
rect 10874 12815 10876 12824
rect 10928 12815 10930 12824
rect 10876 12786 10928 12792
rect 10600 12640 10652 12646
rect 10598 12608 10600 12617
rect 10784 12640 10836 12646
rect 10652 12608 10654 12617
rect 10784 12582 10836 12588
rect 10598 12543 10654 12552
rect 10690 12472 10746 12481
rect 10690 12407 10692 12416
rect 10744 12407 10746 12416
rect 10692 12378 10744 12384
rect 10690 11928 10746 11937
rect 10690 11863 10746 11872
rect 10600 11756 10652 11762
rect 10600 11698 10652 11704
rect 10612 11150 10640 11698
rect 10704 11558 10732 11863
rect 10692 11552 10744 11558
rect 10690 11520 10692 11529
rect 10744 11520 10746 11529
rect 10690 11455 10746 11464
rect 10690 11384 10746 11393
rect 10796 11354 10824 12582
rect 10888 12424 10916 12786
rect 11256 12714 11284 13126
rect 11244 12708 11296 12714
rect 11244 12650 11296 12656
rect 10950 12540 11246 12560
rect 11006 12538 11030 12540
rect 11086 12538 11110 12540
rect 11166 12538 11190 12540
rect 11028 12486 11030 12538
rect 11092 12486 11104 12538
rect 11166 12486 11168 12538
rect 11006 12484 11030 12486
rect 11086 12484 11110 12486
rect 11166 12484 11190 12486
rect 10950 12464 11246 12484
rect 10888 12396 11008 12424
rect 10980 12238 11008 12396
rect 10968 12232 11020 12238
rect 10968 12174 11020 12180
rect 11244 12096 11296 12102
rect 11058 12064 11114 12073
rect 11244 12038 11296 12044
rect 11058 11999 11114 12008
rect 11072 11694 11100 11999
rect 11256 11762 11284 12038
rect 11348 11898 11376 13330
rect 11440 13190 11468 15574
rect 11428 13184 11480 13190
rect 11428 13126 11480 13132
rect 11428 12980 11480 12986
rect 11532 12968 11560 15982
rect 11796 15496 11848 15502
rect 11796 15438 11848 15444
rect 11704 13796 11756 13802
rect 11704 13738 11756 13744
rect 11612 13524 11664 13530
rect 11612 13466 11664 13472
rect 11624 13258 11652 13466
rect 11612 13252 11664 13258
rect 11612 13194 11664 13200
rect 11480 12940 11560 12968
rect 11428 12922 11480 12928
rect 11440 12442 11468 12922
rect 11624 12850 11652 13194
rect 11612 12844 11664 12850
rect 11612 12786 11664 12792
rect 11520 12708 11572 12714
rect 11520 12650 11572 12656
rect 11428 12436 11480 12442
rect 11428 12378 11480 12384
rect 11440 12209 11468 12378
rect 11426 12200 11482 12209
rect 11426 12135 11482 12144
rect 11428 12096 11480 12102
rect 11428 12038 11480 12044
rect 11336 11892 11388 11898
rect 11336 11834 11388 11840
rect 11244 11756 11296 11762
rect 11244 11698 11296 11704
rect 11060 11688 11112 11694
rect 11060 11630 11112 11636
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10690 11319 10746 11328
rect 10784 11348 10836 11354
rect 10704 11286 10732 11319
rect 10784 11290 10836 11296
rect 10888 11286 10916 11494
rect 10950 11452 11246 11472
rect 11006 11450 11030 11452
rect 11086 11450 11110 11452
rect 11166 11450 11190 11452
rect 11028 11398 11030 11450
rect 11092 11398 11104 11450
rect 11166 11398 11168 11450
rect 11006 11396 11030 11398
rect 11086 11396 11110 11398
rect 11166 11396 11190 11398
rect 10950 11376 11246 11396
rect 10692 11280 10744 11286
rect 10692 11222 10744 11228
rect 10876 11280 10928 11286
rect 10876 11222 10928 11228
rect 10968 11280 11020 11286
rect 10968 11222 11020 11228
rect 10600 11144 10652 11150
rect 10600 11086 10652 11092
rect 10876 11144 10928 11150
rect 10876 11086 10928 11092
rect 10784 11008 10836 11014
rect 10784 10950 10836 10956
rect 10692 10804 10744 10810
rect 10692 10746 10744 10752
rect 10600 10736 10652 10742
rect 10600 10678 10652 10684
rect 10508 9988 10560 9994
rect 10508 9930 10560 9936
rect 10612 9926 10640 10678
rect 10600 9920 10652 9926
rect 10600 9862 10652 9868
rect 10508 9648 10560 9654
rect 10508 9590 10560 9596
rect 10520 9353 10548 9590
rect 10506 9344 10562 9353
rect 10506 9279 10562 9288
rect 10506 9208 10562 9217
rect 10506 9143 10562 9152
rect 10520 9042 10548 9143
rect 10508 9036 10560 9042
rect 10508 8978 10560 8984
rect 10612 8974 10640 9862
rect 10704 9217 10732 10746
rect 10796 10198 10824 10950
rect 10888 10674 10916 11086
rect 10876 10668 10928 10674
rect 10876 10610 10928 10616
rect 10888 10577 10916 10610
rect 10874 10568 10930 10577
rect 10874 10503 10930 10512
rect 10980 10452 11008 11222
rect 11060 11212 11112 11218
rect 11060 11154 11112 11160
rect 11072 10810 11100 11154
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 11244 10736 11296 10742
rect 11244 10678 11296 10684
rect 11256 10577 11284 10678
rect 11242 10568 11298 10577
rect 11242 10503 11298 10512
rect 10888 10424 11008 10452
rect 10784 10192 10836 10198
rect 10784 10134 10836 10140
rect 10782 9888 10838 9897
rect 10782 9823 10838 9832
rect 10690 9208 10746 9217
rect 10796 9178 10824 9823
rect 10690 9143 10746 9152
rect 10784 9172 10836 9178
rect 10784 9114 10836 9120
rect 10888 9024 10916 10424
rect 10950 10364 11246 10384
rect 11006 10362 11030 10364
rect 11086 10362 11110 10364
rect 11166 10362 11190 10364
rect 11028 10310 11030 10362
rect 11092 10310 11104 10362
rect 11166 10310 11168 10362
rect 11006 10308 11030 10310
rect 11086 10308 11110 10310
rect 11166 10308 11190 10310
rect 10950 10288 11246 10308
rect 11060 10124 11112 10130
rect 11060 10066 11112 10072
rect 11072 9926 11100 10066
rect 11244 9988 11296 9994
rect 11244 9930 11296 9936
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 11152 9920 11204 9926
rect 11152 9862 11204 9868
rect 11164 9518 11192 9862
rect 11256 9722 11284 9930
rect 11244 9716 11296 9722
rect 11244 9658 11296 9664
rect 11348 9518 11376 11834
rect 11440 11801 11468 12038
rect 11426 11792 11482 11801
rect 11426 11727 11482 11736
rect 11428 11688 11480 11694
rect 11428 11630 11480 11636
rect 11440 10810 11468 11630
rect 11532 11393 11560 12650
rect 11716 11898 11744 13738
rect 11808 12442 11836 15438
rect 11992 12889 12020 16952
rect 12072 16934 12124 16940
rect 11978 12880 12034 12889
rect 11978 12815 12034 12824
rect 11980 12708 12032 12714
rect 12084 12696 12112 16934
rect 12176 16726 12204 19200
rect 12164 16720 12216 16726
rect 12164 16662 12216 16668
rect 12544 16658 12572 19200
rect 12912 17202 12940 19200
rect 12900 17196 12952 17202
rect 12900 17138 12952 17144
rect 12808 17060 12860 17066
rect 12808 17002 12860 17008
rect 12624 16992 12676 16998
rect 12624 16934 12676 16940
rect 12532 16652 12584 16658
rect 12532 16594 12584 16600
rect 12164 16516 12216 16522
rect 12164 16458 12216 16464
rect 12176 12782 12204 16458
rect 12256 14952 12308 14958
rect 12256 14894 12308 14900
rect 12268 12782 12296 14894
rect 12348 13932 12400 13938
rect 12348 13874 12400 13880
rect 12360 13326 12388 13874
rect 12348 13320 12400 13326
rect 12348 13262 12400 13268
rect 12164 12776 12216 12782
rect 12256 12776 12308 12782
rect 12164 12718 12216 12724
rect 12254 12744 12256 12753
rect 12308 12744 12310 12753
rect 12032 12668 12112 12696
rect 12254 12679 12310 12688
rect 11980 12650 12032 12656
rect 11796 12436 11848 12442
rect 11848 12396 11928 12424
rect 11796 12378 11848 12384
rect 11796 12232 11848 12238
rect 11796 12174 11848 12180
rect 11808 12102 11836 12174
rect 11796 12096 11848 12102
rect 11796 12038 11848 12044
rect 11900 11914 11928 12396
rect 11704 11892 11756 11898
rect 11704 11834 11756 11840
rect 11808 11886 11928 11914
rect 11612 11756 11664 11762
rect 11612 11698 11664 11704
rect 11518 11384 11574 11393
rect 11518 11319 11520 11328
rect 11572 11319 11574 11328
rect 11520 11290 11572 11296
rect 11532 11259 11560 11290
rect 11520 11144 11572 11150
rect 11624 11121 11652 11698
rect 11704 11552 11756 11558
rect 11704 11494 11756 11500
rect 11520 11086 11572 11092
rect 11610 11112 11666 11121
rect 11428 10804 11480 10810
rect 11428 10746 11480 10752
rect 11532 10713 11560 11086
rect 11610 11047 11666 11056
rect 11612 11008 11664 11014
rect 11612 10950 11664 10956
rect 11518 10704 11574 10713
rect 11624 10674 11652 10950
rect 11518 10639 11574 10648
rect 11612 10668 11664 10674
rect 11426 9888 11482 9897
rect 11426 9823 11482 9832
rect 11152 9512 11204 9518
rect 11152 9454 11204 9460
rect 11336 9512 11388 9518
rect 11336 9454 11388 9460
rect 10968 9444 11020 9450
rect 11020 9404 11100 9432
rect 10968 9386 11020 9392
rect 11072 9364 11100 9404
rect 11072 9353 11376 9364
rect 11072 9344 11390 9353
rect 11072 9336 11334 9344
rect 10950 9276 11246 9296
rect 11334 9279 11390 9288
rect 11006 9274 11030 9276
rect 11086 9274 11110 9276
rect 11166 9274 11190 9276
rect 11028 9222 11030 9274
rect 11092 9222 11104 9274
rect 11166 9222 11168 9274
rect 11006 9220 11030 9222
rect 11086 9220 11110 9222
rect 11166 9220 11190 9222
rect 10950 9200 11246 9220
rect 11336 9172 11388 9178
rect 11440 9160 11468 9823
rect 11388 9132 11468 9160
rect 11336 9114 11388 9120
rect 11060 9104 11112 9110
rect 11244 9104 11296 9110
rect 11112 9064 11244 9092
rect 11060 9046 11112 9052
rect 11244 9046 11296 9052
rect 10968 9036 11020 9042
rect 10888 8996 10968 9024
rect 10968 8978 11020 8984
rect 10600 8968 10652 8974
rect 10600 8910 10652 8916
rect 10508 8628 10560 8634
rect 10508 8570 10560 8576
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 10416 8356 10468 8362
rect 10416 8298 10468 8304
rect 10322 8256 10378 8265
rect 10322 8191 10378 8200
rect 10428 7478 10456 8298
rect 10520 7886 10548 8570
rect 10612 8090 10640 8570
rect 10980 8378 11008 8978
rect 11532 8974 11560 10639
rect 11612 10610 11664 10616
rect 11624 9722 11652 10610
rect 11716 9722 11744 11494
rect 11612 9716 11664 9722
rect 11612 9658 11664 9664
rect 11704 9716 11756 9722
rect 11704 9658 11756 9664
rect 11702 9616 11758 9625
rect 11702 9551 11758 9560
rect 11716 9217 11744 9551
rect 11702 9208 11758 9217
rect 11702 9143 11758 9152
rect 11704 9036 11756 9042
rect 11704 8978 11756 8984
rect 11336 8968 11388 8974
rect 11336 8910 11388 8916
rect 11520 8968 11572 8974
rect 11520 8910 11572 8916
rect 11348 8634 11376 8910
rect 11716 8786 11744 8978
rect 11532 8758 11744 8786
rect 11532 8673 11560 8758
rect 11518 8664 11574 8673
rect 11336 8628 11388 8634
rect 11518 8599 11574 8608
rect 11336 8570 11388 8576
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 10980 8362 11192 8378
rect 10876 8356 10928 8362
rect 10980 8356 11204 8362
rect 10980 8350 11152 8356
rect 10876 8298 10928 8304
rect 11152 8298 11204 8304
rect 10782 8256 10838 8265
rect 10782 8191 10838 8200
rect 10600 8084 10652 8090
rect 10600 8026 10652 8032
rect 10796 7886 10824 8191
rect 10508 7880 10560 7886
rect 10508 7822 10560 7828
rect 10784 7880 10836 7886
rect 10784 7822 10836 7828
rect 10888 7818 10916 8298
rect 11256 8276 11284 8434
rect 11704 8356 11756 8362
rect 11704 8298 11756 8304
rect 11256 8248 11560 8276
rect 10950 8188 11246 8208
rect 11006 8186 11030 8188
rect 11086 8186 11110 8188
rect 11166 8186 11190 8188
rect 11028 8134 11030 8186
rect 11092 8134 11104 8186
rect 11166 8134 11168 8186
rect 11006 8132 11030 8134
rect 11086 8132 11110 8134
rect 11166 8132 11190 8134
rect 10950 8112 11246 8132
rect 10968 8016 11020 8022
rect 11020 7976 11100 8004
rect 10968 7958 11020 7964
rect 10876 7812 10928 7818
rect 10876 7754 10928 7760
rect 10600 7744 10652 7750
rect 10600 7686 10652 7692
rect 10784 7744 10836 7750
rect 11072 7721 11100 7976
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 11242 7848 11298 7857
rect 10784 7686 10836 7692
rect 10874 7712 10930 7721
rect 10612 7546 10640 7686
rect 10600 7540 10652 7546
rect 10600 7482 10652 7488
rect 10416 7472 10468 7478
rect 10416 7414 10468 7420
rect 10508 7404 10560 7410
rect 10508 7346 10560 7352
rect 10324 7200 10376 7206
rect 10520 7188 10548 7346
rect 10796 7342 10824 7686
rect 10874 7647 10930 7656
rect 11058 7712 11114 7721
rect 11058 7647 11114 7656
rect 10888 7546 10916 7647
rect 10876 7540 10928 7546
rect 10876 7482 10928 7488
rect 10968 7404 11020 7410
rect 11164 7392 11192 7822
rect 11298 7806 11468 7834
rect 11242 7783 11298 7792
rect 11440 7750 11468 7806
rect 11244 7744 11296 7750
rect 11244 7686 11296 7692
rect 11428 7744 11480 7750
rect 11428 7686 11480 7692
rect 11256 7478 11284 7686
rect 11532 7562 11560 8248
rect 11440 7534 11560 7562
rect 11244 7472 11296 7478
rect 11244 7414 11296 7420
rect 11020 7364 11192 7392
rect 10968 7346 11020 7352
rect 10784 7336 10836 7342
rect 10784 7278 10836 7284
rect 10876 7336 10928 7342
rect 10876 7278 10928 7284
rect 11336 7336 11388 7342
rect 11336 7278 11388 7284
rect 10376 7160 10548 7188
rect 10598 7168 10654 7177
rect 10324 7142 10376 7148
rect 10336 6440 10364 7142
rect 10598 7103 10654 7112
rect 10416 6860 10468 6866
rect 10416 6802 10468 6808
rect 10508 6860 10560 6866
rect 10508 6802 10560 6808
rect 10428 6662 10456 6802
rect 10416 6656 10468 6662
rect 10416 6598 10468 6604
rect 10416 6452 10468 6458
rect 10336 6412 10416 6440
rect 10336 6186 10364 6412
rect 10416 6394 10468 6400
rect 10232 6180 10284 6186
rect 10232 6122 10284 6128
rect 10324 6180 10376 6186
rect 10324 6122 10376 6128
rect 10520 6066 10548 6802
rect 10244 6038 10548 6066
rect 10244 5273 10272 6038
rect 10322 5808 10378 5817
rect 10322 5743 10378 5752
rect 10336 5409 10364 5743
rect 10322 5400 10378 5409
rect 10428 5370 10456 6038
rect 10506 5808 10562 5817
rect 10506 5743 10562 5752
rect 10520 5710 10548 5743
rect 10508 5704 10560 5710
rect 10508 5646 10560 5652
rect 10322 5335 10378 5344
rect 10416 5364 10468 5370
rect 10060 5222 10180 5250
rect 10230 5264 10286 5273
rect 10060 4826 10088 5222
rect 10230 5199 10286 5208
rect 10336 5114 10364 5335
rect 10416 5306 10468 5312
rect 10506 5264 10562 5273
rect 10506 5199 10562 5208
rect 10520 5166 10548 5199
rect 10244 5086 10364 5114
rect 10508 5160 10560 5166
rect 10508 5102 10560 5108
rect 10416 5092 10468 5098
rect 10138 4856 10194 4865
rect 10048 4820 10100 4826
rect 10138 4791 10194 4800
rect 10048 4762 10100 4768
rect 10152 4706 10180 4791
rect 10060 4678 10180 4706
rect 9956 4140 10008 4146
rect 9956 4082 10008 4088
rect 10060 3777 10088 4678
rect 10140 4480 10192 4486
rect 10138 4448 10140 4457
rect 10192 4448 10194 4457
rect 10244 4434 10272 5086
rect 10416 5034 10468 5040
rect 10324 4548 10376 4554
rect 10324 4490 10376 4496
rect 10244 4406 10281 4434
rect 10138 4383 10194 4392
rect 10253 4298 10281 4406
rect 10152 4270 10281 4298
rect 10152 4146 10180 4270
rect 10232 4208 10284 4214
rect 10232 4150 10284 4156
rect 10140 4140 10192 4146
rect 10140 4082 10192 4088
rect 10244 4026 10272 4150
rect 10152 3998 10272 4026
rect 10046 3768 10102 3777
rect 10046 3703 10102 3712
rect 9954 3632 10010 3641
rect 9864 3596 9916 3602
rect 9954 3567 10010 3576
rect 9864 3538 9916 3544
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 9968 3176 9996 3567
rect 10048 3460 10100 3466
rect 10048 3402 10100 3408
rect 10060 3369 10088 3402
rect 10046 3360 10102 3369
rect 10046 3295 10102 3304
rect 9784 3148 9996 3176
rect 9680 3120 9732 3126
rect 9680 3062 9732 3068
rect 9784 2990 9812 3148
rect 9862 3088 9918 3097
rect 9862 3023 9918 3032
rect 9876 2990 9904 3023
rect 9772 2984 9824 2990
rect 9772 2926 9824 2932
rect 9864 2984 9916 2990
rect 9864 2926 9916 2932
rect 9680 2848 9732 2854
rect 9876 2825 9904 2926
rect 9956 2848 10008 2854
rect 9680 2790 9732 2796
rect 9862 2816 9918 2825
rect 9496 2644 9548 2650
rect 9496 2586 9548 2592
rect 9588 2644 9640 2650
rect 9588 2586 9640 2592
rect 9128 2576 9180 2582
rect 9128 2518 9180 2524
rect 9220 2576 9272 2582
rect 9220 2518 9272 2524
rect 9404 2508 9456 2514
rect 9404 2450 9456 2456
rect 9310 2408 9366 2417
rect 9128 2372 9180 2378
rect 9310 2343 9366 2352
rect 9128 2314 9180 2320
rect 9140 1426 9168 2314
rect 9128 1420 9180 1426
rect 9128 1362 9180 1368
rect 9324 800 9352 2343
rect 9416 2009 9444 2450
rect 9508 2310 9536 2586
rect 9692 2530 9720 2790
rect 9956 2790 10008 2796
rect 9862 2751 9918 2760
rect 9692 2502 9812 2530
rect 9496 2304 9548 2310
rect 9496 2246 9548 2252
rect 9508 2145 9536 2246
rect 9494 2136 9550 2145
rect 9494 2071 9550 2080
rect 9402 2000 9458 2009
rect 9402 1935 9458 1944
rect 9416 1902 9444 1935
rect 9404 1896 9456 1902
rect 9404 1838 9456 1844
rect 9784 1766 9812 2502
rect 9864 2508 9916 2514
rect 9864 2450 9916 2456
rect 9772 1760 9824 1766
rect 9772 1702 9824 1708
rect 9876 1562 9904 2450
rect 9968 1834 9996 2790
rect 10152 2394 10180 3998
rect 10336 3346 10364 4490
rect 10428 4185 10456 5034
rect 10520 4758 10548 5102
rect 10612 5098 10640 7103
rect 10782 7032 10838 7041
rect 10782 6967 10838 6976
rect 10796 6780 10824 6967
rect 10888 6905 10916 7278
rect 10950 7100 11246 7120
rect 11006 7098 11030 7100
rect 11086 7098 11110 7100
rect 11166 7098 11190 7100
rect 11028 7046 11030 7098
rect 11092 7046 11104 7098
rect 11166 7046 11168 7098
rect 11006 7044 11030 7046
rect 11086 7044 11110 7046
rect 11166 7044 11190 7046
rect 10950 7024 11246 7044
rect 10874 6896 10930 6905
rect 10874 6831 10930 6840
rect 11058 6896 11114 6905
rect 11058 6831 11114 6840
rect 11152 6860 11204 6866
rect 11072 6780 11100 6831
rect 11152 6802 11204 6808
rect 10796 6752 11100 6780
rect 11164 6769 11192 6802
rect 11150 6760 11206 6769
rect 11150 6695 11206 6704
rect 10876 6656 10928 6662
rect 11060 6656 11112 6662
rect 10928 6616 11008 6644
rect 10876 6598 10928 6604
rect 10784 6384 10836 6390
rect 10784 6326 10836 6332
rect 10876 6384 10928 6390
rect 10876 6326 10928 6332
rect 10692 6112 10744 6118
rect 10796 6089 10824 6326
rect 10888 6225 10916 6326
rect 10874 6216 10930 6225
rect 10980 6186 11008 6616
rect 11060 6598 11112 6604
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 11072 6225 11100 6598
rect 11164 6322 11192 6598
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 11058 6216 11114 6225
rect 10874 6151 10930 6160
rect 10968 6180 11020 6186
rect 11058 6151 11114 6160
rect 10968 6122 11020 6128
rect 10876 6112 10928 6118
rect 10692 6054 10744 6060
rect 10782 6080 10838 6089
rect 10704 5914 10732 6054
rect 10876 6054 10928 6060
rect 10782 6015 10838 6024
rect 10888 5930 10916 6054
rect 10950 6012 11246 6032
rect 11006 6010 11030 6012
rect 11086 6010 11110 6012
rect 11166 6010 11190 6012
rect 11028 5958 11030 6010
rect 11092 5958 11104 6010
rect 11166 5958 11168 6010
rect 11006 5956 11030 5958
rect 11086 5956 11110 5958
rect 11166 5956 11190 5958
rect 10950 5936 11246 5956
rect 10692 5908 10744 5914
rect 10692 5850 10744 5856
rect 10796 5902 10916 5930
rect 10600 5092 10652 5098
rect 10600 5034 10652 5040
rect 10598 4992 10654 5001
rect 10598 4927 10654 4936
rect 10508 4752 10560 4758
rect 10508 4694 10560 4700
rect 10612 4570 10640 4927
rect 10704 4690 10732 5850
rect 10796 5386 10824 5902
rect 11348 5896 11376 7278
rect 11440 7206 11468 7534
rect 11716 7528 11744 8298
rect 11808 8265 11836 11886
rect 11992 11830 12020 12650
rect 12256 12640 12308 12646
rect 12256 12582 12308 12588
rect 12268 12442 12296 12582
rect 12256 12436 12308 12442
rect 12256 12378 12308 12384
rect 12360 12238 12388 13262
rect 12440 12844 12492 12850
rect 12440 12786 12492 12792
rect 12348 12232 12400 12238
rect 12348 12174 12400 12180
rect 12072 12096 12124 12102
rect 12072 12038 12124 12044
rect 11980 11824 12032 11830
rect 11980 11766 12032 11772
rect 11992 11354 12020 11766
rect 11980 11348 12032 11354
rect 11980 11290 12032 11296
rect 11980 11212 12032 11218
rect 11980 11154 12032 11160
rect 11888 11144 11940 11150
rect 11888 11086 11940 11092
rect 11900 9897 11928 11086
rect 11992 10130 12020 11154
rect 12084 10985 12112 12038
rect 12452 11830 12480 12786
rect 12636 12424 12664 16934
rect 12820 16658 12848 17002
rect 12808 16652 12860 16658
rect 12808 16594 12860 16600
rect 12808 16448 12860 16454
rect 12808 16390 12860 16396
rect 12820 15552 12848 16390
rect 12912 16182 12940 17138
rect 13084 17128 13136 17134
rect 13084 17070 13136 17076
rect 12900 16176 12952 16182
rect 12900 16118 12952 16124
rect 12820 15524 12940 15552
rect 12808 15428 12860 15434
rect 12808 15370 12860 15376
rect 12716 12436 12768 12442
rect 12636 12396 12716 12424
rect 12716 12378 12768 12384
rect 12530 11928 12586 11937
rect 12530 11863 12532 11872
rect 12584 11863 12586 11872
rect 12532 11834 12584 11840
rect 12440 11824 12492 11830
rect 12440 11766 12492 11772
rect 12438 11656 12494 11665
rect 12438 11591 12494 11600
rect 12256 11280 12308 11286
rect 12254 11248 12256 11257
rect 12308 11248 12310 11257
rect 12254 11183 12310 11192
rect 12452 11082 12480 11591
rect 12544 11286 12572 11834
rect 12716 11756 12768 11762
rect 12716 11698 12768 11704
rect 12624 11620 12676 11626
rect 12624 11562 12676 11568
rect 12532 11280 12584 11286
rect 12532 11222 12584 11228
rect 12164 11076 12216 11082
rect 12164 11018 12216 11024
rect 12440 11076 12492 11082
rect 12440 11018 12492 11024
rect 12070 10976 12126 10985
rect 12070 10911 12126 10920
rect 12072 10804 12124 10810
rect 12072 10746 12124 10752
rect 12084 10441 12112 10746
rect 12070 10432 12126 10441
rect 12070 10367 12126 10376
rect 12084 10198 12112 10367
rect 12072 10192 12124 10198
rect 12072 10134 12124 10140
rect 11980 10124 12032 10130
rect 11980 10066 12032 10072
rect 11886 9888 11942 9897
rect 11886 9823 11942 9832
rect 12070 9888 12126 9897
rect 12070 9823 12126 9832
rect 11980 9716 12032 9722
rect 11980 9658 12032 9664
rect 11888 9376 11940 9382
rect 11886 9344 11888 9353
rect 11940 9344 11942 9353
rect 11886 9279 11942 9288
rect 11992 9178 12020 9658
rect 11980 9172 12032 9178
rect 11980 9114 12032 9120
rect 11888 9036 11940 9042
rect 11888 8978 11940 8984
rect 11794 8256 11850 8265
rect 11794 8191 11850 8200
rect 11794 8120 11850 8129
rect 11794 8055 11796 8064
rect 11848 8055 11850 8064
rect 11796 8026 11848 8032
rect 11900 7857 11928 8978
rect 11992 8809 12020 9114
rect 11978 8800 12034 8809
rect 11978 8735 12034 8744
rect 11978 8664 12034 8673
rect 11978 8599 12034 8608
rect 11992 8430 12020 8599
rect 11980 8424 12032 8430
rect 11980 8366 12032 8372
rect 11980 8288 12032 8294
rect 11980 8230 12032 8236
rect 11992 7886 12020 8230
rect 11980 7880 12032 7886
rect 11886 7848 11942 7857
rect 12084 7857 12112 9823
rect 12176 9586 12204 11018
rect 12254 10976 12310 10985
rect 12254 10911 12310 10920
rect 12268 10538 12296 10911
rect 12636 10810 12664 11562
rect 12728 11150 12756 11698
rect 12716 11144 12768 11150
rect 12714 11112 12716 11121
rect 12768 11112 12770 11121
rect 12714 11047 12770 11056
rect 12820 10810 12848 15370
rect 12912 10826 12940 15524
rect 12992 12436 13044 12442
rect 12992 12378 13044 12384
rect 13004 11914 13032 12378
rect 13096 12345 13124 17070
rect 13280 16674 13308 19200
rect 13648 17626 13676 19200
rect 13648 17598 13860 17626
rect 13449 17436 13745 17456
rect 13505 17434 13529 17436
rect 13585 17434 13609 17436
rect 13665 17434 13689 17436
rect 13527 17382 13529 17434
rect 13591 17382 13603 17434
rect 13665 17382 13667 17434
rect 13505 17380 13529 17382
rect 13585 17380 13609 17382
rect 13665 17380 13689 17382
rect 13449 17360 13745 17380
rect 13832 17338 13860 17598
rect 13820 17332 13872 17338
rect 13820 17274 13872 17280
rect 13832 17134 13860 17274
rect 13820 17128 13872 17134
rect 13820 17070 13872 17076
rect 14016 17082 14044 19200
rect 14384 17134 14412 19200
rect 14648 17332 14700 17338
rect 14648 17274 14700 17280
rect 14096 17128 14148 17134
rect 14016 17076 14096 17082
rect 14016 17070 14148 17076
rect 14372 17128 14424 17134
rect 14372 17070 14424 17076
rect 14016 17054 14136 17070
rect 14016 16794 14044 17054
rect 14096 16992 14148 16998
rect 14096 16934 14148 16940
rect 14004 16788 14056 16794
rect 14004 16730 14056 16736
rect 13360 16720 13412 16726
rect 13280 16668 13360 16674
rect 13280 16662 13412 16668
rect 13280 16646 13400 16662
rect 13268 16516 13320 16522
rect 13268 16458 13320 16464
rect 13176 16448 13228 16454
rect 13176 16390 13228 16396
rect 13082 12336 13138 12345
rect 13082 12271 13138 12280
rect 13004 11886 13124 11914
rect 12992 11824 13044 11830
rect 12992 11766 13044 11772
rect 13004 11286 13032 11766
rect 13096 11558 13124 11886
rect 13188 11626 13216 16390
rect 13280 12442 13308 16458
rect 13372 16250 13400 16646
rect 13912 16516 13964 16522
rect 13912 16458 13964 16464
rect 13449 16348 13745 16368
rect 13505 16346 13529 16348
rect 13585 16346 13609 16348
rect 13665 16346 13689 16348
rect 13527 16294 13529 16346
rect 13591 16294 13603 16346
rect 13665 16294 13667 16346
rect 13505 16292 13529 16294
rect 13585 16292 13609 16294
rect 13665 16292 13689 16294
rect 13449 16272 13745 16292
rect 13360 16244 13412 16250
rect 13360 16186 13412 16192
rect 13820 15972 13872 15978
rect 13820 15914 13872 15920
rect 13449 15260 13745 15280
rect 13505 15258 13529 15260
rect 13585 15258 13609 15260
rect 13665 15258 13689 15260
rect 13527 15206 13529 15258
rect 13591 15206 13603 15258
rect 13665 15206 13667 15258
rect 13505 15204 13529 15206
rect 13585 15204 13609 15206
rect 13665 15204 13689 15206
rect 13449 15184 13745 15204
rect 13449 14172 13745 14192
rect 13505 14170 13529 14172
rect 13585 14170 13609 14172
rect 13665 14170 13689 14172
rect 13527 14118 13529 14170
rect 13591 14118 13603 14170
rect 13665 14118 13667 14170
rect 13505 14116 13529 14118
rect 13585 14116 13609 14118
rect 13665 14116 13689 14118
rect 13449 14096 13745 14116
rect 13449 13084 13745 13104
rect 13505 13082 13529 13084
rect 13585 13082 13609 13084
rect 13665 13082 13689 13084
rect 13527 13030 13529 13082
rect 13591 13030 13603 13082
rect 13665 13030 13667 13082
rect 13505 13028 13529 13030
rect 13585 13028 13609 13030
rect 13665 13028 13689 13030
rect 13449 13008 13745 13028
rect 13268 12436 13320 12442
rect 13320 12396 13400 12424
rect 13268 12378 13320 12384
rect 13372 12102 13400 12396
rect 13360 12096 13412 12102
rect 13360 12038 13412 12044
rect 13372 11898 13400 12038
rect 13449 11996 13745 12016
rect 13505 11994 13529 11996
rect 13585 11994 13609 11996
rect 13665 11994 13689 11996
rect 13527 11942 13529 11994
rect 13591 11942 13603 11994
rect 13665 11942 13667 11994
rect 13505 11940 13529 11942
rect 13585 11940 13609 11942
rect 13665 11940 13689 11942
rect 13449 11920 13745 11940
rect 13360 11892 13412 11898
rect 13360 11834 13412 11840
rect 13176 11620 13228 11626
rect 13176 11562 13228 11568
rect 13084 11552 13136 11558
rect 13084 11494 13136 11500
rect 12992 11280 13044 11286
rect 12992 11222 13044 11228
rect 13176 11280 13228 11286
rect 13176 11222 13228 11228
rect 12624 10804 12676 10810
rect 12624 10746 12676 10752
rect 12808 10804 12860 10810
rect 12912 10798 13032 10826
rect 12808 10746 12860 10752
rect 12900 10736 12952 10742
rect 12900 10678 12952 10684
rect 12624 10668 12676 10674
rect 12624 10610 12676 10616
rect 12256 10532 12308 10538
rect 12256 10474 12308 10480
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12254 10296 12310 10305
rect 12452 10282 12480 10406
rect 12452 10266 12572 10282
rect 12452 10260 12584 10266
rect 12452 10254 12532 10260
rect 12254 10231 12256 10240
rect 12308 10231 12310 10240
rect 12256 10202 12308 10208
rect 12532 10202 12584 10208
rect 12348 10124 12400 10130
rect 12348 10066 12400 10072
rect 12360 9674 12388 10066
rect 12440 10056 12492 10062
rect 12440 9998 12492 10004
rect 12452 9897 12480 9998
rect 12438 9888 12494 9897
rect 12438 9823 12494 9832
rect 12636 9704 12664 10610
rect 12808 10464 12860 10470
rect 12808 10406 12860 10412
rect 12716 9988 12768 9994
rect 12716 9930 12768 9936
rect 12268 9646 12388 9674
rect 12452 9676 12664 9704
rect 12164 9580 12216 9586
rect 12164 9522 12216 9528
rect 12268 9518 12296 9646
rect 12348 9580 12400 9586
rect 12452 9568 12480 9676
rect 12622 9616 12678 9625
rect 12400 9540 12480 9568
rect 12532 9580 12584 9586
rect 12348 9522 12400 9528
rect 12728 9586 12756 9930
rect 12820 9625 12848 10406
rect 12912 9722 12940 10678
rect 12900 9716 12952 9722
rect 12900 9658 12952 9664
rect 12806 9616 12862 9625
rect 12622 9551 12678 9560
rect 12716 9580 12768 9586
rect 12532 9522 12584 9528
rect 12256 9512 12308 9518
rect 12256 9454 12308 9460
rect 12162 9208 12218 9217
rect 12162 9143 12218 9152
rect 12176 8634 12204 9143
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 12360 8634 12388 8910
rect 12544 8838 12572 9522
rect 12636 9178 12664 9551
rect 12806 9551 12862 9560
rect 12716 9522 12768 9528
rect 12808 9512 12860 9518
rect 12806 9480 12808 9489
rect 13004 9500 13032 10798
rect 13084 10804 13136 10810
rect 13084 10746 13136 10752
rect 12860 9480 13032 9500
rect 12862 9472 13032 9480
rect 12806 9415 12862 9424
rect 12900 9376 12952 9382
rect 12900 9318 12952 9324
rect 12912 9217 12940 9318
rect 12898 9208 12954 9217
rect 12624 9172 12676 9178
rect 12808 9172 12860 9178
rect 12624 9114 12676 9120
rect 12728 9132 12808 9160
rect 12728 9081 12756 9132
rect 12898 9143 12954 9152
rect 12808 9114 12860 9120
rect 12714 9072 12770 9081
rect 13096 9058 13124 10746
rect 13188 10169 13216 11222
rect 13268 11144 13320 11150
rect 13268 11086 13320 11092
rect 13280 10849 13308 11086
rect 13360 11008 13412 11014
rect 13360 10950 13412 10956
rect 13266 10840 13322 10849
rect 13266 10775 13322 10784
rect 13372 10538 13400 10950
rect 13449 10908 13745 10928
rect 13505 10906 13529 10908
rect 13585 10906 13609 10908
rect 13665 10906 13689 10908
rect 13527 10854 13529 10906
rect 13591 10854 13603 10906
rect 13665 10854 13667 10906
rect 13505 10852 13529 10854
rect 13585 10852 13609 10854
rect 13665 10852 13689 10854
rect 13449 10832 13745 10852
rect 13450 10704 13506 10713
rect 13450 10639 13506 10648
rect 13268 10532 13320 10538
rect 13268 10474 13320 10480
rect 13360 10532 13412 10538
rect 13360 10474 13412 10480
rect 13280 10266 13308 10474
rect 13268 10260 13320 10266
rect 13268 10202 13320 10208
rect 13174 10160 13230 10169
rect 13174 10095 13230 10104
rect 13268 10124 13320 10130
rect 12714 9007 12770 9016
rect 12820 9030 13124 9058
rect 12716 8968 12768 8974
rect 12716 8910 12768 8916
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 12164 8628 12216 8634
rect 12164 8570 12216 8576
rect 12348 8628 12400 8634
rect 12348 8570 12400 8576
rect 12532 8560 12584 8566
rect 12530 8528 12532 8537
rect 12584 8528 12586 8537
rect 12440 8492 12492 8498
rect 12530 8463 12586 8472
rect 12440 8434 12492 8440
rect 12164 8424 12216 8430
rect 12164 8366 12216 8372
rect 12176 8265 12204 8366
rect 12348 8288 12400 8294
rect 12162 8256 12218 8265
rect 12162 8191 12218 8200
rect 12268 8248 12348 8276
rect 11980 7822 12032 7828
rect 12070 7848 12126 7857
rect 11886 7783 11942 7792
rect 11716 7500 11836 7528
rect 11702 7440 11758 7449
rect 11702 7375 11758 7384
rect 11716 7206 11744 7375
rect 11428 7200 11480 7206
rect 11428 7142 11480 7148
rect 11704 7200 11756 7206
rect 11704 7142 11756 7148
rect 11808 6934 11836 7500
rect 11992 7449 12020 7822
rect 12070 7783 12126 7792
rect 12176 7721 12204 8191
rect 12268 8090 12296 8248
rect 12348 8230 12400 8236
rect 12256 8084 12308 8090
rect 12256 8026 12308 8032
rect 12348 8084 12400 8090
rect 12348 8026 12400 8032
rect 12254 7984 12310 7993
rect 12254 7919 12310 7928
rect 12268 7818 12296 7919
rect 12256 7812 12308 7818
rect 12256 7754 12308 7760
rect 12360 7750 12388 8026
rect 12452 7993 12480 8434
rect 12532 8424 12584 8430
rect 12532 8366 12584 8372
rect 12624 8424 12676 8430
rect 12624 8366 12676 8372
rect 12438 7984 12494 7993
rect 12544 7954 12572 8366
rect 12636 8265 12664 8366
rect 12622 8256 12678 8265
rect 12622 8191 12678 8200
rect 12438 7919 12494 7928
rect 12532 7948 12584 7954
rect 12532 7890 12584 7896
rect 12440 7880 12492 7886
rect 12440 7822 12492 7828
rect 12348 7744 12400 7750
rect 12162 7712 12218 7721
rect 12348 7686 12400 7692
rect 12162 7647 12218 7656
rect 11978 7440 12034 7449
rect 11978 7375 12034 7384
rect 11980 7336 12032 7342
rect 12176 7290 12204 7647
rect 11980 7278 12032 7284
rect 11886 7168 11942 7177
rect 11886 7103 11942 7112
rect 11612 6928 11664 6934
rect 11796 6928 11848 6934
rect 11612 6870 11664 6876
rect 11702 6896 11758 6905
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 11428 6180 11480 6186
rect 11428 6122 11480 6128
rect 11256 5868 11376 5896
rect 10876 5840 10928 5846
rect 10928 5800 11100 5828
rect 10876 5782 10928 5788
rect 10888 5710 10916 5782
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 10966 5672 11022 5681
rect 10966 5607 11022 5616
rect 10796 5358 10916 5386
rect 10782 5264 10838 5273
rect 10782 5199 10838 5208
rect 10796 5098 10824 5199
rect 10784 5092 10836 5098
rect 10784 5034 10836 5040
rect 10796 4865 10824 5034
rect 10782 4856 10838 4865
rect 10782 4791 10838 4800
rect 10692 4684 10744 4690
rect 10692 4626 10744 4632
rect 10612 4542 10824 4570
rect 10796 4486 10824 4542
rect 10508 4480 10560 4486
rect 10508 4422 10560 4428
rect 10692 4480 10744 4486
rect 10692 4422 10744 4428
rect 10784 4480 10836 4486
rect 10784 4422 10836 4428
rect 10414 4176 10470 4185
rect 10414 4111 10470 4120
rect 10428 4010 10456 4111
rect 10416 4004 10468 4010
rect 10416 3946 10468 3952
rect 10414 3768 10470 3777
rect 10414 3703 10470 3712
rect 10428 3670 10456 3703
rect 10416 3664 10468 3670
rect 10416 3606 10468 3612
rect 10520 3602 10548 4422
rect 10508 3596 10560 3602
rect 10508 3538 10560 3544
rect 10508 3460 10560 3466
rect 10508 3402 10560 3408
rect 10244 3318 10364 3346
rect 10416 3392 10468 3398
rect 10416 3334 10468 3340
rect 10244 2990 10272 3318
rect 10322 3224 10378 3233
rect 10322 3159 10378 3168
rect 10232 2984 10284 2990
rect 10232 2926 10284 2932
rect 10232 2848 10284 2854
rect 10232 2790 10284 2796
rect 10060 2366 10180 2394
rect 9956 1828 10008 1834
rect 9956 1770 10008 1776
rect 10060 1698 10088 2366
rect 10140 2304 10192 2310
rect 10140 2246 10192 2252
rect 10152 1970 10180 2246
rect 10140 1964 10192 1970
rect 10140 1906 10192 1912
rect 10048 1692 10100 1698
rect 10048 1634 10100 1640
rect 9864 1556 9916 1562
rect 9864 1498 9916 1504
rect 9680 1488 9732 1494
rect 9680 1430 9732 1436
rect 9692 800 9720 1430
rect 10244 1426 10272 2790
rect 10336 2650 10364 3159
rect 10428 2650 10456 3334
rect 10520 3097 10548 3402
rect 10600 3392 10652 3398
rect 10704 3380 10732 4422
rect 10888 4214 10916 5358
rect 10980 5166 11008 5607
rect 11072 5574 11100 5800
rect 11060 5568 11112 5574
rect 11060 5510 11112 5516
rect 11256 5250 11284 5868
rect 11334 5672 11390 5681
rect 11334 5607 11390 5616
rect 11348 5370 11376 5607
rect 11440 5370 11468 6122
rect 11532 5710 11560 6734
rect 11520 5704 11572 5710
rect 11520 5646 11572 5652
rect 11336 5364 11388 5370
rect 11336 5306 11388 5312
rect 11428 5364 11480 5370
rect 11428 5306 11480 5312
rect 11256 5222 11376 5250
rect 10968 5160 11020 5166
rect 10968 5102 11020 5108
rect 11058 5128 11114 5137
rect 11058 5063 11060 5072
rect 11112 5063 11114 5072
rect 11060 5034 11112 5040
rect 10950 4924 11246 4944
rect 11006 4922 11030 4924
rect 11086 4922 11110 4924
rect 11166 4922 11190 4924
rect 11028 4870 11030 4922
rect 11092 4870 11104 4922
rect 11166 4870 11168 4922
rect 11006 4868 11030 4870
rect 11086 4868 11110 4870
rect 11166 4868 11190 4870
rect 10950 4848 11246 4868
rect 11348 4808 11376 5222
rect 11520 5228 11572 5234
rect 11520 5170 11572 5176
rect 11532 5137 11560 5170
rect 11518 5128 11574 5137
rect 11518 5063 11574 5072
rect 11520 5024 11572 5030
rect 11426 4992 11482 5001
rect 11520 4966 11572 4972
rect 11426 4927 11482 4936
rect 11164 4780 11376 4808
rect 11060 4752 11112 4758
rect 11060 4694 11112 4700
rect 11072 4554 11100 4694
rect 11060 4548 11112 4554
rect 11060 4490 11112 4496
rect 11164 4214 11192 4780
rect 11440 4740 11468 4927
rect 11348 4712 11468 4740
rect 11348 4554 11376 4712
rect 11532 4604 11560 4966
rect 11440 4576 11560 4604
rect 11336 4548 11388 4554
rect 11336 4490 11388 4496
rect 10876 4208 10928 4214
rect 10876 4150 10928 4156
rect 11152 4208 11204 4214
rect 11152 4150 11204 4156
rect 11244 4140 11296 4146
rect 11244 4082 11296 4088
rect 10784 4072 10836 4078
rect 10784 4014 10836 4020
rect 10796 3913 10824 4014
rect 11060 4004 11112 4010
rect 11256 3992 11284 4082
rect 11112 3964 11284 3992
rect 11060 3946 11112 3952
rect 10876 3936 10928 3942
rect 10782 3904 10838 3913
rect 10876 3878 10928 3884
rect 11336 3936 11388 3942
rect 11336 3878 11388 3884
rect 10782 3839 10838 3848
rect 10888 3738 10916 3878
rect 10950 3836 11246 3856
rect 11006 3834 11030 3836
rect 11086 3834 11110 3836
rect 11166 3834 11190 3836
rect 11028 3782 11030 3834
rect 11092 3782 11104 3834
rect 11166 3782 11168 3834
rect 11006 3780 11030 3782
rect 11086 3780 11110 3782
rect 11166 3780 11190 3782
rect 10950 3760 11246 3780
rect 10784 3732 10836 3738
rect 10784 3674 10836 3680
rect 10876 3732 10928 3738
rect 10876 3674 10928 3680
rect 10796 3482 10824 3674
rect 11348 3618 11376 3878
rect 10980 3590 11376 3618
rect 10796 3454 10892 3482
rect 10864 3448 10892 3454
rect 10864 3420 10916 3448
rect 10784 3392 10836 3398
rect 10704 3352 10784 3380
rect 10600 3334 10652 3340
rect 10784 3334 10836 3340
rect 10506 3088 10562 3097
rect 10506 3023 10562 3032
rect 10520 2990 10548 3023
rect 10517 2984 10569 2990
rect 10517 2926 10569 2932
rect 10324 2644 10376 2650
rect 10324 2586 10376 2592
rect 10416 2644 10468 2650
rect 10416 2586 10468 2592
rect 10506 2544 10562 2553
rect 10324 2508 10376 2514
rect 10324 2450 10376 2456
rect 10416 2508 10468 2514
rect 10612 2514 10640 3334
rect 10796 2689 10824 3334
rect 10888 2938 10916 3420
rect 10980 3233 11008 3590
rect 11440 3584 11468 4576
rect 11520 4208 11572 4214
rect 11520 4150 11572 4156
rect 11532 3913 11560 4150
rect 11518 3904 11574 3913
rect 11518 3839 11574 3848
rect 11518 3768 11574 3777
rect 11518 3703 11520 3712
rect 11572 3703 11574 3712
rect 11520 3674 11572 3680
rect 11440 3556 11560 3584
rect 11428 3460 11480 3466
rect 11428 3402 11480 3408
rect 11060 3392 11112 3398
rect 11060 3334 11112 3340
rect 10966 3224 11022 3233
rect 10966 3159 11022 3168
rect 11072 3126 11100 3334
rect 11060 3120 11112 3126
rect 11060 3062 11112 3068
rect 11242 3088 11298 3097
rect 11242 3023 11298 3032
rect 11152 2984 11204 2990
rect 10888 2910 11008 2938
rect 11256 2972 11284 3023
rect 11204 2944 11284 2972
rect 11353 2984 11405 2990
rect 11152 2926 11204 2932
rect 11440 2972 11468 3402
rect 11405 2944 11468 2972
rect 11353 2926 11405 2932
rect 10876 2848 10928 2854
rect 10980 2836 11008 2910
rect 11532 2904 11560 3556
rect 11624 3505 11652 6870
rect 11796 6870 11848 6876
rect 11702 6831 11758 6840
rect 11716 6798 11744 6831
rect 11704 6792 11756 6798
rect 11704 6734 11756 6740
rect 11796 6792 11848 6798
rect 11796 6734 11848 6740
rect 11716 6202 11744 6734
rect 11808 6458 11836 6734
rect 11796 6452 11848 6458
rect 11796 6394 11848 6400
rect 11900 6390 11928 7103
rect 11992 7002 12020 7278
rect 12084 7262 12204 7290
rect 11980 6996 12032 7002
rect 11980 6938 12032 6944
rect 11980 6860 12032 6866
rect 11980 6802 12032 6808
rect 11888 6384 11940 6390
rect 11992 6361 12020 6802
rect 11888 6326 11940 6332
rect 11978 6352 12034 6361
rect 11716 6174 11836 6202
rect 11704 6112 11756 6118
rect 11704 6054 11756 6060
rect 11716 5817 11744 6054
rect 11808 5953 11836 6174
rect 11794 5944 11850 5953
rect 11900 5914 11928 6326
rect 11978 6287 12034 6296
rect 11980 6180 12032 6186
rect 11980 6122 12032 6128
rect 11794 5879 11850 5888
rect 11888 5908 11940 5914
rect 11702 5808 11758 5817
rect 11702 5743 11758 5752
rect 11704 5636 11756 5642
rect 11704 5578 11756 5584
rect 11716 5545 11744 5578
rect 11702 5536 11758 5545
rect 11702 5471 11758 5480
rect 11808 5234 11836 5879
rect 11888 5850 11940 5856
rect 11888 5772 11940 5778
rect 11888 5714 11940 5720
rect 11796 5228 11848 5234
rect 11796 5170 11848 5176
rect 11796 5024 11848 5030
rect 11796 4966 11848 4972
rect 11702 4856 11758 4865
rect 11702 4791 11704 4800
rect 11756 4791 11758 4800
rect 11704 4762 11756 4768
rect 11702 4720 11758 4729
rect 11702 4655 11704 4664
rect 11756 4655 11758 4664
rect 11704 4626 11756 4632
rect 11716 4457 11744 4626
rect 11808 4554 11836 4966
rect 11900 4865 11928 5714
rect 11992 5001 12020 6122
rect 11978 4992 12034 5001
rect 11978 4927 12034 4936
rect 11886 4856 11942 4865
rect 11886 4791 11942 4800
rect 11888 4684 11940 4690
rect 11888 4626 11940 4632
rect 11796 4548 11848 4554
rect 11796 4490 11848 4496
rect 11702 4448 11758 4457
rect 11900 4434 11928 4626
rect 11978 4584 12034 4593
rect 11978 4519 11980 4528
rect 12032 4519 12034 4528
rect 11980 4490 12032 4496
rect 11702 4383 11758 4392
rect 11808 4406 11928 4434
rect 11808 4078 11836 4406
rect 12084 4321 12112 7262
rect 12164 7200 12216 7206
rect 12164 7142 12216 7148
rect 12348 7200 12400 7206
rect 12348 7142 12400 7148
rect 12176 6905 12204 7142
rect 12360 7041 12388 7142
rect 12346 7032 12402 7041
rect 12256 6996 12308 7002
rect 12346 6967 12402 6976
rect 12256 6938 12308 6944
rect 12162 6896 12218 6905
rect 12162 6831 12218 6840
rect 12268 6730 12296 6938
rect 12348 6928 12400 6934
rect 12452 6916 12480 7822
rect 12532 7744 12584 7750
rect 12532 7686 12584 7692
rect 12544 7546 12572 7686
rect 12728 7546 12756 8910
rect 12532 7540 12584 7546
rect 12532 7482 12584 7488
rect 12716 7540 12768 7546
rect 12716 7482 12768 7488
rect 12400 6888 12480 6916
rect 12348 6870 12400 6876
rect 12256 6724 12308 6730
rect 12256 6666 12308 6672
rect 12268 6372 12296 6666
rect 12176 6344 12296 6372
rect 12176 6089 12204 6344
rect 12360 6304 12388 6870
rect 12438 6488 12494 6497
rect 12438 6423 12494 6432
rect 12268 6276 12388 6304
rect 12162 6080 12218 6089
rect 12162 6015 12218 6024
rect 11886 4312 11942 4321
rect 11886 4247 11942 4256
rect 12070 4312 12126 4321
rect 12070 4247 12126 4256
rect 11796 4072 11848 4078
rect 11796 4014 11848 4020
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 11716 3534 11744 3878
rect 11796 3664 11848 3670
rect 11796 3606 11848 3612
rect 11704 3528 11756 3534
rect 11610 3496 11666 3505
rect 11808 3505 11836 3606
rect 11704 3470 11756 3476
rect 11794 3496 11850 3505
rect 11610 3431 11666 3440
rect 11900 3482 11928 4247
rect 11980 4208 12032 4214
rect 11980 4150 12032 4156
rect 11992 3641 12020 4150
rect 12072 4072 12124 4078
rect 12072 4014 12124 4020
rect 11978 3632 12034 3641
rect 12084 3602 12112 4014
rect 11978 3567 12034 3576
rect 12072 3596 12124 3602
rect 12072 3538 12124 3544
rect 11900 3454 12112 3482
rect 11794 3431 11850 3440
rect 11612 3392 11664 3398
rect 11980 3392 12032 3398
rect 11664 3352 11980 3380
rect 11612 3334 11664 3340
rect 11980 3334 12032 3340
rect 11796 3188 11848 3194
rect 11624 3148 11796 3176
rect 11624 3058 11652 3148
rect 11796 3130 11848 3136
rect 11980 3188 12032 3194
rect 12084 3176 12112 3454
rect 12032 3148 12112 3176
rect 11980 3130 12032 3136
rect 11612 3052 11664 3058
rect 11612 2994 11664 3000
rect 11796 3052 11848 3058
rect 11796 2994 11848 3000
rect 11704 2984 11756 2990
rect 11704 2926 11756 2932
rect 11440 2876 11560 2904
rect 11612 2916 11664 2922
rect 10980 2808 11376 2836
rect 10876 2790 10928 2796
rect 10782 2680 10838 2689
rect 10782 2615 10838 2624
rect 10506 2479 10562 2488
rect 10600 2508 10652 2514
rect 10416 2450 10468 2456
rect 10336 1902 10364 2450
rect 10428 2310 10456 2450
rect 10520 2446 10548 2479
rect 10600 2450 10652 2456
rect 10508 2440 10560 2446
rect 10508 2382 10560 2388
rect 10416 2304 10468 2310
rect 10416 2246 10468 2252
rect 10612 1986 10640 2450
rect 10428 1958 10640 1986
rect 10324 1896 10376 1902
rect 10324 1838 10376 1844
rect 10232 1420 10284 1426
rect 10232 1362 10284 1368
rect 10336 1306 10364 1838
rect 10060 1278 10364 1306
rect 10060 800 10088 1278
rect 10428 800 10456 1958
rect 10796 1834 10824 2615
rect 10888 2582 10916 2790
rect 10950 2748 11246 2768
rect 11006 2746 11030 2748
rect 11086 2746 11110 2748
rect 11166 2746 11190 2748
rect 11028 2694 11030 2746
rect 11092 2694 11104 2746
rect 11166 2694 11168 2746
rect 11006 2692 11030 2694
rect 11086 2692 11110 2694
rect 11166 2692 11190 2694
rect 10950 2672 11246 2692
rect 11348 2632 11376 2808
rect 11256 2604 11376 2632
rect 10876 2576 10928 2582
rect 11060 2576 11112 2582
rect 10876 2518 10928 2524
rect 10966 2544 11022 2553
rect 11152 2576 11204 2582
rect 11112 2536 11152 2564
rect 11060 2518 11112 2524
rect 11152 2518 11204 2524
rect 11256 2514 11284 2604
rect 10966 2479 11022 2488
rect 11244 2508 11296 2514
rect 10980 2310 11008 2479
rect 11244 2450 11296 2456
rect 10968 2304 11020 2310
rect 10968 2246 11020 2252
rect 11244 2304 11296 2310
rect 11244 2246 11296 2252
rect 11256 2106 11284 2246
rect 11244 2100 11296 2106
rect 11244 2042 11296 2048
rect 10784 1828 10836 1834
rect 10784 1770 10836 1776
rect 10692 1760 10744 1766
rect 10692 1702 10744 1708
rect 11058 1728 11114 1737
rect 10704 800 10732 1702
rect 11058 1663 11114 1672
rect 11072 800 11100 1663
rect 11440 1630 11468 2876
rect 11612 2858 11664 2864
rect 11518 2816 11574 2825
rect 11518 2751 11574 2760
rect 11532 2650 11560 2751
rect 11520 2644 11572 2650
rect 11520 2586 11572 2592
rect 11520 2508 11572 2514
rect 11520 2450 11572 2456
rect 11532 1766 11560 2450
rect 11624 2417 11652 2858
rect 11716 2689 11744 2926
rect 11702 2680 11758 2689
rect 11808 2650 11836 2994
rect 12072 2984 12124 2990
rect 11886 2952 11942 2961
rect 12072 2926 12124 2932
rect 11886 2887 11942 2896
rect 11702 2615 11758 2624
rect 11796 2644 11848 2650
rect 11610 2408 11666 2417
rect 11610 2343 11666 2352
rect 11520 1760 11572 1766
rect 11520 1702 11572 1708
rect 11428 1624 11480 1630
rect 11428 1566 11480 1572
rect 11716 1476 11744 2615
rect 11796 2586 11848 2592
rect 11796 2508 11848 2514
rect 11796 2450 11848 2456
rect 11440 1448 11744 1476
rect 11440 800 11468 1448
rect 11808 800 11836 2450
rect 11900 2360 11928 2887
rect 11980 2848 12032 2854
rect 11978 2816 11980 2825
rect 12032 2816 12034 2825
rect 11978 2751 12034 2760
rect 11980 2644 12032 2650
rect 11980 2586 12032 2592
rect 11992 2553 12020 2586
rect 11978 2544 12034 2553
rect 11978 2479 12034 2488
rect 11980 2372 12032 2378
rect 11900 2332 11980 2360
rect 11980 2314 12032 2320
rect 12084 800 12112 2926
rect 12176 1970 12204 6015
rect 12268 5681 12296 6276
rect 12452 6118 12480 6423
rect 12348 6112 12400 6118
rect 12346 6080 12348 6089
rect 12440 6112 12492 6118
rect 12400 6080 12402 6089
rect 12440 6054 12492 6060
rect 12346 6015 12402 6024
rect 12254 5672 12310 5681
rect 12254 5607 12310 5616
rect 12256 5364 12308 5370
rect 12256 5306 12308 5312
rect 12268 4282 12296 5306
rect 12360 4690 12388 6015
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 12452 5778 12480 5850
rect 12440 5772 12492 5778
rect 12440 5714 12492 5720
rect 12440 5636 12492 5642
rect 12440 5578 12492 5584
rect 12452 5409 12480 5578
rect 12438 5400 12494 5409
rect 12438 5335 12494 5344
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 12452 4826 12480 5102
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 12348 4684 12400 4690
rect 12348 4626 12400 4632
rect 12348 4548 12400 4554
rect 12348 4490 12400 4496
rect 12256 4276 12308 4282
rect 12256 4218 12308 4224
rect 12268 3738 12296 4218
rect 12360 4010 12388 4490
rect 12438 4312 12494 4321
rect 12544 4282 12572 7482
rect 12624 7268 12676 7274
rect 12624 7210 12676 7216
rect 12636 7041 12664 7210
rect 12622 7032 12678 7041
rect 12820 7018 12848 9030
rect 12900 8968 12952 8974
rect 13188 8956 13216 10095
rect 13268 10066 13320 10072
rect 12900 8910 12952 8916
rect 13096 8928 13216 8956
rect 12912 8498 12940 8910
rect 12992 8900 13044 8906
rect 12992 8842 13044 8848
rect 12900 8492 12952 8498
rect 12900 8434 12952 8440
rect 12898 7984 12954 7993
rect 12898 7919 12954 7928
rect 12912 7886 12940 7919
rect 12900 7880 12952 7886
rect 12900 7822 12952 7828
rect 12912 7342 12940 7822
rect 13004 7750 13032 8842
rect 13096 7954 13124 8928
rect 13280 8786 13308 10066
rect 13464 10062 13492 10639
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13740 10305 13768 10406
rect 13726 10296 13782 10305
rect 13832 10266 13860 15914
rect 13924 10742 13952 16458
rect 14108 14822 14136 16934
rect 14384 16658 14412 17070
rect 14556 16720 14608 16726
rect 14556 16662 14608 16668
rect 14372 16652 14424 16658
rect 14372 16594 14424 16600
rect 14464 16448 14516 16454
rect 14464 16390 14516 16396
rect 14372 14884 14424 14890
rect 14372 14826 14424 14832
rect 14096 14816 14148 14822
rect 14096 14758 14148 14764
rect 14188 14000 14240 14006
rect 14188 13942 14240 13948
rect 14096 12776 14148 12782
rect 14096 12718 14148 12724
rect 14004 12096 14056 12102
rect 14004 12038 14056 12044
rect 14016 11762 14044 12038
rect 14004 11756 14056 11762
rect 14004 11698 14056 11704
rect 14004 11076 14056 11082
rect 14004 11018 14056 11024
rect 13912 10736 13964 10742
rect 13912 10678 13964 10684
rect 14016 10606 14044 11018
rect 14108 10606 14136 12718
rect 14200 10810 14228 13942
rect 14280 13864 14332 13870
rect 14280 13806 14332 13812
rect 14188 10804 14240 10810
rect 14188 10746 14240 10752
rect 14004 10600 14056 10606
rect 14004 10542 14056 10548
rect 14096 10600 14148 10606
rect 14096 10542 14148 10548
rect 13910 10432 13966 10441
rect 13910 10367 13966 10376
rect 13726 10231 13782 10240
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 13452 10056 13504 10062
rect 13452 9998 13504 10004
rect 13449 9820 13745 9840
rect 13505 9818 13529 9820
rect 13585 9818 13609 9820
rect 13665 9818 13689 9820
rect 13527 9766 13529 9818
rect 13591 9766 13603 9818
rect 13665 9766 13667 9818
rect 13505 9764 13529 9766
rect 13585 9764 13609 9766
rect 13665 9764 13689 9766
rect 13449 9744 13745 9764
rect 13832 9704 13860 10202
rect 13924 10130 13952 10367
rect 13912 10124 13964 10130
rect 13912 10066 13964 10072
rect 14016 10010 14044 10542
rect 14096 10464 14148 10470
rect 14096 10406 14148 10412
rect 14108 10266 14136 10406
rect 14096 10260 14148 10266
rect 14096 10202 14148 10208
rect 14292 10198 14320 13806
rect 14384 11354 14412 14826
rect 14476 13870 14504 16390
rect 14568 16250 14596 16662
rect 14556 16244 14608 16250
rect 14556 16186 14608 16192
rect 14556 14816 14608 14822
rect 14556 14758 14608 14764
rect 14464 13864 14516 13870
rect 14464 13806 14516 13812
rect 14464 13728 14516 13734
rect 14464 13670 14516 13676
rect 14476 12918 14504 13670
rect 14464 12912 14516 12918
rect 14464 12854 14516 12860
rect 14476 11778 14504 12854
rect 14568 11880 14596 14758
rect 14660 12102 14688 17274
rect 14752 17202 14780 19200
rect 14740 17196 14792 17202
rect 14740 17138 14792 17144
rect 14752 16250 14780 17138
rect 14832 17060 14884 17066
rect 14832 17002 14884 17008
rect 14740 16244 14792 16250
rect 14740 16186 14792 16192
rect 14844 13734 14872 17002
rect 14922 16688 14978 16697
rect 15120 16674 15148 19200
rect 15292 17060 15344 17066
rect 15292 17002 15344 17008
rect 15200 16720 15252 16726
rect 15120 16668 15200 16674
rect 15120 16662 15252 16668
rect 15120 16646 15240 16662
rect 14922 16623 14978 16632
rect 14936 16250 14964 16623
rect 15108 16516 15160 16522
rect 15108 16458 15160 16464
rect 14924 16244 14976 16250
rect 14924 16186 14976 16192
rect 14832 13728 14884 13734
rect 14832 13670 14884 13676
rect 14648 12096 14700 12102
rect 14648 12038 14700 12044
rect 14568 11852 15056 11880
rect 14476 11750 14964 11778
rect 14740 11688 14792 11694
rect 14740 11630 14792 11636
rect 14648 11620 14700 11626
rect 14648 11562 14700 11568
rect 14464 11552 14516 11558
rect 14464 11494 14516 11500
rect 14372 11348 14424 11354
rect 14372 11290 14424 11296
rect 14280 10192 14332 10198
rect 14280 10134 14332 10140
rect 14188 10124 14240 10130
rect 14188 10066 14240 10072
rect 14016 9982 14136 10010
rect 14004 9920 14056 9926
rect 14004 9862 14056 9868
rect 13556 9676 13860 9704
rect 13452 9172 13504 9178
rect 13452 9114 13504 9120
rect 13360 8968 13412 8974
rect 13360 8910 13412 8916
rect 13372 8838 13400 8910
rect 13464 8906 13492 9114
rect 13556 9081 13584 9676
rect 14016 9625 14044 9862
rect 14002 9616 14058 9625
rect 14002 9551 14058 9560
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 13740 9217 13768 9318
rect 13726 9208 13782 9217
rect 13726 9143 13782 9152
rect 13912 9172 13964 9178
rect 13912 9114 13964 9120
rect 13542 9072 13598 9081
rect 13542 9007 13598 9016
rect 13820 8968 13872 8974
rect 13924 8945 13952 9114
rect 13820 8910 13872 8916
rect 13910 8936 13966 8945
rect 13452 8900 13504 8906
rect 13452 8842 13504 8848
rect 13188 8758 13308 8786
rect 13360 8832 13412 8838
rect 13360 8774 13412 8780
rect 13188 7954 13216 8758
rect 13449 8732 13745 8752
rect 13505 8730 13529 8732
rect 13585 8730 13609 8732
rect 13665 8730 13689 8732
rect 13527 8678 13529 8730
rect 13591 8678 13603 8730
rect 13665 8678 13667 8730
rect 13505 8676 13529 8678
rect 13585 8676 13609 8678
rect 13665 8676 13689 8678
rect 13449 8656 13745 8676
rect 13360 8560 13412 8566
rect 13360 8502 13412 8508
rect 13544 8560 13596 8566
rect 13544 8502 13596 8508
rect 13372 8401 13400 8502
rect 13556 8430 13584 8502
rect 13832 8498 13860 8910
rect 13910 8871 13966 8880
rect 13912 8628 13964 8634
rect 13912 8570 13964 8576
rect 13636 8492 13688 8498
rect 13636 8434 13688 8440
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 13544 8424 13596 8430
rect 13358 8392 13414 8401
rect 13544 8366 13596 8372
rect 13358 8327 13414 8336
rect 13452 8356 13504 8362
rect 13452 8298 13504 8304
rect 13268 8288 13320 8294
rect 13266 8256 13268 8265
rect 13320 8256 13322 8265
rect 13464 8242 13492 8298
rect 13266 8191 13322 8200
rect 13372 8214 13492 8242
rect 13084 7948 13136 7954
rect 13084 7890 13136 7896
rect 13176 7948 13228 7954
rect 13176 7890 13228 7896
rect 12992 7744 13044 7750
rect 12992 7686 13044 7692
rect 13084 7744 13136 7750
rect 13084 7686 13136 7692
rect 13096 7585 13124 7686
rect 13082 7576 13138 7585
rect 13082 7511 13138 7520
rect 12992 7472 13044 7478
rect 12992 7414 13044 7420
rect 13082 7440 13138 7449
rect 12900 7336 12952 7342
rect 12900 7278 12952 7284
rect 13004 7290 13032 7414
rect 13138 7384 13308 7392
rect 13082 7375 13084 7384
rect 13136 7364 13308 7384
rect 13084 7346 13136 7352
rect 13004 7262 13124 7290
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 12992 7200 13044 7206
rect 12992 7142 13044 7148
rect 12728 7002 12848 7018
rect 12622 6967 12678 6976
rect 12716 6996 12848 7002
rect 12768 6990 12848 6996
rect 12716 6938 12768 6944
rect 12808 6860 12860 6866
rect 12808 6802 12860 6808
rect 12624 6792 12676 6798
rect 12624 6734 12676 6740
rect 12636 6390 12664 6734
rect 12624 6384 12676 6390
rect 12624 6326 12676 6332
rect 12716 6316 12768 6322
rect 12716 6258 12768 6264
rect 12624 6248 12676 6254
rect 12624 6190 12676 6196
rect 12636 5914 12664 6190
rect 12728 5953 12756 6258
rect 12820 6118 12848 6802
rect 12808 6112 12860 6118
rect 12808 6054 12860 6060
rect 12714 5944 12770 5953
rect 12624 5908 12676 5914
rect 12714 5879 12770 5888
rect 12624 5850 12676 5856
rect 12820 5846 12848 6054
rect 12716 5840 12768 5846
rect 12714 5808 12716 5817
rect 12808 5840 12860 5846
rect 12768 5808 12770 5817
rect 12808 5782 12860 5788
rect 12714 5743 12770 5752
rect 12716 5704 12768 5710
rect 12716 5646 12768 5652
rect 12728 5370 12756 5646
rect 12716 5364 12768 5370
rect 12636 5324 12716 5352
rect 12438 4247 12494 4256
rect 12532 4276 12584 4282
rect 12452 4162 12480 4247
rect 12532 4218 12584 4224
rect 12452 4134 12572 4162
rect 12440 4072 12492 4078
rect 12440 4014 12492 4020
rect 12348 4004 12400 4010
rect 12348 3946 12400 3952
rect 12346 3904 12402 3913
rect 12346 3839 12402 3848
rect 12256 3732 12308 3738
rect 12256 3674 12308 3680
rect 12256 3596 12308 3602
rect 12256 3538 12308 3544
rect 12164 1964 12216 1970
rect 12164 1906 12216 1912
rect 12268 1494 12296 3538
rect 12360 3194 12388 3839
rect 12452 3670 12480 4014
rect 12440 3664 12492 3670
rect 12440 3606 12492 3612
rect 12440 3528 12492 3534
rect 12438 3496 12440 3505
rect 12492 3496 12494 3505
rect 12438 3431 12494 3440
rect 12348 3188 12400 3194
rect 12348 3130 12400 3136
rect 12348 3052 12400 3058
rect 12348 2994 12400 3000
rect 12360 2514 12388 2994
rect 12440 2984 12492 2990
rect 12440 2926 12492 2932
rect 12348 2508 12400 2514
rect 12348 2450 12400 2456
rect 12348 2304 12400 2310
rect 12348 2246 12400 2252
rect 12360 2038 12388 2246
rect 12348 2032 12400 2038
rect 12348 1974 12400 1980
rect 12256 1488 12308 1494
rect 12256 1430 12308 1436
rect 12452 800 12480 2926
rect 12544 2650 12572 4134
rect 12636 3505 12664 5324
rect 12716 5306 12768 5312
rect 12808 5296 12860 5302
rect 12912 5284 12940 7142
rect 13004 6633 13032 7142
rect 12990 6624 13046 6633
rect 12990 6559 13046 6568
rect 12992 6452 13044 6458
rect 12992 6394 13044 6400
rect 13004 6254 13032 6394
rect 13096 6322 13124 7262
rect 13176 6996 13228 7002
rect 13176 6938 13228 6944
rect 13084 6316 13136 6322
rect 13084 6258 13136 6264
rect 12992 6248 13044 6254
rect 12992 6190 13044 6196
rect 12992 5840 13044 5846
rect 12992 5782 13044 5788
rect 12860 5256 12940 5284
rect 12808 5238 12860 5244
rect 12716 5228 12768 5234
rect 12716 5170 12768 5176
rect 12728 4146 12756 5170
rect 13004 5098 13032 5782
rect 13082 5536 13138 5545
rect 13082 5471 13138 5480
rect 13096 5370 13124 5471
rect 13084 5364 13136 5370
rect 13084 5306 13136 5312
rect 13188 5137 13216 6938
rect 13280 6798 13308 7364
rect 13268 6792 13320 6798
rect 13268 6734 13320 6740
rect 13372 6474 13400 8214
rect 13648 7886 13676 8434
rect 13728 8288 13780 8294
rect 13728 8230 13780 8236
rect 13740 8022 13768 8230
rect 13728 8016 13780 8022
rect 13728 7958 13780 7964
rect 13820 7948 13872 7954
rect 13820 7890 13872 7896
rect 13636 7880 13688 7886
rect 13636 7822 13688 7828
rect 13449 7644 13745 7664
rect 13505 7642 13529 7644
rect 13585 7642 13609 7644
rect 13665 7642 13689 7644
rect 13527 7590 13529 7642
rect 13591 7590 13603 7642
rect 13665 7590 13667 7642
rect 13505 7588 13529 7590
rect 13585 7588 13609 7590
rect 13665 7588 13689 7590
rect 13449 7568 13745 7588
rect 13832 7528 13860 7890
rect 13740 7500 13860 7528
rect 13740 7018 13768 7500
rect 13820 7200 13872 7206
rect 13818 7168 13820 7177
rect 13872 7168 13874 7177
rect 13818 7103 13874 7112
rect 13740 6990 13860 7018
rect 13449 6556 13745 6576
rect 13505 6554 13529 6556
rect 13585 6554 13609 6556
rect 13665 6554 13689 6556
rect 13527 6502 13529 6554
rect 13591 6502 13603 6554
rect 13665 6502 13667 6554
rect 13505 6500 13529 6502
rect 13585 6500 13609 6502
rect 13665 6500 13689 6502
rect 13449 6480 13745 6500
rect 13280 6446 13400 6474
rect 13174 5128 13230 5137
rect 12992 5092 13044 5098
rect 13174 5063 13230 5072
rect 12992 5034 13044 5040
rect 13084 5024 13136 5030
rect 12806 4992 12862 5001
rect 12806 4927 12862 4936
rect 13082 4992 13084 5001
rect 13280 5012 13308 6446
rect 13358 6216 13414 6225
rect 13358 6151 13414 6160
rect 13544 6180 13596 6186
rect 13372 6118 13400 6151
rect 13544 6122 13596 6128
rect 13636 6180 13688 6186
rect 13636 6122 13688 6128
rect 13360 6112 13412 6118
rect 13360 6054 13412 6060
rect 13556 5846 13584 6122
rect 13648 6089 13676 6122
rect 13832 6118 13860 6990
rect 13820 6112 13872 6118
rect 13634 6080 13690 6089
rect 13820 6054 13872 6060
rect 13634 6015 13690 6024
rect 13544 5840 13596 5846
rect 13372 5800 13544 5828
rect 13372 5574 13400 5800
rect 13544 5782 13596 5788
rect 13360 5568 13412 5574
rect 13360 5510 13412 5516
rect 13136 4992 13138 5001
rect 13082 4927 13138 4936
rect 13188 4984 13308 5012
rect 12820 4282 12848 4927
rect 13096 4826 13124 4927
rect 13084 4820 13136 4826
rect 13084 4762 13136 4768
rect 13084 4684 13136 4690
rect 13084 4626 13136 4632
rect 12992 4548 13044 4554
rect 12992 4490 13044 4496
rect 12900 4480 12952 4486
rect 12900 4422 12952 4428
rect 12808 4276 12860 4282
rect 12808 4218 12860 4224
rect 12716 4140 12768 4146
rect 12716 4082 12768 4088
rect 12808 4004 12860 4010
rect 12808 3946 12860 3952
rect 12622 3496 12678 3505
rect 12622 3431 12678 3440
rect 12624 3392 12676 3398
rect 12624 3334 12676 3340
rect 12636 2854 12664 3334
rect 12716 3188 12768 3194
rect 12716 3130 12768 3136
rect 12624 2848 12676 2854
rect 12624 2790 12676 2796
rect 12532 2644 12584 2650
rect 12532 2586 12584 2592
rect 12728 1873 12756 3130
rect 12820 3108 12848 3946
rect 12912 3398 12940 4422
rect 13004 4214 13032 4490
rect 12992 4208 13044 4214
rect 12992 4150 13044 4156
rect 12990 4040 13046 4049
rect 12990 3975 12992 3984
rect 13044 3975 13046 3984
rect 12992 3946 13044 3952
rect 13096 3738 13124 4626
rect 13084 3732 13136 3738
rect 13084 3674 13136 3680
rect 12992 3528 13044 3534
rect 12992 3470 13044 3476
rect 12900 3392 12952 3398
rect 12900 3334 12952 3340
rect 12912 3233 12940 3334
rect 12898 3224 12954 3233
rect 12898 3159 12954 3168
rect 12820 3080 12940 3108
rect 12808 2848 12860 2854
rect 12808 2790 12860 2796
rect 12820 2514 12848 2790
rect 12808 2508 12860 2514
rect 12808 2450 12860 2456
rect 12714 1864 12770 1873
rect 12714 1799 12770 1808
rect 12820 800 12848 2450
rect 12912 1834 12940 3080
rect 13004 1902 13032 3470
rect 13084 3392 13136 3398
rect 13188 3380 13216 4984
rect 13268 4820 13320 4826
rect 13268 4762 13320 4768
rect 13280 3670 13308 4762
rect 13372 4282 13400 5510
rect 13449 5468 13745 5488
rect 13505 5466 13529 5468
rect 13585 5466 13609 5468
rect 13665 5466 13689 5468
rect 13527 5414 13529 5466
rect 13591 5414 13603 5466
rect 13665 5414 13667 5466
rect 13505 5412 13529 5414
rect 13585 5412 13609 5414
rect 13665 5412 13689 5414
rect 13449 5392 13745 5412
rect 13452 5296 13504 5302
rect 13544 5296 13596 5302
rect 13452 5238 13504 5244
rect 13542 5264 13544 5273
rect 13596 5264 13598 5273
rect 13464 4826 13492 5238
rect 13542 5199 13598 5208
rect 13636 5024 13688 5030
rect 13636 4966 13688 4972
rect 13648 4865 13676 4966
rect 13634 4856 13690 4865
rect 13452 4820 13504 4826
rect 13634 4791 13690 4800
rect 13452 4762 13504 4768
rect 13634 4720 13690 4729
rect 13634 4655 13636 4664
rect 13688 4655 13690 4664
rect 13636 4626 13688 4632
rect 13449 4380 13745 4400
rect 13505 4378 13529 4380
rect 13585 4378 13609 4380
rect 13665 4378 13689 4380
rect 13527 4326 13529 4378
rect 13591 4326 13603 4378
rect 13665 4326 13667 4378
rect 13505 4324 13529 4326
rect 13585 4324 13609 4326
rect 13665 4324 13689 4326
rect 13449 4304 13745 4324
rect 13360 4276 13412 4282
rect 13832 4264 13860 6054
rect 13360 4218 13412 4224
rect 13740 4236 13860 4264
rect 13740 4185 13768 4236
rect 13726 4176 13782 4185
rect 13726 4111 13782 4120
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 13268 3664 13320 3670
rect 13268 3606 13320 3612
rect 13358 3632 13414 3641
rect 13832 3602 13860 4082
rect 13924 3652 13952 8570
rect 14016 8430 14044 9551
rect 14108 8945 14136 9982
rect 14094 8936 14150 8945
rect 14094 8871 14150 8880
rect 14096 8832 14148 8838
rect 14096 8774 14148 8780
rect 14004 8424 14056 8430
rect 14004 8366 14056 8372
rect 14016 7546 14044 8366
rect 14108 8362 14136 8774
rect 14096 8356 14148 8362
rect 14096 8298 14148 8304
rect 14200 7954 14228 10066
rect 14370 10024 14426 10033
rect 14370 9959 14372 9968
rect 14424 9959 14426 9968
rect 14372 9930 14424 9936
rect 14280 9580 14332 9586
rect 14280 9522 14332 9528
rect 14292 8498 14320 9522
rect 14476 9382 14504 11494
rect 14556 11076 14608 11082
rect 14556 11018 14608 11024
rect 14568 10470 14596 11018
rect 14556 10464 14608 10470
rect 14556 10406 14608 10412
rect 14464 9376 14516 9382
rect 14464 9318 14516 9324
rect 14372 8900 14424 8906
rect 14372 8842 14424 8848
rect 14280 8492 14332 8498
rect 14280 8434 14332 8440
rect 14280 8356 14332 8362
rect 14280 8298 14332 8304
rect 14292 8129 14320 8298
rect 14278 8120 14334 8129
rect 14278 8055 14334 8064
rect 14188 7948 14240 7954
rect 14188 7890 14240 7896
rect 14096 7812 14148 7818
rect 14096 7754 14148 7760
rect 14004 7540 14056 7546
rect 14004 7482 14056 7488
rect 14004 7336 14056 7342
rect 14004 7278 14056 7284
rect 14016 5574 14044 7278
rect 14108 7002 14136 7754
rect 14188 7744 14240 7750
rect 14292 7732 14320 8055
rect 14240 7704 14320 7732
rect 14188 7686 14240 7692
rect 14096 6996 14148 7002
rect 14096 6938 14148 6944
rect 14108 6769 14136 6938
rect 14094 6760 14150 6769
rect 14094 6695 14150 6704
rect 14108 5914 14136 6695
rect 14096 5908 14148 5914
rect 14096 5850 14148 5856
rect 14004 5568 14056 5574
rect 14004 5510 14056 5516
rect 14016 5030 14044 5510
rect 14096 5160 14148 5166
rect 14096 5102 14148 5108
rect 14004 5024 14056 5030
rect 14004 4966 14056 4972
rect 14004 4684 14056 4690
rect 14004 4626 14056 4632
rect 14016 4282 14044 4626
rect 14004 4276 14056 4282
rect 14004 4218 14056 4224
rect 14004 3664 14056 3670
rect 13924 3624 14004 3652
rect 14004 3606 14056 3612
rect 13358 3567 13360 3576
rect 13412 3567 13414 3576
rect 13820 3596 13872 3602
rect 13360 3538 13412 3544
rect 13820 3538 13872 3544
rect 13136 3352 13216 3380
rect 13084 3334 13136 3340
rect 13096 2145 13124 3334
rect 13449 3292 13745 3312
rect 13505 3290 13529 3292
rect 13585 3290 13609 3292
rect 13665 3290 13689 3292
rect 13527 3238 13529 3290
rect 13591 3238 13603 3290
rect 13665 3238 13667 3290
rect 13505 3236 13529 3238
rect 13585 3236 13609 3238
rect 13665 3236 13689 3238
rect 13449 3216 13745 3236
rect 13832 3126 13860 3538
rect 14108 3194 14136 5102
rect 14096 3188 14148 3194
rect 14016 3148 14096 3176
rect 13820 3120 13872 3126
rect 13820 3062 13872 3068
rect 13176 2984 13228 2990
rect 13176 2926 13228 2932
rect 13188 2514 13216 2926
rect 13452 2916 13504 2922
rect 13452 2858 13504 2864
rect 13464 2514 13492 2858
rect 13820 2848 13872 2854
rect 13820 2790 13872 2796
rect 13832 2514 13860 2790
rect 14016 2514 14044 3148
rect 14096 3130 14148 3136
rect 14200 3074 14228 7686
rect 14280 7540 14332 7546
rect 14280 7482 14332 7488
rect 14292 6662 14320 7482
rect 14384 7206 14412 8842
rect 14476 7274 14504 9318
rect 14464 7268 14516 7274
rect 14464 7210 14516 7216
rect 14372 7200 14424 7206
rect 14372 7142 14424 7148
rect 14384 6905 14412 7142
rect 14370 6896 14426 6905
rect 14370 6831 14426 6840
rect 14280 6656 14332 6662
rect 14280 6598 14332 6604
rect 14292 4554 14320 6598
rect 14370 6352 14426 6361
rect 14370 6287 14372 6296
rect 14424 6287 14426 6296
rect 14372 6258 14424 6264
rect 14280 4548 14332 4554
rect 14280 4490 14332 4496
rect 14384 4214 14412 6258
rect 14464 5296 14516 5302
rect 14568 5284 14596 10406
rect 14660 7342 14688 11562
rect 14752 11354 14780 11630
rect 14740 11348 14792 11354
rect 14740 11290 14792 11296
rect 14740 11212 14792 11218
rect 14740 11154 14792 11160
rect 14752 10674 14780 11154
rect 14740 10668 14792 10674
rect 14792 10628 14872 10656
rect 14740 10610 14792 10616
rect 14844 10062 14872 10628
rect 14832 10056 14884 10062
rect 14832 9998 14884 10004
rect 14740 9376 14792 9382
rect 14740 9318 14792 9324
rect 14752 9178 14780 9318
rect 14740 9172 14792 9178
rect 14740 9114 14792 9120
rect 14832 8968 14884 8974
rect 14832 8910 14884 8916
rect 14844 8634 14872 8910
rect 14832 8628 14884 8634
rect 14832 8570 14884 8576
rect 14832 8288 14884 8294
rect 14936 8276 14964 11750
rect 14884 8248 14964 8276
rect 14832 8230 14884 8236
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 14752 7546 14780 7686
rect 14740 7540 14792 7546
rect 14740 7482 14792 7488
rect 14648 7336 14700 7342
rect 14648 7278 14700 7284
rect 14738 7032 14794 7041
rect 14738 6967 14794 6976
rect 14752 6662 14780 6967
rect 14740 6656 14792 6662
rect 14740 6598 14792 6604
rect 14516 5256 14596 5284
rect 14464 5238 14516 5244
rect 14476 4282 14504 5238
rect 14752 4826 14780 6598
rect 14844 5234 14872 8230
rect 15028 8022 15056 11852
rect 15120 11014 15148 16458
rect 15212 15638 15240 16646
rect 15200 15632 15252 15638
rect 15200 15574 15252 15580
rect 15304 11354 15332 17002
rect 15488 16658 15516 19200
rect 15658 16688 15714 16697
rect 15476 16652 15528 16658
rect 15658 16623 15660 16632
rect 15476 16594 15528 16600
rect 15712 16623 15714 16632
rect 15660 16594 15712 16600
rect 15384 15904 15436 15910
rect 15384 15846 15436 15852
rect 15396 15570 15424 15846
rect 15384 15564 15436 15570
rect 15384 15506 15436 15512
rect 15488 15502 15516 16594
rect 15856 16046 15884 19200
rect 16224 16794 16252 19200
rect 16592 16998 16620 19200
rect 16580 16992 16632 16998
rect 16580 16934 16632 16940
rect 16212 16788 16264 16794
rect 16212 16730 16264 16736
rect 15844 16040 15896 16046
rect 15844 15982 15896 15988
rect 15856 15706 15884 15982
rect 16960 15978 16988 19200
rect 16948 15972 17000 15978
rect 16948 15914 17000 15920
rect 15844 15700 15896 15706
rect 15844 15642 15896 15648
rect 15476 15496 15528 15502
rect 15476 15438 15528 15444
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 15108 11008 15160 11014
rect 15108 10950 15160 10956
rect 15108 9512 15160 9518
rect 15108 9454 15160 9460
rect 15120 9382 15148 9454
rect 15108 9376 15160 9382
rect 15106 9344 15108 9353
rect 15160 9344 15162 9353
rect 15106 9279 15162 9288
rect 15016 8016 15068 8022
rect 15016 7958 15068 7964
rect 14924 7744 14976 7750
rect 14924 7686 14976 7692
rect 14936 6934 14964 7686
rect 14924 6928 14976 6934
rect 14924 6870 14976 6876
rect 14832 5228 14884 5234
rect 14832 5170 14884 5176
rect 14740 4820 14792 4826
rect 14740 4762 14792 4768
rect 15016 4752 15068 4758
rect 15016 4694 15068 4700
rect 14556 4616 14608 4622
rect 14556 4558 14608 4564
rect 14464 4276 14516 4282
rect 14464 4218 14516 4224
rect 14372 4208 14424 4214
rect 14372 4150 14424 4156
rect 14464 3596 14516 3602
rect 14464 3538 14516 3544
rect 14476 3398 14504 3538
rect 14568 3466 14596 4558
rect 14648 3732 14700 3738
rect 14648 3674 14700 3680
rect 14556 3460 14608 3466
rect 14556 3402 14608 3408
rect 14464 3392 14516 3398
rect 14464 3334 14516 3340
rect 14108 3046 14228 3074
rect 14108 2650 14136 3046
rect 14188 2916 14240 2922
rect 14188 2858 14240 2864
rect 14096 2644 14148 2650
rect 14096 2586 14148 2592
rect 13176 2508 13228 2514
rect 13452 2508 13504 2514
rect 13176 2450 13228 2456
rect 13372 2468 13452 2496
rect 13082 2136 13138 2145
rect 13082 2071 13138 2080
rect 12992 1896 13044 1902
rect 12992 1838 13044 1844
rect 12900 1828 12952 1834
rect 12900 1770 12952 1776
rect 13188 800 13216 2450
rect 13372 1986 13400 2468
rect 13452 2450 13504 2456
rect 13820 2508 13872 2514
rect 13820 2450 13872 2456
rect 14004 2508 14056 2514
rect 14004 2450 14056 2456
rect 13449 2204 13745 2224
rect 13505 2202 13529 2204
rect 13585 2202 13609 2204
rect 13665 2202 13689 2204
rect 13527 2150 13529 2202
rect 13591 2150 13603 2202
rect 13665 2150 13667 2202
rect 13505 2148 13529 2150
rect 13585 2148 13609 2150
rect 13665 2148 13689 2150
rect 13449 2128 13745 2148
rect 13372 1958 13492 1986
rect 13464 800 13492 1958
rect 13832 800 13860 2450
rect 14200 800 14228 2858
rect 14476 2360 14504 3334
rect 14568 3058 14596 3402
rect 14556 3052 14608 3058
rect 14556 2994 14608 3000
rect 14660 2990 14688 3674
rect 14832 3596 14884 3602
rect 14832 3538 14884 3544
rect 14648 2984 14700 2990
rect 14648 2926 14700 2932
rect 14556 2848 14608 2854
rect 14556 2790 14608 2796
rect 14568 2514 14596 2790
rect 14556 2508 14608 2514
rect 14556 2450 14608 2456
rect 14476 2332 14596 2360
rect 14568 800 14596 2332
rect 14844 800 14872 3538
rect 15028 3466 15056 4694
rect 15120 4026 15148 9279
rect 15200 9036 15252 9042
rect 15200 8978 15252 8984
rect 15212 8537 15240 8978
rect 15198 8528 15254 8537
rect 15198 8463 15200 8472
rect 15252 8463 15254 8472
rect 15200 8434 15252 8440
rect 15212 5846 15240 8434
rect 15200 5840 15252 5846
rect 15200 5782 15252 5788
rect 15304 4146 15332 11290
rect 15476 10124 15528 10130
rect 15476 10066 15528 10072
rect 15488 9722 15516 10066
rect 15658 10024 15714 10033
rect 15658 9959 15660 9968
rect 15712 9959 15714 9968
rect 15660 9930 15712 9936
rect 15476 9716 15528 9722
rect 15476 9658 15528 9664
rect 15474 9480 15530 9489
rect 15474 9415 15476 9424
rect 15528 9415 15530 9424
rect 15476 9386 15528 9392
rect 15292 4140 15344 4146
rect 15292 4082 15344 4088
rect 15120 3998 15240 4026
rect 15108 3936 15160 3942
rect 15108 3878 15160 3884
rect 15120 3602 15148 3878
rect 15108 3596 15160 3602
rect 15108 3538 15160 3544
rect 15212 3482 15240 3998
rect 15292 3936 15344 3942
rect 15292 3878 15344 3884
rect 16212 3936 16264 3942
rect 16212 3878 16264 3884
rect 15304 3602 15332 3878
rect 15292 3596 15344 3602
rect 15292 3538 15344 3544
rect 15016 3460 15068 3466
rect 15016 3402 15068 3408
rect 15120 3454 15240 3482
rect 15028 2990 15056 3402
rect 15016 2984 15068 2990
rect 15016 2926 15068 2932
rect 14924 2848 14976 2854
rect 14924 2790 14976 2796
rect 14936 2582 14964 2790
rect 14924 2576 14976 2582
rect 14924 2518 14976 2524
rect 15120 2378 15148 3454
rect 15304 2774 15332 3538
rect 15660 3460 15712 3466
rect 15660 3402 15712 3408
rect 15672 3369 15700 3402
rect 15658 3360 15714 3369
rect 15658 3295 15714 3304
rect 15212 2746 15332 2774
rect 15108 2372 15160 2378
rect 15108 2314 15160 2320
rect 15212 800 15240 2746
rect 15936 2372 15988 2378
rect 15936 2314 15988 2320
rect 15568 2304 15620 2310
rect 15568 2246 15620 2252
rect 15580 800 15608 2246
rect 15948 800 15976 2314
rect 16224 800 16252 3878
rect 16948 2916 17000 2922
rect 16948 2858 17000 2864
rect 16580 2440 16632 2446
rect 16580 2382 16632 2388
rect 16592 800 16620 2382
rect 16960 800 16988 2858
rect 1674 504 1730 513
rect 1674 439 1730 448
rect 1766 0 1822 800
rect 2134 0 2190 800
rect 2502 0 2558 800
rect 2778 0 2834 800
rect 3146 0 3202 800
rect 3514 0 3570 800
rect 3882 0 3938 800
rect 4158 0 4214 800
rect 4526 0 4582 800
rect 4894 0 4950 800
rect 5262 0 5318 800
rect 5538 0 5594 800
rect 5906 0 5962 800
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 6918 0 6974 800
rect 7286 0 7342 800
rect 7654 0 7710 800
rect 8022 0 8078 800
rect 8298 0 8354 800
rect 8666 0 8722 800
rect 9034 0 9090 800
rect 9310 0 9366 800
rect 9678 0 9734 800
rect 10046 0 10102 800
rect 10414 0 10470 800
rect 10690 0 10746 800
rect 11058 0 11114 800
rect 11426 0 11482 800
rect 11794 0 11850 800
rect 12070 0 12126 800
rect 12438 0 12494 800
rect 12806 0 12862 800
rect 13174 0 13230 800
rect 13450 0 13506 800
rect 13818 0 13874 800
rect 14186 0 14242 800
rect 14554 0 14610 800
rect 14830 0 14886 800
rect 15198 0 15254 800
rect 15566 0 15622 800
rect 15934 0 15990 800
rect 16210 0 16266 800
rect 16578 0 16634 800
rect 16946 0 17002 800
<< via2 >>
rect 1398 19352 1454 19408
rect 1950 17312 2006 17368
rect 1490 16360 1546 16416
rect 2778 18400 2834 18456
rect 3454 17434 3510 17436
rect 3534 17434 3590 17436
rect 3614 17434 3670 17436
rect 3694 17434 3750 17436
rect 3454 17382 3480 17434
rect 3480 17382 3510 17434
rect 3534 17382 3544 17434
rect 3544 17382 3590 17434
rect 3614 17382 3660 17434
rect 3660 17382 3670 17434
rect 3694 17382 3724 17434
rect 3724 17382 3750 17434
rect 3454 17380 3510 17382
rect 3534 17380 3590 17382
rect 3614 17380 3670 17382
rect 3694 17380 3750 17382
rect 1398 15428 1454 15464
rect 1398 15408 1400 15428
rect 1400 15408 1452 15428
rect 1452 15408 1454 15428
rect 1398 14340 1454 14376
rect 1398 14320 1400 14340
rect 1400 14320 1452 14340
rect 1452 14320 1454 14340
rect 1398 13388 1454 13424
rect 1398 13368 1400 13388
rect 1400 13368 1452 13388
rect 1452 13368 1454 13388
rect 1398 12416 1454 12472
rect 2410 12552 2466 12608
rect 1950 11620 2006 11656
rect 1950 11600 1952 11620
rect 1952 11600 2004 11620
rect 2004 11600 2006 11620
rect 2410 11736 2466 11792
rect 3146 13368 3202 13424
rect 1490 11348 1546 11384
rect 1490 11328 1492 11348
rect 1492 11328 1544 11348
rect 1544 11328 1546 11348
rect 1490 10412 1492 10432
rect 1492 10412 1544 10432
rect 1544 10412 1546 10432
rect 1490 10376 1546 10412
rect 1398 9460 1400 9480
rect 1400 9460 1452 9480
rect 1452 9460 1454 9480
rect 1398 9424 1454 9460
rect 1490 9288 1546 9344
rect 1398 8356 1454 8392
rect 1398 8336 1400 8356
rect 1400 8336 1452 8356
rect 1452 8336 1454 8356
rect 1398 7404 1454 7440
rect 1398 7384 1400 7404
rect 1400 7384 1452 7404
rect 1452 7384 1454 7404
rect 1490 6452 1546 6488
rect 1490 6432 1492 6452
rect 1492 6432 1544 6452
rect 1544 6432 1546 6452
rect 1490 5364 1546 5400
rect 1490 5344 1492 5364
rect 1492 5344 1544 5364
rect 1544 5344 1546 5364
rect 1490 4428 1492 4448
rect 1492 4428 1544 4448
rect 1544 4428 1546 4448
rect 1490 4392 1546 4428
rect 1490 2352 1546 2408
rect 2226 9968 2282 10024
rect 2686 10512 2742 10568
rect 2594 9424 2650 9480
rect 2502 9152 2558 9208
rect 2410 9036 2466 9072
rect 2410 9016 2412 9036
rect 2412 9016 2464 9036
rect 2464 9016 2466 9036
rect 2870 12280 2926 12336
rect 3882 16360 3938 16416
rect 3454 16346 3510 16348
rect 3534 16346 3590 16348
rect 3614 16346 3670 16348
rect 3694 16346 3750 16348
rect 3454 16294 3480 16346
rect 3480 16294 3510 16346
rect 3534 16294 3544 16346
rect 3544 16294 3590 16346
rect 3614 16294 3660 16346
rect 3660 16294 3670 16346
rect 3694 16294 3724 16346
rect 3724 16294 3750 16346
rect 3454 16292 3510 16294
rect 3534 16292 3590 16294
rect 3614 16292 3670 16294
rect 3694 16292 3750 16294
rect 3454 15258 3510 15260
rect 3534 15258 3590 15260
rect 3614 15258 3670 15260
rect 3694 15258 3750 15260
rect 3454 15206 3480 15258
rect 3480 15206 3510 15258
rect 3534 15206 3544 15258
rect 3544 15206 3590 15258
rect 3614 15206 3660 15258
rect 3660 15206 3670 15258
rect 3694 15206 3724 15258
rect 3724 15206 3750 15258
rect 3454 15204 3510 15206
rect 3534 15204 3590 15206
rect 3614 15204 3670 15206
rect 3694 15204 3750 15206
rect 3238 12280 3294 12336
rect 3238 12180 3240 12200
rect 3240 12180 3292 12200
rect 3292 12180 3294 12200
rect 3238 12144 3294 12180
rect 3454 14170 3510 14172
rect 3534 14170 3590 14172
rect 3614 14170 3670 14172
rect 3694 14170 3750 14172
rect 3454 14118 3480 14170
rect 3480 14118 3510 14170
rect 3534 14118 3544 14170
rect 3544 14118 3590 14170
rect 3614 14118 3660 14170
rect 3660 14118 3670 14170
rect 3694 14118 3724 14170
rect 3724 14118 3750 14170
rect 3454 14116 3510 14118
rect 3534 14116 3590 14118
rect 3614 14116 3670 14118
rect 3694 14116 3750 14118
rect 3422 13776 3478 13832
rect 3454 13082 3510 13084
rect 3534 13082 3590 13084
rect 3614 13082 3670 13084
rect 3694 13082 3750 13084
rect 3454 13030 3480 13082
rect 3480 13030 3510 13082
rect 3534 13030 3544 13082
rect 3544 13030 3590 13082
rect 3614 13030 3660 13082
rect 3660 13030 3670 13082
rect 3694 13030 3724 13082
rect 3724 13030 3750 13082
rect 3454 13028 3510 13030
rect 3534 13028 3590 13030
rect 3614 13028 3670 13030
rect 3694 13028 3750 13030
rect 3514 12824 3570 12880
rect 3454 11994 3510 11996
rect 3534 11994 3590 11996
rect 3614 11994 3670 11996
rect 3694 11994 3750 11996
rect 3454 11942 3480 11994
rect 3480 11942 3510 11994
rect 3534 11942 3544 11994
rect 3544 11942 3590 11994
rect 3614 11942 3660 11994
rect 3660 11942 3670 11994
rect 3694 11942 3724 11994
rect 3724 11942 3750 11994
rect 3454 11940 3510 11942
rect 3534 11940 3590 11942
rect 3614 11940 3670 11942
rect 3694 11940 3750 11942
rect 8452 17434 8508 17436
rect 8532 17434 8588 17436
rect 8612 17434 8668 17436
rect 8692 17434 8748 17436
rect 8452 17382 8478 17434
rect 8478 17382 8508 17434
rect 8532 17382 8542 17434
rect 8542 17382 8588 17434
rect 8612 17382 8658 17434
rect 8658 17382 8668 17434
rect 8692 17382 8722 17434
rect 8722 17382 8748 17434
rect 8452 17380 8508 17382
rect 8532 17380 8588 17382
rect 8612 17380 8668 17382
rect 8692 17380 8748 17382
rect 5953 16890 6009 16892
rect 6033 16890 6089 16892
rect 6113 16890 6169 16892
rect 6193 16890 6249 16892
rect 5953 16838 5979 16890
rect 5979 16838 6009 16890
rect 6033 16838 6043 16890
rect 6043 16838 6089 16890
rect 6113 16838 6159 16890
rect 6159 16838 6169 16890
rect 6193 16838 6223 16890
rect 6223 16838 6249 16890
rect 5953 16836 6009 16838
rect 6033 16836 6089 16838
rect 6113 16836 6169 16838
rect 6193 16836 6249 16838
rect 5953 15802 6009 15804
rect 6033 15802 6089 15804
rect 6113 15802 6169 15804
rect 6193 15802 6249 15804
rect 5953 15750 5979 15802
rect 5979 15750 6009 15802
rect 6033 15750 6043 15802
rect 6043 15750 6089 15802
rect 6113 15750 6159 15802
rect 6159 15750 6169 15802
rect 6193 15750 6223 15802
rect 6223 15750 6249 15802
rect 5953 15748 6009 15750
rect 6033 15748 6089 15750
rect 6113 15748 6169 15750
rect 6193 15748 6249 15750
rect 4618 15000 4674 15056
rect 4066 13096 4122 13152
rect 3454 10906 3510 10908
rect 3534 10906 3590 10908
rect 3614 10906 3670 10908
rect 3694 10906 3750 10908
rect 3454 10854 3480 10906
rect 3480 10854 3510 10906
rect 3534 10854 3544 10906
rect 3544 10854 3590 10906
rect 3614 10854 3660 10906
rect 3660 10854 3670 10906
rect 3694 10854 3724 10906
rect 3724 10854 3750 10906
rect 3454 10852 3510 10854
rect 3534 10852 3590 10854
rect 3614 10852 3670 10854
rect 3694 10852 3750 10854
rect 2686 8880 2742 8936
rect 2686 8336 2742 8392
rect 2502 8200 2558 8256
rect 3054 9560 3110 9616
rect 2410 7948 2466 7984
rect 2410 7928 2412 7948
rect 2412 7928 2464 7948
rect 2464 7928 2466 7948
rect 2962 8236 2964 8256
rect 2964 8236 3016 8256
rect 3016 8236 3018 8256
rect 2962 8200 3018 8236
rect 2962 7948 3018 7984
rect 2962 7928 2964 7948
rect 2964 7928 3016 7948
rect 3016 7928 3018 7948
rect 2502 6876 2504 6896
rect 2504 6876 2556 6896
rect 2556 6876 2558 6896
rect 2502 6840 2558 6876
rect 2226 6160 2282 6216
rect 2134 6024 2190 6080
rect 2134 5888 2190 5944
rect 2410 5752 2466 5808
rect 1950 4936 2006 4992
rect 1858 3440 1914 3496
rect 2410 4020 2412 4040
rect 2412 4020 2464 4040
rect 2464 4020 2466 4040
rect 2410 3984 2466 4020
rect 2502 3848 2558 3904
rect 2226 3032 2282 3088
rect 1858 1400 1914 1456
rect 2226 2624 2282 2680
rect 2686 4800 2742 4856
rect 4066 12280 4122 12336
rect 4526 12552 4582 12608
rect 4342 11872 4398 11928
rect 4710 13232 4766 13288
rect 4802 12688 4858 12744
rect 3454 9818 3510 9820
rect 3534 9818 3590 9820
rect 3614 9818 3670 9820
rect 3694 9818 3750 9820
rect 3454 9766 3480 9818
rect 3480 9766 3510 9818
rect 3534 9766 3544 9818
rect 3544 9766 3590 9818
rect 3614 9766 3660 9818
rect 3660 9766 3670 9818
rect 3694 9766 3724 9818
rect 3724 9766 3750 9818
rect 3454 9764 3510 9766
rect 3534 9764 3590 9766
rect 3614 9764 3670 9766
rect 3694 9764 3750 9766
rect 3238 9580 3294 9616
rect 3238 9560 3240 9580
rect 3240 9560 3292 9580
rect 3292 9560 3294 9580
rect 3454 8730 3510 8732
rect 3534 8730 3590 8732
rect 3614 8730 3670 8732
rect 3694 8730 3750 8732
rect 3454 8678 3480 8730
rect 3480 8678 3510 8730
rect 3534 8678 3544 8730
rect 3544 8678 3590 8730
rect 3614 8678 3660 8730
rect 3660 8678 3670 8730
rect 3694 8678 3724 8730
rect 3724 8678 3750 8730
rect 3454 8676 3510 8678
rect 3534 8676 3590 8678
rect 3614 8676 3670 8678
rect 3694 8676 3750 8678
rect 3146 7792 3202 7848
rect 3698 7928 3754 7984
rect 3454 7642 3510 7644
rect 3534 7642 3590 7644
rect 3614 7642 3670 7644
rect 3694 7642 3750 7644
rect 3454 7590 3480 7642
rect 3480 7590 3510 7642
rect 3534 7590 3544 7642
rect 3544 7590 3590 7642
rect 3614 7590 3660 7642
rect 3660 7590 3670 7642
rect 3694 7590 3724 7642
rect 3724 7590 3750 7642
rect 3454 7588 3510 7590
rect 3534 7588 3590 7590
rect 3614 7588 3670 7590
rect 3694 7588 3750 7590
rect 2870 6704 2926 6760
rect 2778 4664 2834 4720
rect 4158 9696 4214 9752
rect 4342 10512 4398 10568
rect 3882 8472 3938 8528
rect 3882 7928 3938 7984
rect 3790 7248 3846 7304
rect 3606 7112 3662 7168
rect 3330 6976 3386 7032
rect 3882 6840 3938 6896
rect 3454 6554 3510 6556
rect 3534 6554 3590 6556
rect 3614 6554 3670 6556
rect 3694 6554 3750 6556
rect 3454 6502 3480 6554
rect 3480 6502 3510 6554
rect 3534 6502 3544 6554
rect 3544 6502 3590 6554
rect 3614 6502 3660 6554
rect 3660 6502 3670 6554
rect 3694 6502 3724 6554
rect 3724 6502 3750 6554
rect 3454 6500 3510 6502
rect 3534 6500 3590 6502
rect 3614 6500 3670 6502
rect 3694 6500 3750 6502
rect 4066 7792 4122 7848
rect 4158 7656 4214 7712
rect 4066 6840 4122 6896
rect 3882 6432 3938 6488
rect 2962 4120 3018 4176
rect 2318 2388 2320 2408
rect 2320 2388 2372 2408
rect 2372 2388 2374 2408
rect 2318 2352 2374 2388
rect 2778 3440 2834 3496
rect 2686 2624 2742 2680
rect 3146 4972 3148 4992
rect 3148 4972 3200 4992
rect 3200 4972 3202 4992
rect 3146 4936 3202 4972
rect 4526 10124 4582 10160
rect 4526 10104 4528 10124
rect 4528 10104 4580 10124
rect 4580 10104 4582 10124
rect 4342 8608 4398 8664
rect 5446 11872 5502 11928
rect 5262 11212 5318 11248
rect 5262 11192 5264 11212
rect 5264 11192 5316 11212
rect 5316 11192 5318 11212
rect 5170 11056 5226 11112
rect 5953 14714 6009 14716
rect 6033 14714 6089 14716
rect 6113 14714 6169 14716
rect 6193 14714 6249 14716
rect 5953 14662 5979 14714
rect 5979 14662 6009 14714
rect 6033 14662 6043 14714
rect 6043 14662 6089 14714
rect 6113 14662 6159 14714
rect 6159 14662 6169 14714
rect 6193 14662 6223 14714
rect 6223 14662 6249 14714
rect 5953 14660 6009 14662
rect 6033 14660 6089 14662
rect 6113 14660 6169 14662
rect 6193 14660 6249 14662
rect 5814 13912 5870 13968
rect 5953 13626 6009 13628
rect 6033 13626 6089 13628
rect 6113 13626 6169 13628
rect 6193 13626 6249 13628
rect 5953 13574 5979 13626
rect 5979 13574 6009 13626
rect 6033 13574 6043 13626
rect 6043 13574 6089 13626
rect 6113 13574 6159 13626
rect 6159 13574 6169 13626
rect 6193 13574 6223 13626
rect 6223 13574 6249 13626
rect 5953 13572 6009 13574
rect 6033 13572 6089 13574
rect 6113 13572 6169 13574
rect 6193 13572 6249 13574
rect 5722 12824 5778 12880
rect 5953 12538 6009 12540
rect 6033 12538 6089 12540
rect 6113 12538 6169 12540
rect 6193 12538 6249 12540
rect 5953 12486 5979 12538
rect 5979 12486 6009 12538
rect 6033 12486 6043 12538
rect 6043 12486 6089 12538
rect 6113 12486 6159 12538
rect 6159 12486 6169 12538
rect 6193 12486 6223 12538
rect 6223 12486 6249 12538
rect 5953 12484 6009 12486
rect 6033 12484 6089 12486
rect 6113 12484 6169 12486
rect 6193 12484 6249 12486
rect 5953 11450 6009 11452
rect 6033 11450 6089 11452
rect 6113 11450 6169 11452
rect 6193 11450 6249 11452
rect 5953 11398 5979 11450
rect 5979 11398 6009 11450
rect 6033 11398 6043 11450
rect 6043 11398 6089 11450
rect 6113 11398 6159 11450
rect 6159 11398 6169 11450
rect 6193 11398 6223 11450
rect 6223 11398 6249 11450
rect 5953 11396 6009 11398
rect 6033 11396 6089 11398
rect 6113 11396 6169 11398
rect 6193 11396 6249 11398
rect 6734 15700 6790 15736
rect 6734 15680 6736 15700
rect 6736 15680 6788 15700
rect 6788 15680 6790 15700
rect 6366 12552 6422 12608
rect 5953 10362 6009 10364
rect 6033 10362 6089 10364
rect 6113 10362 6169 10364
rect 6193 10362 6249 10364
rect 5953 10310 5979 10362
rect 5979 10310 6009 10362
rect 6033 10310 6043 10362
rect 6043 10310 6089 10362
rect 6113 10310 6159 10362
rect 6159 10310 6169 10362
rect 6193 10310 6223 10362
rect 6223 10310 6249 10362
rect 5953 10308 6009 10310
rect 6033 10308 6089 10310
rect 6113 10308 6169 10310
rect 6193 10308 6249 10310
rect 4526 7928 4582 7984
rect 4710 7928 4766 7984
rect 4158 6568 4214 6624
rect 4342 5652 4344 5672
rect 4344 5652 4396 5672
rect 4396 5652 4398 5672
rect 3882 5480 3938 5536
rect 3454 5466 3510 5468
rect 3534 5466 3590 5468
rect 3614 5466 3670 5468
rect 3694 5466 3750 5468
rect 3454 5414 3480 5466
rect 3480 5414 3510 5466
rect 3534 5414 3544 5466
rect 3544 5414 3590 5466
rect 3614 5414 3660 5466
rect 3660 5414 3670 5466
rect 3694 5414 3724 5466
rect 3724 5414 3750 5466
rect 3454 5412 3510 5414
rect 3534 5412 3590 5414
rect 3614 5412 3670 5414
rect 3694 5412 3750 5414
rect 3882 5344 3938 5400
rect 4342 5616 4398 5652
rect 3514 4936 3570 4992
rect 3422 4564 3424 4584
rect 3424 4564 3476 4584
rect 3476 4564 3478 4584
rect 3422 4528 3478 4564
rect 3454 4378 3510 4380
rect 3534 4378 3590 4380
rect 3614 4378 3670 4380
rect 3694 4378 3750 4380
rect 3454 4326 3480 4378
rect 3480 4326 3510 4378
rect 3534 4326 3544 4378
rect 3544 4326 3590 4378
rect 3614 4326 3660 4378
rect 3660 4326 3670 4378
rect 3694 4326 3724 4378
rect 3724 4326 3750 4378
rect 3454 4324 3510 4326
rect 3534 4324 3590 4326
rect 3614 4324 3670 4326
rect 3694 4324 3750 4326
rect 3330 3712 3386 3768
rect 3698 3596 3754 3632
rect 3698 3576 3700 3596
rect 3700 3576 3752 3596
rect 3752 3576 3754 3596
rect 3238 2896 3294 2952
rect 3454 3290 3510 3292
rect 3534 3290 3590 3292
rect 3614 3290 3670 3292
rect 3694 3290 3750 3292
rect 3454 3238 3480 3290
rect 3480 3238 3510 3290
rect 3534 3238 3544 3290
rect 3544 3238 3590 3290
rect 3614 3238 3660 3290
rect 3660 3238 3670 3290
rect 3694 3238 3724 3290
rect 3724 3238 3750 3290
rect 3454 3236 3510 3238
rect 3534 3236 3590 3238
rect 3614 3236 3670 3238
rect 3694 3236 3750 3238
rect 4066 4528 4122 4584
rect 4434 4256 4490 4312
rect 4618 4936 4674 4992
rect 4342 3848 4398 3904
rect 4526 3168 4582 3224
rect 3454 2202 3510 2204
rect 3534 2202 3590 2204
rect 3614 2202 3670 2204
rect 3694 2202 3750 2204
rect 3454 2150 3480 2202
rect 3480 2150 3510 2202
rect 3534 2150 3544 2202
rect 3544 2150 3590 2202
rect 3614 2150 3660 2202
rect 3660 2150 3670 2202
rect 3694 2150 3724 2202
rect 3724 2150 3750 2202
rect 3454 2148 3510 2150
rect 3534 2148 3590 2150
rect 3614 2148 3670 2150
rect 3694 2148 3750 2150
rect 6366 10104 6422 10160
rect 5630 9560 5686 9616
rect 5538 9324 5540 9344
rect 5540 9324 5592 9344
rect 5592 9324 5594 9344
rect 5078 8744 5134 8800
rect 5538 9288 5594 9324
rect 5953 9274 6009 9276
rect 6033 9274 6089 9276
rect 6113 9274 6169 9276
rect 6193 9274 6249 9276
rect 5953 9222 5979 9274
rect 5979 9222 6009 9274
rect 6033 9222 6043 9274
rect 6043 9222 6089 9274
rect 6113 9222 6159 9274
rect 6159 9222 6169 9274
rect 6193 9222 6223 9274
rect 6223 9222 6249 9274
rect 5953 9220 6009 9222
rect 6033 9220 6089 9222
rect 6113 9220 6169 9222
rect 6193 9220 6249 9222
rect 5630 9016 5686 9072
rect 6550 8608 6606 8664
rect 6734 14320 6790 14376
rect 7194 13776 7250 13832
rect 7010 12824 7066 12880
rect 6918 12688 6974 12744
rect 6734 11464 6790 11520
rect 7194 10240 7250 10296
rect 6826 10104 6882 10160
rect 7194 9696 7250 9752
rect 5814 8200 5870 8256
rect 5170 7928 5226 7984
rect 4802 4936 4858 4992
rect 4710 4800 4766 4856
rect 4710 4256 4766 4312
rect 5262 6976 5318 7032
rect 5953 8186 6009 8188
rect 6033 8186 6089 8188
rect 6113 8186 6169 8188
rect 6193 8186 6249 8188
rect 5953 8134 5979 8186
rect 5979 8134 6009 8186
rect 6033 8134 6043 8186
rect 6043 8134 6089 8186
rect 6113 8134 6159 8186
rect 6159 8134 6169 8186
rect 6193 8134 6223 8186
rect 6223 8134 6249 8186
rect 5953 8132 6009 8134
rect 6033 8132 6089 8134
rect 6113 8132 6169 8134
rect 6193 8132 6249 8134
rect 8206 15680 8262 15736
rect 8452 16346 8508 16348
rect 8532 16346 8588 16348
rect 8612 16346 8668 16348
rect 8692 16346 8748 16348
rect 8452 16294 8478 16346
rect 8478 16294 8508 16346
rect 8532 16294 8542 16346
rect 8542 16294 8588 16346
rect 8612 16294 8658 16346
rect 8658 16294 8668 16346
rect 8692 16294 8722 16346
rect 8722 16294 8748 16346
rect 8452 16292 8508 16294
rect 8532 16292 8588 16294
rect 8612 16292 8668 16294
rect 8692 16292 8748 16294
rect 7470 13504 7526 13560
rect 7378 13096 7434 13152
rect 8206 15408 8262 15464
rect 7838 14340 7894 14376
rect 7838 14320 7840 14340
rect 7840 14320 7892 14340
rect 7892 14320 7894 14340
rect 8022 13232 8078 13288
rect 8206 13640 8262 13696
rect 7930 12144 7986 12200
rect 8452 15258 8508 15260
rect 8532 15258 8588 15260
rect 8612 15258 8668 15260
rect 8692 15258 8748 15260
rect 8452 15206 8478 15258
rect 8478 15206 8508 15258
rect 8532 15206 8542 15258
rect 8542 15206 8588 15258
rect 8612 15206 8658 15258
rect 8658 15206 8668 15258
rect 8692 15206 8722 15258
rect 8722 15206 8748 15258
rect 8452 15204 8508 15206
rect 8532 15204 8588 15206
rect 8612 15204 8668 15206
rect 8692 15204 8748 15206
rect 8758 15020 8814 15056
rect 8758 15000 8760 15020
rect 8760 15000 8812 15020
rect 8812 15000 8814 15020
rect 8452 14170 8508 14172
rect 8532 14170 8588 14172
rect 8612 14170 8668 14172
rect 8692 14170 8748 14172
rect 8452 14118 8478 14170
rect 8478 14118 8508 14170
rect 8532 14118 8542 14170
rect 8542 14118 8588 14170
rect 8612 14118 8658 14170
rect 8658 14118 8668 14170
rect 8692 14118 8722 14170
rect 8722 14118 8748 14170
rect 8452 14116 8508 14118
rect 8532 14116 8588 14118
rect 8612 14116 8668 14118
rect 8692 14116 8748 14118
rect 8482 13776 8538 13832
rect 9494 15852 9496 15872
rect 9496 15852 9548 15872
rect 9548 15852 9550 15872
rect 9494 15816 9550 15852
rect 9126 13912 9182 13968
rect 9310 13776 9366 13832
rect 9034 13640 9090 13696
rect 9126 13504 9182 13560
rect 8452 13082 8508 13084
rect 8532 13082 8588 13084
rect 8612 13082 8668 13084
rect 8692 13082 8748 13084
rect 8452 13030 8478 13082
rect 8478 13030 8508 13082
rect 8532 13030 8542 13082
rect 8542 13030 8588 13082
rect 8612 13030 8658 13082
rect 8658 13030 8668 13082
rect 8692 13030 8722 13082
rect 8722 13030 8748 13082
rect 8452 13028 8508 13030
rect 8532 13028 8588 13030
rect 8612 13028 8668 13030
rect 8692 13028 8748 13030
rect 8758 12416 8814 12472
rect 9770 16532 9772 16552
rect 9772 16532 9824 16552
rect 9824 16532 9826 16552
rect 9770 16496 9826 16532
rect 9770 15000 9826 15056
rect 9678 14340 9734 14376
rect 9678 14320 9680 14340
rect 9680 14320 9732 14340
rect 9732 14320 9734 14340
rect 9678 13912 9734 13968
rect 9494 13776 9550 13832
rect 9310 13232 9366 13288
rect 9126 12860 9128 12880
rect 9128 12860 9180 12880
rect 9180 12860 9182 12880
rect 9126 12824 9182 12860
rect 8942 12552 8998 12608
rect 8452 11994 8508 11996
rect 8532 11994 8588 11996
rect 8612 11994 8668 11996
rect 8692 11994 8748 11996
rect 8452 11942 8478 11994
rect 8478 11942 8508 11994
rect 8532 11942 8542 11994
rect 8542 11942 8588 11994
rect 8612 11942 8658 11994
rect 8658 11942 8668 11994
rect 8692 11942 8722 11994
rect 8722 11942 8748 11994
rect 8452 11940 8508 11942
rect 8532 11940 8588 11942
rect 8612 11940 8668 11942
rect 8692 11940 8748 11942
rect 8114 11056 8170 11112
rect 7746 10376 7802 10432
rect 7286 8880 7342 8936
rect 8452 10906 8508 10908
rect 8532 10906 8588 10908
rect 8612 10906 8668 10908
rect 8692 10906 8748 10908
rect 8452 10854 8478 10906
rect 8478 10854 8508 10906
rect 8532 10854 8542 10906
rect 8542 10854 8588 10906
rect 8612 10854 8658 10906
rect 8658 10854 8668 10906
rect 8692 10854 8722 10906
rect 8722 10854 8748 10906
rect 8452 10852 8508 10854
rect 8532 10852 8588 10854
rect 8612 10852 8668 10854
rect 8692 10852 8748 10854
rect 8850 10412 8852 10432
rect 8852 10412 8904 10432
rect 8904 10412 8906 10432
rect 8850 10376 8906 10412
rect 8850 10240 8906 10296
rect 9126 12552 9182 12608
rect 9034 11464 9090 11520
rect 9678 13676 9680 13696
rect 9680 13676 9732 13696
rect 9732 13676 9734 13696
rect 9678 13640 9734 13676
rect 8452 9818 8508 9820
rect 8532 9818 8588 9820
rect 8612 9818 8668 9820
rect 8692 9818 8748 9820
rect 8452 9766 8478 9818
rect 8478 9766 8508 9818
rect 8532 9766 8542 9818
rect 8542 9766 8588 9818
rect 8612 9766 8658 9818
rect 8658 9766 8668 9818
rect 8692 9766 8722 9818
rect 8722 9766 8748 9818
rect 8452 9764 8508 9766
rect 8532 9764 8588 9766
rect 8612 9764 8668 9766
rect 8692 9764 8748 9766
rect 8114 9424 8170 9480
rect 8114 9152 8170 9208
rect 7470 8744 7526 8800
rect 7286 8336 7342 8392
rect 5722 7112 5778 7168
rect 6366 7112 6422 7168
rect 5953 7098 6009 7100
rect 6033 7098 6089 7100
rect 6113 7098 6169 7100
rect 6193 7098 6249 7100
rect 5953 7046 5979 7098
rect 5979 7046 6009 7098
rect 6033 7046 6043 7098
rect 6043 7046 6089 7098
rect 6113 7046 6159 7098
rect 6159 7046 6169 7098
rect 6193 7046 6223 7098
rect 6223 7046 6249 7098
rect 5953 7044 6009 7046
rect 6033 7044 6089 7046
rect 6113 7044 6169 7046
rect 6193 7044 6249 7046
rect 6458 6976 6514 7032
rect 5953 6010 6009 6012
rect 6033 6010 6089 6012
rect 6113 6010 6169 6012
rect 6193 6010 6249 6012
rect 5953 5958 5979 6010
rect 5979 5958 6009 6010
rect 6033 5958 6043 6010
rect 6043 5958 6089 6010
rect 6113 5958 6159 6010
rect 6159 5958 6169 6010
rect 6193 5958 6223 6010
rect 6223 5958 6249 6010
rect 5953 5956 6009 5958
rect 6033 5956 6089 5958
rect 6113 5956 6169 5958
rect 6193 5956 6249 5958
rect 5814 5888 5870 5944
rect 5354 4936 5410 4992
rect 5078 3884 5080 3904
rect 5080 3884 5132 3904
rect 5132 3884 5134 3904
rect 5078 3848 5134 3884
rect 5170 3712 5226 3768
rect 5354 3848 5410 3904
rect 5630 5480 5686 5536
rect 5814 5480 5870 5536
rect 5538 4392 5594 4448
rect 5170 3304 5226 3360
rect 5446 3304 5502 3360
rect 5078 2916 5134 2952
rect 5953 4922 6009 4924
rect 6033 4922 6089 4924
rect 6113 4922 6169 4924
rect 6193 4922 6249 4924
rect 5953 4870 5979 4922
rect 5979 4870 6009 4922
rect 6033 4870 6043 4922
rect 6043 4870 6089 4922
rect 6113 4870 6159 4922
rect 6159 4870 6169 4922
rect 6193 4870 6223 4922
rect 6223 4870 6249 4922
rect 5953 4868 6009 4870
rect 6033 4868 6089 4870
rect 6113 4868 6169 4870
rect 6193 4868 6249 4870
rect 5814 4392 5870 4448
rect 6918 6024 6974 6080
rect 6550 5344 6606 5400
rect 6734 5480 6790 5536
rect 5953 3834 6009 3836
rect 6033 3834 6089 3836
rect 6113 3834 6169 3836
rect 6193 3834 6249 3836
rect 5953 3782 5979 3834
rect 5979 3782 6009 3834
rect 6033 3782 6043 3834
rect 6043 3782 6089 3834
rect 6113 3782 6159 3834
rect 6159 3782 6169 3834
rect 6193 3782 6223 3834
rect 6223 3782 6249 3834
rect 5953 3780 6009 3782
rect 6033 3780 6089 3782
rect 6113 3780 6169 3782
rect 6193 3780 6249 3782
rect 6458 4256 6514 4312
rect 5078 2896 5080 2916
rect 5080 2896 5132 2916
rect 5132 2896 5134 2916
rect 4710 2352 4766 2408
rect 6458 3884 6460 3904
rect 6460 3884 6512 3904
rect 6512 3884 6514 3904
rect 6458 3848 6514 3884
rect 6550 3712 6606 3768
rect 6274 2896 6330 2952
rect 5953 2746 6009 2748
rect 6033 2746 6089 2748
rect 6113 2746 6169 2748
rect 6193 2746 6249 2748
rect 5953 2694 5979 2746
rect 5979 2694 6009 2746
rect 6033 2694 6043 2746
rect 6043 2694 6089 2746
rect 6113 2694 6159 2746
rect 6159 2694 6169 2746
rect 6193 2694 6223 2746
rect 6223 2694 6249 2746
rect 5953 2692 6009 2694
rect 6033 2692 6089 2694
rect 6113 2692 6169 2694
rect 6193 2692 6249 2694
rect 6550 3304 6606 3360
rect 6550 2760 6606 2816
rect 6550 2488 6606 2544
rect 6090 2388 6092 2408
rect 6092 2388 6144 2408
rect 6144 2388 6146 2408
rect 6090 2352 6146 2388
rect 7010 2760 7066 2816
rect 7378 6432 7434 6488
rect 7378 5888 7434 5944
rect 7286 3032 7342 3088
rect 8114 8064 8170 8120
rect 8298 8744 8354 8800
rect 8452 8730 8508 8732
rect 8532 8730 8588 8732
rect 8612 8730 8668 8732
rect 8692 8730 8748 8732
rect 8452 8678 8478 8730
rect 8478 8678 8508 8730
rect 8532 8678 8542 8730
rect 8542 8678 8588 8730
rect 8612 8678 8658 8730
rect 8658 8678 8668 8730
rect 8692 8678 8722 8730
rect 8722 8678 8748 8730
rect 8452 8676 8508 8678
rect 8532 8676 8588 8678
rect 8612 8676 8668 8678
rect 8692 8676 8748 8678
rect 8850 7656 8906 7712
rect 8452 7642 8508 7644
rect 8532 7642 8588 7644
rect 8612 7642 8668 7644
rect 8692 7642 8748 7644
rect 8452 7590 8478 7642
rect 8478 7590 8508 7642
rect 8532 7590 8542 7642
rect 8542 7590 8588 7642
rect 8612 7590 8658 7642
rect 8658 7590 8668 7642
rect 8692 7590 8722 7642
rect 8722 7590 8748 7642
rect 8452 7588 8508 7590
rect 8532 7588 8588 7590
rect 8612 7588 8668 7590
rect 8692 7588 8748 7590
rect 8206 7520 8262 7576
rect 8850 7520 8906 7576
rect 8114 7112 8170 7168
rect 8298 6568 8354 6624
rect 8850 6568 8906 6624
rect 8452 6554 8508 6556
rect 8532 6554 8588 6556
rect 8612 6554 8668 6556
rect 8692 6554 8748 6556
rect 8452 6502 8478 6554
rect 8478 6502 8508 6554
rect 8532 6502 8542 6554
rect 8542 6502 8588 6554
rect 8612 6502 8658 6554
rect 8658 6502 8668 6554
rect 8692 6502 8722 6554
rect 8722 6502 8748 6554
rect 8452 6500 8508 6502
rect 8532 6500 8588 6502
rect 8612 6500 8668 6502
rect 8692 6500 8748 6502
rect 8206 6296 8262 6352
rect 8206 5788 8208 5808
rect 8208 5788 8260 5808
rect 8260 5788 8262 5808
rect 8206 5752 8262 5788
rect 8390 5752 8446 5808
rect 8666 6160 8722 6216
rect 8850 5752 8906 5808
rect 8298 5480 8354 5536
rect 8452 5466 8508 5468
rect 8532 5466 8588 5468
rect 8612 5466 8668 5468
rect 8692 5466 8748 5468
rect 8452 5414 8478 5466
rect 8478 5414 8508 5466
rect 8532 5414 8542 5466
rect 8542 5414 8588 5466
rect 8612 5414 8658 5466
rect 8658 5414 8668 5466
rect 8692 5414 8722 5466
rect 8722 5414 8748 5466
rect 8452 5412 8508 5414
rect 8532 5412 8588 5414
rect 8612 5412 8668 5414
rect 8692 5412 8748 5414
rect 8114 4392 8170 4448
rect 8452 4378 8508 4380
rect 8532 4378 8588 4380
rect 8612 4378 8668 4380
rect 8692 4378 8748 4380
rect 8452 4326 8478 4378
rect 8478 4326 8508 4378
rect 8532 4326 8542 4378
rect 8542 4326 8588 4378
rect 8612 4326 8658 4378
rect 8658 4326 8668 4378
rect 8692 4326 8722 4378
rect 8722 4326 8748 4378
rect 8452 4324 8508 4326
rect 8532 4324 8588 4326
rect 8612 4324 8668 4326
rect 8692 4324 8748 4326
rect 8022 3848 8078 3904
rect 8114 3168 8170 3224
rect 7930 3032 7986 3088
rect 8114 2896 8170 2952
rect 7654 2624 7710 2680
rect 7746 1944 7802 2000
rect 8206 2488 8262 2544
rect 8114 2216 8170 2272
rect 8452 3290 8508 3292
rect 8532 3290 8588 3292
rect 8612 3290 8668 3292
rect 8692 3290 8748 3292
rect 8452 3238 8478 3290
rect 8478 3238 8508 3290
rect 8532 3238 8542 3290
rect 8542 3238 8588 3290
rect 8612 3238 8658 3290
rect 8658 3238 8668 3290
rect 8692 3238 8722 3290
rect 8722 3238 8748 3290
rect 8452 3236 8508 3238
rect 8532 3236 8588 3238
rect 8612 3236 8668 3238
rect 8692 3236 8748 3238
rect 9126 9696 9182 9752
rect 9126 9288 9182 9344
rect 9310 10684 9312 10704
rect 9312 10684 9364 10704
rect 9364 10684 9366 10704
rect 9310 10648 9366 10684
rect 9770 13232 9826 13288
rect 9862 12824 9918 12880
rect 9862 12708 9918 12744
rect 9862 12688 9864 12708
rect 9864 12688 9916 12708
rect 9916 12688 9918 12708
rect 9862 12280 9918 12336
rect 9494 11056 9550 11112
rect 9770 10784 9826 10840
rect 9402 10104 9458 10160
rect 9494 9152 9550 9208
rect 9678 9288 9734 9344
rect 9218 8608 9274 8664
rect 10046 12144 10102 12200
rect 9954 11328 10010 11384
rect 10322 15408 10378 15464
rect 10414 13776 10470 13832
rect 10414 10920 10470 10976
rect 9770 6704 9826 6760
rect 9494 6568 9550 6624
rect 9770 6160 9826 6216
rect 9494 5364 9550 5400
rect 9494 5344 9496 5364
rect 9496 5344 9548 5364
rect 9548 5344 9550 5364
rect 9310 5208 9366 5264
rect 9494 5228 9550 5264
rect 9494 5208 9496 5228
rect 9496 5208 9548 5228
rect 9548 5208 9550 5228
rect 9310 4800 9366 4856
rect 9126 4528 9182 4584
rect 9310 4392 9366 4448
rect 9126 4276 9182 4312
rect 9126 4256 9128 4276
rect 9128 4256 9180 4276
rect 9180 4256 9182 4276
rect 8666 2796 8668 2816
rect 8668 2796 8720 2816
rect 8720 2796 8722 2816
rect 8666 2760 8722 2796
rect 8452 2202 8508 2204
rect 8532 2202 8588 2204
rect 8612 2202 8668 2204
rect 8692 2202 8748 2204
rect 8452 2150 8478 2202
rect 8478 2150 8508 2202
rect 8532 2150 8542 2202
rect 8542 2150 8588 2202
rect 8612 2150 8658 2202
rect 8658 2150 8668 2202
rect 8692 2150 8722 2202
rect 8722 2150 8748 2202
rect 8452 2148 8508 2150
rect 8532 2148 8588 2150
rect 8612 2148 8668 2150
rect 8692 2148 8748 2150
rect 9494 4120 9550 4176
rect 10138 8744 10194 8800
rect 10046 7112 10102 7168
rect 10046 6568 10102 6624
rect 10046 6160 10102 6216
rect 9770 4392 9826 4448
rect 9586 3304 9642 3360
rect 9494 3168 9550 3224
rect 10046 5364 10102 5400
rect 10046 5344 10048 5364
rect 10048 5344 10100 5364
rect 10100 5344 10102 5364
rect 10230 8608 10286 8664
rect 10414 10376 10470 10432
rect 10950 16890 11006 16892
rect 11030 16890 11086 16892
rect 11110 16890 11166 16892
rect 11190 16890 11246 16892
rect 10950 16838 10976 16890
rect 10976 16838 11006 16890
rect 11030 16838 11040 16890
rect 11040 16838 11086 16890
rect 11110 16838 11156 16890
rect 11156 16838 11166 16890
rect 11190 16838 11220 16890
rect 11220 16838 11246 16890
rect 10950 16836 11006 16838
rect 11030 16836 11086 16838
rect 11110 16836 11166 16838
rect 11190 16836 11246 16838
rect 10950 15802 11006 15804
rect 11030 15802 11086 15804
rect 11110 15802 11166 15804
rect 11190 15802 11246 15804
rect 10950 15750 10976 15802
rect 10976 15750 11006 15802
rect 11030 15750 11040 15802
rect 11040 15750 11086 15802
rect 11110 15750 11156 15802
rect 11156 15750 11166 15802
rect 11190 15750 11220 15802
rect 11220 15750 11246 15802
rect 10950 15748 11006 15750
rect 11030 15748 11086 15750
rect 11110 15748 11166 15750
rect 11190 15748 11246 15750
rect 10950 14714 11006 14716
rect 11030 14714 11086 14716
rect 11110 14714 11166 14716
rect 11190 14714 11246 14716
rect 10950 14662 10976 14714
rect 10976 14662 11006 14714
rect 11030 14662 11040 14714
rect 11040 14662 11086 14714
rect 11110 14662 11156 14714
rect 11156 14662 11166 14714
rect 11190 14662 11220 14714
rect 11220 14662 11246 14714
rect 10950 14660 11006 14662
rect 11030 14660 11086 14662
rect 11110 14660 11166 14662
rect 11190 14660 11246 14662
rect 10950 13626 11006 13628
rect 11030 13626 11086 13628
rect 11110 13626 11166 13628
rect 11190 13626 11246 13628
rect 10950 13574 10976 13626
rect 10976 13574 11006 13626
rect 11030 13574 11040 13626
rect 11040 13574 11086 13626
rect 11110 13574 11156 13626
rect 11156 13574 11166 13626
rect 11190 13574 11220 13626
rect 11220 13574 11246 13626
rect 10950 13572 11006 13574
rect 11030 13572 11086 13574
rect 11110 13572 11166 13574
rect 11190 13572 11246 13574
rect 10690 12960 10746 13016
rect 11150 13132 11152 13152
rect 11152 13132 11204 13152
rect 11204 13132 11206 13152
rect 11150 13096 11206 13132
rect 10874 12844 10930 12880
rect 10874 12824 10876 12844
rect 10876 12824 10928 12844
rect 10928 12824 10930 12844
rect 10598 12588 10600 12608
rect 10600 12588 10652 12608
rect 10652 12588 10654 12608
rect 10598 12552 10654 12588
rect 10690 12436 10746 12472
rect 10690 12416 10692 12436
rect 10692 12416 10744 12436
rect 10744 12416 10746 12436
rect 10690 11872 10746 11928
rect 10690 11500 10692 11520
rect 10692 11500 10744 11520
rect 10744 11500 10746 11520
rect 10690 11464 10746 11500
rect 10690 11328 10746 11384
rect 10950 12538 11006 12540
rect 11030 12538 11086 12540
rect 11110 12538 11166 12540
rect 11190 12538 11246 12540
rect 10950 12486 10976 12538
rect 10976 12486 11006 12538
rect 11030 12486 11040 12538
rect 11040 12486 11086 12538
rect 11110 12486 11156 12538
rect 11156 12486 11166 12538
rect 11190 12486 11220 12538
rect 11220 12486 11246 12538
rect 10950 12484 11006 12486
rect 11030 12484 11086 12486
rect 11110 12484 11166 12486
rect 11190 12484 11246 12486
rect 11058 12008 11114 12064
rect 11426 12144 11482 12200
rect 10950 11450 11006 11452
rect 11030 11450 11086 11452
rect 11110 11450 11166 11452
rect 11190 11450 11246 11452
rect 10950 11398 10976 11450
rect 10976 11398 11006 11450
rect 11030 11398 11040 11450
rect 11040 11398 11086 11450
rect 11110 11398 11156 11450
rect 11156 11398 11166 11450
rect 11190 11398 11220 11450
rect 11220 11398 11246 11450
rect 10950 11396 11006 11398
rect 11030 11396 11086 11398
rect 11110 11396 11166 11398
rect 11190 11396 11246 11398
rect 10506 9288 10562 9344
rect 10506 9152 10562 9208
rect 10874 10512 10930 10568
rect 11242 10512 11298 10568
rect 10782 9832 10838 9888
rect 10690 9152 10746 9208
rect 10950 10362 11006 10364
rect 11030 10362 11086 10364
rect 11110 10362 11166 10364
rect 11190 10362 11246 10364
rect 10950 10310 10976 10362
rect 10976 10310 11006 10362
rect 11030 10310 11040 10362
rect 11040 10310 11086 10362
rect 11110 10310 11156 10362
rect 11156 10310 11166 10362
rect 11190 10310 11220 10362
rect 11220 10310 11246 10362
rect 10950 10308 11006 10310
rect 11030 10308 11086 10310
rect 11110 10308 11166 10310
rect 11190 10308 11246 10310
rect 11426 11736 11482 11792
rect 11978 12824 12034 12880
rect 12254 12724 12256 12744
rect 12256 12724 12308 12744
rect 12308 12724 12310 12744
rect 12254 12688 12310 12724
rect 11518 11348 11574 11384
rect 11518 11328 11520 11348
rect 11520 11328 11572 11348
rect 11572 11328 11574 11348
rect 11610 11056 11666 11112
rect 11518 10648 11574 10704
rect 11426 9832 11482 9888
rect 11334 9288 11390 9344
rect 10950 9274 11006 9276
rect 11030 9274 11086 9276
rect 11110 9274 11166 9276
rect 11190 9274 11246 9276
rect 10950 9222 10976 9274
rect 10976 9222 11006 9274
rect 11030 9222 11040 9274
rect 11040 9222 11086 9274
rect 11110 9222 11156 9274
rect 11156 9222 11166 9274
rect 11190 9222 11220 9274
rect 11220 9222 11246 9274
rect 10950 9220 11006 9222
rect 11030 9220 11086 9222
rect 11110 9220 11166 9222
rect 11190 9220 11246 9222
rect 10322 8200 10378 8256
rect 11702 9560 11758 9616
rect 11702 9152 11758 9208
rect 11518 8608 11574 8664
rect 10782 8200 10838 8256
rect 10950 8186 11006 8188
rect 11030 8186 11086 8188
rect 11110 8186 11166 8188
rect 11190 8186 11246 8188
rect 10950 8134 10976 8186
rect 10976 8134 11006 8186
rect 11030 8134 11040 8186
rect 11040 8134 11086 8186
rect 11110 8134 11156 8186
rect 11156 8134 11166 8186
rect 11190 8134 11220 8186
rect 11220 8134 11246 8186
rect 10950 8132 11006 8134
rect 11030 8132 11086 8134
rect 11110 8132 11166 8134
rect 11190 8132 11246 8134
rect 10874 7656 10930 7712
rect 11058 7656 11114 7712
rect 11242 7792 11298 7848
rect 10598 7112 10654 7168
rect 10322 5752 10378 5808
rect 10322 5344 10378 5400
rect 10506 5752 10562 5808
rect 10230 5208 10286 5264
rect 10506 5208 10562 5264
rect 10138 4800 10194 4856
rect 10138 4428 10140 4448
rect 10140 4428 10192 4448
rect 10192 4428 10194 4448
rect 10138 4392 10194 4428
rect 10046 3712 10102 3768
rect 9954 3576 10010 3632
rect 10046 3304 10102 3360
rect 9862 3032 9918 3088
rect 9310 2352 9366 2408
rect 9862 2760 9918 2816
rect 9494 2080 9550 2136
rect 9402 1944 9458 2000
rect 10782 6976 10838 7032
rect 10950 7098 11006 7100
rect 11030 7098 11086 7100
rect 11110 7098 11166 7100
rect 11190 7098 11246 7100
rect 10950 7046 10976 7098
rect 10976 7046 11006 7098
rect 11030 7046 11040 7098
rect 11040 7046 11086 7098
rect 11110 7046 11156 7098
rect 11156 7046 11166 7098
rect 11190 7046 11220 7098
rect 11220 7046 11246 7098
rect 10950 7044 11006 7046
rect 11030 7044 11086 7046
rect 11110 7044 11166 7046
rect 11190 7044 11246 7046
rect 10874 6840 10930 6896
rect 11058 6840 11114 6896
rect 11150 6704 11206 6760
rect 10874 6160 10930 6216
rect 11058 6160 11114 6216
rect 10782 6024 10838 6080
rect 10950 6010 11006 6012
rect 11030 6010 11086 6012
rect 11110 6010 11166 6012
rect 11190 6010 11246 6012
rect 10950 5958 10976 6010
rect 10976 5958 11006 6010
rect 11030 5958 11040 6010
rect 11040 5958 11086 6010
rect 11110 5958 11156 6010
rect 11156 5958 11166 6010
rect 11190 5958 11220 6010
rect 11220 5958 11246 6010
rect 10950 5956 11006 5958
rect 11030 5956 11086 5958
rect 11110 5956 11166 5958
rect 11190 5956 11246 5958
rect 10598 4936 10654 4992
rect 12530 11892 12586 11928
rect 12530 11872 12532 11892
rect 12532 11872 12584 11892
rect 12584 11872 12586 11892
rect 12438 11600 12494 11656
rect 12254 11228 12256 11248
rect 12256 11228 12308 11248
rect 12308 11228 12310 11248
rect 12254 11192 12310 11228
rect 12070 10920 12126 10976
rect 12070 10376 12126 10432
rect 11886 9832 11942 9888
rect 12070 9832 12126 9888
rect 11886 9324 11888 9344
rect 11888 9324 11940 9344
rect 11940 9324 11942 9344
rect 11886 9288 11942 9324
rect 11794 8200 11850 8256
rect 11794 8084 11850 8120
rect 11794 8064 11796 8084
rect 11796 8064 11848 8084
rect 11848 8064 11850 8084
rect 11978 8744 12034 8800
rect 11978 8608 12034 8664
rect 11886 7792 11942 7848
rect 12254 10920 12310 10976
rect 12714 11092 12716 11112
rect 12716 11092 12768 11112
rect 12768 11092 12770 11112
rect 12714 11056 12770 11092
rect 13449 17434 13505 17436
rect 13529 17434 13585 17436
rect 13609 17434 13665 17436
rect 13689 17434 13745 17436
rect 13449 17382 13475 17434
rect 13475 17382 13505 17434
rect 13529 17382 13539 17434
rect 13539 17382 13585 17434
rect 13609 17382 13655 17434
rect 13655 17382 13665 17434
rect 13689 17382 13719 17434
rect 13719 17382 13745 17434
rect 13449 17380 13505 17382
rect 13529 17380 13585 17382
rect 13609 17380 13665 17382
rect 13689 17380 13745 17382
rect 13082 12280 13138 12336
rect 13449 16346 13505 16348
rect 13529 16346 13585 16348
rect 13609 16346 13665 16348
rect 13689 16346 13745 16348
rect 13449 16294 13475 16346
rect 13475 16294 13505 16346
rect 13529 16294 13539 16346
rect 13539 16294 13585 16346
rect 13609 16294 13655 16346
rect 13655 16294 13665 16346
rect 13689 16294 13719 16346
rect 13719 16294 13745 16346
rect 13449 16292 13505 16294
rect 13529 16292 13585 16294
rect 13609 16292 13665 16294
rect 13689 16292 13745 16294
rect 13449 15258 13505 15260
rect 13529 15258 13585 15260
rect 13609 15258 13665 15260
rect 13689 15258 13745 15260
rect 13449 15206 13475 15258
rect 13475 15206 13505 15258
rect 13529 15206 13539 15258
rect 13539 15206 13585 15258
rect 13609 15206 13655 15258
rect 13655 15206 13665 15258
rect 13689 15206 13719 15258
rect 13719 15206 13745 15258
rect 13449 15204 13505 15206
rect 13529 15204 13585 15206
rect 13609 15204 13665 15206
rect 13689 15204 13745 15206
rect 13449 14170 13505 14172
rect 13529 14170 13585 14172
rect 13609 14170 13665 14172
rect 13689 14170 13745 14172
rect 13449 14118 13475 14170
rect 13475 14118 13505 14170
rect 13529 14118 13539 14170
rect 13539 14118 13585 14170
rect 13609 14118 13655 14170
rect 13655 14118 13665 14170
rect 13689 14118 13719 14170
rect 13719 14118 13745 14170
rect 13449 14116 13505 14118
rect 13529 14116 13585 14118
rect 13609 14116 13665 14118
rect 13689 14116 13745 14118
rect 13449 13082 13505 13084
rect 13529 13082 13585 13084
rect 13609 13082 13665 13084
rect 13689 13082 13745 13084
rect 13449 13030 13475 13082
rect 13475 13030 13505 13082
rect 13529 13030 13539 13082
rect 13539 13030 13585 13082
rect 13609 13030 13655 13082
rect 13655 13030 13665 13082
rect 13689 13030 13719 13082
rect 13719 13030 13745 13082
rect 13449 13028 13505 13030
rect 13529 13028 13585 13030
rect 13609 13028 13665 13030
rect 13689 13028 13745 13030
rect 13449 11994 13505 11996
rect 13529 11994 13585 11996
rect 13609 11994 13665 11996
rect 13689 11994 13745 11996
rect 13449 11942 13475 11994
rect 13475 11942 13505 11994
rect 13529 11942 13539 11994
rect 13539 11942 13585 11994
rect 13609 11942 13655 11994
rect 13655 11942 13665 11994
rect 13689 11942 13719 11994
rect 13719 11942 13745 11994
rect 13449 11940 13505 11942
rect 13529 11940 13585 11942
rect 13609 11940 13665 11942
rect 13689 11940 13745 11942
rect 12254 10260 12310 10296
rect 12254 10240 12256 10260
rect 12256 10240 12308 10260
rect 12308 10240 12310 10260
rect 12438 9832 12494 9888
rect 12622 9560 12678 9616
rect 12162 9152 12218 9208
rect 12806 9560 12862 9616
rect 12806 9460 12808 9480
rect 12808 9460 12860 9480
rect 12860 9460 12862 9480
rect 12806 9424 12862 9460
rect 12898 9152 12954 9208
rect 12714 9016 12770 9072
rect 13266 10784 13322 10840
rect 13449 10906 13505 10908
rect 13529 10906 13585 10908
rect 13609 10906 13665 10908
rect 13689 10906 13745 10908
rect 13449 10854 13475 10906
rect 13475 10854 13505 10906
rect 13529 10854 13539 10906
rect 13539 10854 13585 10906
rect 13609 10854 13655 10906
rect 13655 10854 13665 10906
rect 13689 10854 13719 10906
rect 13719 10854 13745 10906
rect 13449 10852 13505 10854
rect 13529 10852 13585 10854
rect 13609 10852 13665 10854
rect 13689 10852 13745 10854
rect 13450 10648 13506 10704
rect 13174 10104 13230 10160
rect 12530 8508 12532 8528
rect 12532 8508 12584 8528
rect 12584 8508 12586 8528
rect 12530 8472 12586 8508
rect 12162 8200 12218 8256
rect 11702 7384 11758 7440
rect 12070 7792 12126 7848
rect 12254 7928 12310 7984
rect 12438 7928 12494 7984
rect 12622 8200 12678 8256
rect 12162 7656 12218 7712
rect 11978 7384 12034 7440
rect 11886 7112 11942 7168
rect 10966 5616 11022 5672
rect 10782 5208 10838 5264
rect 10782 4800 10838 4856
rect 10414 4120 10470 4176
rect 10414 3712 10470 3768
rect 10322 3168 10378 3224
rect 11334 5616 11390 5672
rect 11058 5092 11114 5128
rect 11058 5072 11060 5092
rect 11060 5072 11112 5092
rect 11112 5072 11114 5092
rect 10950 4922 11006 4924
rect 11030 4922 11086 4924
rect 11110 4922 11166 4924
rect 11190 4922 11246 4924
rect 10950 4870 10976 4922
rect 10976 4870 11006 4922
rect 11030 4870 11040 4922
rect 11040 4870 11086 4922
rect 11110 4870 11156 4922
rect 11156 4870 11166 4922
rect 11190 4870 11220 4922
rect 11220 4870 11246 4922
rect 10950 4868 11006 4870
rect 11030 4868 11086 4870
rect 11110 4868 11166 4870
rect 11190 4868 11246 4870
rect 11518 5072 11574 5128
rect 11426 4936 11482 4992
rect 10782 3848 10838 3904
rect 10950 3834 11006 3836
rect 11030 3834 11086 3836
rect 11110 3834 11166 3836
rect 11190 3834 11246 3836
rect 10950 3782 10976 3834
rect 10976 3782 11006 3834
rect 11030 3782 11040 3834
rect 11040 3782 11086 3834
rect 11110 3782 11156 3834
rect 11156 3782 11166 3834
rect 11190 3782 11220 3834
rect 11220 3782 11246 3834
rect 10950 3780 11006 3782
rect 11030 3780 11086 3782
rect 11110 3780 11166 3782
rect 11190 3780 11246 3782
rect 10506 3032 10562 3088
rect 10506 2488 10562 2544
rect 11518 3848 11574 3904
rect 11518 3732 11574 3768
rect 11518 3712 11520 3732
rect 11520 3712 11572 3732
rect 11572 3712 11574 3732
rect 10966 3168 11022 3224
rect 11242 3032 11298 3088
rect 11702 6840 11758 6896
rect 11794 5888 11850 5944
rect 11978 6296 12034 6352
rect 11702 5752 11758 5808
rect 11702 5480 11758 5536
rect 11702 4820 11758 4856
rect 11702 4800 11704 4820
rect 11704 4800 11756 4820
rect 11756 4800 11758 4820
rect 11702 4684 11758 4720
rect 11702 4664 11704 4684
rect 11704 4664 11756 4684
rect 11756 4664 11758 4684
rect 11978 4936 12034 4992
rect 11886 4800 11942 4856
rect 11702 4392 11758 4448
rect 11978 4548 12034 4584
rect 11978 4528 11980 4548
rect 11980 4528 12032 4548
rect 12032 4528 12034 4548
rect 12346 6976 12402 7032
rect 12162 6840 12218 6896
rect 12438 6432 12494 6488
rect 12162 6024 12218 6080
rect 11886 4256 11942 4312
rect 12070 4256 12126 4312
rect 11610 3440 11666 3496
rect 11794 3440 11850 3496
rect 11978 3576 12034 3632
rect 10782 2624 10838 2680
rect 10950 2746 11006 2748
rect 11030 2746 11086 2748
rect 11110 2746 11166 2748
rect 11190 2746 11246 2748
rect 10950 2694 10976 2746
rect 10976 2694 11006 2746
rect 11030 2694 11040 2746
rect 11040 2694 11086 2746
rect 11110 2694 11156 2746
rect 11156 2694 11166 2746
rect 11190 2694 11220 2746
rect 11220 2694 11246 2746
rect 10950 2692 11006 2694
rect 11030 2692 11086 2694
rect 11110 2692 11166 2694
rect 11190 2692 11246 2694
rect 10966 2488 11022 2544
rect 11058 1672 11114 1728
rect 11518 2760 11574 2816
rect 11702 2624 11758 2680
rect 11886 2896 11942 2952
rect 11610 2352 11666 2408
rect 11978 2796 11980 2816
rect 11980 2796 12032 2816
rect 12032 2796 12034 2816
rect 11978 2760 12034 2796
rect 11978 2488 12034 2544
rect 12346 6060 12348 6080
rect 12348 6060 12400 6080
rect 12400 6060 12402 6080
rect 12346 6024 12402 6060
rect 12254 5616 12310 5672
rect 12438 5344 12494 5400
rect 12438 4256 12494 4312
rect 12622 6976 12678 7032
rect 12898 7928 12954 7984
rect 13726 10240 13782 10296
rect 13910 10376 13966 10432
rect 13449 9818 13505 9820
rect 13529 9818 13585 9820
rect 13609 9818 13665 9820
rect 13689 9818 13745 9820
rect 13449 9766 13475 9818
rect 13475 9766 13505 9818
rect 13529 9766 13539 9818
rect 13539 9766 13585 9818
rect 13609 9766 13655 9818
rect 13655 9766 13665 9818
rect 13689 9766 13719 9818
rect 13719 9766 13745 9818
rect 13449 9764 13505 9766
rect 13529 9764 13585 9766
rect 13609 9764 13665 9766
rect 13689 9764 13745 9766
rect 14922 16632 14978 16688
rect 14002 9560 14058 9616
rect 13726 9152 13782 9208
rect 13542 9016 13598 9072
rect 13449 8730 13505 8732
rect 13529 8730 13585 8732
rect 13609 8730 13665 8732
rect 13689 8730 13745 8732
rect 13449 8678 13475 8730
rect 13475 8678 13505 8730
rect 13529 8678 13539 8730
rect 13539 8678 13585 8730
rect 13609 8678 13655 8730
rect 13655 8678 13665 8730
rect 13689 8678 13719 8730
rect 13719 8678 13745 8730
rect 13449 8676 13505 8678
rect 13529 8676 13585 8678
rect 13609 8676 13665 8678
rect 13689 8676 13745 8678
rect 13910 8880 13966 8936
rect 13358 8336 13414 8392
rect 13266 8236 13268 8256
rect 13268 8236 13320 8256
rect 13320 8236 13322 8256
rect 13266 8200 13322 8236
rect 13082 7520 13138 7576
rect 13082 7404 13138 7440
rect 13082 7384 13084 7404
rect 13084 7384 13136 7404
rect 13136 7384 13138 7404
rect 12714 5888 12770 5944
rect 12714 5788 12716 5808
rect 12716 5788 12768 5808
rect 12768 5788 12770 5808
rect 12714 5752 12770 5788
rect 12346 3848 12402 3904
rect 12438 3476 12440 3496
rect 12440 3476 12492 3496
rect 12492 3476 12494 3496
rect 12438 3440 12494 3476
rect 12990 6568 13046 6624
rect 13082 5480 13138 5536
rect 13449 7642 13505 7644
rect 13529 7642 13585 7644
rect 13609 7642 13665 7644
rect 13689 7642 13745 7644
rect 13449 7590 13475 7642
rect 13475 7590 13505 7642
rect 13529 7590 13539 7642
rect 13539 7590 13585 7642
rect 13609 7590 13655 7642
rect 13655 7590 13665 7642
rect 13689 7590 13719 7642
rect 13719 7590 13745 7642
rect 13449 7588 13505 7590
rect 13529 7588 13585 7590
rect 13609 7588 13665 7590
rect 13689 7588 13745 7590
rect 13818 7148 13820 7168
rect 13820 7148 13872 7168
rect 13872 7148 13874 7168
rect 13818 7112 13874 7148
rect 13449 6554 13505 6556
rect 13529 6554 13585 6556
rect 13609 6554 13665 6556
rect 13689 6554 13745 6556
rect 13449 6502 13475 6554
rect 13475 6502 13505 6554
rect 13529 6502 13539 6554
rect 13539 6502 13585 6554
rect 13609 6502 13655 6554
rect 13655 6502 13665 6554
rect 13689 6502 13719 6554
rect 13719 6502 13745 6554
rect 13449 6500 13505 6502
rect 13529 6500 13585 6502
rect 13609 6500 13665 6502
rect 13689 6500 13745 6502
rect 13174 5072 13230 5128
rect 12806 4936 12862 4992
rect 13358 6160 13414 6216
rect 13634 6024 13690 6080
rect 13082 4972 13084 4992
rect 13084 4972 13136 4992
rect 13136 4972 13138 4992
rect 13082 4936 13138 4972
rect 12622 3440 12678 3496
rect 12990 4004 13046 4040
rect 12990 3984 12992 4004
rect 12992 3984 13044 4004
rect 13044 3984 13046 4004
rect 12898 3168 12954 3224
rect 12714 1808 12770 1864
rect 13449 5466 13505 5468
rect 13529 5466 13585 5468
rect 13609 5466 13665 5468
rect 13689 5466 13745 5468
rect 13449 5414 13475 5466
rect 13475 5414 13505 5466
rect 13529 5414 13539 5466
rect 13539 5414 13585 5466
rect 13609 5414 13655 5466
rect 13655 5414 13665 5466
rect 13689 5414 13719 5466
rect 13719 5414 13745 5466
rect 13449 5412 13505 5414
rect 13529 5412 13585 5414
rect 13609 5412 13665 5414
rect 13689 5412 13745 5414
rect 13542 5244 13544 5264
rect 13544 5244 13596 5264
rect 13596 5244 13598 5264
rect 13542 5208 13598 5244
rect 13634 4800 13690 4856
rect 13634 4684 13690 4720
rect 13634 4664 13636 4684
rect 13636 4664 13688 4684
rect 13688 4664 13690 4684
rect 13449 4378 13505 4380
rect 13529 4378 13585 4380
rect 13609 4378 13665 4380
rect 13689 4378 13745 4380
rect 13449 4326 13475 4378
rect 13475 4326 13505 4378
rect 13529 4326 13539 4378
rect 13539 4326 13585 4378
rect 13609 4326 13655 4378
rect 13655 4326 13665 4378
rect 13689 4326 13719 4378
rect 13719 4326 13745 4378
rect 13449 4324 13505 4326
rect 13529 4324 13585 4326
rect 13609 4324 13665 4326
rect 13689 4324 13745 4326
rect 13726 4120 13782 4176
rect 13358 3596 13414 3632
rect 14094 8880 14150 8936
rect 14370 9988 14426 10024
rect 14370 9968 14372 9988
rect 14372 9968 14424 9988
rect 14424 9968 14426 9988
rect 14278 8064 14334 8120
rect 14094 6704 14150 6760
rect 13358 3576 13360 3596
rect 13360 3576 13412 3596
rect 13412 3576 13414 3596
rect 13449 3290 13505 3292
rect 13529 3290 13585 3292
rect 13609 3290 13665 3292
rect 13689 3290 13745 3292
rect 13449 3238 13475 3290
rect 13475 3238 13505 3290
rect 13529 3238 13539 3290
rect 13539 3238 13585 3290
rect 13609 3238 13655 3290
rect 13655 3238 13665 3290
rect 13689 3238 13719 3290
rect 13719 3238 13745 3290
rect 13449 3236 13505 3238
rect 13529 3236 13585 3238
rect 13609 3236 13665 3238
rect 13689 3236 13745 3238
rect 14370 6840 14426 6896
rect 14370 6316 14426 6352
rect 14370 6296 14372 6316
rect 14372 6296 14424 6316
rect 14424 6296 14426 6316
rect 14738 6976 14794 7032
rect 15658 16652 15714 16688
rect 15658 16632 15660 16652
rect 15660 16632 15712 16652
rect 15712 16632 15714 16652
rect 15106 9324 15108 9344
rect 15108 9324 15160 9344
rect 15160 9324 15162 9344
rect 15106 9288 15162 9324
rect 13082 2080 13138 2136
rect 13449 2202 13505 2204
rect 13529 2202 13585 2204
rect 13609 2202 13665 2204
rect 13689 2202 13745 2204
rect 13449 2150 13475 2202
rect 13475 2150 13505 2202
rect 13529 2150 13539 2202
rect 13539 2150 13585 2202
rect 13609 2150 13655 2202
rect 13655 2150 13665 2202
rect 13689 2150 13719 2202
rect 13719 2150 13745 2202
rect 13449 2148 13505 2150
rect 13529 2148 13585 2150
rect 13609 2148 13665 2150
rect 13689 2148 13745 2150
rect 15198 8492 15254 8528
rect 15198 8472 15200 8492
rect 15200 8472 15252 8492
rect 15252 8472 15254 8492
rect 15658 9988 15714 10024
rect 15658 9968 15660 9988
rect 15660 9968 15712 9988
rect 15712 9968 15714 9988
rect 15474 9444 15530 9480
rect 15474 9424 15476 9444
rect 15476 9424 15528 9444
rect 15528 9424 15530 9444
rect 15658 3304 15714 3360
rect 1674 448 1730 504
<< metal3 >>
rect 0 19410 800 19440
rect 1393 19410 1459 19413
rect 0 19408 1459 19410
rect 0 19352 1398 19408
rect 1454 19352 1459 19408
rect 0 19350 1459 19352
rect 0 19320 800 19350
rect 1393 19347 1459 19350
rect 0 18458 800 18488
rect 2773 18458 2839 18461
rect 0 18456 2839 18458
rect 0 18400 2778 18456
rect 2834 18400 2839 18456
rect 0 18398 2839 18400
rect 0 18368 800 18398
rect 2773 18395 2839 18398
rect 3442 17440 3762 17441
rect 0 17370 800 17400
rect 3442 17376 3450 17440
rect 3514 17376 3530 17440
rect 3594 17376 3610 17440
rect 3674 17376 3690 17440
rect 3754 17376 3762 17440
rect 3442 17375 3762 17376
rect 8440 17440 8760 17441
rect 8440 17376 8448 17440
rect 8512 17376 8528 17440
rect 8592 17376 8608 17440
rect 8672 17376 8688 17440
rect 8752 17376 8760 17440
rect 8440 17375 8760 17376
rect 13437 17440 13757 17441
rect 13437 17376 13445 17440
rect 13509 17376 13525 17440
rect 13589 17376 13605 17440
rect 13669 17376 13685 17440
rect 13749 17376 13757 17440
rect 13437 17375 13757 17376
rect 1945 17370 2011 17373
rect 0 17368 2011 17370
rect 0 17312 1950 17368
rect 2006 17312 2011 17368
rect 0 17310 2011 17312
rect 0 17280 800 17310
rect 1945 17307 2011 17310
rect 5941 16896 6261 16897
rect 5941 16832 5949 16896
rect 6013 16832 6029 16896
rect 6093 16832 6109 16896
rect 6173 16832 6189 16896
rect 6253 16832 6261 16896
rect 5941 16831 6261 16832
rect 10938 16896 11258 16897
rect 10938 16832 10946 16896
rect 11010 16832 11026 16896
rect 11090 16832 11106 16896
rect 11170 16832 11186 16896
rect 11250 16832 11258 16896
rect 10938 16831 11258 16832
rect 14917 16690 14983 16693
rect 15653 16690 15719 16693
rect 16400 16690 17200 16720
rect 14917 16688 17200 16690
rect 14917 16632 14922 16688
rect 14978 16632 15658 16688
rect 15714 16632 17200 16688
rect 14917 16630 17200 16632
rect 14917 16627 14983 16630
rect 15653 16627 15719 16630
rect 16400 16600 17200 16630
rect 9765 16554 9831 16557
rect 9990 16554 9996 16556
rect 9765 16552 9996 16554
rect 9765 16496 9770 16552
rect 9826 16496 9996 16552
rect 9765 16494 9996 16496
rect 9765 16491 9831 16494
rect 9990 16492 9996 16494
rect 10060 16492 10066 16556
rect 0 16418 800 16448
rect 1485 16418 1551 16421
rect 0 16416 1551 16418
rect 0 16360 1490 16416
rect 1546 16360 1551 16416
rect 0 16358 1551 16360
rect 0 16328 800 16358
rect 1485 16355 1551 16358
rect 3877 16418 3943 16421
rect 6494 16418 6500 16420
rect 3877 16416 6500 16418
rect 3877 16360 3882 16416
rect 3938 16360 6500 16416
rect 3877 16358 6500 16360
rect 3877 16355 3943 16358
rect 6494 16356 6500 16358
rect 6564 16356 6570 16420
rect 3442 16352 3762 16353
rect 3442 16288 3450 16352
rect 3514 16288 3530 16352
rect 3594 16288 3610 16352
rect 3674 16288 3690 16352
rect 3754 16288 3762 16352
rect 3442 16287 3762 16288
rect 8440 16352 8760 16353
rect 8440 16288 8448 16352
rect 8512 16288 8528 16352
rect 8592 16288 8608 16352
rect 8672 16288 8688 16352
rect 8752 16288 8760 16352
rect 8440 16287 8760 16288
rect 13437 16352 13757 16353
rect 13437 16288 13445 16352
rect 13509 16288 13525 16352
rect 13589 16288 13605 16352
rect 13669 16288 13685 16352
rect 13749 16288 13757 16352
rect 13437 16287 13757 16288
rect 9489 15874 9555 15877
rect 9622 15874 9628 15876
rect 9489 15872 9628 15874
rect 9489 15816 9494 15872
rect 9550 15816 9628 15872
rect 9489 15814 9628 15816
rect 9489 15811 9555 15814
rect 9622 15812 9628 15814
rect 9692 15812 9698 15876
rect 5941 15808 6261 15809
rect 5941 15744 5949 15808
rect 6013 15744 6029 15808
rect 6093 15744 6109 15808
rect 6173 15744 6189 15808
rect 6253 15744 6261 15808
rect 5941 15743 6261 15744
rect 10938 15808 11258 15809
rect 10938 15744 10946 15808
rect 11010 15744 11026 15808
rect 11090 15744 11106 15808
rect 11170 15744 11186 15808
rect 11250 15744 11258 15808
rect 10938 15743 11258 15744
rect 6729 15738 6795 15741
rect 8201 15738 8267 15741
rect 6729 15736 8267 15738
rect 6729 15680 6734 15736
rect 6790 15680 8206 15736
rect 8262 15680 8267 15736
rect 6729 15678 8267 15680
rect 6729 15675 6795 15678
rect 8201 15675 8267 15678
rect 0 15466 800 15496
rect 1393 15466 1459 15469
rect 0 15464 1459 15466
rect 0 15408 1398 15464
rect 1454 15408 1459 15464
rect 0 15406 1459 15408
rect 0 15376 800 15406
rect 1393 15403 1459 15406
rect 8201 15466 8267 15469
rect 10317 15466 10383 15469
rect 8201 15464 10383 15466
rect 8201 15408 8206 15464
rect 8262 15408 10322 15464
rect 10378 15408 10383 15464
rect 8201 15406 10383 15408
rect 8201 15403 8267 15406
rect 10317 15403 10383 15406
rect 3442 15264 3762 15265
rect 3442 15200 3450 15264
rect 3514 15200 3530 15264
rect 3594 15200 3610 15264
rect 3674 15200 3690 15264
rect 3754 15200 3762 15264
rect 3442 15199 3762 15200
rect 8440 15264 8760 15265
rect 8440 15200 8448 15264
rect 8512 15200 8528 15264
rect 8592 15200 8608 15264
rect 8672 15200 8688 15264
rect 8752 15200 8760 15264
rect 8440 15199 8760 15200
rect 13437 15264 13757 15265
rect 13437 15200 13445 15264
rect 13509 15200 13525 15264
rect 13589 15200 13605 15264
rect 13669 15200 13685 15264
rect 13749 15200 13757 15264
rect 13437 15199 13757 15200
rect 4613 15058 4679 15061
rect 8753 15058 8819 15061
rect 4613 15056 8819 15058
rect 4613 15000 4618 15056
rect 4674 15000 8758 15056
rect 8814 15000 8819 15056
rect 4613 14998 8819 15000
rect 4613 14995 4679 14998
rect 8753 14995 8819 14998
rect 9765 15058 9831 15061
rect 10358 15058 10364 15060
rect 9765 15056 10364 15058
rect 9765 15000 9770 15056
rect 9826 15000 10364 15056
rect 9765 14998 10364 15000
rect 9765 14995 9831 14998
rect 10358 14996 10364 14998
rect 10428 14996 10434 15060
rect 5941 14720 6261 14721
rect 5941 14656 5949 14720
rect 6013 14656 6029 14720
rect 6093 14656 6109 14720
rect 6173 14656 6189 14720
rect 6253 14656 6261 14720
rect 5941 14655 6261 14656
rect 10938 14720 11258 14721
rect 10938 14656 10946 14720
rect 11010 14656 11026 14720
rect 11090 14656 11106 14720
rect 11170 14656 11186 14720
rect 11250 14656 11258 14720
rect 10938 14655 11258 14656
rect 0 14378 800 14408
rect 1393 14378 1459 14381
rect 0 14376 1459 14378
rect 0 14320 1398 14376
rect 1454 14320 1459 14376
rect 0 14318 1459 14320
rect 0 14288 800 14318
rect 1393 14315 1459 14318
rect 6729 14378 6795 14381
rect 7833 14378 7899 14381
rect 9673 14378 9739 14381
rect 6729 14376 9739 14378
rect 6729 14320 6734 14376
rect 6790 14320 7838 14376
rect 7894 14320 9678 14376
rect 9734 14320 9739 14376
rect 6729 14318 9739 14320
rect 6729 14315 6795 14318
rect 7833 14315 7899 14318
rect 9673 14315 9739 14318
rect 3442 14176 3762 14177
rect 3442 14112 3450 14176
rect 3514 14112 3530 14176
rect 3594 14112 3610 14176
rect 3674 14112 3690 14176
rect 3754 14112 3762 14176
rect 3442 14111 3762 14112
rect 8440 14176 8760 14177
rect 8440 14112 8448 14176
rect 8512 14112 8528 14176
rect 8592 14112 8608 14176
rect 8672 14112 8688 14176
rect 8752 14112 8760 14176
rect 8440 14111 8760 14112
rect 13437 14176 13757 14177
rect 13437 14112 13445 14176
rect 13509 14112 13525 14176
rect 13589 14112 13605 14176
rect 13669 14112 13685 14176
rect 13749 14112 13757 14176
rect 13437 14111 13757 14112
rect 5809 13972 5875 13973
rect 5758 13970 5764 13972
rect 5682 13910 5764 13970
rect 5828 13970 5875 13972
rect 9121 13970 9187 13973
rect 9673 13970 9739 13973
rect 9806 13970 9812 13972
rect 5828 13968 9552 13970
rect 5870 13912 9126 13968
rect 9182 13912 9552 13968
rect 5758 13908 5764 13910
rect 5828 13910 9552 13912
rect 5828 13908 5875 13910
rect 5809 13907 5875 13908
rect 9121 13907 9187 13910
rect 9492 13837 9552 13910
rect 9673 13968 9812 13970
rect 9673 13912 9678 13968
rect 9734 13912 9812 13968
rect 9673 13910 9812 13912
rect 9673 13907 9739 13910
rect 9806 13908 9812 13910
rect 9876 13908 9882 13972
rect 3417 13834 3483 13837
rect 7189 13834 7255 13837
rect 3417 13832 7255 13834
rect 3417 13776 3422 13832
rect 3478 13776 7194 13832
rect 7250 13776 7255 13832
rect 3417 13774 7255 13776
rect 3417 13771 3483 13774
rect 7189 13771 7255 13774
rect 8477 13834 8543 13837
rect 9305 13834 9371 13837
rect 8477 13832 9371 13834
rect 8477 13776 8482 13832
rect 8538 13776 9310 13832
rect 9366 13776 9371 13832
rect 8477 13774 9371 13776
rect 8477 13771 8543 13774
rect 9305 13771 9371 13774
rect 9489 13834 9555 13837
rect 10409 13834 10475 13837
rect 9489 13832 10475 13834
rect 9489 13776 9494 13832
rect 9550 13776 10414 13832
rect 10470 13776 10475 13832
rect 9489 13774 10475 13776
rect 9489 13771 9555 13774
rect 10409 13771 10475 13774
rect 8201 13700 8267 13701
rect 8150 13636 8156 13700
rect 8220 13698 8267 13700
rect 9029 13698 9095 13701
rect 9673 13698 9739 13701
rect 8220 13696 8312 13698
rect 8262 13640 8312 13696
rect 8220 13638 8312 13640
rect 9029 13696 9739 13698
rect 9029 13640 9034 13696
rect 9090 13640 9678 13696
rect 9734 13640 9739 13696
rect 9029 13638 9739 13640
rect 8220 13636 8267 13638
rect 8201 13635 8267 13636
rect 9029 13635 9095 13638
rect 9673 13635 9739 13638
rect 5941 13632 6261 13633
rect 5941 13568 5949 13632
rect 6013 13568 6029 13632
rect 6093 13568 6109 13632
rect 6173 13568 6189 13632
rect 6253 13568 6261 13632
rect 5941 13567 6261 13568
rect 10938 13632 11258 13633
rect 10938 13568 10946 13632
rect 11010 13568 11026 13632
rect 11090 13568 11106 13632
rect 11170 13568 11186 13632
rect 11250 13568 11258 13632
rect 10938 13567 11258 13568
rect 7465 13562 7531 13565
rect 9121 13562 9187 13565
rect 7465 13560 9187 13562
rect 7465 13504 7470 13560
rect 7526 13504 9126 13560
rect 9182 13504 9187 13560
rect 7465 13502 9187 13504
rect 7465 13499 7531 13502
rect 9121 13499 9187 13502
rect 0 13426 800 13456
rect 1393 13426 1459 13429
rect 0 13424 1459 13426
rect 0 13368 1398 13424
rect 1454 13368 1459 13424
rect 0 13366 1459 13368
rect 0 13336 800 13366
rect 1393 13363 1459 13366
rect 3141 13426 3207 13429
rect 3141 13424 8218 13426
rect 3141 13368 3146 13424
rect 3202 13368 8218 13424
rect 3141 13366 8218 13368
rect 3141 13363 3207 13366
rect 4705 13290 4771 13293
rect 8017 13290 8083 13293
rect 4705 13288 8083 13290
rect 4705 13232 4710 13288
rect 4766 13232 8022 13288
rect 8078 13232 8083 13288
rect 4705 13230 8083 13232
rect 8158 13290 8218 13366
rect 9305 13290 9371 13293
rect 8158 13288 9371 13290
rect 8158 13232 9310 13288
rect 9366 13232 9371 13288
rect 8158 13230 9371 13232
rect 4705 13227 4771 13230
rect 8017 13227 8083 13230
rect 9305 13227 9371 13230
rect 9765 13290 9831 13293
rect 14038 13290 14044 13292
rect 9765 13288 14044 13290
rect 9765 13232 9770 13288
rect 9826 13232 14044 13288
rect 9765 13230 14044 13232
rect 9765 13227 9831 13230
rect 14038 13228 14044 13230
rect 14108 13228 14114 13292
rect 4061 13154 4127 13157
rect 7373 13154 7439 13157
rect 4061 13152 7439 13154
rect 4061 13096 4066 13152
rect 4122 13096 7378 13152
rect 7434 13096 7439 13152
rect 4061 13094 7439 13096
rect 4061 13091 4127 13094
rect 7373 13091 7439 13094
rect 11145 13154 11211 13157
rect 11462 13154 11468 13156
rect 11145 13152 11468 13154
rect 11145 13096 11150 13152
rect 11206 13096 11468 13152
rect 11145 13094 11468 13096
rect 11145 13091 11211 13094
rect 11462 13092 11468 13094
rect 11532 13092 11538 13156
rect 3442 13088 3762 13089
rect 3442 13024 3450 13088
rect 3514 13024 3530 13088
rect 3594 13024 3610 13088
rect 3674 13024 3690 13088
rect 3754 13024 3762 13088
rect 3442 13023 3762 13024
rect 8440 13088 8760 13089
rect 8440 13024 8448 13088
rect 8512 13024 8528 13088
rect 8592 13024 8608 13088
rect 8672 13024 8688 13088
rect 8752 13024 8760 13088
rect 8440 13023 8760 13024
rect 13437 13088 13757 13089
rect 13437 13024 13445 13088
rect 13509 13024 13525 13088
rect 13589 13024 13605 13088
rect 13669 13024 13685 13088
rect 13749 13024 13757 13088
rect 13437 13023 13757 13024
rect 10685 13018 10751 13021
rect 11646 13018 11652 13020
rect 10685 13016 11652 13018
rect 10685 12960 10690 13016
rect 10746 12960 11652 13016
rect 10685 12958 11652 12960
rect 10685 12955 10751 12958
rect 11646 12956 11652 12958
rect 11716 12956 11722 13020
rect 3509 12882 3575 12885
rect 5717 12882 5783 12885
rect 3509 12880 5783 12882
rect 3509 12824 3514 12880
rect 3570 12824 5722 12880
rect 5778 12824 5783 12880
rect 3509 12822 5783 12824
rect 3509 12819 3575 12822
rect 5717 12819 5783 12822
rect 7005 12882 7071 12885
rect 9121 12882 9187 12885
rect 7005 12880 9187 12882
rect 7005 12824 7010 12880
rect 7066 12824 9126 12880
rect 9182 12824 9187 12880
rect 7005 12822 9187 12824
rect 7005 12819 7071 12822
rect 9121 12819 9187 12822
rect 9857 12882 9923 12885
rect 10869 12882 10935 12885
rect 9857 12880 10935 12882
rect 9857 12824 9862 12880
rect 9918 12824 10874 12880
rect 10930 12824 10935 12880
rect 9857 12822 10935 12824
rect 9857 12819 9923 12822
rect 10869 12819 10935 12822
rect 11973 12884 12039 12885
rect 11973 12880 12020 12884
rect 12084 12882 12090 12884
rect 11973 12824 11978 12880
rect 11973 12820 12020 12824
rect 12084 12822 12130 12882
rect 12084 12820 12090 12822
rect 11973 12819 12039 12820
rect 4797 12746 4863 12749
rect 6913 12746 6979 12749
rect 9857 12746 9923 12749
rect 4797 12744 6979 12746
rect 4797 12688 4802 12744
rect 4858 12688 6918 12744
rect 6974 12688 6979 12744
rect 4797 12686 6979 12688
rect 4797 12683 4863 12686
rect 6913 12683 6979 12686
rect 8940 12744 9923 12746
rect 8940 12688 9862 12744
rect 9918 12688 9923 12744
rect 8940 12686 9923 12688
rect 8940 12613 9000 12686
rect 9857 12683 9923 12686
rect 10542 12684 10548 12748
rect 10612 12746 10618 12748
rect 12249 12746 12315 12749
rect 10612 12744 12315 12746
rect 10612 12688 12254 12744
rect 12310 12688 12315 12744
rect 10612 12686 12315 12688
rect 10612 12684 10618 12686
rect 12249 12683 12315 12686
rect 2405 12610 2471 12613
rect 4521 12610 4587 12613
rect 2405 12608 4587 12610
rect 2405 12552 2410 12608
rect 2466 12552 4526 12608
rect 4582 12552 4587 12608
rect 2405 12550 4587 12552
rect 2405 12547 2471 12550
rect 4521 12547 4587 12550
rect 6361 12610 6427 12613
rect 8937 12610 9003 12613
rect 6361 12608 9003 12610
rect 6361 12552 6366 12608
rect 6422 12552 8942 12608
rect 8998 12552 9003 12608
rect 6361 12550 9003 12552
rect 6361 12547 6427 12550
rect 8937 12547 9003 12550
rect 9121 12610 9187 12613
rect 9806 12610 9812 12612
rect 9121 12608 9812 12610
rect 9121 12552 9126 12608
rect 9182 12552 9812 12608
rect 9121 12550 9812 12552
rect 9121 12547 9187 12550
rect 9806 12548 9812 12550
rect 9876 12610 9882 12612
rect 10593 12610 10659 12613
rect 9876 12608 10659 12610
rect 9876 12552 10598 12608
rect 10654 12552 10659 12608
rect 9876 12550 10659 12552
rect 9876 12548 9882 12550
rect 10593 12547 10659 12550
rect 5941 12544 6261 12545
rect 0 12474 800 12504
rect 5941 12480 5949 12544
rect 6013 12480 6029 12544
rect 6093 12480 6109 12544
rect 6173 12480 6189 12544
rect 6253 12480 6261 12544
rect 5941 12479 6261 12480
rect 10938 12544 11258 12545
rect 10938 12480 10946 12544
rect 11010 12480 11026 12544
rect 11090 12480 11106 12544
rect 11170 12480 11186 12544
rect 11250 12480 11258 12544
rect 10938 12479 11258 12480
rect 1393 12474 1459 12477
rect 0 12472 1459 12474
rect 0 12416 1398 12472
rect 1454 12416 1459 12472
rect 0 12414 1459 12416
rect 0 12384 800 12414
rect 1393 12411 1459 12414
rect 8753 12474 8819 12477
rect 10685 12474 10751 12477
rect 8753 12472 10751 12474
rect 8753 12416 8758 12472
rect 8814 12416 10690 12472
rect 10746 12416 10751 12472
rect 8753 12414 10751 12416
rect 8753 12411 8819 12414
rect 10685 12411 10751 12414
rect 2865 12338 2931 12341
rect 3233 12338 3299 12341
rect 2865 12336 3299 12338
rect 2865 12280 2870 12336
rect 2926 12280 3238 12336
rect 3294 12280 3299 12336
rect 2865 12278 3299 12280
rect 2865 12275 2931 12278
rect 3233 12275 3299 12278
rect 4061 12338 4127 12341
rect 9857 12338 9923 12341
rect 9990 12338 9996 12340
rect 4061 12336 8908 12338
rect 4061 12280 4066 12336
rect 4122 12280 8908 12336
rect 4061 12278 8908 12280
rect 4061 12275 4127 12278
rect 3233 12202 3299 12205
rect 7925 12202 7991 12205
rect 3233 12200 7991 12202
rect 3233 12144 3238 12200
rect 3294 12144 7930 12200
rect 7986 12144 7991 12200
rect 3233 12142 7991 12144
rect 3233 12139 3299 12142
rect 7925 12139 7991 12142
rect 8848 12066 8908 12278
rect 9857 12336 9996 12338
rect 9857 12280 9862 12336
rect 9918 12280 9996 12336
rect 9857 12278 9996 12280
rect 9857 12275 9923 12278
rect 9990 12276 9996 12278
rect 10060 12276 10066 12340
rect 12934 12276 12940 12340
rect 13004 12338 13010 12340
rect 13077 12338 13143 12341
rect 13004 12336 13143 12338
rect 13004 12280 13082 12336
rect 13138 12280 13143 12336
rect 13004 12278 13143 12280
rect 13004 12276 13010 12278
rect 13077 12275 13143 12278
rect 10041 12202 10107 12205
rect 11421 12202 11487 12205
rect 10041 12200 11487 12202
rect 10041 12144 10046 12200
rect 10102 12144 11426 12200
rect 11482 12144 11487 12200
rect 10041 12142 11487 12144
rect 10041 12139 10107 12142
rect 11421 12139 11487 12142
rect 11053 12066 11119 12069
rect 8848 12064 11119 12066
rect 8848 12008 11058 12064
rect 11114 12008 11119 12064
rect 8848 12006 11119 12008
rect 11053 12003 11119 12006
rect 3442 12000 3762 12001
rect 3442 11936 3450 12000
rect 3514 11936 3530 12000
rect 3594 11936 3610 12000
rect 3674 11936 3690 12000
rect 3754 11936 3762 12000
rect 3442 11935 3762 11936
rect 8440 12000 8760 12001
rect 8440 11936 8448 12000
rect 8512 11936 8528 12000
rect 8592 11936 8608 12000
rect 8672 11936 8688 12000
rect 8752 11936 8760 12000
rect 8440 11935 8760 11936
rect 13437 12000 13757 12001
rect 13437 11936 13445 12000
rect 13509 11936 13525 12000
rect 13589 11936 13605 12000
rect 13669 11936 13685 12000
rect 13749 11936 13757 12000
rect 13437 11935 13757 11936
rect 4337 11930 4403 11933
rect 5441 11930 5507 11933
rect 4337 11928 5507 11930
rect 4337 11872 4342 11928
rect 4398 11872 5446 11928
rect 5502 11872 5507 11928
rect 4337 11870 5507 11872
rect 4337 11867 4403 11870
rect 5441 11867 5507 11870
rect 10685 11930 10751 11933
rect 12525 11930 12591 11933
rect 10685 11928 12591 11930
rect 10685 11872 10690 11928
rect 10746 11872 12530 11928
rect 12586 11872 12591 11928
rect 10685 11870 12591 11872
rect 10685 11867 10751 11870
rect 12525 11867 12591 11870
rect 2405 11794 2471 11797
rect 11421 11794 11487 11797
rect 2405 11792 11487 11794
rect 2405 11736 2410 11792
rect 2466 11736 11426 11792
rect 11482 11736 11487 11792
rect 2405 11734 11487 11736
rect 2405 11731 2471 11734
rect 11421 11731 11487 11734
rect 1945 11658 2011 11661
rect 12433 11658 12499 11661
rect 1945 11656 12499 11658
rect 1945 11600 1950 11656
rect 2006 11600 12438 11656
rect 12494 11600 12499 11656
rect 1945 11598 12499 11600
rect 1945 11595 2011 11598
rect 12433 11595 12499 11598
rect 6729 11522 6795 11525
rect 9029 11522 9095 11525
rect 6729 11520 9095 11522
rect 6729 11464 6734 11520
rect 6790 11464 9034 11520
rect 9090 11464 9095 11520
rect 6729 11462 9095 11464
rect 6729 11459 6795 11462
rect 9029 11459 9095 11462
rect 10358 11460 10364 11524
rect 10428 11522 10434 11524
rect 10685 11522 10751 11525
rect 10428 11520 10751 11522
rect 10428 11464 10690 11520
rect 10746 11464 10751 11520
rect 10428 11462 10751 11464
rect 10428 11460 10434 11462
rect 10685 11459 10751 11462
rect 5941 11456 6261 11457
rect 0 11386 800 11416
rect 5941 11392 5949 11456
rect 6013 11392 6029 11456
rect 6093 11392 6109 11456
rect 6173 11392 6189 11456
rect 6253 11392 6261 11456
rect 5941 11391 6261 11392
rect 10938 11456 11258 11457
rect 10938 11392 10946 11456
rect 11010 11392 11026 11456
rect 11090 11392 11106 11456
rect 11170 11392 11186 11456
rect 11250 11392 11258 11456
rect 10938 11391 11258 11392
rect 1485 11386 1551 11389
rect 0 11384 1551 11386
rect 0 11328 1490 11384
rect 1546 11328 1551 11384
rect 0 11326 1551 11328
rect 0 11296 800 11326
rect 1485 11323 1551 11326
rect 9949 11386 10015 11389
rect 10685 11386 10751 11389
rect 9949 11384 10751 11386
rect 9949 11328 9954 11384
rect 10010 11328 10690 11384
rect 10746 11328 10751 11384
rect 9949 11326 10751 11328
rect 9949 11323 10015 11326
rect 10685 11323 10751 11326
rect 11513 11386 11579 11389
rect 12198 11386 12204 11388
rect 11513 11384 12204 11386
rect 11513 11328 11518 11384
rect 11574 11328 12204 11384
rect 11513 11326 12204 11328
rect 11513 11323 11579 11326
rect 12198 11324 12204 11326
rect 12268 11324 12274 11388
rect 5257 11250 5323 11253
rect 12249 11250 12315 11253
rect 5257 11248 12315 11250
rect 5257 11192 5262 11248
rect 5318 11192 12254 11248
rect 12310 11192 12315 11248
rect 5257 11190 12315 11192
rect 5257 11187 5323 11190
rect 12249 11187 12315 11190
rect 5165 11114 5231 11117
rect 8109 11114 8175 11117
rect 5165 11112 8175 11114
rect 5165 11056 5170 11112
rect 5226 11056 8114 11112
rect 8170 11056 8175 11112
rect 5165 11054 8175 11056
rect 5165 11051 5231 11054
rect 8109 11051 8175 11054
rect 9489 11112 9555 11117
rect 9489 11056 9494 11112
rect 9550 11056 9555 11112
rect 9489 11051 9555 11056
rect 10726 11052 10732 11116
rect 10796 11114 10802 11116
rect 11605 11114 11671 11117
rect 10796 11112 11671 11114
rect 10796 11056 11610 11112
rect 11666 11056 11671 11112
rect 10796 11054 11671 11056
rect 10796 11052 10802 11054
rect 11605 11051 11671 11054
rect 12709 11116 12775 11117
rect 12709 11112 12756 11116
rect 12820 11114 12826 11116
rect 12709 11056 12714 11112
rect 12709 11052 12756 11056
rect 12820 11054 12866 11114
rect 12820 11052 12826 11054
rect 12709 11051 12775 11052
rect 9492 10978 9552 11051
rect 10409 10978 10475 10981
rect 11830 10978 11836 10980
rect 9492 10918 10288 10978
rect 3442 10912 3762 10913
rect 3442 10848 3450 10912
rect 3514 10848 3530 10912
rect 3594 10848 3610 10912
rect 3674 10848 3690 10912
rect 3754 10848 3762 10912
rect 3442 10847 3762 10848
rect 8440 10912 8760 10913
rect 8440 10848 8448 10912
rect 8512 10848 8528 10912
rect 8592 10848 8608 10912
rect 8672 10848 8688 10912
rect 8752 10848 8760 10912
rect 8440 10847 8760 10848
rect 9622 10780 9628 10844
rect 9692 10842 9698 10844
rect 9765 10842 9831 10845
rect 9692 10840 9831 10842
rect 9692 10784 9770 10840
rect 9826 10784 9831 10840
rect 9692 10782 9831 10784
rect 10228 10842 10288 10918
rect 10409 10976 11836 10978
rect 10409 10920 10414 10976
rect 10470 10920 11836 10976
rect 10409 10918 11836 10920
rect 10409 10915 10475 10918
rect 11830 10916 11836 10918
rect 11900 10916 11906 10980
rect 12065 10978 12131 10981
rect 12249 10978 12315 10981
rect 12065 10976 12315 10978
rect 12065 10920 12070 10976
rect 12126 10920 12254 10976
rect 12310 10920 12315 10976
rect 12065 10918 12315 10920
rect 12065 10915 12131 10918
rect 12249 10915 12315 10918
rect 13437 10912 13757 10913
rect 13437 10848 13445 10912
rect 13509 10848 13525 10912
rect 13589 10848 13605 10912
rect 13669 10848 13685 10912
rect 13749 10848 13757 10912
rect 13437 10847 13757 10848
rect 13118 10842 13124 10844
rect 10228 10782 13124 10842
rect 9692 10780 9698 10782
rect 9765 10779 9831 10782
rect 13118 10780 13124 10782
rect 13188 10842 13194 10844
rect 13261 10842 13327 10845
rect 13188 10840 13327 10842
rect 13188 10784 13266 10840
rect 13322 10784 13327 10840
rect 13188 10782 13327 10784
rect 13188 10780 13194 10782
rect 13261 10779 13327 10782
rect 9305 10706 9371 10709
rect 11513 10706 11579 10709
rect 13445 10706 13511 10709
rect 9305 10704 13511 10706
rect 9305 10648 9310 10704
rect 9366 10648 11518 10704
rect 11574 10648 13450 10704
rect 13506 10648 13511 10704
rect 9305 10646 13511 10648
rect 9305 10643 9371 10646
rect 11513 10643 11579 10646
rect 13445 10643 13511 10646
rect 2681 10570 2747 10573
rect 4337 10570 4403 10573
rect 10869 10570 10935 10573
rect 2681 10568 4403 10570
rect 2681 10512 2686 10568
rect 2742 10512 4342 10568
rect 4398 10512 4403 10568
rect 2681 10510 4403 10512
rect 2681 10507 2747 10510
rect 4337 10507 4403 10510
rect 10412 10568 10935 10570
rect 10412 10512 10874 10568
rect 10930 10512 10935 10568
rect 10412 10510 10935 10512
rect 0 10434 800 10464
rect 10412 10437 10472 10510
rect 10869 10507 10935 10510
rect 11237 10570 11303 10573
rect 11462 10570 11468 10572
rect 11237 10568 11468 10570
rect 11237 10512 11242 10568
rect 11298 10512 11468 10568
rect 11237 10510 11468 10512
rect 11237 10507 11303 10510
rect 11462 10508 11468 10510
rect 11532 10508 11538 10572
rect 1485 10434 1551 10437
rect 0 10432 1551 10434
rect 0 10376 1490 10432
rect 1546 10376 1551 10432
rect 0 10374 1551 10376
rect 0 10344 800 10374
rect 1485 10371 1551 10374
rect 7741 10434 7807 10437
rect 8845 10434 8911 10437
rect 7741 10432 8911 10434
rect 7741 10376 7746 10432
rect 7802 10376 8850 10432
rect 8906 10376 8911 10432
rect 7741 10374 8911 10376
rect 7741 10371 7807 10374
rect 8845 10371 8911 10374
rect 10409 10432 10475 10437
rect 10409 10376 10414 10432
rect 10470 10376 10475 10432
rect 10409 10371 10475 10376
rect 12065 10434 12131 10437
rect 13905 10434 13971 10437
rect 12065 10432 13971 10434
rect 12065 10376 12070 10432
rect 12126 10376 13910 10432
rect 13966 10376 13971 10432
rect 12065 10374 13971 10376
rect 12065 10371 12131 10374
rect 13905 10371 13971 10374
rect 5941 10368 6261 10369
rect 5941 10304 5949 10368
rect 6013 10304 6029 10368
rect 6093 10304 6109 10368
rect 6173 10304 6189 10368
rect 6253 10304 6261 10368
rect 5941 10303 6261 10304
rect 10938 10368 11258 10369
rect 10938 10304 10946 10368
rect 11010 10304 11026 10368
rect 11090 10304 11106 10368
rect 11170 10304 11186 10368
rect 11250 10304 11258 10368
rect 10938 10303 11258 10304
rect 7189 10298 7255 10301
rect 8845 10298 8911 10301
rect 7189 10296 8911 10298
rect 7189 10240 7194 10296
rect 7250 10240 8850 10296
rect 8906 10240 8911 10296
rect 7189 10238 8911 10240
rect 7189 10235 7255 10238
rect 8845 10235 8911 10238
rect 12249 10298 12315 10301
rect 12249 10296 12588 10298
rect 12249 10240 12254 10296
rect 12310 10240 12588 10296
rect 12249 10238 12588 10240
rect 12249 10235 12315 10238
rect 4521 10162 4587 10165
rect 6361 10162 6427 10165
rect 4521 10160 6427 10162
rect 4521 10104 4526 10160
rect 4582 10104 6366 10160
rect 6422 10104 6427 10160
rect 4521 10102 6427 10104
rect 4521 10099 4587 10102
rect 6361 10099 6427 10102
rect 6821 10162 6887 10165
rect 8150 10162 8156 10164
rect 6821 10160 8156 10162
rect 6821 10104 6826 10160
rect 6882 10104 8156 10160
rect 6821 10102 8156 10104
rect 6821 10099 6887 10102
rect 8150 10100 8156 10102
rect 8220 10162 8226 10164
rect 9397 10162 9463 10165
rect 12382 10162 12388 10164
rect 8220 10160 12388 10162
rect 8220 10104 9402 10160
rect 9458 10104 12388 10160
rect 8220 10102 12388 10104
rect 8220 10100 8226 10102
rect 9397 10099 9463 10102
rect 12382 10100 12388 10102
rect 12452 10100 12458 10164
rect 12528 10162 12588 10238
rect 12934 10236 12940 10300
rect 13004 10298 13010 10300
rect 13721 10298 13787 10301
rect 13004 10296 13787 10298
rect 13004 10240 13726 10296
rect 13782 10240 13787 10296
rect 13004 10238 13787 10240
rect 13004 10236 13010 10238
rect 13721 10235 13787 10238
rect 13169 10162 13235 10165
rect 12528 10160 13235 10162
rect 12528 10104 13174 10160
rect 13230 10104 13235 10160
rect 12528 10102 13235 10104
rect 13169 10099 13235 10102
rect 2221 10026 2287 10029
rect 14365 10026 14431 10029
rect 2221 10024 14431 10026
rect 2221 9968 2226 10024
rect 2282 9968 14370 10024
rect 14426 9968 14431 10024
rect 2221 9966 14431 9968
rect 2221 9963 2287 9966
rect 14365 9963 14431 9966
rect 15653 10026 15719 10029
rect 16400 10026 17200 10056
rect 15653 10024 17200 10026
rect 15653 9968 15658 10024
rect 15714 9968 17200 10024
rect 15653 9966 17200 9968
rect 15653 9963 15719 9966
rect 16400 9936 17200 9966
rect 10777 9892 10843 9893
rect 10726 9890 10732 9892
rect 10686 9830 10732 9890
rect 10796 9888 10843 9892
rect 10838 9832 10843 9888
rect 10726 9828 10732 9830
rect 10796 9828 10843 9832
rect 10777 9827 10843 9828
rect 11421 9890 11487 9893
rect 11881 9890 11947 9893
rect 11421 9888 11947 9890
rect 11421 9832 11426 9888
rect 11482 9832 11886 9888
rect 11942 9832 11947 9888
rect 11421 9830 11947 9832
rect 11421 9827 11487 9830
rect 11881 9827 11947 9830
rect 12065 9890 12131 9893
rect 12198 9890 12204 9892
rect 12065 9888 12204 9890
rect 12065 9832 12070 9888
rect 12126 9832 12204 9888
rect 12065 9830 12204 9832
rect 12065 9827 12131 9830
rect 12198 9828 12204 9830
rect 12268 9890 12274 9892
rect 12433 9890 12499 9893
rect 12268 9888 12499 9890
rect 12268 9832 12438 9888
rect 12494 9832 12499 9888
rect 12268 9830 12499 9832
rect 12268 9828 12274 9830
rect 12433 9827 12499 9830
rect 3442 9824 3762 9825
rect 3442 9760 3450 9824
rect 3514 9760 3530 9824
rect 3594 9760 3610 9824
rect 3674 9760 3690 9824
rect 3754 9760 3762 9824
rect 3442 9759 3762 9760
rect 8440 9824 8760 9825
rect 8440 9760 8448 9824
rect 8512 9760 8528 9824
rect 8592 9760 8608 9824
rect 8672 9760 8688 9824
rect 8752 9760 8760 9824
rect 8440 9759 8760 9760
rect 13437 9824 13757 9825
rect 13437 9760 13445 9824
rect 13509 9760 13525 9824
rect 13589 9760 13605 9824
rect 13669 9760 13685 9824
rect 13749 9760 13757 9824
rect 13437 9759 13757 9760
rect 4153 9754 4219 9757
rect 7189 9754 7255 9757
rect 3880 9752 7255 9754
rect 3880 9696 4158 9752
rect 4214 9696 7194 9752
rect 7250 9696 7255 9752
rect 3880 9694 7255 9696
rect 3049 9620 3115 9621
rect 2998 9618 3004 9620
rect 2958 9558 3004 9618
rect 3068 9616 3115 9620
rect 3110 9560 3115 9616
rect 2998 9556 3004 9558
rect 3068 9556 3115 9560
rect 3049 9555 3115 9556
rect 3233 9618 3299 9621
rect 3880 9618 3940 9694
rect 4153 9691 4219 9694
rect 7189 9691 7255 9694
rect 9121 9754 9187 9757
rect 9121 9752 13370 9754
rect 9121 9696 9126 9752
rect 9182 9696 13370 9752
rect 9121 9694 13370 9696
rect 9121 9691 9187 9694
rect 3233 9616 3940 9618
rect 3233 9560 3238 9616
rect 3294 9560 3940 9616
rect 3233 9558 3940 9560
rect 5625 9618 5691 9621
rect 11697 9618 11763 9621
rect 5625 9616 11763 9618
rect 5625 9560 5630 9616
rect 5686 9560 11702 9616
rect 11758 9560 11763 9616
rect 5625 9558 11763 9560
rect 3233 9555 3299 9558
rect 5625 9555 5691 9558
rect 11697 9555 11763 9558
rect 12617 9618 12683 9621
rect 12801 9618 12867 9621
rect 12617 9616 12867 9618
rect 12617 9560 12622 9616
rect 12678 9560 12806 9616
rect 12862 9560 12867 9616
rect 12617 9558 12867 9560
rect 13310 9618 13370 9694
rect 13997 9618 14063 9621
rect 13310 9616 14063 9618
rect 13310 9560 14002 9616
rect 14058 9560 14063 9616
rect 13310 9558 14063 9560
rect 12617 9555 12683 9558
rect 12801 9555 12867 9558
rect 13997 9555 14063 9558
rect 0 9482 800 9512
rect 1393 9482 1459 9485
rect 0 9480 1459 9482
rect 0 9424 1398 9480
rect 1454 9424 1459 9480
rect 0 9422 1459 9424
rect 0 9392 800 9422
rect 1393 9419 1459 9422
rect 2589 9482 2655 9485
rect 8109 9482 8175 9485
rect 2589 9480 8034 9482
rect 2589 9424 2594 9480
rect 2650 9424 8034 9480
rect 2589 9422 8034 9424
rect 2589 9419 2655 9422
rect 1485 9346 1551 9349
rect 5533 9346 5599 9349
rect 1485 9344 5599 9346
rect 1485 9288 1490 9344
rect 1546 9288 5538 9344
rect 5594 9288 5599 9344
rect 1485 9286 5599 9288
rect 1485 9283 1551 9286
rect 5533 9283 5599 9286
rect 5941 9280 6261 9281
rect 5941 9216 5949 9280
rect 6013 9216 6029 9280
rect 6093 9216 6109 9280
rect 6173 9216 6189 9280
rect 6253 9216 6261 9280
rect 5941 9215 6261 9216
rect 2497 9210 2563 9213
rect 2497 9208 5826 9210
rect 2497 9152 2502 9208
rect 2558 9152 5826 9208
rect 2497 9150 5826 9152
rect 2497 9147 2563 9150
rect 2405 9074 2471 9077
rect 5625 9074 5691 9077
rect 2405 9072 5691 9074
rect 2405 9016 2410 9072
rect 2466 9016 5630 9072
rect 5686 9016 5691 9072
rect 2405 9014 5691 9016
rect 5766 9074 5826 9150
rect 7974 9074 8034 9422
rect 8109 9480 12450 9482
rect 8109 9424 8114 9480
rect 8170 9424 12450 9480
rect 8109 9422 12450 9424
rect 8109 9419 8175 9422
rect 9121 9346 9187 9349
rect 9673 9346 9739 9349
rect 10501 9346 10567 9349
rect 9121 9344 10567 9346
rect 9121 9288 9126 9344
rect 9182 9288 9678 9344
rect 9734 9288 10506 9344
rect 10562 9288 10567 9344
rect 9121 9286 10567 9288
rect 9121 9283 9187 9286
rect 9673 9283 9739 9286
rect 10501 9283 10567 9286
rect 11329 9346 11395 9349
rect 11881 9346 11947 9349
rect 11329 9344 11947 9346
rect 11329 9288 11334 9344
rect 11390 9288 11886 9344
rect 11942 9288 11947 9344
rect 11329 9286 11947 9288
rect 12390 9346 12450 9422
rect 12566 9420 12572 9484
rect 12636 9482 12642 9484
rect 12801 9482 12867 9485
rect 15469 9482 15535 9485
rect 12636 9480 15535 9482
rect 12636 9424 12806 9480
rect 12862 9424 15474 9480
rect 15530 9424 15535 9480
rect 12636 9422 15535 9424
rect 12636 9420 12642 9422
rect 12801 9419 12867 9422
rect 15469 9419 15535 9422
rect 15101 9346 15167 9349
rect 12390 9344 15167 9346
rect 12390 9288 15106 9344
rect 15162 9288 15167 9344
rect 12390 9286 15167 9288
rect 11329 9283 11395 9286
rect 11881 9283 11947 9286
rect 15101 9283 15167 9286
rect 10938 9280 11258 9281
rect 10938 9216 10946 9280
rect 11010 9216 11026 9280
rect 11090 9216 11106 9280
rect 11170 9216 11186 9280
rect 11250 9216 11258 9280
rect 10938 9215 11258 9216
rect 8109 9210 8175 9213
rect 9489 9210 9555 9213
rect 8109 9208 9555 9210
rect 8109 9152 8114 9208
rect 8170 9152 9494 9208
rect 9550 9152 9555 9208
rect 8109 9150 9555 9152
rect 8109 9147 8175 9150
rect 9489 9147 9555 9150
rect 9806 9148 9812 9212
rect 9876 9210 9882 9212
rect 10501 9210 10567 9213
rect 10685 9210 10751 9213
rect 9876 9208 10751 9210
rect 9876 9152 10506 9208
rect 10562 9152 10690 9208
rect 10746 9152 10751 9208
rect 9876 9150 10751 9152
rect 9876 9148 9882 9150
rect 10501 9147 10567 9150
rect 10685 9147 10751 9150
rect 11697 9210 11763 9213
rect 12157 9210 12223 9213
rect 12893 9212 12959 9213
rect 12893 9210 12940 9212
rect 11697 9208 12223 9210
rect 11697 9152 11702 9208
rect 11758 9152 12162 9208
rect 12218 9152 12223 9208
rect 11697 9150 12223 9152
rect 12848 9208 12940 9210
rect 12848 9152 12898 9208
rect 12848 9150 12940 9152
rect 11697 9147 11763 9150
rect 12157 9147 12223 9150
rect 12893 9148 12940 9150
rect 13004 9148 13010 9212
rect 13721 9210 13787 9213
rect 14038 9210 14044 9212
rect 13721 9208 14044 9210
rect 13721 9152 13726 9208
rect 13782 9152 14044 9208
rect 13721 9150 14044 9152
rect 12893 9147 12959 9148
rect 13721 9147 13787 9150
rect 14038 9148 14044 9150
rect 14108 9148 14114 9212
rect 12709 9074 12775 9077
rect 5766 9014 7850 9074
rect 7974 9072 12775 9074
rect 7974 9016 12714 9072
rect 12770 9016 12775 9072
rect 7974 9014 12775 9016
rect 2405 9011 2471 9014
rect 5625 9011 5691 9014
rect 2681 8938 2747 8941
rect 7281 8938 7347 8941
rect 2681 8936 7347 8938
rect 2681 8880 2686 8936
rect 2742 8880 7286 8936
rect 7342 8880 7347 8936
rect 2681 8878 7347 8880
rect 7790 8938 7850 9014
rect 12709 9011 12775 9014
rect 13537 9074 13603 9077
rect 13854 9074 13860 9076
rect 13537 9072 13860 9074
rect 13537 9016 13542 9072
rect 13598 9016 13860 9072
rect 13537 9014 13860 9016
rect 13537 9011 13603 9014
rect 13854 9012 13860 9014
rect 13924 9012 13930 9076
rect 13905 8938 13971 8941
rect 7790 8936 13971 8938
rect 7790 8880 13910 8936
rect 13966 8880 13971 8936
rect 7790 8878 13971 8880
rect 2681 8875 2747 8878
rect 7281 8875 7347 8878
rect 13905 8875 13971 8878
rect 14089 8936 14155 8941
rect 14089 8880 14094 8936
rect 14150 8880 14155 8936
rect 14089 8875 14155 8880
rect 5073 8802 5139 8805
rect 7465 8802 7531 8805
rect 8293 8802 8359 8805
rect 5073 8800 8359 8802
rect 5073 8744 5078 8800
rect 5134 8744 7470 8800
rect 7526 8744 8298 8800
rect 8354 8744 8359 8800
rect 5073 8742 8359 8744
rect 5073 8739 5139 8742
rect 7465 8739 7531 8742
rect 8293 8739 8359 8742
rect 10133 8802 10199 8805
rect 11973 8802 12039 8805
rect 10133 8800 12039 8802
rect 10133 8744 10138 8800
rect 10194 8744 11978 8800
rect 12034 8744 12039 8800
rect 10133 8742 12039 8744
rect 10133 8739 10199 8742
rect 11973 8739 12039 8742
rect 3442 8736 3762 8737
rect 3442 8672 3450 8736
rect 3514 8672 3530 8736
rect 3594 8672 3610 8736
rect 3674 8672 3690 8736
rect 3754 8672 3762 8736
rect 3442 8671 3762 8672
rect 8440 8736 8760 8737
rect 8440 8672 8448 8736
rect 8512 8672 8528 8736
rect 8592 8672 8608 8736
rect 8672 8672 8688 8736
rect 8752 8672 8760 8736
rect 8440 8671 8760 8672
rect 13437 8736 13757 8737
rect 13437 8672 13445 8736
rect 13509 8672 13525 8736
rect 13589 8672 13605 8736
rect 13669 8672 13685 8736
rect 13749 8672 13757 8736
rect 13437 8671 13757 8672
rect 4337 8666 4403 8669
rect 6545 8666 6611 8669
rect 4337 8664 6611 8666
rect 4337 8608 4342 8664
rect 4398 8608 6550 8664
rect 6606 8608 6611 8664
rect 4337 8606 6611 8608
rect 4337 8603 4403 8606
rect 6545 8603 6611 8606
rect 9213 8666 9279 8669
rect 9622 8666 9628 8668
rect 9213 8664 9628 8666
rect 9213 8608 9218 8664
rect 9274 8608 9628 8664
rect 9213 8606 9628 8608
rect 9213 8603 9279 8606
rect 9622 8604 9628 8606
rect 9692 8604 9698 8668
rect 10225 8666 10291 8669
rect 11513 8666 11579 8669
rect 10225 8664 11579 8666
rect 10225 8608 10230 8664
rect 10286 8608 11518 8664
rect 11574 8608 11579 8664
rect 10225 8606 11579 8608
rect 10225 8603 10291 8606
rect 11513 8603 11579 8606
rect 11973 8666 12039 8669
rect 11973 8664 13370 8666
rect 11973 8608 11978 8664
rect 12034 8608 13370 8664
rect 11973 8606 13370 8608
rect 11973 8603 12039 8606
rect 3877 8530 3943 8533
rect 12525 8530 12591 8533
rect 3877 8528 12591 8530
rect 3877 8472 3882 8528
rect 3938 8472 12530 8528
rect 12586 8472 12591 8528
rect 3877 8470 12591 8472
rect 13310 8530 13370 8606
rect 14092 8530 14152 8875
rect 15193 8530 15259 8533
rect 13310 8528 15259 8530
rect 13310 8472 15198 8528
rect 15254 8472 15259 8528
rect 13310 8470 15259 8472
rect 3877 8467 3943 8470
rect 12525 8467 12591 8470
rect 15193 8467 15259 8470
rect 0 8394 800 8424
rect 1393 8394 1459 8397
rect 0 8392 1459 8394
rect 0 8336 1398 8392
rect 1454 8336 1459 8392
rect 0 8334 1459 8336
rect 0 8304 800 8334
rect 1393 8331 1459 8334
rect 2681 8394 2747 8397
rect 7281 8394 7347 8397
rect 13353 8394 13419 8397
rect 2681 8392 6562 8394
rect 2681 8336 2686 8392
rect 2742 8336 6562 8392
rect 2681 8334 6562 8336
rect 2681 8331 2747 8334
rect 2497 8258 2563 8261
rect 2957 8258 3023 8261
rect 5809 8258 5875 8261
rect 2497 8256 2790 8258
rect 2497 8200 2502 8256
rect 2558 8200 2790 8256
rect 2497 8198 2790 8200
rect 2497 8195 2563 8198
rect 2730 8122 2790 8198
rect 2957 8256 5875 8258
rect 2957 8200 2962 8256
rect 3018 8200 5814 8256
rect 5870 8200 5875 8256
rect 2957 8198 5875 8200
rect 6502 8258 6562 8334
rect 7281 8392 13419 8394
rect 7281 8336 7286 8392
rect 7342 8336 13358 8392
rect 13414 8336 13419 8392
rect 7281 8334 13419 8336
rect 7281 8331 7347 8334
rect 13353 8331 13419 8334
rect 10317 8258 10383 8261
rect 10777 8258 10843 8261
rect 6502 8256 10843 8258
rect 6502 8200 10322 8256
rect 10378 8200 10782 8256
rect 10838 8200 10843 8256
rect 6502 8198 10843 8200
rect 2957 8195 3023 8198
rect 5809 8195 5875 8198
rect 10317 8195 10383 8198
rect 10777 8195 10843 8198
rect 11789 8258 11855 8261
rect 12157 8258 12223 8261
rect 11789 8256 12223 8258
rect 11789 8200 11794 8256
rect 11850 8200 12162 8256
rect 12218 8200 12223 8256
rect 11789 8198 12223 8200
rect 11789 8195 11855 8198
rect 12157 8195 12223 8198
rect 12617 8258 12683 8261
rect 13261 8260 13327 8261
rect 12750 8258 12756 8260
rect 12617 8256 12756 8258
rect 12617 8200 12622 8256
rect 12678 8200 12756 8256
rect 12617 8198 12756 8200
rect 12617 8195 12683 8198
rect 12750 8196 12756 8198
rect 12820 8196 12826 8260
rect 13261 8258 13308 8260
rect 13216 8256 13308 8258
rect 13216 8200 13266 8256
rect 13216 8198 13308 8200
rect 13261 8196 13308 8198
rect 13372 8196 13378 8260
rect 13261 8195 13327 8196
rect 5941 8192 6261 8193
rect 5941 8128 5949 8192
rect 6013 8128 6029 8192
rect 6093 8128 6109 8192
rect 6173 8128 6189 8192
rect 6253 8128 6261 8192
rect 5941 8127 6261 8128
rect 10938 8192 11258 8193
rect 10938 8128 10946 8192
rect 11010 8128 11026 8192
rect 11090 8128 11106 8192
rect 11170 8128 11186 8192
rect 11250 8128 11258 8192
rect 10938 8127 11258 8128
rect 8109 8122 8175 8125
rect 10726 8122 10732 8124
rect 2730 8062 5826 8122
rect 2405 7986 2471 7989
rect 2957 7986 3023 7989
rect 3693 7986 3759 7989
rect 2405 7984 2790 7986
rect 2405 7928 2410 7984
rect 2466 7928 2790 7984
rect 2405 7926 2790 7928
rect 2405 7923 2471 7926
rect 0 7442 800 7472
rect 1393 7442 1459 7445
rect 0 7440 1459 7442
rect 0 7384 1398 7440
rect 1454 7384 1459 7440
rect 0 7382 1459 7384
rect 2730 7442 2790 7926
rect 2957 7984 3759 7986
rect 2957 7928 2962 7984
rect 3018 7928 3698 7984
rect 3754 7928 3759 7984
rect 2957 7926 3759 7928
rect 2957 7923 3023 7926
rect 3693 7923 3759 7926
rect 3877 7986 3943 7989
rect 4286 7986 4292 7988
rect 3877 7984 4292 7986
rect 3877 7928 3882 7984
rect 3938 7928 4292 7984
rect 3877 7926 4292 7928
rect 3877 7923 3943 7926
rect 4286 7924 4292 7926
rect 4356 7924 4362 7988
rect 4521 7986 4587 7989
rect 4705 7986 4771 7989
rect 5165 7986 5231 7989
rect 4521 7984 5231 7986
rect 4521 7928 4526 7984
rect 4582 7928 4710 7984
rect 4766 7928 5170 7984
rect 5226 7928 5231 7984
rect 4521 7926 5231 7928
rect 5766 7986 5826 8062
rect 8109 8120 10732 8122
rect 8109 8064 8114 8120
rect 8170 8064 10732 8120
rect 8109 8062 10732 8064
rect 8109 8059 8175 8062
rect 10726 8060 10732 8062
rect 10796 8060 10802 8124
rect 11646 8060 11652 8124
rect 11716 8122 11722 8124
rect 11789 8122 11855 8125
rect 14273 8122 14339 8125
rect 11716 8120 14339 8122
rect 11716 8064 11794 8120
rect 11850 8064 14278 8120
rect 14334 8064 14339 8120
rect 11716 8062 14339 8064
rect 11716 8060 11722 8062
rect 11789 8059 11855 8062
rect 14273 8059 14339 8062
rect 12249 7986 12315 7989
rect 5766 7984 12315 7986
rect 5766 7928 12254 7984
rect 12310 7928 12315 7984
rect 5766 7926 12315 7928
rect 4521 7923 4587 7926
rect 4705 7923 4771 7926
rect 5165 7923 5231 7926
rect 12249 7923 12315 7926
rect 12433 7986 12499 7989
rect 12893 7986 12959 7989
rect 12433 7984 12959 7986
rect 12433 7928 12438 7984
rect 12494 7928 12898 7984
rect 12954 7928 12959 7984
rect 12433 7926 12959 7928
rect 12433 7923 12499 7926
rect 12893 7923 12959 7926
rect 3141 7850 3207 7853
rect 4061 7850 4127 7853
rect 11237 7850 11303 7853
rect 11881 7852 11947 7853
rect 3141 7848 3940 7850
rect 3141 7792 3146 7848
rect 3202 7792 3940 7848
rect 3141 7790 3940 7792
rect 3141 7787 3207 7790
rect 3442 7648 3762 7649
rect 3442 7584 3450 7648
rect 3514 7584 3530 7648
rect 3594 7584 3610 7648
rect 3674 7584 3690 7648
rect 3754 7584 3762 7648
rect 3442 7583 3762 7584
rect 3880 7578 3940 7790
rect 4061 7848 11303 7850
rect 4061 7792 4066 7848
rect 4122 7792 11242 7848
rect 11298 7792 11303 7848
rect 4061 7790 11303 7792
rect 4061 7787 4127 7790
rect 11237 7787 11303 7790
rect 11830 7788 11836 7852
rect 11900 7850 11947 7852
rect 12065 7850 12131 7853
rect 12198 7850 12204 7852
rect 11900 7848 11992 7850
rect 11942 7792 11992 7848
rect 11900 7790 11992 7792
rect 12065 7848 12204 7850
rect 12065 7792 12070 7848
rect 12126 7792 12204 7848
rect 12065 7790 12204 7792
rect 11900 7788 11947 7790
rect 11881 7787 11947 7788
rect 12065 7787 12131 7790
rect 12198 7788 12204 7790
rect 12268 7788 12274 7852
rect 4153 7714 4219 7717
rect 5758 7714 5764 7716
rect 4153 7712 5764 7714
rect 4153 7656 4158 7712
rect 4214 7656 5764 7712
rect 4153 7654 5764 7656
rect 4153 7651 4219 7654
rect 5758 7652 5764 7654
rect 5828 7652 5834 7716
rect 8845 7714 8911 7717
rect 10869 7714 10935 7717
rect 8845 7712 10935 7714
rect 8845 7656 8850 7712
rect 8906 7656 10874 7712
rect 10930 7656 10935 7712
rect 8845 7654 10935 7656
rect 8845 7651 8911 7654
rect 10869 7651 10935 7654
rect 11053 7714 11119 7717
rect 12157 7714 12223 7717
rect 11053 7712 12223 7714
rect 11053 7656 11058 7712
rect 11114 7656 12162 7712
rect 12218 7656 12223 7712
rect 11053 7654 12223 7656
rect 11053 7651 11119 7654
rect 12157 7651 12223 7654
rect 8440 7648 8760 7649
rect 8440 7584 8448 7648
rect 8512 7584 8528 7648
rect 8592 7584 8608 7648
rect 8672 7584 8688 7648
rect 8752 7584 8760 7648
rect 8440 7583 8760 7584
rect 13437 7648 13757 7649
rect 13437 7584 13445 7648
rect 13509 7584 13525 7648
rect 13589 7584 13605 7648
rect 13669 7584 13685 7648
rect 13749 7584 13757 7648
rect 13437 7583 13757 7584
rect 8201 7578 8267 7581
rect 3880 7576 8267 7578
rect 3880 7520 8206 7576
rect 8262 7520 8267 7576
rect 3880 7518 8267 7520
rect 8201 7515 8267 7518
rect 8845 7578 8911 7581
rect 13077 7578 13143 7581
rect 8845 7576 13143 7578
rect 8845 7520 8850 7576
rect 8906 7520 13082 7576
rect 13138 7520 13143 7576
rect 8845 7518 13143 7520
rect 8845 7515 8911 7518
rect 13077 7515 13143 7518
rect 11697 7442 11763 7445
rect 2730 7440 11763 7442
rect 2730 7384 11702 7440
rect 11758 7384 11763 7440
rect 2730 7382 11763 7384
rect 0 7352 800 7382
rect 1393 7379 1459 7382
rect 11697 7379 11763 7382
rect 11973 7442 12039 7445
rect 13077 7442 13143 7445
rect 11973 7440 13143 7442
rect 11973 7384 11978 7440
rect 12034 7384 13082 7440
rect 13138 7384 13143 7440
rect 11973 7382 13143 7384
rect 11973 7379 12039 7382
rect 13077 7379 13143 7382
rect 3785 7306 3851 7309
rect 3785 7304 11484 7306
rect 3785 7248 3790 7304
rect 3846 7248 11484 7304
rect 3785 7246 11484 7248
rect 3785 7243 3851 7246
rect 3601 7170 3667 7173
rect 5717 7170 5783 7173
rect 3601 7168 5783 7170
rect 3601 7112 3606 7168
rect 3662 7112 5722 7168
rect 5778 7112 5783 7168
rect 3601 7110 5783 7112
rect 3601 7107 3667 7110
rect 5717 7107 5783 7110
rect 6361 7170 6427 7173
rect 6678 7170 6684 7172
rect 6361 7168 6684 7170
rect 6361 7112 6366 7168
rect 6422 7112 6684 7168
rect 6361 7110 6684 7112
rect 6361 7107 6427 7110
rect 6678 7108 6684 7110
rect 6748 7108 6754 7172
rect 8109 7170 8175 7173
rect 10041 7170 10107 7173
rect 10593 7172 10659 7173
rect 8109 7168 10107 7170
rect 8109 7112 8114 7168
rect 8170 7112 10046 7168
rect 10102 7112 10107 7168
rect 8109 7110 10107 7112
rect 8109 7107 8175 7110
rect 10041 7107 10107 7110
rect 10542 7108 10548 7172
rect 10612 7170 10659 7172
rect 10612 7168 10704 7170
rect 10654 7112 10704 7168
rect 10612 7110 10704 7112
rect 10612 7108 10659 7110
rect 10593 7107 10659 7108
rect 5941 7104 6261 7105
rect 5941 7040 5949 7104
rect 6013 7040 6029 7104
rect 6093 7040 6109 7104
rect 6173 7040 6189 7104
rect 6253 7040 6261 7104
rect 5941 7039 6261 7040
rect 10938 7104 11258 7105
rect 10938 7040 10946 7104
rect 11010 7040 11026 7104
rect 11090 7040 11106 7104
rect 11170 7040 11186 7104
rect 11250 7040 11258 7104
rect 10938 7039 11258 7040
rect 3325 7034 3391 7037
rect 5257 7034 5323 7037
rect 3325 7032 5323 7034
rect 3325 6976 3330 7032
rect 3386 6976 5262 7032
rect 5318 6976 5323 7032
rect 3325 6974 5323 6976
rect 3325 6971 3391 6974
rect 5257 6971 5323 6974
rect 6453 7034 6519 7037
rect 10777 7034 10843 7037
rect 6453 7032 10843 7034
rect 6453 6976 6458 7032
rect 6514 6976 10782 7032
rect 10838 6976 10843 7032
rect 6453 6974 10843 6976
rect 11424 7034 11484 7246
rect 11881 7170 11947 7173
rect 13813 7170 13879 7173
rect 11881 7168 13879 7170
rect 11881 7112 11886 7168
rect 11942 7112 13818 7168
rect 13874 7112 13879 7168
rect 11881 7110 13879 7112
rect 11881 7107 11947 7110
rect 13813 7107 13879 7110
rect 12341 7034 12407 7037
rect 11424 7032 12407 7034
rect 11424 6976 12346 7032
rect 12402 6976 12407 7032
rect 11424 6974 12407 6976
rect 6453 6971 6519 6974
rect 10777 6971 10843 6974
rect 12341 6971 12407 6974
rect 12617 7034 12683 7037
rect 14733 7034 14799 7037
rect 12617 7032 14799 7034
rect 12617 6976 12622 7032
rect 12678 6976 14738 7032
rect 14794 6976 14799 7032
rect 12617 6974 14799 6976
rect 12617 6971 12683 6974
rect 14733 6971 14799 6974
rect 2497 6898 2563 6901
rect 3877 6898 3943 6901
rect 2497 6896 3943 6898
rect 2497 6840 2502 6896
rect 2558 6840 3882 6896
rect 3938 6840 3943 6896
rect 2497 6838 3943 6840
rect 2497 6835 2563 6838
rect 3877 6835 3943 6838
rect 4061 6898 4127 6901
rect 10869 6898 10935 6901
rect 4061 6896 10935 6898
rect 4061 6840 4066 6896
rect 4122 6840 10874 6896
rect 10930 6840 10935 6896
rect 4061 6838 10935 6840
rect 4061 6835 4127 6838
rect 10869 6835 10935 6838
rect 11053 6898 11119 6901
rect 11697 6898 11763 6901
rect 11053 6896 11763 6898
rect 11053 6840 11058 6896
rect 11114 6840 11702 6896
rect 11758 6840 11763 6896
rect 11053 6838 11763 6840
rect 11053 6835 11119 6838
rect 11697 6835 11763 6838
rect 12157 6898 12223 6901
rect 12382 6898 12388 6900
rect 12157 6896 12388 6898
rect 12157 6840 12162 6896
rect 12218 6840 12388 6896
rect 12157 6838 12388 6840
rect 12157 6835 12223 6838
rect 12382 6836 12388 6838
rect 12452 6898 12458 6900
rect 14365 6898 14431 6901
rect 12452 6896 14431 6898
rect 12452 6840 14370 6896
rect 14426 6840 14431 6896
rect 12452 6838 14431 6840
rect 12452 6836 12458 6838
rect 14365 6835 14431 6838
rect 2865 6762 2931 6765
rect 9765 6762 9831 6765
rect 11145 6762 11211 6765
rect 14089 6762 14155 6765
rect 2865 6760 9690 6762
rect 2865 6704 2870 6760
rect 2926 6704 9690 6760
rect 2865 6702 9690 6704
rect 2865 6699 2931 6702
rect 4153 6626 4219 6629
rect 8293 6626 8359 6629
rect 4153 6624 8359 6626
rect 4153 6568 4158 6624
rect 4214 6568 8298 6624
rect 8354 6568 8359 6624
rect 4153 6566 8359 6568
rect 4153 6563 4219 6566
rect 8293 6563 8359 6566
rect 8845 6626 8911 6629
rect 9489 6626 9555 6629
rect 8845 6624 9555 6626
rect 8845 6568 8850 6624
rect 8906 6568 9494 6624
rect 9550 6568 9555 6624
rect 8845 6566 9555 6568
rect 8845 6563 8911 6566
rect 9489 6563 9555 6566
rect 3442 6560 3762 6561
rect 0 6490 800 6520
rect 3442 6496 3450 6560
rect 3514 6496 3530 6560
rect 3594 6496 3610 6560
rect 3674 6496 3690 6560
rect 3754 6496 3762 6560
rect 3442 6495 3762 6496
rect 8440 6560 8760 6561
rect 8440 6496 8448 6560
rect 8512 6496 8528 6560
rect 8592 6496 8608 6560
rect 8672 6496 8688 6560
rect 8752 6496 8760 6560
rect 8440 6495 8760 6496
rect 1485 6490 1551 6493
rect 0 6488 1551 6490
rect 0 6432 1490 6488
rect 1546 6432 1551 6488
rect 0 6430 1551 6432
rect 0 6400 800 6430
rect 1485 6427 1551 6430
rect 3877 6490 3943 6493
rect 7373 6490 7439 6493
rect 3877 6488 7439 6490
rect 3877 6432 3882 6488
rect 3938 6432 7378 6488
rect 7434 6432 7439 6488
rect 3877 6430 7439 6432
rect 9630 6490 9690 6702
rect 9765 6760 14155 6762
rect 9765 6704 9770 6760
rect 9826 6704 11150 6760
rect 11206 6704 14094 6760
rect 14150 6704 14155 6760
rect 9765 6702 14155 6704
rect 9765 6699 9831 6702
rect 11145 6699 11211 6702
rect 14089 6699 14155 6702
rect 10041 6628 10107 6629
rect 9990 6626 9996 6628
rect 9950 6566 9996 6626
rect 10060 6624 10107 6628
rect 10102 6568 10107 6624
rect 9990 6564 9996 6566
rect 10060 6564 10107 6568
rect 10174 6564 10180 6628
rect 10244 6626 10250 6628
rect 12985 6626 13051 6629
rect 10244 6624 13051 6626
rect 10244 6568 12990 6624
rect 13046 6568 13051 6624
rect 10244 6566 13051 6568
rect 10244 6564 10250 6566
rect 10041 6563 10107 6564
rect 12985 6563 13051 6566
rect 13437 6560 13757 6561
rect 13437 6496 13445 6560
rect 13509 6496 13525 6560
rect 13589 6496 13605 6560
rect 13669 6496 13685 6560
rect 13749 6496 13757 6560
rect 13437 6495 13757 6496
rect 12433 6490 12499 6493
rect 9630 6488 12499 6490
rect 9630 6432 12438 6488
rect 12494 6432 12499 6488
rect 9630 6430 12499 6432
rect 3877 6427 3943 6430
rect 7373 6427 7439 6430
rect 12433 6427 12499 6430
rect 8201 6354 8267 6357
rect 11973 6354 12039 6357
rect 12934 6354 12940 6356
rect 2224 6352 8267 6354
rect 2224 6296 8206 6352
rect 8262 6296 8267 6352
rect 2224 6294 8267 6296
rect 2224 6221 2284 6294
rect 8201 6291 8267 6294
rect 8526 6294 11668 6354
rect 8526 6252 8586 6294
rect 2221 6216 2287 6221
rect 8342 6218 8586 6252
rect 2221 6160 2226 6216
rect 2282 6160 2287 6216
rect 2221 6155 2287 6160
rect 5766 6192 8586 6218
rect 8661 6218 8727 6221
rect 8886 6218 8892 6220
rect 8661 6216 8892 6218
rect 5766 6158 8402 6192
rect 8661 6160 8666 6216
rect 8722 6160 8892 6216
rect 8661 6158 8892 6160
rect 2129 6082 2195 6085
rect 5766 6082 5826 6158
rect 8661 6155 8727 6158
rect 8886 6156 8892 6158
rect 8956 6218 8962 6220
rect 9765 6218 9831 6221
rect 8956 6216 9831 6218
rect 8956 6160 9770 6216
rect 9826 6160 9831 6216
rect 8956 6158 9831 6160
rect 8956 6156 8962 6158
rect 9765 6155 9831 6158
rect 10041 6218 10107 6221
rect 10542 6218 10548 6220
rect 10041 6216 10548 6218
rect 10041 6160 10046 6216
rect 10102 6160 10548 6216
rect 10041 6158 10548 6160
rect 10041 6155 10107 6158
rect 10542 6156 10548 6158
rect 10612 6156 10618 6220
rect 10726 6156 10732 6220
rect 10796 6218 10802 6220
rect 10869 6218 10935 6221
rect 10796 6216 10935 6218
rect 10796 6160 10874 6216
rect 10930 6160 10935 6216
rect 10796 6158 10935 6160
rect 10796 6156 10802 6158
rect 10869 6155 10935 6158
rect 11053 6218 11119 6221
rect 11462 6218 11468 6220
rect 11053 6216 11468 6218
rect 11053 6160 11058 6216
rect 11114 6160 11468 6216
rect 11053 6158 11468 6160
rect 11053 6155 11119 6158
rect 11462 6156 11468 6158
rect 11532 6156 11538 6220
rect 11608 6218 11668 6294
rect 11973 6352 12940 6354
rect 11973 6296 11978 6352
rect 12034 6296 12940 6352
rect 11973 6294 12940 6296
rect 11973 6291 12039 6294
rect 12934 6292 12940 6294
rect 13004 6354 13010 6356
rect 14365 6354 14431 6357
rect 13004 6352 14431 6354
rect 13004 6296 14370 6352
rect 14426 6296 14431 6352
rect 13004 6294 14431 6296
rect 13004 6292 13010 6294
rect 14365 6291 14431 6294
rect 13353 6218 13419 6221
rect 11608 6216 13419 6218
rect 11608 6160 13358 6216
rect 13414 6160 13419 6216
rect 11608 6158 13419 6160
rect 13353 6155 13419 6158
rect 2129 6080 5826 6082
rect 2129 6024 2134 6080
rect 2190 6024 5826 6080
rect 2129 6022 5826 6024
rect 6913 6082 6979 6085
rect 10777 6082 10843 6085
rect 6913 6080 10843 6082
rect 6913 6024 6918 6080
rect 6974 6024 10782 6080
rect 10838 6024 10843 6080
rect 6913 6022 10843 6024
rect 2129 6019 2195 6022
rect 6913 6019 6979 6022
rect 10777 6019 10843 6022
rect 11646 6020 11652 6084
rect 11716 6082 11722 6084
rect 12157 6082 12223 6085
rect 11716 6080 12223 6082
rect 11716 6024 12162 6080
rect 12218 6024 12223 6080
rect 11716 6022 12223 6024
rect 11716 6020 11722 6022
rect 12157 6019 12223 6022
rect 12341 6082 12407 6085
rect 12566 6082 12572 6084
rect 12341 6080 12572 6082
rect 12341 6024 12346 6080
rect 12402 6024 12572 6080
rect 12341 6022 12572 6024
rect 12341 6019 12407 6022
rect 12566 6020 12572 6022
rect 12636 6082 12642 6084
rect 13629 6082 13695 6085
rect 12636 6080 13695 6082
rect 12636 6024 13634 6080
rect 13690 6024 13695 6080
rect 12636 6022 13695 6024
rect 12636 6020 12642 6022
rect 13629 6019 13695 6022
rect 5941 6016 6261 6017
rect 5941 5952 5949 6016
rect 6013 5952 6029 6016
rect 6093 5952 6109 6016
rect 6173 5952 6189 6016
rect 6253 5952 6261 6016
rect 5941 5951 6261 5952
rect 10938 6016 11258 6017
rect 10938 5952 10946 6016
rect 11010 5952 11026 6016
rect 11090 5952 11106 6016
rect 11170 5952 11186 6016
rect 11250 5952 11258 6016
rect 10938 5951 11258 5952
rect 2129 5946 2195 5949
rect 5809 5946 5875 5949
rect 2129 5944 5875 5946
rect 2129 5888 2134 5944
rect 2190 5888 5814 5944
rect 5870 5888 5875 5944
rect 2129 5886 5875 5888
rect 2129 5883 2195 5886
rect 5809 5883 5875 5886
rect 7373 5946 7439 5949
rect 11789 5946 11855 5949
rect 12709 5946 12775 5949
rect 7373 5944 10840 5946
rect 7373 5888 7378 5944
rect 7434 5888 10840 5944
rect 7373 5886 10840 5888
rect 7373 5883 7439 5886
rect 2405 5810 2471 5813
rect 8201 5810 8267 5813
rect 2405 5808 8267 5810
rect 2405 5752 2410 5808
rect 2466 5752 8206 5808
rect 8262 5752 8267 5808
rect 2405 5750 8267 5752
rect 2405 5747 2471 5750
rect 8201 5747 8267 5750
rect 8385 5810 8451 5813
rect 8845 5810 8911 5813
rect 10317 5810 10383 5813
rect 10501 5812 10567 5813
rect 10501 5810 10548 5812
rect 8385 5808 10383 5810
rect 8385 5752 8390 5808
rect 8446 5752 8850 5808
rect 8906 5752 10322 5808
rect 10378 5752 10383 5808
rect 8385 5750 10383 5752
rect 10456 5808 10548 5810
rect 10456 5752 10506 5808
rect 10456 5750 10548 5752
rect 8385 5747 8451 5750
rect 8845 5747 8911 5750
rect 10317 5747 10383 5750
rect 10501 5748 10548 5750
rect 10612 5748 10618 5812
rect 10780 5810 10840 5886
rect 11789 5944 12775 5946
rect 11789 5888 11794 5944
rect 11850 5888 12714 5944
rect 12770 5888 12775 5944
rect 11789 5886 12775 5888
rect 11789 5883 11855 5886
rect 12709 5883 12775 5886
rect 11697 5810 11763 5813
rect 10780 5808 11763 5810
rect 10780 5752 11702 5808
rect 11758 5752 11763 5808
rect 10780 5750 11763 5752
rect 10501 5747 10567 5748
rect 11697 5747 11763 5750
rect 12566 5748 12572 5812
rect 12636 5810 12642 5812
rect 12709 5810 12775 5813
rect 13854 5810 13860 5812
rect 12636 5808 13860 5810
rect 12636 5752 12714 5808
rect 12770 5752 13860 5808
rect 12636 5750 13860 5752
rect 12636 5748 12642 5750
rect 12709 5747 12775 5750
rect 13854 5748 13860 5750
rect 13924 5748 13930 5812
rect 4337 5674 4403 5677
rect 10961 5674 11027 5677
rect 4337 5672 11027 5674
rect 4337 5616 4342 5672
rect 4398 5616 10966 5672
rect 11022 5616 11027 5672
rect 4337 5614 11027 5616
rect 4337 5611 4403 5614
rect 10961 5611 11027 5614
rect 11329 5674 11395 5677
rect 12249 5674 12315 5677
rect 11329 5672 12315 5674
rect 11329 5616 11334 5672
rect 11390 5616 12254 5672
rect 12310 5616 12315 5672
rect 11329 5614 12315 5616
rect 11329 5611 11395 5614
rect 12249 5611 12315 5614
rect 3877 5538 3943 5541
rect 5625 5538 5691 5541
rect 3877 5536 5691 5538
rect 3877 5480 3882 5536
rect 3938 5480 5630 5536
rect 5686 5480 5691 5536
rect 3877 5478 5691 5480
rect 3877 5475 3943 5478
rect 5625 5475 5691 5478
rect 5809 5538 5875 5541
rect 6729 5538 6795 5541
rect 8293 5538 8359 5541
rect 5809 5536 8359 5538
rect 5809 5480 5814 5536
rect 5870 5480 6734 5536
rect 6790 5480 8298 5536
rect 8354 5480 8359 5536
rect 5809 5478 8359 5480
rect 5809 5475 5875 5478
rect 6729 5475 6795 5478
rect 8293 5475 8359 5478
rect 9070 5476 9076 5540
rect 9140 5538 9146 5540
rect 11697 5538 11763 5541
rect 9140 5536 11763 5538
rect 9140 5480 11702 5536
rect 11758 5480 11763 5536
rect 9140 5478 11763 5480
rect 12252 5538 12312 5611
rect 13077 5538 13143 5541
rect 12252 5536 13143 5538
rect 12252 5480 13082 5536
rect 13138 5480 13143 5536
rect 12252 5478 13143 5480
rect 9140 5476 9146 5478
rect 11697 5475 11763 5478
rect 13077 5475 13143 5478
rect 3442 5472 3762 5473
rect 0 5402 800 5432
rect 3442 5408 3450 5472
rect 3514 5408 3530 5472
rect 3594 5408 3610 5472
rect 3674 5408 3690 5472
rect 3754 5408 3762 5472
rect 3442 5407 3762 5408
rect 8440 5472 8760 5473
rect 8440 5408 8448 5472
rect 8512 5408 8528 5472
rect 8592 5408 8608 5472
rect 8672 5408 8688 5472
rect 8752 5408 8760 5472
rect 8440 5407 8760 5408
rect 13437 5472 13757 5473
rect 13437 5408 13445 5472
rect 13509 5408 13525 5472
rect 13589 5408 13605 5472
rect 13669 5408 13685 5472
rect 13749 5408 13757 5472
rect 13437 5407 13757 5408
rect 1485 5402 1551 5405
rect 0 5400 1551 5402
rect 0 5344 1490 5400
rect 1546 5344 1551 5400
rect 0 5342 1551 5344
rect 0 5312 800 5342
rect 1485 5339 1551 5342
rect 3877 5402 3943 5405
rect 6545 5402 6611 5405
rect 3877 5400 6611 5402
rect 3877 5344 3882 5400
rect 3938 5344 6550 5400
rect 6606 5344 6611 5400
rect 3877 5342 6611 5344
rect 3877 5339 3943 5342
rect 6545 5339 6611 5342
rect 9489 5402 9555 5405
rect 10041 5402 10107 5405
rect 9489 5400 10107 5402
rect 9489 5344 9494 5400
rect 9550 5344 10046 5400
rect 10102 5344 10107 5400
rect 9489 5342 10107 5344
rect 9489 5339 9555 5342
rect 10041 5339 10107 5342
rect 10317 5402 10383 5405
rect 12433 5402 12499 5405
rect 10317 5400 12499 5402
rect 10317 5344 10322 5400
rect 10378 5344 12438 5400
rect 12494 5344 12499 5400
rect 10317 5342 12499 5344
rect 10317 5339 10383 5342
rect 12433 5339 12499 5342
rect 2998 5204 3004 5268
rect 3068 5266 3074 5268
rect 9305 5266 9371 5269
rect 3068 5264 9371 5266
rect 3068 5208 9310 5264
rect 9366 5208 9371 5264
rect 3068 5206 9371 5208
rect 3068 5204 3074 5206
rect 9305 5203 9371 5206
rect 9489 5266 9555 5269
rect 10225 5266 10291 5269
rect 9489 5264 10291 5266
rect 9489 5208 9494 5264
rect 9550 5208 10230 5264
rect 10286 5208 10291 5264
rect 9489 5206 10291 5208
rect 9489 5203 9555 5206
rect 10225 5203 10291 5206
rect 10358 5204 10364 5268
rect 10428 5266 10434 5268
rect 10501 5266 10567 5269
rect 10428 5264 10567 5266
rect 10428 5208 10506 5264
rect 10562 5208 10567 5264
rect 10428 5206 10567 5208
rect 10428 5204 10434 5206
rect 10501 5203 10567 5206
rect 10777 5266 10843 5269
rect 13537 5266 13603 5269
rect 10777 5264 13603 5266
rect 10777 5208 10782 5264
rect 10838 5208 13542 5264
rect 13598 5208 13603 5264
rect 10777 5206 13603 5208
rect 10777 5203 10843 5206
rect 13537 5203 13603 5206
rect 11053 5130 11119 5133
rect 2730 5128 11119 5130
rect 2730 5072 11058 5128
rect 11114 5072 11119 5128
rect 2730 5070 11119 5072
rect 1945 4994 2011 4997
rect 2730 4994 2790 5070
rect 11053 5067 11119 5070
rect 11513 5130 11579 5133
rect 11646 5130 11652 5132
rect 11513 5128 11652 5130
rect 11513 5072 11518 5128
rect 11574 5072 11652 5128
rect 11513 5070 11652 5072
rect 11513 5067 11579 5070
rect 11646 5068 11652 5070
rect 11716 5130 11722 5132
rect 13169 5130 13235 5133
rect 11716 5128 13235 5130
rect 11716 5072 13174 5128
rect 13230 5072 13235 5128
rect 11716 5070 13235 5072
rect 11716 5068 11722 5070
rect 13169 5067 13235 5070
rect 3141 4996 3207 4997
rect 3141 4994 3188 4996
rect 1945 4992 2790 4994
rect 1945 4936 1950 4992
rect 2006 4936 2790 4992
rect 1945 4934 2790 4936
rect 3096 4992 3188 4994
rect 3096 4936 3146 4992
rect 3096 4934 3188 4936
rect 1945 4931 2011 4934
rect 3141 4932 3188 4934
rect 3252 4932 3258 4996
rect 3509 4994 3575 4997
rect 4613 4994 4679 4997
rect 3509 4992 4679 4994
rect 3509 4936 3514 4992
rect 3570 4936 4618 4992
rect 4674 4936 4679 4992
rect 3509 4934 4679 4936
rect 3141 4931 3207 4932
rect 3509 4931 3575 4934
rect 4613 4931 4679 4934
rect 4797 4994 4863 4997
rect 5349 4994 5415 4997
rect 4797 4992 5415 4994
rect 4797 4936 4802 4992
rect 4858 4936 5354 4992
rect 5410 4936 5415 4992
rect 4797 4934 5415 4936
rect 4797 4931 4863 4934
rect 5349 4931 5415 4934
rect 6494 4932 6500 4996
rect 6564 4994 6570 4996
rect 10593 4994 10659 4997
rect 6564 4992 10659 4994
rect 6564 4936 10598 4992
rect 10654 4936 10659 4992
rect 6564 4934 10659 4936
rect 6564 4932 6570 4934
rect 10593 4931 10659 4934
rect 11421 4994 11487 4997
rect 11973 4994 12039 4997
rect 11421 4992 12039 4994
rect 11421 4936 11426 4992
rect 11482 4936 11978 4992
rect 12034 4936 12039 4992
rect 11421 4934 12039 4936
rect 11421 4931 11487 4934
rect 11973 4931 12039 4934
rect 12382 4932 12388 4996
rect 12452 4994 12458 4996
rect 12801 4994 12867 4997
rect 13077 4996 13143 4997
rect 13077 4994 13124 4996
rect 12452 4992 12867 4994
rect 12452 4936 12806 4992
rect 12862 4936 12867 4992
rect 12452 4934 12867 4936
rect 13032 4992 13124 4994
rect 13032 4936 13082 4992
rect 13032 4934 13124 4936
rect 12452 4932 12458 4934
rect 12801 4931 12867 4934
rect 13077 4932 13124 4934
rect 13188 4932 13194 4996
rect 13077 4931 13143 4932
rect 5941 4928 6261 4929
rect 5941 4864 5949 4928
rect 6013 4864 6029 4928
rect 6093 4864 6109 4928
rect 6173 4864 6189 4928
rect 6253 4864 6261 4928
rect 5941 4863 6261 4864
rect 10938 4928 11258 4929
rect 10938 4864 10946 4928
rect 11010 4864 11026 4928
rect 11090 4864 11106 4928
rect 11170 4864 11186 4928
rect 11250 4864 11258 4928
rect 10938 4863 11258 4864
rect 2681 4858 2747 4861
rect 4705 4858 4771 4861
rect 2681 4856 4771 4858
rect 2681 4800 2686 4856
rect 2742 4800 4710 4856
rect 4766 4800 4771 4856
rect 2681 4798 4771 4800
rect 2681 4795 2747 4798
rect 4705 4795 4771 4798
rect 9305 4858 9371 4861
rect 10133 4858 10199 4861
rect 10777 4858 10843 4861
rect 11697 4858 11763 4861
rect 9305 4856 9644 4858
rect 9305 4800 9310 4856
rect 9366 4800 9644 4856
rect 9305 4798 9644 4800
rect 9305 4795 9371 4798
rect 2773 4722 2839 4725
rect 9584 4722 9644 4798
rect 10133 4856 10843 4858
rect 10133 4800 10138 4856
rect 10194 4800 10782 4856
rect 10838 4800 10843 4856
rect 10133 4798 10843 4800
rect 10133 4795 10199 4798
rect 10777 4795 10843 4798
rect 11516 4856 11763 4858
rect 11516 4800 11702 4856
rect 11758 4800 11763 4856
rect 11516 4798 11763 4800
rect 11516 4722 11576 4798
rect 11697 4795 11763 4798
rect 11881 4858 11947 4861
rect 13629 4858 13695 4861
rect 11881 4856 13695 4858
rect 11881 4800 11886 4856
rect 11942 4800 13634 4856
rect 13690 4800 13695 4856
rect 11881 4798 13695 4800
rect 11881 4795 11947 4798
rect 13629 4795 13695 4798
rect 2773 4720 9506 4722
rect 2773 4664 2778 4720
rect 2834 4664 9506 4720
rect 2773 4662 9506 4664
rect 9584 4662 11576 4722
rect 11697 4722 11763 4725
rect 12014 4722 12020 4724
rect 11697 4720 12020 4722
rect 11697 4664 11702 4720
rect 11758 4664 12020 4720
rect 11697 4662 12020 4664
rect 2773 4659 2839 4662
rect 3417 4586 3483 4589
rect 4061 4586 4127 4589
rect 9121 4586 9187 4589
rect 3417 4584 3986 4586
rect 3417 4528 3422 4584
rect 3478 4528 3986 4584
rect 3417 4526 3986 4528
rect 3417 4523 3483 4526
rect 0 4450 800 4480
rect 1485 4450 1551 4453
rect 0 4448 1551 4450
rect 0 4392 1490 4448
rect 1546 4392 1551 4448
rect 0 4390 1551 4392
rect 3926 4450 3986 4526
rect 4061 4584 9187 4586
rect 4061 4528 4066 4584
rect 4122 4528 9126 4584
rect 9182 4528 9187 4584
rect 4061 4526 9187 4528
rect 9446 4586 9506 4662
rect 11697 4659 11763 4662
rect 12014 4660 12020 4662
rect 12084 4722 12090 4724
rect 13629 4722 13695 4725
rect 12084 4720 13695 4722
rect 12084 4664 13634 4720
rect 13690 4664 13695 4720
rect 12084 4662 13695 4664
rect 12084 4660 12090 4662
rect 13629 4659 13695 4662
rect 11973 4586 12039 4589
rect 9446 4584 12039 4586
rect 9446 4528 11978 4584
rect 12034 4528 12039 4584
rect 9446 4526 12039 4528
rect 4061 4523 4127 4526
rect 9121 4523 9187 4526
rect 11973 4523 12039 4526
rect 5533 4450 5599 4453
rect 3926 4448 5599 4450
rect 3926 4392 5538 4448
rect 5594 4392 5599 4448
rect 3926 4390 5599 4392
rect 0 4360 800 4390
rect 1485 4387 1551 4390
rect 5533 4387 5599 4390
rect 5809 4450 5875 4453
rect 8109 4450 8175 4453
rect 9305 4452 9371 4453
rect 9254 4450 9260 4452
rect 5809 4448 8175 4450
rect 5809 4392 5814 4448
rect 5870 4392 8114 4448
rect 8170 4392 8175 4448
rect 5809 4390 8175 4392
rect 9214 4390 9260 4450
rect 9324 4448 9371 4452
rect 9366 4392 9371 4448
rect 5809 4387 5875 4390
rect 8109 4387 8175 4390
rect 9254 4388 9260 4390
rect 9324 4388 9371 4392
rect 9305 4387 9371 4388
rect 9765 4452 9831 4453
rect 10133 4452 10199 4453
rect 9765 4448 9812 4452
rect 9876 4450 9882 4452
rect 10133 4450 10180 4452
rect 9765 4392 9770 4448
rect 9765 4388 9812 4392
rect 9876 4390 9922 4450
rect 10088 4448 10180 4450
rect 10088 4392 10138 4448
rect 10088 4390 10180 4392
rect 9876 4388 9882 4390
rect 10133 4388 10180 4390
rect 10244 4388 10250 4452
rect 11697 4450 11763 4453
rect 10320 4448 11763 4450
rect 10320 4392 11702 4448
rect 11758 4392 11763 4448
rect 10320 4390 11763 4392
rect 9765 4387 9831 4388
rect 10133 4387 10199 4388
rect 3442 4384 3762 4385
rect 3442 4320 3450 4384
rect 3514 4320 3530 4384
rect 3594 4320 3610 4384
rect 3674 4320 3690 4384
rect 3754 4320 3762 4384
rect 3442 4319 3762 4320
rect 8440 4384 8760 4385
rect 8440 4320 8448 4384
rect 8512 4320 8528 4384
rect 8592 4320 8608 4384
rect 8672 4320 8688 4384
rect 8752 4320 8760 4384
rect 8440 4319 8760 4320
rect 4429 4316 4495 4317
rect 4429 4312 4476 4316
rect 4540 4314 4546 4316
rect 4705 4314 4771 4317
rect 6453 4314 6519 4317
rect 4429 4256 4434 4312
rect 4429 4252 4476 4256
rect 4540 4254 4586 4314
rect 4705 4312 6519 4314
rect 4705 4256 4710 4312
rect 4766 4256 6458 4312
rect 6514 4256 6519 4312
rect 4705 4254 6519 4256
rect 4540 4252 4546 4254
rect 4429 4251 4495 4252
rect 4705 4251 4771 4254
rect 6453 4251 6519 4254
rect 9121 4314 9187 4317
rect 10320 4314 10380 4390
rect 11697 4387 11763 4390
rect 13437 4384 13757 4385
rect 13437 4320 13445 4384
rect 13509 4320 13525 4384
rect 13589 4320 13605 4384
rect 13669 4320 13685 4384
rect 13749 4320 13757 4384
rect 13437 4319 13757 4320
rect 11881 4314 11947 4317
rect 9121 4312 10380 4314
rect 9121 4256 9126 4312
rect 9182 4256 10380 4312
rect 9121 4254 10380 4256
rect 10596 4312 11947 4314
rect 10596 4256 11886 4312
rect 11942 4256 11947 4312
rect 10596 4254 11947 4256
rect 9121 4251 9187 4254
rect 2957 4178 3023 4181
rect 9489 4178 9555 4181
rect 2957 4176 9555 4178
rect 2957 4120 2962 4176
rect 3018 4120 9494 4176
rect 9550 4120 9555 4176
rect 2957 4118 9555 4120
rect 2957 4115 3023 4118
rect 9489 4115 9555 4118
rect 10409 4178 10475 4181
rect 10596 4178 10656 4254
rect 11881 4251 11947 4254
rect 12065 4314 12131 4317
rect 12433 4314 12499 4317
rect 12065 4312 12499 4314
rect 12065 4256 12070 4312
rect 12126 4256 12438 4312
rect 12494 4256 12499 4312
rect 12065 4254 12499 4256
rect 12065 4251 12131 4254
rect 12433 4251 12499 4254
rect 10409 4176 10656 4178
rect 10409 4120 10414 4176
rect 10470 4120 10656 4176
rect 10409 4118 10656 4120
rect 10409 4115 10475 4118
rect 10726 4116 10732 4180
rect 10796 4178 10802 4180
rect 13721 4178 13787 4181
rect 10796 4176 13787 4178
rect 10796 4120 13726 4176
rect 13782 4120 13787 4176
rect 10796 4118 13787 4120
rect 10796 4116 10802 4118
rect 13721 4115 13787 4118
rect 2405 4042 2471 4045
rect 9630 4042 10196 4076
rect 12750 4042 12756 4044
rect 2405 4040 12756 4042
rect 2405 3984 2410 4040
rect 2466 4016 12756 4040
rect 2466 3984 9690 4016
rect 2405 3982 9690 3984
rect 10136 3982 12756 4016
rect 2405 3979 2471 3982
rect 12750 3980 12756 3982
rect 12820 4042 12826 4044
rect 12985 4042 13051 4045
rect 12820 4040 13051 4042
rect 12820 3984 12990 4040
rect 13046 3984 13051 4040
rect 12820 3982 13051 3984
rect 12820 3980 12826 3982
rect 12985 3979 13051 3982
rect 2497 3906 2563 3909
rect 4337 3906 4403 3909
rect 2497 3904 4403 3906
rect 2497 3848 2502 3904
rect 2558 3848 4342 3904
rect 4398 3848 4403 3904
rect 2497 3846 4403 3848
rect 2497 3843 2563 3846
rect 4337 3843 4403 3846
rect 5073 3906 5139 3909
rect 5349 3906 5415 3909
rect 6453 3908 6519 3909
rect 6453 3906 6500 3908
rect 5073 3904 5415 3906
rect 5073 3848 5078 3904
rect 5134 3848 5354 3904
rect 5410 3848 5415 3904
rect 5073 3846 5415 3848
rect 6408 3904 6500 3906
rect 6408 3848 6458 3904
rect 6408 3846 6500 3848
rect 5073 3843 5139 3846
rect 5349 3843 5415 3846
rect 6453 3844 6500 3846
rect 6564 3844 6570 3908
rect 8017 3906 8083 3909
rect 9438 3906 9444 3908
rect 8017 3904 9444 3906
rect 8017 3848 8022 3904
rect 8078 3848 9444 3904
rect 8017 3846 9444 3848
rect 6453 3843 6519 3844
rect 8017 3843 8083 3846
rect 9438 3844 9444 3846
rect 9508 3844 9514 3908
rect 10777 3906 10843 3909
rect 9584 3904 10843 3906
rect 9584 3848 10782 3904
rect 10838 3848 10843 3904
rect 9584 3846 10843 3848
rect 5941 3840 6261 3841
rect 5941 3776 5949 3840
rect 6013 3776 6029 3840
rect 6093 3776 6109 3840
rect 6173 3776 6189 3840
rect 6253 3776 6261 3840
rect 5941 3775 6261 3776
rect 3325 3770 3391 3773
rect 5165 3770 5231 3773
rect 3325 3768 5231 3770
rect 3325 3712 3330 3768
rect 3386 3712 5170 3768
rect 5226 3712 5231 3768
rect 3325 3710 5231 3712
rect 3325 3707 3391 3710
rect 5165 3707 5231 3710
rect 6545 3770 6611 3773
rect 9584 3770 9644 3846
rect 10777 3843 10843 3846
rect 11513 3906 11579 3909
rect 12014 3906 12020 3908
rect 11513 3904 12020 3906
rect 11513 3848 11518 3904
rect 11574 3848 12020 3904
rect 11513 3846 12020 3848
rect 11513 3843 11579 3846
rect 12014 3844 12020 3846
rect 12084 3844 12090 3908
rect 12198 3844 12204 3908
rect 12268 3906 12274 3908
rect 12341 3906 12407 3909
rect 12268 3904 12407 3906
rect 12268 3848 12346 3904
rect 12402 3848 12407 3904
rect 12268 3846 12407 3848
rect 12268 3844 12274 3846
rect 12341 3843 12407 3846
rect 10938 3840 11258 3841
rect 10938 3776 10946 3840
rect 11010 3776 11026 3840
rect 11090 3776 11106 3840
rect 11170 3776 11186 3840
rect 11250 3776 11258 3840
rect 10938 3775 11258 3776
rect 10041 3770 10107 3773
rect 6545 3768 9644 3770
rect 6545 3712 6550 3768
rect 6606 3712 9644 3768
rect 6545 3710 9644 3712
rect 9814 3768 10107 3770
rect 9814 3712 10046 3768
rect 10102 3712 10107 3768
rect 9814 3710 10107 3712
rect 6545 3707 6611 3710
rect 3693 3634 3759 3637
rect 9814 3634 9874 3710
rect 10041 3707 10107 3710
rect 10409 3770 10475 3773
rect 10726 3770 10732 3772
rect 10409 3768 10732 3770
rect 10409 3712 10414 3768
rect 10470 3712 10732 3768
rect 10409 3710 10732 3712
rect 10409 3707 10475 3710
rect 10726 3708 10732 3710
rect 10796 3708 10802 3772
rect 11513 3770 11579 3773
rect 12382 3770 12388 3772
rect 11513 3768 12388 3770
rect 11513 3712 11518 3768
rect 11574 3712 12388 3768
rect 11513 3710 12388 3712
rect 11513 3707 11579 3710
rect 12382 3708 12388 3710
rect 12452 3708 12458 3772
rect 3693 3632 9874 3634
rect 3693 3576 3698 3632
rect 3754 3576 9874 3632
rect 3693 3574 9874 3576
rect 9949 3634 10015 3637
rect 11973 3634 12039 3637
rect 13353 3636 13419 3637
rect 9949 3632 12039 3634
rect 9949 3576 9954 3632
rect 10010 3576 11978 3632
rect 12034 3576 12039 3632
rect 9949 3574 12039 3576
rect 3693 3571 3759 3574
rect 9949 3571 10015 3574
rect 11973 3571 12039 3574
rect 13302 3572 13308 3636
rect 13372 3634 13419 3636
rect 13372 3632 13464 3634
rect 13414 3576 13464 3632
rect 13372 3574 13464 3576
rect 13372 3572 13419 3574
rect 13310 3571 13419 3572
rect 0 3498 800 3528
rect 1853 3498 1919 3501
rect 0 3496 1919 3498
rect 0 3440 1858 3496
rect 1914 3440 1919 3496
rect 0 3438 1919 3440
rect 0 3408 800 3438
rect 1853 3435 1919 3438
rect 2773 3498 2839 3501
rect 11605 3498 11671 3501
rect 2773 3496 11671 3498
rect 2773 3440 2778 3496
rect 2834 3440 11610 3496
rect 11666 3440 11671 3496
rect 2773 3438 11671 3440
rect 2773 3435 2839 3438
rect 11605 3435 11671 3438
rect 11789 3498 11855 3501
rect 12014 3498 12020 3500
rect 11789 3496 12020 3498
rect 11789 3440 11794 3496
rect 11850 3440 12020 3496
rect 11789 3438 12020 3440
rect 11789 3435 11855 3438
rect 12014 3436 12020 3438
rect 12084 3498 12090 3500
rect 12433 3498 12499 3501
rect 12084 3496 12499 3498
rect 12084 3440 12438 3496
rect 12494 3440 12499 3496
rect 12084 3438 12499 3440
rect 12084 3436 12090 3438
rect 12433 3435 12499 3438
rect 12617 3498 12683 3501
rect 12750 3498 12756 3500
rect 12617 3496 12756 3498
rect 12617 3440 12622 3496
rect 12678 3440 12756 3496
rect 12617 3438 12756 3440
rect 12617 3435 12683 3438
rect 12750 3436 12756 3438
rect 12820 3436 12826 3500
rect 4286 3300 4292 3364
rect 4356 3362 4362 3364
rect 5165 3362 5231 3365
rect 4356 3360 5231 3362
rect 4356 3304 5170 3360
rect 5226 3304 5231 3360
rect 4356 3302 5231 3304
rect 4356 3300 4362 3302
rect 5165 3299 5231 3302
rect 5441 3362 5507 3365
rect 6545 3362 6611 3365
rect 5441 3360 6611 3362
rect 5441 3304 5446 3360
rect 5502 3304 6550 3360
rect 6606 3304 6611 3360
rect 5441 3302 6611 3304
rect 5441 3299 5507 3302
rect 6545 3299 6611 3302
rect 8886 3300 8892 3364
rect 8956 3362 8962 3364
rect 9581 3362 9647 3365
rect 8956 3360 9647 3362
rect 8956 3304 9586 3360
rect 9642 3304 9647 3360
rect 8956 3302 9647 3304
rect 8956 3300 8962 3302
rect 9581 3299 9647 3302
rect 9806 3300 9812 3364
rect 9876 3362 9882 3364
rect 10041 3362 10107 3365
rect 9876 3360 10107 3362
rect 9876 3304 10046 3360
rect 10102 3304 10107 3360
rect 9876 3302 10107 3304
rect 9876 3300 9882 3302
rect 10041 3299 10107 3302
rect 10174 3300 10180 3364
rect 10244 3362 10250 3364
rect 13310 3362 13370 3571
rect 10244 3302 13370 3362
rect 15653 3362 15719 3365
rect 16400 3362 17200 3392
rect 15653 3360 17200 3362
rect 15653 3304 15658 3360
rect 15714 3304 17200 3360
rect 15653 3302 17200 3304
rect 10244 3300 10250 3302
rect 15653 3299 15719 3302
rect 3442 3296 3762 3297
rect 3442 3232 3450 3296
rect 3514 3232 3530 3296
rect 3594 3232 3610 3296
rect 3674 3232 3690 3296
rect 3754 3232 3762 3296
rect 3442 3231 3762 3232
rect 8440 3296 8760 3297
rect 8440 3232 8448 3296
rect 8512 3232 8528 3296
rect 8592 3232 8608 3296
rect 8672 3232 8688 3296
rect 8752 3232 8760 3296
rect 8440 3231 8760 3232
rect 13437 3296 13757 3297
rect 13437 3232 13445 3296
rect 13509 3232 13525 3296
rect 13589 3232 13605 3296
rect 13669 3232 13685 3296
rect 13749 3232 13757 3296
rect 16400 3272 17200 3302
rect 13437 3231 13757 3232
rect 4521 3226 4587 3229
rect 8109 3226 8175 3229
rect 4521 3224 8175 3226
rect 4521 3168 4526 3224
rect 4582 3168 8114 3224
rect 8170 3168 8175 3224
rect 4521 3166 8175 3168
rect 4521 3163 4587 3166
rect 8109 3163 8175 3166
rect 9489 3226 9555 3229
rect 10317 3226 10383 3229
rect 10961 3226 11027 3229
rect 12893 3226 12959 3229
rect 9489 3224 10196 3226
rect 9489 3168 9494 3224
rect 9550 3168 10196 3224
rect 9489 3166 10196 3168
rect 9489 3163 9555 3166
rect 2221 3090 2287 3093
rect 7281 3090 7347 3093
rect 2221 3088 7347 3090
rect 2221 3032 2226 3088
rect 2282 3032 7286 3088
rect 7342 3032 7347 3088
rect 2221 3030 7347 3032
rect 2221 3027 2287 3030
rect 7281 3027 7347 3030
rect 7925 3090 7991 3093
rect 9857 3090 9923 3093
rect 7925 3088 9923 3090
rect 7925 3032 7930 3088
rect 7986 3032 9862 3088
rect 9918 3032 9923 3088
rect 7925 3030 9923 3032
rect 7925 3027 7991 3030
rect 9857 3027 9923 3030
rect 3233 2954 3299 2957
rect 5073 2954 5139 2957
rect 3233 2952 5139 2954
rect 3233 2896 3238 2952
rect 3294 2896 5078 2952
rect 5134 2896 5139 2952
rect 3233 2894 5139 2896
rect 3233 2891 3299 2894
rect 5073 2891 5139 2894
rect 6269 2954 6335 2957
rect 6678 2954 6684 2956
rect 6269 2952 6684 2954
rect 6269 2896 6274 2952
rect 6330 2896 6684 2952
rect 6269 2894 6684 2896
rect 6269 2891 6335 2894
rect 6678 2892 6684 2894
rect 6748 2892 6754 2956
rect 8109 2954 8175 2957
rect 9622 2954 9628 2956
rect 8109 2952 9628 2954
rect 8109 2896 8114 2952
rect 8170 2896 9628 2952
rect 8109 2894 9628 2896
rect 8109 2891 8175 2894
rect 9622 2892 9628 2894
rect 9692 2892 9698 2956
rect 10136 2954 10196 3166
rect 10317 3224 11027 3226
rect 10317 3168 10322 3224
rect 10378 3168 10966 3224
rect 11022 3168 11027 3224
rect 10317 3166 11027 3168
rect 10317 3163 10383 3166
rect 10961 3163 11027 3166
rect 11102 3224 12959 3226
rect 11102 3168 12898 3224
rect 12954 3168 12959 3224
rect 11102 3166 12959 3168
rect 10501 3090 10567 3093
rect 11102 3090 11162 3166
rect 12893 3163 12959 3166
rect 10501 3088 11162 3090
rect 10501 3032 10506 3088
rect 10562 3032 11162 3088
rect 10501 3030 11162 3032
rect 11237 3090 11303 3093
rect 12566 3090 12572 3092
rect 11237 3088 12572 3090
rect 11237 3032 11242 3088
rect 11298 3032 12572 3088
rect 11237 3030 12572 3032
rect 10501 3027 10567 3030
rect 11237 3027 11303 3030
rect 12566 3028 12572 3030
rect 12636 3028 12642 3092
rect 11881 2954 11947 2957
rect 10136 2952 11947 2954
rect 10136 2896 11886 2952
rect 11942 2896 11947 2952
rect 10136 2894 11947 2896
rect 11881 2891 11947 2894
rect 6545 2820 6611 2821
rect 6494 2818 6500 2820
rect 6454 2758 6500 2818
rect 6564 2816 6611 2820
rect 6606 2760 6611 2816
rect 6494 2756 6500 2758
rect 6564 2756 6611 2760
rect 6545 2755 6611 2756
rect 7005 2818 7071 2821
rect 8661 2818 8727 2821
rect 7005 2816 8727 2818
rect 7005 2760 7010 2816
rect 7066 2760 8666 2816
rect 8722 2760 8727 2816
rect 7005 2758 8727 2760
rect 7005 2755 7071 2758
rect 8661 2755 8727 2758
rect 9857 2818 9923 2821
rect 10174 2818 10180 2820
rect 9857 2816 10180 2818
rect 9857 2760 9862 2816
rect 9918 2760 10180 2816
rect 9857 2758 10180 2760
rect 9857 2755 9923 2758
rect 10174 2756 10180 2758
rect 10244 2756 10250 2820
rect 11513 2818 11579 2821
rect 11830 2818 11836 2820
rect 11513 2816 11836 2818
rect 11513 2760 11518 2816
rect 11574 2760 11836 2816
rect 11513 2758 11836 2760
rect 11513 2755 11579 2758
rect 11830 2756 11836 2758
rect 11900 2756 11906 2820
rect 11973 2818 12039 2821
rect 14038 2818 14044 2820
rect 11973 2816 14044 2818
rect 11973 2760 11978 2816
rect 12034 2760 14044 2816
rect 11973 2758 14044 2760
rect 11973 2755 12039 2758
rect 14038 2756 14044 2758
rect 14108 2756 14114 2820
rect 5941 2752 6261 2753
rect 5941 2688 5949 2752
rect 6013 2688 6029 2752
rect 6093 2688 6109 2752
rect 6173 2688 6189 2752
rect 6253 2688 6261 2752
rect 5941 2687 6261 2688
rect 10938 2752 11258 2753
rect 10938 2688 10946 2752
rect 11010 2688 11026 2752
rect 11090 2688 11106 2752
rect 11170 2688 11186 2752
rect 11250 2688 11258 2752
rect 10938 2687 11258 2688
rect 2221 2682 2287 2685
rect 2681 2682 2747 2685
rect 2221 2680 2747 2682
rect 2221 2624 2226 2680
rect 2282 2624 2686 2680
rect 2742 2624 2747 2680
rect 2221 2622 2747 2624
rect 2221 2619 2287 2622
rect 2681 2619 2747 2622
rect 7649 2682 7715 2685
rect 10777 2682 10843 2685
rect 7649 2680 10843 2682
rect 7649 2624 7654 2680
rect 7710 2624 10782 2680
rect 10838 2624 10843 2680
rect 7649 2622 10843 2624
rect 7649 2619 7715 2622
rect 10777 2619 10843 2622
rect 11697 2682 11763 2685
rect 12382 2682 12388 2684
rect 11697 2680 12388 2682
rect 11697 2624 11702 2680
rect 11758 2624 12388 2680
rect 11697 2622 12388 2624
rect 11697 2619 11763 2622
rect 12382 2620 12388 2622
rect 12452 2620 12458 2684
rect 3182 2484 3188 2548
rect 3252 2546 3258 2548
rect 6545 2546 6611 2549
rect 3252 2544 6611 2546
rect 3252 2488 6550 2544
rect 6606 2488 6611 2544
rect 3252 2486 6611 2488
rect 3252 2484 3258 2486
rect 6545 2483 6611 2486
rect 8201 2546 8267 2549
rect 9254 2546 9260 2548
rect 8201 2544 9260 2546
rect 8201 2488 8206 2544
rect 8262 2488 9260 2544
rect 8201 2486 9260 2488
rect 8201 2483 8267 2486
rect 9254 2484 9260 2486
rect 9324 2484 9330 2548
rect 9990 2484 9996 2548
rect 10060 2546 10066 2548
rect 10501 2546 10567 2549
rect 10060 2544 10567 2546
rect 10060 2488 10506 2544
rect 10562 2488 10567 2544
rect 10060 2486 10567 2488
rect 10060 2484 10066 2486
rect 10501 2483 10567 2486
rect 10961 2546 11027 2549
rect 11646 2546 11652 2548
rect 10961 2544 11652 2546
rect 10961 2488 10966 2544
rect 11022 2488 11652 2544
rect 10961 2486 11652 2488
rect 10961 2483 11027 2486
rect 11646 2484 11652 2486
rect 11716 2484 11722 2548
rect 11973 2546 12039 2549
rect 12750 2546 12756 2548
rect 11973 2544 12756 2546
rect 11973 2488 11978 2544
rect 12034 2488 12756 2544
rect 11973 2486 12756 2488
rect 11973 2483 12039 2486
rect 12750 2484 12756 2486
rect 12820 2484 12826 2548
rect 0 2410 800 2440
rect 1485 2410 1551 2413
rect 0 2408 1551 2410
rect 0 2352 1490 2408
rect 1546 2352 1551 2408
rect 0 2350 1551 2352
rect 0 2320 800 2350
rect 1485 2347 1551 2350
rect 2313 2410 2379 2413
rect 4705 2410 4771 2413
rect 2313 2408 4771 2410
rect 2313 2352 2318 2408
rect 2374 2352 4710 2408
rect 4766 2352 4771 2408
rect 2313 2350 4771 2352
rect 2313 2347 2379 2350
rect 4705 2347 4771 2350
rect 6085 2410 6151 2413
rect 9305 2410 9371 2413
rect 11605 2410 11671 2413
rect 6085 2408 8954 2410
rect 6085 2352 6090 2408
rect 6146 2352 8954 2408
rect 6085 2350 8954 2352
rect 6085 2347 6151 2350
rect 4470 2212 4476 2276
rect 4540 2274 4546 2276
rect 8109 2274 8175 2277
rect 4540 2272 8175 2274
rect 4540 2216 8114 2272
rect 8170 2216 8175 2272
rect 4540 2214 8175 2216
rect 8894 2274 8954 2350
rect 9305 2408 11671 2410
rect 9305 2352 9310 2408
rect 9366 2352 11610 2408
rect 11666 2352 11671 2408
rect 9305 2350 11671 2352
rect 9305 2347 9371 2350
rect 11605 2347 11671 2350
rect 11462 2274 11468 2276
rect 8894 2214 11468 2274
rect 4540 2212 4546 2214
rect 8109 2211 8175 2214
rect 11462 2212 11468 2214
rect 11532 2212 11538 2276
rect 3442 2208 3762 2209
rect 3442 2144 3450 2208
rect 3514 2144 3530 2208
rect 3594 2144 3610 2208
rect 3674 2144 3690 2208
rect 3754 2144 3762 2208
rect 3442 2143 3762 2144
rect 8440 2208 8760 2209
rect 8440 2144 8448 2208
rect 8512 2144 8528 2208
rect 8592 2144 8608 2208
rect 8672 2144 8688 2208
rect 8752 2144 8760 2208
rect 8440 2143 8760 2144
rect 13437 2208 13757 2209
rect 13437 2144 13445 2208
rect 13509 2144 13525 2208
rect 13589 2144 13605 2208
rect 13669 2144 13685 2208
rect 13749 2144 13757 2208
rect 13437 2143 13757 2144
rect 9489 2138 9555 2141
rect 13077 2138 13143 2141
rect 9489 2136 13143 2138
rect 9489 2080 9494 2136
rect 9550 2080 13082 2136
rect 13138 2080 13143 2136
rect 9489 2078 13143 2080
rect 9489 2075 9555 2078
rect 13077 2075 13143 2078
rect 7741 2002 7807 2005
rect 9070 2002 9076 2004
rect 7741 2000 9076 2002
rect 7741 1944 7746 2000
rect 7802 1944 9076 2000
rect 7741 1942 9076 1944
rect 7741 1939 7807 1942
rect 9070 1940 9076 1942
rect 9140 1940 9146 2004
rect 9397 2002 9463 2005
rect 12198 2002 12204 2004
rect 9397 2000 12204 2002
rect 9397 1944 9402 2000
rect 9458 1944 12204 2000
rect 9397 1942 12204 1944
rect 9397 1939 9463 1942
rect 12198 1940 12204 1942
rect 12268 1940 12274 2004
rect 9438 1804 9444 1868
rect 9508 1866 9514 1868
rect 12709 1866 12775 1869
rect 9508 1864 12775 1866
rect 9508 1808 12714 1864
rect 12770 1808 12775 1864
rect 9508 1806 12775 1808
rect 9508 1804 9514 1806
rect 12709 1803 12775 1806
rect 11053 1730 11119 1733
rect 12014 1730 12020 1732
rect 11053 1728 12020 1730
rect 11053 1672 11058 1728
rect 11114 1672 12020 1728
rect 11053 1670 12020 1672
rect 11053 1667 11119 1670
rect 12014 1668 12020 1670
rect 12084 1668 12090 1732
rect 0 1458 800 1488
rect 1853 1458 1919 1461
rect 0 1456 1919 1458
rect 0 1400 1858 1456
rect 1914 1400 1919 1456
rect 0 1398 1919 1400
rect 0 1368 800 1398
rect 1853 1395 1919 1398
rect 0 506 800 536
rect 1669 506 1735 509
rect 0 504 1735 506
rect 0 448 1674 504
rect 1730 448 1735 504
rect 0 446 1735 448
rect 0 416 800 446
rect 1669 443 1735 446
<< via3 >>
rect 3450 17436 3514 17440
rect 3450 17380 3454 17436
rect 3454 17380 3510 17436
rect 3510 17380 3514 17436
rect 3450 17376 3514 17380
rect 3530 17436 3594 17440
rect 3530 17380 3534 17436
rect 3534 17380 3590 17436
rect 3590 17380 3594 17436
rect 3530 17376 3594 17380
rect 3610 17436 3674 17440
rect 3610 17380 3614 17436
rect 3614 17380 3670 17436
rect 3670 17380 3674 17436
rect 3610 17376 3674 17380
rect 3690 17436 3754 17440
rect 3690 17380 3694 17436
rect 3694 17380 3750 17436
rect 3750 17380 3754 17436
rect 3690 17376 3754 17380
rect 8448 17436 8512 17440
rect 8448 17380 8452 17436
rect 8452 17380 8508 17436
rect 8508 17380 8512 17436
rect 8448 17376 8512 17380
rect 8528 17436 8592 17440
rect 8528 17380 8532 17436
rect 8532 17380 8588 17436
rect 8588 17380 8592 17436
rect 8528 17376 8592 17380
rect 8608 17436 8672 17440
rect 8608 17380 8612 17436
rect 8612 17380 8668 17436
rect 8668 17380 8672 17436
rect 8608 17376 8672 17380
rect 8688 17436 8752 17440
rect 8688 17380 8692 17436
rect 8692 17380 8748 17436
rect 8748 17380 8752 17436
rect 8688 17376 8752 17380
rect 13445 17436 13509 17440
rect 13445 17380 13449 17436
rect 13449 17380 13505 17436
rect 13505 17380 13509 17436
rect 13445 17376 13509 17380
rect 13525 17436 13589 17440
rect 13525 17380 13529 17436
rect 13529 17380 13585 17436
rect 13585 17380 13589 17436
rect 13525 17376 13589 17380
rect 13605 17436 13669 17440
rect 13605 17380 13609 17436
rect 13609 17380 13665 17436
rect 13665 17380 13669 17436
rect 13605 17376 13669 17380
rect 13685 17436 13749 17440
rect 13685 17380 13689 17436
rect 13689 17380 13745 17436
rect 13745 17380 13749 17436
rect 13685 17376 13749 17380
rect 5949 16892 6013 16896
rect 5949 16836 5953 16892
rect 5953 16836 6009 16892
rect 6009 16836 6013 16892
rect 5949 16832 6013 16836
rect 6029 16892 6093 16896
rect 6029 16836 6033 16892
rect 6033 16836 6089 16892
rect 6089 16836 6093 16892
rect 6029 16832 6093 16836
rect 6109 16892 6173 16896
rect 6109 16836 6113 16892
rect 6113 16836 6169 16892
rect 6169 16836 6173 16892
rect 6109 16832 6173 16836
rect 6189 16892 6253 16896
rect 6189 16836 6193 16892
rect 6193 16836 6249 16892
rect 6249 16836 6253 16892
rect 6189 16832 6253 16836
rect 10946 16892 11010 16896
rect 10946 16836 10950 16892
rect 10950 16836 11006 16892
rect 11006 16836 11010 16892
rect 10946 16832 11010 16836
rect 11026 16892 11090 16896
rect 11026 16836 11030 16892
rect 11030 16836 11086 16892
rect 11086 16836 11090 16892
rect 11026 16832 11090 16836
rect 11106 16892 11170 16896
rect 11106 16836 11110 16892
rect 11110 16836 11166 16892
rect 11166 16836 11170 16892
rect 11106 16832 11170 16836
rect 11186 16892 11250 16896
rect 11186 16836 11190 16892
rect 11190 16836 11246 16892
rect 11246 16836 11250 16892
rect 11186 16832 11250 16836
rect 9996 16492 10060 16556
rect 6500 16356 6564 16420
rect 3450 16348 3514 16352
rect 3450 16292 3454 16348
rect 3454 16292 3510 16348
rect 3510 16292 3514 16348
rect 3450 16288 3514 16292
rect 3530 16348 3594 16352
rect 3530 16292 3534 16348
rect 3534 16292 3590 16348
rect 3590 16292 3594 16348
rect 3530 16288 3594 16292
rect 3610 16348 3674 16352
rect 3610 16292 3614 16348
rect 3614 16292 3670 16348
rect 3670 16292 3674 16348
rect 3610 16288 3674 16292
rect 3690 16348 3754 16352
rect 3690 16292 3694 16348
rect 3694 16292 3750 16348
rect 3750 16292 3754 16348
rect 3690 16288 3754 16292
rect 8448 16348 8512 16352
rect 8448 16292 8452 16348
rect 8452 16292 8508 16348
rect 8508 16292 8512 16348
rect 8448 16288 8512 16292
rect 8528 16348 8592 16352
rect 8528 16292 8532 16348
rect 8532 16292 8588 16348
rect 8588 16292 8592 16348
rect 8528 16288 8592 16292
rect 8608 16348 8672 16352
rect 8608 16292 8612 16348
rect 8612 16292 8668 16348
rect 8668 16292 8672 16348
rect 8608 16288 8672 16292
rect 8688 16348 8752 16352
rect 8688 16292 8692 16348
rect 8692 16292 8748 16348
rect 8748 16292 8752 16348
rect 8688 16288 8752 16292
rect 13445 16348 13509 16352
rect 13445 16292 13449 16348
rect 13449 16292 13505 16348
rect 13505 16292 13509 16348
rect 13445 16288 13509 16292
rect 13525 16348 13589 16352
rect 13525 16292 13529 16348
rect 13529 16292 13585 16348
rect 13585 16292 13589 16348
rect 13525 16288 13589 16292
rect 13605 16348 13669 16352
rect 13605 16292 13609 16348
rect 13609 16292 13665 16348
rect 13665 16292 13669 16348
rect 13605 16288 13669 16292
rect 13685 16348 13749 16352
rect 13685 16292 13689 16348
rect 13689 16292 13745 16348
rect 13745 16292 13749 16348
rect 13685 16288 13749 16292
rect 9628 15812 9692 15876
rect 5949 15804 6013 15808
rect 5949 15748 5953 15804
rect 5953 15748 6009 15804
rect 6009 15748 6013 15804
rect 5949 15744 6013 15748
rect 6029 15804 6093 15808
rect 6029 15748 6033 15804
rect 6033 15748 6089 15804
rect 6089 15748 6093 15804
rect 6029 15744 6093 15748
rect 6109 15804 6173 15808
rect 6109 15748 6113 15804
rect 6113 15748 6169 15804
rect 6169 15748 6173 15804
rect 6109 15744 6173 15748
rect 6189 15804 6253 15808
rect 6189 15748 6193 15804
rect 6193 15748 6249 15804
rect 6249 15748 6253 15804
rect 6189 15744 6253 15748
rect 10946 15804 11010 15808
rect 10946 15748 10950 15804
rect 10950 15748 11006 15804
rect 11006 15748 11010 15804
rect 10946 15744 11010 15748
rect 11026 15804 11090 15808
rect 11026 15748 11030 15804
rect 11030 15748 11086 15804
rect 11086 15748 11090 15804
rect 11026 15744 11090 15748
rect 11106 15804 11170 15808
rect 11106 15748 11110 15804
rect 11110 15748 11166 15804
rect 11166 15748 11170 15804
rect 11106 15744 11170 15748
rect 11186 15804 11250 15808
rect 11186 15748 11190 15804
rect 11190 15748 11246 15804
rect 11246 15748 11250 15804
rect 11186 15744 11250 15748
rect 3450 15260 3514 15264
rect 3450 15204 3454 15260
rect 3454 15204 3510 15260
rect 3510 15204 3514 15260
rect 3450 15200 3514 15204
rect 3530 15260 3594 15264
rect 3530 15204 3534 15260
rect 3534 15204 3590 15260
rect 3590 15204 3594 15260
rect 3530 15200 3594 15204
rect 3610 15260 3674 15264
rect 3610 15204 3614 15260
rect 3614 15204 3670 15260
rect 3670 15204 3674 15260
rect 3610 15200 3674 15204
rect 3690 15260 3754 15264
rect 3690 15204 3694 15260
rect 3694 15204 3750 15260
rect 3750 15204 3754 15260
rect 3690 15200 3754 15204
rect 8448 15260 8512 15264
rect 8448 15204 8452 15260
rect 8452 15204 8508 15260
rect 8508 15204 8512 15260
rect 8448 15200 8512 15204
rect 8528 15260 8592 15264
rect 8528 15204 8532 15260
rect 8532 15204 8588 15260
rect 8588 15204 8592 15260
rect 8528 15200 8592 15204
rect 8608 15260 8672 15264
rect 8608 15204 8612 15260
rect 8612 15204 8668 15260
rect 8668 15204 8672 15260
rect 8608 15200 8672 15204
rect 8688 15260 8752 15264
rect 8688 15204 8692 15260
rect 8692 15204 8748 15260
rect 8748 15204 8752 15260
rect 8688 15200 8752 15204
rect 13445 15260 13509 15264
rect 13445 15204 13449 15260
rect 13449 15204 13505 15260
rect 13505 15204 13509 15260
rect 13445 15200 13509 15204
rect 13525 15260 13589 15264
rect 13525 15204 13529 15260
rect 13529 15204 13585 15260
rect 13585 15204 13589 15260
rect 13525 15200 13589 15204
rect 13605 15260 13669 15264
rect 13605 15204 13609 15260
rect 13609 15204 13665 15260
rect 13665 15204 13669 15260
rect 13605 15200 13669 15204
rect 13685 15260 13749 15264
rect 13685 15204 13689 15260
rect 13689 15204 13745 15260
rect 13745 15204 13749 15260
rect 13685 15200 13749 15204
rect 10364 14996 10428 15060
rect 5949 14716 6013 14720
rect 5949 14660 5953 14716
rect 5953 14660 6009 14716
rect 6009 14660 6013 14716
rect 5949 14656 6013 14660
rect 6029 14716 6093 14720
rect 6029 14660 6033 14716
rect 6033 14660 6089 14716
rect 6089 14660 6093 14716
rect 6029 14656 6093 14660
rect 6109 14716 6173 14720
rect 6109 14660 6113 14716
rect 6113 14660 6169 14716
rect 6169 14660 6173 14716
rect 6109 14656 6173 14660
rect 6189 14716 6253 14720
rect 6189 14660 6193 14716
rect 6193 14660 6249 14716
rect 6249 14660 6253 14716
rect 6189 14656 6253 14660
rect 10946 14716 11010 14720
rect 10946 14660 10950 14716
rect 10950 14660 11006 14716
rect 11006 14660 11010 14716
rect 10946 14656 11010 14660
rect 11026 14716 11090 14720
rect 11026 14660 11030 14716
rect 11030 14660 11086 14716
rect 11086 14660 11090 14716
rect 11026 14656 11090 14660
rect 11106 14716 11170 14720
rect 11106 14660 11110 14716
rect 11110 14660 11166 14716
rect 11166 14660 11170 14716
rect 11106 14656 11170 14660
rect 11186 14716 11250 14720
rect 11186 14660 11190 14716
rect 11190 14660 11246 14716
rect 11246 14660 11250 14716
rect 11186 14656 11250 14660
rect 3450 14172 3514 14176
rect 3450 14116 3454 14172
rect 3454 14116 3510 14172
rect 3510 14116 3514 14172
rect 3450 14112 3514 14116
rect 3530 14172 3594 14176
rect 3530 14116 3534 14172
rect 3534 14116 3590 14172
rect 3590 14116 3594 14172
rect 3530 14112 3594 14116
rect 3610 14172 3674 14176
rect 3610 14116 3614 14172
rect 3614 14116 3670 14172
rect 3670 14116 3674 14172
rect 3610 14112 3674 14116
rect 3690 14172 3754 14176
rect 3690 14116 3694 14172
rect 3694 14116 3750 14172
rect 3750 14116 3754 14172
rect 3690 14112 3754 14116
rect 8448 14172 8512 14176
rect 8448 14116 8452 14172
rect 8452 14116 8508 14172
rect 8508 14116 8512 14172
rect 8448 14112 8512 14116
rect 8528 14172 8592 14176
rect 8528 14116 8532 14172
rect 8532 14116 8588 14172
rect 8588 14116 8592 14172
rect 8528 14112 8592 14116
rect 8608 14172 8672 14176
rect 8608 14116 8612 14172
rect 8612 14116 8668 14172
rect 8668 14116 8672 14172
rect 8608 14112 8672 14116
rect 8688 14172 8752 14176
rect 8688 14116 8692 14172
rect 8692 14116 8748 14172
rect 8748 14116 8752 14172
rect 8688 14112 8752 14116
rect 13445 14172 13509 14176
rect 13445 14116 13449 14172
rect 13449 14116 13505 14172
rect 13505 14116 13509 14172
rect 13445 14112 13509 14116
rect 13525 14172 13589 14176
rect 13525 14116 13529 14172
rect 13529 14116 13585 14172
rect 13585 14116 13589 14172
rect 13525 14112 13589 14116
rect 13605 14172 13669 14176
rect 13605 14116 13609 14172
rect 13609 14116 13665 14172
rect 13665 14116 13669 14172
rect 13605 14112 13669 14116
rect 13685 14172 13749 14176
rect 13685 14116 13689 14172
rect 13689 14116 13745 14172
rect 13745 14116 13749 14172
rect 13685 14112 13749 14116
rect 5764 13968 5828 13972
rect 5764 13912 5814 13968
rect 5814 13912 5828 13968
rect 5764 13908 5828 13912
rect 9812 13908 9876 13972
rect 8156 13696 8220 13700
rect 8156 13640 8206 13696
rect 8206 13640 8220 13696
rect 8156 13636 8220 13640
rect 5949 13628 6013 13632
rect 5949 13572 5953 13628
rect 5953 13572 6009 13628
rect 6009 13572 6013 13628
rect 5949 13568 6013 13572
rect 6029 13628 6093 13632
rect 6029 13572 6033 13628
rect 6033 13572 6089 13628
rect 6089 13572 6093 13628
rect 6029 13568 6093 13572
rect 6109 13628 6173 13632
rect 6109 13572 6113 13628
rect 6113 13572 6169 13628
rect 6169 13572 6173 13628
rect 6109 13568 6173 13572
rect 6189 13628 6253 13632
rect 6189 13572 6193 13628
rect 6193 13572 6249 13628
rect 6249 13572 6253 13628
rect 6189 13568 6253 13572
rect 10946 13628 11010 13632
rect 10946 13572 10950 13628
rect 10950 13572 11006 13628
rect 11006 13572 11010 13628
rect 10946 13568 11010 13572
rect 11026 13628 11090 13632
rect 11026 13572 11030 13628
rect 11030 13572 11086 13628
rect 11086 13572 11090 13628
rect 11026 13568 11090 13572
rect 11106 13628 11170 13632
rect 11106 13572 11110 13628
rect 11110 13572 11166 13628
rect 11166 13572 11170 13628
rect 11106 13568 11170 13572
rect 11186 13628 11250 13632
rect 11186 13572 11190 13628
rect 11190 13572 11246 13628
rect 11246 13572 11250 13628
rect 11186 13568 11250 13572
rect 14044 13228 14108 13292
rect 11468 13092 11532 13156
rect 3450 13084 3514 13088
rect 3450 13028 3454 13084
rect 3454 13028 3510 13084
rect 3510 13028 3514 13084
rect 3450 13024 3514 13028
rect 3530 13084 3594 13088
rect 3530 13028 3534 13084
rect 3534 13028 3590 13084
rect 3590 13028 3594 13084
rect 3530 13024 3594 13028
rect 3610 13084 3674 13088
rect 3610 13028 3614 13084
rect 3614 13028 3670 13084
rect 3670 13028 3674 13084
rect 3610 13024 3674 13028
rect 3690 13084 3754 13088
rect 3690 13028 3694 13084
rect 3694 13028 3750 13084
rect 3750 13028 3754 13084
rect 3690 13024 3754 13028
rect 8448 13084 8512 13088
rect 8448 13028 8452 13084
rect 8452 13028 8508 13084
rect 8508 13028 8512 13084
rect 8448 13024 8512 13028
rect 8528 13084 8592 13088
rect 8528 13028 8532 13084
rect 8532 13028 8588 13084
rect 8588 13028 8592 13084
rect 8528 13024 8592 13028
rect 8608 13084 8672 13088
rect 8608 13028 8612 13084
rect 8612 13028 8668 13084
rect 8668 13028 8672 13084
rect 8608 13024 8672 13028
rect 8688 13084 8752 13088
rect 8688 13028 8692 13084
rect 8692 13028 8748 13084
rect 8748 13028 8752 13084
rect 8688 13024 8752 13028
rect 13445 13084 13509 13088
rect 13445 13028 13449 13084
rect 13449 13028 13505 13084
rect 13505 13028 13509 13084
rect 13445 13024 13509 13028
rect 13525 13084 13589 13088
rect 13525 13028 13529 13084
rect 13529 13028 13585 13084
rect 13585 13028 13589 13084
rect 13525 13024 13589 13028
rect 13605 13084 13669 13088
rect 13605 13028 13609 13084
rect 13609 13028 13665 13084
rect 13665 13028 13669 13084
rect 13605 13024 13669 13028
rect 13685 13084 13749 13088
rect 13685 13028 13689 13084
rect 13689 13028 13745 13084
rect 13745 13028 13749 13084
rect 13685 13024 13749 13028
rect 11652 12956 11716 13020
rect 12020 12880 12084 12884
rect 12020 12824 12034 12880
rect 12034 12824 12084 12880
rect 12020 12820 12084 12824
rect 10548 12684 10612 12748
rect 9812 12548 9876 12612
rect 5949 12540 6013 12544
rect 5949 12484 5953 12540
rect 5953 12484 6009 12540
rect 6009 12484 6013 12540
rect 5949 12480 6013 12484
rect 6029 12540 6093 12544
rect 6029 12484 6033 12540
rect 6033 12484 6089 12540
rect 6089 12484 6093 12540
rect 6029 12480 6093 12484
rect 6109 12540 6173 12544
rect 6109 12484 6113 12540
rect 6113 12484 6169 12540
rect 6169 12484 6173 12540
rect 6109 12480 6173 12484
rect 6189 12540 6253 12544
rect 6189 12484 6193 12540
rect 6193 12484 6249 12540
rect 6249 12484 6253 12540
rect 6189 12480 6253 12484
rect 10946 12540 11010 12544
rect 10946 12484 10950 12540
rect 10950 12484 11006 12540
rect 11006 12484 11010 12540
rect 10946 12480 11010 12484
rect 11026 12540 11090 12544
rect 11026 12484 11030 12540
rect 11030 12484 11086 12540
rect 11086 12484 11090 12540
rect 11026 12480 11090 12484
rect 11106 12540 11170 12544
rect 11106 12484 11110 12540
rect 11110 12484 11166 12540
rect 11166 12484 11170 12540
rect 11106 12480 11170 12484
rect 11186 12540 11250 12544
rect 11186 12484 11190 12540
rect 11190 12484 11246 12540
rect 11246 12484 11250 12540
rect 11186 12480 11250 12484
rect 9996 12276 10060 12340
rect 12940 12276 13004 12340
rect 3450 11996 3514 12000
rect 3450 11940 3454 11996
rect 3454 11940 3510 11996
rect 3510 11940 3514 11996
rect 3450 11936 3514 11940
rect 3530 11996 3594 12000
rect 3530 11940 3534 11996
rect 3534 11940 3590 11996
rect 3590 11940 3594 11996
rect 3530 11936 3594 11940
rect 3610 11996 3674 12000
rect 3610 11940 3614 11996
rect 3614 11940 3670 11996
rect 3670 11940 3674 11996
rect 3610 11936 3674 11940
rect 3690 11996 3754 12000
rect 3690 11940 3694 11996
rect 3694 11940 3750 11996
rect 3750 11940 3754 11996
rect 3690 11936 3754 11940
rect 8448 11996 8512 12000
rect 8448 11940 8452 11996
rect 8452 11940 8508 11996
rect 8508 11940 8512 11996
rect 8448 11936 8512 11940
rect 8528 11996 8592 12000
rect 8528 11940 8532 11996
rect 8532 11940 8588 11996
rect 8588 11940 8592 11996
rect 8528 11936 8592 11940
rect 8608 11996 8672 12000
rect 8608 11940 8612 11996
rect 8612 11940 8668 11996
rect 8668 11940 8672 11996
rect 8608 11936 8672 11940
rect 8688 11996 8752 12000
rect 8688 11940 8692 11996
rect 8692 11940 8748 11996
rect 8748 11940 8752 11996
rect 8688 11936 8752 11940
rect 13445 11996 13509 12000
rect 13445 11940 13449 11996
rect 13449 11940 13505 11996
rect 13505 11940 13509 11996
rect 13445 11936 13509 11940
rect 13525 11996 13589 12000
rect 13525 11940 13529 11996
rect 13529 11940 13585 11996
rect 13585 11940 13589 11996
rect 13525 11936 13589 11940
rect 13605 11996 13669 12000
rect 13605 11940 13609 11996
rect 13609 11940 13665 11996
rect 13665 11940 13669 11996
rect 13605 11936 13669 11940
rect 13685 11996 13749 12000
rect 13685 11940 13689 11996
rect 13689 11940 13745 11996
rect 13745 11940 13749 11996
rect 13685 11936 13749 11940
rect 10364 11460 10428 11524
rect 5949 11452 6013 11456
rect 5949 11396 5953 11452
rect 5953 11396 6009 11452
rect 6009 11396 6013 11452
rect 5949 11392 6013 11396
rect 6029 11452 6093 11456
rect 6029 11396 6033 11452
rect 6033 11396 6089 11452
rect 6089 11396 6093 11452
rect 6029 11392 6093 11396
rect 6109 11452 6173 11456
rect 6109 11396 6113 11452
rect 6113 11396 6169 11452
rect 6169 11396 6173 11452
rect 6109 11392 6173 11396
rect 6189 11452 6253 11456
rect 6189 11396 6193 11452
rect 6193 11396 6249 11452
rect 6249 11396 6253 11452
rect 6189 11392 6253 11396
rect 10946 11452 11010 11456
rect 10946 11396 10950 11452
rect 10950 11396 11006 11452
rect 11006 11396 11010 11452
rect 10946 11392 11010 11396
rect 11026 11452 11090 11456
rect 11026 11396 11030 11452
rect 11030 11396 11086 11452
rect 11086 11396 11090 11452
rect 11026 11392 11090 11396
rect 11106 11452 11170 11456
rect 11106 11396 11110 11452
rect 11110 11396 11166 11452
rect 11166 11396 11170 11452
rect 11106 11392 11170 11396
rect 11186 11452 11250 11456
rect 11186 11396 11190 11452
rect 11190 11396 11246 11452
rect 11246 11396 11250 11452
rect 11186 11392 11250 11396
rect 12204 11324 12268 11388
rect 10732 11052 10796 11116
rect 12756 11112 12820 11116
rect 12756 11056 12770 11112
rect 12770 11056 12820 11112
rect 12756 11052 12820 11056
rect 3450 10908 3514 10912
rect 3450 10852 3454 10908
rect 3454 10852 3510 10908
rect 3510 10852 3514 10908
rect 3450 10848 3514 10852
rect 3530 10908 3594 10912
rect 3530 10852 3534 10908
rect 3534 10852 3590 10908
rect 3590 10852 3594 10908
rect 3530 10848 3594 10852
rect 3610 10908 3674 10912
rect 3610 10852 3614 10908
rect 3614 10852 3670 10908
rect 3670 10852 3674 10908
rect 3610 10848 3674 10852
rect 3690 10908 3754 10912
rect 3690 10852 3694 10908
rect 3694 10852 3750 10908
rect 3750 10852 3754 10908
rect 3690 10848 3754 10852
rect 8448 10908 8512 10912
rect 8448 10852 8452 10908
rect 8452 10852 8508 10908
rect 8508 10852 8512 10908
rect 8448 10848 8512 10852
rect 8528 10908 8592 10912
rect 8528 10852 8532 10908
rect 8532 10852 8588 10908
rect 8588 10852 8592 10908
rect 8528 10848 8592 10852
rect 8608 10908 8672 10912
rect 8608 10852 8612 10908
rect 8612 10852 8668 10908
rect 8668 10852 8672 10908
rect 8608 10848 8672 10852
rect 8688 10908 8752 10912
rect 8688 10852 8692 10908
rect 8692 10852 8748 10908
rect 8748 10852 8752 10908
rect 8688 10848 8752 10852
rect 9628 10780 9692 10844
rect 11836 10916 11900 10980
rect 13445 10908 13509 10912
rect 13445 10852 13449 10908
rect 13449 10852 13505 10908
rect 13505 10852 13509 10908
rect 13445 10848 13509 10852
rect 13525 10908 13589 10912
rect 13525 10852 13529 10908
rect 13529 10852 13585 10908
rect 13585 10852 13589 10908
rect 13525 10848 13589 10852
rect 13605 10908 13669 10912
rect 13605 10852 13609 10908
rect 13609 10852 13665 10908
rect 13665 10852 13669 10908
rect 13605 10848 13669 10852
rect 13685 10908 13749 10912
rect 13685 10852 13689 10908
rect 13689 10852 13745 10908
rect 13745 10852 13749 10908
rect 13685 10848 13749 10852
rect 13124 10780 13188 10844
rect 11468 10508 11532 10572
rect 5949 10364 6013 10368
rect 5949 10308 5953 10364
rect 5953 10308 6009 10364
rect 6009 10308 6013 10364
rect 5949 10304 6013 10308
rect 6029 10364 6093 10368
rect 6029 10308 6033 10364
rect 6033 10308 6089 10364
rect 6089 10308 6093 10364
rect 6029 10304 6093 10308
rect 6109 10364 6173 10368
rect 6109 10308 6113 10364
rect 6113 10308 6169 10364
rect 6169 10308 6173 10364
rect 6109 10304 6173 10308
rect 6189 10364 6253 10368
rect 6189 10308 6193 10364
rect 6193 10308 6249 10364
rect 6249 10308 6253 10364
rect 6189 10304 6253 10308
rect 10946 10364 11010 10368
rect 10946 10308 10950 10364
rect 10950 10308 11006 10364
rect 11006 10308 11010 10364
rect 10946 10304 11010 10308
rect 11026 10364 11090 10368
rect 11026 10308 11030 10364
rect 11030 10308 11086 10364
rect 11086 10308 11090 10364
rect 11026 10304 11090 10308
rect 11106 10364 11170 10368
rect 11106 10308 11110 10364
rect 11110 10308 11166 10364
rect 11166 10308 11170 10364
rect 11106 10304 11170 10308
rect 11186 10364 11250 10368
rect 11186 10308 11190 10364
rect 11190 10308 11246 10364
rect 11246 10308 11250 10364
rect 11186 10304 11250 10308
rect 8156 10100 8220 10164
rect 12388 10100 12452 10164
rect 12940 10236 13004 10300
rect 10732 9888 10796 9892
rect 10732 9832 10782 9888
rect 10782 9832 10796 9888
rect 10732 9828 10796 9832
rect 12204 9828 12268 9892
rect 3450 9820 3514 9824
rect 3450 9764 3454 9820
rect 3454 9764 3510 9820
rect 3510 9764 3514 9820
rect 3450 9760 3514 9764
rect 3530 9820 3594 9824
rect 3530 9764 3534 9820
rect 3534 9764 3590 9820
rect 3590 9764 3594 9820
rect 3530 9760 3594 9764
rect 3610 9820 3674 9824
rect 3610 9764 3614 9820
rect 3614 9764 3670 9820
rect 3670 9764 3674 9820
rect 3610 9760 3674 9764
rect 3690 9820 3754 9824
rect 3690 9764 3694 9820
rect 3694 9764 3750 9820
rect 3750 9764 3754 9820
rect 3690 9760 3754 9764
rect 8448 9820 8512 9824
rect 8448 9764 8452 9820
rect 8452 9764 8508 9820
rect 8508 9764 8512 9820
rect 8448 9760 8512 9764
rect 8528 9820 8592 9824
rect 8528 9764 8532 9820
rect 8532 9764 8588 9820
rect 8588 9764 8592 9820
rect 8528 9760 8592 9764
rect 8608 9820 8672 9824
rect 8608 9764 8612 9820
rect 8612 9764 8668 9820
rect 8668 9764 8672 9820
rect 8608 9760 8672 9764
rect 8688 9820 8752 9824
rect 8688 9764 8692 9820
rect 8692 9764 8748 9820
rect 8748 9764 8752 9820
rect 8688 9760 8752 9764
rect 13445 9820 13509 9824
rect 13445 9764 13449 9820
rect 13449 9764 13505 9820
rect 13505 9764 13509 9820
rect 13445 9760 13509 9764
rect 13525 9820 13589 9824
rect 13525 9764 13529 9820
rect 13529 9764 13585 9820
rect 13585 9764 13589 9820
rect 13525 9760 13589 9764
rect 13605 9820 13669 9824
rect 13605 9764 13609 9820
rect 13609 9764 13665 9820
rect 13665 9764 13669 9820
rect 13605 9760 13669 9764
rect 13685 9820 13749 9824
rect 13685 9764 13689 9820
rect 13689 9764 13745 9820
rect 13745 9764 13749 9820
rect 13685 9760 13749 9764
rect 3004 9616 3068 9620
rect 3004 9560 3054 9616
rect 3054 9560 3068 9616
rect 3004 9556 3068 9560
rect 5949 9276 6013 9280
rect 5949 9220 5953 9276
rect 5953 9220 6009 9276
rect 6009 9220 6013 9276
rect 5949 9216 6013 9220
rect 6029 9276 6093 9280
rect 6029 9220 6033 9276
rect 6033 9220 6089 9276
rect 6089 9220 6093 9276
rect 6029 9216 6093 9220
rect 6109 9276 6173 9280
rect 6109 9220 6113 9276
rect 6113 9220 6169 9276
rect 6169 9220 6173 9276
rect 6109 9216 6173 9220
rect 6189 9276 6253 9280
rect 6189 9220 6193 9276
rect 6193 9220 6249 9276
rect 6249 9220 6253 9276
rect 6189 9216 6253 9220
rect 12572 9420 12636 9484
rect 10946 9276 11010 9280
rect 10946 9220 10950 9276
rect 10950 9220 11006 9276
rect 11006 9220 11010 9276
rect 10946 9216 11010 9220
rect 11026 9276 11090 9280
rect 11026 9220 11030 9276
rect 11030 9220 11086 9276
rect 11086 9220 11090 9276
rect 11026 9216 11090 9220
rect 11106 9276 11170 9280
rect 11106 9220 11110 9276
rect 11110 9220 11166 9276
rect 11166 9220 11170 9276
rect 11106 9216 11170 9220
rect 11186 9276 11250 9280
rect 11186 9220 11190 9276
rect 11190 9220 11246 9276
rect 11246 9220 11250 9276
rect 11186 9216 11250 9220
rect 9812 9148 9876 9212
rect 12940 9208 13004 9212
rect 12940 9152 12954 9208
rect 12954 9152 13004 9208
rect 12940 9148 13004 9152
rect 14044 9148 14108 9212
rect 13860 9012 13924 9076
rect 3450 8732 3514 8736
rect 3450 8676 3454 8732
rect 3454 8676 3510 8732
rect 3510 8676 3514 8732
rect 3450 8672 3514 8676
rect 3530 8732 3594 8736
rect 3530 8676 3534 8732
rect 3534 8676 3590 8732
rect 3590 8676 3594 8732
rect 3530 8672 3594 8676
rect 3610 8732 3674 8736
rect 3610 8676 3614 8732
rect 3614 8676 3670 8732
rect 3670 8676 3674 8732
rect 3610 8672 3674 8676
rect 3690 8732 3754 8736
rect 3690 8676 3694 8732
rect 3694 8676 3750 8732
rect 3750 8676 3754 8732
rect 3690 8672 3754 8676
rect 8448 8732 8512 8736
rect 8448 8676 8452 8732
rect 8452 8676 8508 8732
rect 8508 8676 8512 8732
rect 8448 8672 8512 8676
rect 8528 8732 8592 8736
rect 8528 8676 8532 8732
rect 8532 8676 8588 8732
rect 8588 8676 8592 8732
rect 8528 8672 8592 8676
rect 8608 8732 8672 8736
rect 8608 8676 8612 8732
rect 8612 8676 8668 8732
rect 8668 8676 8672 8732
rect 8608 8672 8672 8676
rect 8688 8732 8752 8736
rect 8688 8676 8692 8732
rect 8692 8676 8748 8732
rect 8748 8676 8752 8732
rect 8688 8672 8752 8676
rect 13445 8732 13509 8736
rect 13445 8676 13449 8732
rect 13449 8676 13505 8732
rect 13505 8676 13509 8732
rect 13445 8672 13509 8676
rect 13525 8732 13589 8736
rect 13525 8676 13529 8732
rect 13529 8676 13585 8732
rect 13585 8676 13589 8732
rect 13525 8672 13589 8676
rect 13605 8732 13669 8736
rect 13605 8676 13609 8732
rect 13609 8676 13665 8732
rect 13665 8676 13669 8732
rect 13605 8672 13669 8676
rect 13685 8732 13749 8736
rect 13685 8676 13689 8732
rect 13689 8676 13745 8732
rect 13745 8676 13749 8732
rect 13685 8672 13749 8676
rect 9628 8604 9692 8668
rect 12756 8196 12820 8260
rect 13308 8256 13372 8260
rect 13308 8200 13322 8256
rect 13322 8200 13372 8256
rect 13308 8196 13372 8200
rect 5949 8188 6013 8192
rect 5949 8132 5953 8188
rect 5953 8132 6009 8188
rect 6009 8132 6013 8188
rect 5949 8128 6013 8132
rect 6029 8188 6093 8192
rect 6029 8132 6033 8188
rect 6033 8132 6089 8188
rect 6089 8132 6093 8188
rect 6029 8128 6093 8132
rect 6109 8188 6173 8192
rect 6109 8132 6113 8188
rect 6113 8132 6169 8188
rect 6169 8132 6173 8188
rect 6109 8128 6173 8132
rect 6189 8188 6253 8192
rect 6189 8132 6193 8188
rect 6193 8132 6249 8188
rect 6249 8132 6253 8188
rect 6189 8128 6253 8132
rect 10946 8188 11010 8192
rect 10946 8132 10950 8188
rect 10950 8132 11006 8188
rect 11006 8132 11010 8188
rect 10946 8128 11010 8132
rect 11026 8188 11090 8192
rect 11026 8132 11030 8188
rect 11030 8132 11086 8188
rect 11086 8132 11090 8188
rect 11026 8128 11090 8132
rect 11106 8188 11170 8192
rect 11106 8132 11110 8188
rect 11110 8132 11166 8188
rect 11166 8132 11170 8188
rect 11106 8128 11170 8132
rect 11186 8188 11250 8192
rect 11186 8132 11190 8188
rect 11190 8132 11246 8188
rect 11246 8132 11250 8188
rect 11186 8128 11250 8132
rect 4292 7924 4356 7988
rect 10732 8060 10796 8124
rect 11652 8060 11716 8124
rect 3450 7644 3514 7648
rect 3450 7588 3454 7644
rect 3454 7588 3510 7644
rect 3510 7588 3514 7644
rect 3450 7584 3514 7588
rect 3530 7644 3594 7648
rect 3530 7588 3534 7644
rect 3534 7588 3590 7644
rect 3590 7588 3594 7644
rect 3530 7584 3594 7588
rect 3610 7644 3674 7648
rect 3610 7588 3614 7644
rect 3614 7588 3670 7644
rect 3670 7588 3674 7644
rect 3610 7584 3674 7588
rect 3690 7644 3754 7648
rect 3690 7588 3694 7644
rect 3694 7588 3750 7644
rect 3750 7588 3754 7644
rect 3690 7584 3754 7588
rect 11836 7848 11900 7852
rect 11836 7792 11886 7848
rect 11886 7792 11900 7848
rect 11836 7788 11900 7792
rect 12204 7788 12268 7852
rect 5764 7652 5828 7716
rect 8448 7644 8512 7648
rect 8448 7588 8452 7644
rect 8452 7588 8508 7644
rect 8508 7588 8512 7644
rect 8448 7584 8512 7588
rect 8528 7644 8592 7648
rect 8528 7588 8532 7644
rect 8532 7588 8588 7644
rect 8588 7588 8592 7644
rect 8528 7584 8592 7588
rect 8608 7644 8672 7648
rect 8608 7588 8612 7644
rect 8612 7588 8668 7644
rect 8668 7588 8672 7644
rect 8608 7584 8672 7588
rect 8688 7644 8752 7648
rect 8688 7588 8692 7644
rect 8692 7588 8748 7644
rect 8748 7588 8752 7644
rect 8688 7584 8752 7588
rect 13445 7644 13509 7648
rect 13445 7588 13449 7644
rect 13449 7588 13505 7644
rect 13505 7588 13509 7644
rect 13445 7584 13509 7588
rect 13525 7644 13589 7648
rect 13525 7588 13529 7644
rect 13529 7588 13585 7644
rect 13585 7588 13589 7644
rect 13525 7584 13589 7588
rect 13605 7644 13669 7648
rect 13605 7588 13609 7644
rect 13609 7588 13665 7644
rect 13665 7588 13669 7644
rect 13605 7584 13669 7588
rect 13685 7644 13749 7648
rect 13685 7588 13689 7644
rect 13689 7588 13745 7644
rect 13745 7588 13749 7644
rect 13685 7584 13749 7588
rect 6684 7108 6748 7172
rect 10548 7168 10612 7172
rect 10548 7112 10598 7168
rect 10598 7112 10612 7168
rect 10548 7108 10612 7112
rect 5949 7100 6013 7104
rect 5949 7044 5953 7100
rect 5953 7044 6009 7100
rect 6009 7044 6013 7100
rect 5949 7040 6013 7044
rect 6029 7100 6093 7104
rect 6029 7044 6033 7100
rect 6033 7044 6089 7100
rect 6089 7044 6093 7100
rect 6029 7040 6093 7044
rect 6109 7100 6173 7104
rect 6109 7044 6113 7100
rect 6113 7044 6169 7100
rect 6169 7044 6173 7100
rect 6109 7040 6173 7044
rect 6189 7100 6253 7104
rect 6189 7044 6193 7100
rect 6193 7044 6249 7100
rect 6249 7044 6253 7100
rect 6189 7040 6253 7044
rect 10946 7100 11010 7104
rect 10946 7044 10950 7100
rect 10950 7044 11006 7100
rect 11006 7044 11010 7100
rect 10946 7040 11010 7044
rect 11026 7100 11090 7104
rect 11026 7044 11030 7100
rect 11030 7044 11086 7100
rect 11086 7044 11090 7100
rect 11026 7040 11090 7044
rect 11106 7100 11170 7104
rect 11106 7044 11110 7100
rect 11110 7044 11166 7100
rect 11166 7044 11170 7100
rect 11106 7040 11170 7044
rect 11186 7100 11250 7104
rect 11186 7044 11190 7100
rect 11190 7044 11246 7100
rect 11246 7044 11250 7100
rect 11186 7040 11250 7044
rect 12388 6836 12452 6900
rect 3450 6556 3514 6560
rect 3450 6500 3454 6556
rect 3454 6500 3510 6556
rect 3510 6500 3514 6556
rect 3450 6496 3514 6500
rect 3530 6556 3594 6560
rect 3530 6500 3534 6556
rect 3534 6500 3590 6556
rect 3590 6500 3594 6556
rect 3530 6496 3594 6500
rect 3610 6556 3674 6560
rect 3610 6500 3614 6556
rect 3614 6500 3670 6556
rect 3670 6500 3674 6556
rect 3610 6496 3674 6500
rect 3690 6556 3754 6560
rect 3690 6500 3694 6556
rect 3694 6500 3750 6556
rect 3750 6500 3754 6556
rect 3690 6496 3754 6500
rect 8448 6556 8512 6560
rect 8448 6500 8452 6556
rect 8452 6500 8508 6556
rect 8508 6500 8512 6556
rect 8448 6496 8512 6500
rect 8528 6556 8592 6560
rect 8528 6500 8532 6556
rect 8532 6500 8588 6556
rect 8588 6500 8592 6556
rect 8528 6496 8592 6500
rect 8608 6556 8672 6560
rect 8608 6500 8612 6556
rect 8612 6500 8668 6556
rect 8668 6500 8672 6556
rect 8608 6496 8672 6500
rect 8688 6556 8752 6560
rect 8688 6500 8692 6556
rect 8692 6500 8748 6556
rect 8748 6500 8752 6556
rect 8688 6496 8752 6500
rect 9996 6624 10060 6628
rect 9996 6568 10046 6624
rect 10046 6568 10060 6624
rect 9996 6564 10060 6568
rect 10180 6564 10244 6628
rect 13445 6556 13509 6560
rect 13445 6500 13449 6556
rect 13449 6500 13505 6556
rect 13505 6500 13509 6556
rect 13445 6496 13509 6500
rect 13525 6556 13589 6560
rect 13525 6500 13529 6556
rect 13529 6500 13585 6556
rect 13585 6500 13589 6556
rect 13525 6496 13589 6500
rect 13605 6556 13669 6560
rect 13605 6500 13609 6556
rect 13609 6500 13665 6556
rect 13665 6500 13669 6556
rect 13605 6496 13669 6500
rect 13685 6556 13749 6560
rect 13685 6500 13689 6556
rect 13689 6500 13745 6556
rect 13745 6500 13749 6556
rect 13685 6496 13749 6500
rect 8892 6156 8956 6220
rect 10548 6156 10612 6220
rect 10732 6156 10796 6220
rect 11468 6156 11532 6220
rect 12940 6292 13004 6356
rect 11652 6020 11716 6084
rect 12572 6020 12636 6084
rect 5949 6012 6013 6016
rect 5949 5956 5953 6012
rect 5953 5956 6009 6012
rect 6009 5956 6013 6012
rect 5949 5952 6013 5956
rect 6029 6012 6093 6016
rect 6029 5956 6033 6012
rect 6033 5956 6089 6012
rect 6089 5956 6093 6012
rect 6029 5952 6093 5956
rect 6109 6012 6173 6016
rect 6109 5956 6113 6012
rect 6113 5956 6169 6012
rect 6169 5956 6173 6012
rect 6109 5952 6173 5956
rect 6189 6012 6253 6016
rect 6189 5956 6193 6012
rect 6193 5956 6249 6012
rect 6249 5956 6253 6012
rect 6189 5952 6253 5956
rect 10946 6012 11010 6016
rect 10946 5956 10950 6012
rect 10950 5956 11006 6012
rect 11006 5956 11010 6012
rect 10946 5952 11010 5956
rect 11026 6012 11090 6016
rect 11026 5956 11030 6012
rect 11030 5956 11086 6012
rect 11086 5956 11090 6012
rect 11026 5952 11090 5956
rect 11106 6012 11170 6016
rect 11106 5956 11110 6012
rect 11110 5956 11166 6012
rect 11166 5956 11170 6012
rect 11106 5952 11170 5956
rect 11186 6012 11250 6016
rect 11186 5956 11190 6012
rect 11190 5956 11246 6012
rect 11246 5956 11250 6012
rect 11186 5952 11250 5956
rect 10548 5808 10612 5812
rect 10548 5752 10562 5808
rect 10562 5752 10612 5808
rect 10548 5748 10612 5752
rect 12572 5748 12636 5812
rect 13860 5748 13924 5812
rect 9076 5476 9140 5540
rect 3450 5468 3514 5472
rect 3450 5412 3454 5468
rect 3454 5412 3510 5468
rect 3510 5412 3514 5468
rect 3450 5408 3514 5412
rect 3530 5468 3594 5472
rect 3530 5412 3534 5468
rect 3534 5412 3590 5468
rect 3590 5412 3594 5468
rect 3530 5408 3594 5412
rect 3610 5468 3674 5472
rect 3610 5412 3614 5468
rect 3614 5412 3670 5468
rect 3670 5412 3674 5468
rect 3610 5408 3674 5412
rect 3690 5468 3754 5472
rect 3690 5412 3694 5468
rect 3694 5412 3750 5468
rect 3750 5412 3754 5468
rect 3690 5408 3754 5412
rect 8448 5468 8512 5472
rect 8448 5412 8452 5468
rect 8452 5412 8508 5468
rect 8508 5412 8512 5468
rect 8448 5408 8512 5412
rect 8528 5468 8592 5472
rect 8528 5412 8532 5468
rect 8532 5412 8588 5468
rect 8588 5412 8592 5468
rect 8528 5408 8592 5412
rect 8608 5468 8672 5472
rect 8608 5412 8612 5468
rect 8612 5412 8668 5468
rect 8668 5412 8672 5468
rect 8608 5408 8672 5412
rect 8688 5468 8752 5472
rect 8688 5412 8692 5468
rect 8692 5412 8748 5468
rect 8748 5412 8752 5468
rect 8688 5408 8752 5412
rect 13445 5468 13509 5472
rect 13445 5412 13449 5468
rect 13449 5412 13505 5468
rect 13505 5412 13509 5468
rect 13445 5408 13509 5412
rect 13525 5468 13589 5472
rect 13525 5412 13529 5468
rect 13529 5412 13585 5468
rect 13585 5412 13589 5468
rect 13525 5408 13589 5412
rect 13605 5468 13669 5472
rect 13605 5412 13609 5468
rect 13609 5412 13665 5468
rect 13665 5412 13669 5468
rect 13605 5408 13669 5412
rect 13685 5468 13749 5472
rect 13685 5412 13689 5468
rect 13689 5412 13745 5468
rect 13745 5412 13749 5468
rect 13685 5408 13749 5412
rect 3004 5204 3068 5268
rect 10364 5204 10428 5268
rect 11652 5068 11716 5132
rect 3188 4992 3252 4996
rect 3188 4936 3202 4992
rect 3202 4936 3252 4992
rect 3188 4932 3252 4936
rect 6500 4932 6564 4996
rect 12388 4932 12452 4996
rect 13124 4992 13188 4996
rect 13124 4936 13138 4992
rect 13138 4936 13188 4992
rect 13124 4932 13188 4936
rect 5949 4924 6013 4928
rect 5949 4868 5953 4924
rect 5953 4868 6009 4924
rect 6009 4868 6013 4924
rect 5949 4864 6013 4868
rect 6029 4924 6093 4928
rect 6029 4868 6033 4924
rect 6033 4868 6089 4924
rect 6089 4868 6093 4924
rect 6029 4864 6093 4868
rect 6109 4924 6173 4928
rect 6109 4868 6113 4924
rect 6113 4868 6169 4924
rect 6169 4868 6173 4924
rect 6109 4864 6173 4868
rect 6189 4924 6253 4928
rect 6189 4868 6193 4924
rect 6193 4868 6249 4924
rect 6249 4868 6253 4924
rect 6189 4864 6253 4868
rect 10946 4924 11010 4928
rect 10946 4868 10950 4924
rect 10950 4868 11006 4924
rect 11006 4868 11010 4924
rect 10946 4864 11010 4868
rect 11026 4924 11090 4928
rect 11026 4868 11030 4924
rect 11030 4868 11086 4924
rect 11086 4868 11090 4924
rect 11026 4864 11090 4868
rect 11106 4924 11170 4928
rect 11106 4868 11110 4924
rect 11110 4868 11166 4924
rect 11166 4868 11170 4924
rect 11106 4864 11170 4868
rect 11186 4924 11250 4928
rect 11186 4868 11190 4924
rect 11190 4868 11246 4924
rect 11246 4868 11250 4924
rect 11186 4864 11250 4868
rect 12020 4660 12084 4724
rect 9260 4448 9324 4452
rect 9260 4392 9310 4448
rect 9310 4392 9324 4448
rect 9260 4388 9324 4392
rect 9812 4448 9876 4452
rect 9812 4392 9826 4448
rect 9826 4392 9876 4448
rect 9812 4388 9876 4392
rect 10180 4448 10244 4452
rect 10180 4392 10194 4448
rect 10194 4392 10244 4448
rect 10180 4388 10244 4392
rect 3450 4380 3514 4384
rect 3450 4324 3454 4380
rect 3454 4324 3510 4380
rect 3510 4324 3514 4380
rect 3450 4320 3514 4324
rect 3530 4380 3594 4384
rect 3530 4324 3534 4380
rect 3534 4324 3590 4380
rect 3590 4324 3594 4380
rect 3530 4320 3594 4324
rect 3610 4380 3674 4384
rect 3610 4324 3614 4380
rect 3614 4324 3670 4380
rect 3670 4324 3674 4380
rect 3610 4320 3674 4324
rect 3690 4380 3754 4384
rect 3690 4324 3694 4380
rect 3694 4324 3750 4380
rect 3750 4324 3754 4380
rect 3690 4320 3754 4324
rect 8448 4380 8512 4384
rect 8448 4324 8452 4380
rect 8452 4324 8508 4380
rect 8508 4324 8512 4380
rect 8448 4320 8512 4324
rect 8528 4380 8592 4384
rect 8528 4324 8532 4380
rect 8532 4324 8588 4380
rect 8588 4324 8592 4380
rect 8528 4320 8592 4324
rect 8608 4380 8672 4384
rect 8608 4324 8612 4380
rect 8612 4324 8668 4380
rect 8668 4324 8672 4380
rect 8608 4320 8672 4324
rect 8688 4380 8752 4384
rect 8688 4324 8692 4380
rect 8692 4324 8748 4380
rect 8748 4324 8752 4380
rect 8688 4320 8752 4324
rect 4476 4312 4540 4316
rect 4476 4256 4490 4312
rect 4490 4256 4540 4312
rect 4476 4252 4540 4256
rect 13445 4380 13509 4384
rect 13445 4324 13449 4380
rect 13449 4324 13505 4380
rect 13505 4324 13509 4380
rect 13445 4320 13509 4324
rect 13525 4380 13589 4384
rect 13525 4324 13529 4380
rect 13529 4324 13585 4380
rect 13585 4324 13589 4380
rect 13525 4320 13589 4324
rect 13605 4380 13669 4384
rect 13605 4324 13609 4380
rect 13609 4324 13665 4380
rect 13665 4324 13669 4380
rect 13605 4320 13669 4324
rect 13685 4380 13749 4384
rect 13685 4324 13689 4380
rect 13689 4324 13745 4380
rect 13745 4324 13749 4380
rect 13685 4320 13749 4324
rect 10732 4116 10796 4180
rect 12756 3980 12820 4044
rect 6500 3904 6564 3908
rect 6500 3848 6514 3904
rect 6514 3848 6564 3904
rect 6500 3844 6564 3848
rect 9444 3844 9508 3908
rect 5949 3836 6013 3840
rect 5949 3780 5953 3836
rect 5953 3780 6009 3836
rect 6009 3780 6013 3836
rect 5949 3776 6013 3780
rect 6029 3836 6093 3840
rect 6029 3780 6033 3836
rect 6033 3780 6089 3836
rect 6089 3780 6093 3836
rect 6029 3776 6093 3780
rect 6109 3836 6173 3840
rect 6109 3780 6113 3836
rect 6113 3780 6169 3836
rect 6169 3780 6173 3836
rect 6109 3776 6173 3780
rect 6189 3836 6253 3840
rect 6189 3780 6193 3836
rect 6193 3780 6249 3836
rect 6249 3780 6253 3836
rect 6189 3776 6253 3780
rect 12020 3844 12084 3908
rect 12204 3844 12268 3908
rect 10946 3836 11010 3840
rect 10946 3780 10950 3836
rect 10950 3780 11006 3836
rect 11006 3780 11010 3836
rect 10946 3776 11010 3780
rect 11026 3836 11090 3840
rect 11026 3780 11030 3836
rect 11030 3780 11086 3836
rect 11086 3780 11090 3836
rect 11026 3776 11090 3780
rect 11106 3836 11170 3840
rect 11106 3780 11110 3836
rect 11110 3780 11166 3836
rect 11166 3780 11170 3836
rect 11106 3776 11170 3780
rect 11186 3836 11250 3840
rect 11186 3780 11190 3836
rect 11190 3780 11246 3836
rect 11246 3780 11250 3836
rect 11186 3776 11250 3780
rect 10732 3708 10796 3772
rect 12388 3708 12452 3772
rect 13308 3632 13372 3636
rect 13308 3576 13358 3632
rect 13358 3576 13372 3632
rect 13308 3572 13372 3576
rect 12020 3436 12084 3500
rect 12756 3436 12820 3500
rect 4292 3300 4356 3364
rect 8892 3300 8956 3364
rect 9812 3300 9876 3364
rect 10180 3300 10244 3364
rect 3450 3292 3514 3296
rect 3450 3236 3454 3292
rect 3454 3236 3510 3292
rect 3510 3236 3514 3292
rect 3450 3232 3514 3236
rect 3530 3292 3594 3296
rect 3530 3236 3534 3292
rect 3534 3236 3590 3292
rect 3590 3236 3594 3292
rect 3530 3232 3594 3236
rect 3610 3292 3674 3296
rect 3610 3236 3614 3292
rect 3614 3236 3670 3292
rect 3670 3236 3674 3292
rect 3610 3232 3674 3236
rect 3690 3292 3754 3296
rect 3690 3236 3694 3292
rect 3694 3236 3750 3292
rect 3750 3236 3754 3292
rect 3690 3232 3754 3236
rect 8448 3292 8512 3296
rect 8448 3236 8452 3292
rect 8452 3236 8508 3292
rect 8508 3236 8512 3292
rect 8448 3232 8512 3236
rect 8528 3292 8592 3296
rect 8528 3236 8532 3292
rect 8532 3236 8588 3292
rect 8588 3236 8592 3292
rect 8528 3232 8592 3236
rect 8608 3292 8672 3296
rect 8608 3236 8612 3292
rect 8612 3236 8668 3292
rect 8668 3236 8672 3292
rect 8608 3232 8672 3236
rect 8688 3292 8752 3296
rect 8688 3236 8692 3292
rect 8692 3236 8748 3292
rect 8748 3236 8752 3292
rect 8688 3232 8752 3236
rect 13445 3292 13509 3296
rect 13445 3236 13449 3292
rect 13449 3236 13505 3292
rect 13505 3236 13509 3292
rect 13445 3232 13509 3236
rect 13525 3292 13589 3296
rect 13525 3236 13529 3292
rect 13529 3236 13585 3292
rect 13585 3236 13589 3292
rect 13525 3232 13589 3236
rect 13605 3292 13669 3296
rect 13605 3236 13609 3292
rect 13609 3236 13665 3292
rect 13665 3236 13669 3292
rect 13605 3232 13669 3236
rect 13685 3292 13749 3296
rect 13685 3236 13689 3292
rect 13689 3236 13745 3292
rect 13745 3236 13749 3292
rect 13685 3232 13749 3236
rect 6684 2892 6748 2956
rect 9628 2892 9692 2956
rect 12572 3028 12636 3092
rect 6500 2816 6564 2820
rect 6500 2760 6550 2816
rect 6550 2760 6564 2816
rect 6500 2756 6564 2760
rect 10180 2756 10244 2820
rect 11836 2756 11900 2820
rect 14044 2756 14108 2820
rect 5949 2748 6013 2752
rect 5949 2692 5953 2748
rect 5953 2692 6009 2748
rect 6009 2692 6013 2748
rect 5949 2688 6013 2692
rect 6029 2748 6093 2752
rect 6029 2692 6033 2748
rect 6033 2692 6089 2748
rect 6089 2692 6093 2748
rect 6029 2688 6093 2692
rect 6109 2748 6173 2752
rect 6109 2692 6113 2748
rect 6113 2692 6169 2748
rect 6169 2692 6173 2748
rect 6109 2688 6173 2692
rect 6189 2748 6253 2752
rect 6189 2692 6193 2748
rect 6193 2692 6249 2748
rect 6249 2692 6253 2748
rect 6189 2688 6253 2692
rect 10946 2748 11010 2752
rect 10946 2692 10950 2748
rect 10950 2692 11006 2748
rect 11006 2692 11010 2748
rect 10946 2688 11010 2692
rect 11026 2748 11090 2752
rect 11026 2692 11030 2748
rect 11030 2692 11086 2748
rect 11086 2692 11090 2748
rect 11026 2688 11090 2692
rect 11106 2748 11170 2752
rect 11106 2692 11110 2748
rect 11110 2692 11166 2748
rect 11166 2692 11170 2748
rect 11106 2688 11170 2692
rect 11186 2748 11250 2752
rect 11186 2692 11190 2748
rect 11190 2692 11246 2748
rect 11246 2692 11250 2748
rect 11186 2688 11250 2692
rect 12388 2620 12452 2684
rect 3188 2484 3252 2548
rect 9260 2484 9324 2548
rect 9996 2484 10060 2548
rect 11652 2484 11716 2548
rect 12756 2484 12820 2548
rect 4476 2212 4540 2276
rect 11468 2212 11532 2276
rect 3450 2204 3514 2208
rect 3450 2148 3454 2204
rect 3454 2148 3510 2204
rect 3510 2148 3514 2204
rect 3450 2144 3514 2148
rect 3530 2204 3594 2208
rect 3530 2148 3534 2204
rect 3534 2148 3590 2204
rect 3590 2148 3594 2204
rect 3530 2144 3594 2148
rect 3610 2204 3674 2208
rect 3610 2148 3614 2204
rect 3614 2148 3670 2204
rect 3670 2148 3674 2204
rect 3610 2144 3674 2148
rect 3690 2204 3754 2208
rect 3690 2148 3694 2204
rect 3694 2148 3750 2204
rect 3750 2148 3754 2204
rect 3690 2144 3754 2148
rect 8448 2204 8512 2208
rect 8448 2148 8452 2204
rect 8452 2148 8508 2204
rect 8508 2148 8512 2204
rect 8448 2144 8512 2148
rect 8528 2204 8592 2208
rect 8528 2148 8532 2204
rect 8532 2148 8588 2204
rect 8588 2148 8592 2204
rect 8528 2144 8592 2148
rect 8608 2204 8672 2208
rect 8608 2148 8612 2204
rect 8612 2148 8668 2204
rect 8668 2148 8672 2204
rect 8608 2144 8672 2148
rect 8688 2204 8752 2208
rect 8688 2148 8692 2204
rect 8692 2148 8748 2204
rect 8748 2148 8752 2204
rect 8688 2144 8752 2148
rect 13445 2204 13509 2208
rect 13445 2148 13449 2204
rect 13449 2148 13505 2204
rect 13505 2148 13509 2204
rect 13445 2144 13509 2148
rect 13525 2204 13589 2208
rect 13525 2148 13529 2204
rect 13529 2148 13585 2204
rect 13585 2148 13589 2204
rect 13525 2144 13589 2148
rect 13605 2204 13669 2208
rect 13605 2148 13609 2204
rect 13609 2148 13665 2204
rect 13665 2148 13669 2204
rect 13605 2144 13669 2148
rect 13685 2204 13749 2208
rect 13685 2148 13689 2204
rect 13689 2148 13745 2204
rect 13745 2148 13749 2204
rect 13685 2144 13749 2148
rect 9076 1940 9140 2004
rect 12204 1940 12268 2004
rect 9444 1804 9508 1868
rect 12020 1668 12084 1732
<< metal4 >>
rect 3442 17440 3763 17456
rect 3442 17376 3450 17440
rect 3514 17376 3530 17440
rect 3594 17376 3610 17440
rect 3674 17376 3690 17440
rect 3754 17376 3763 17440
rect 3442 16352 3763 17376
rect 3442 16288 3450 16352
rect 3514 16288 3530 16352
rect 3594 16288 3610 16352
rect 3674 16288 3690 16352
rect 3754 16288 3763 16352
rect 3442 15264 3763 16288
rect 3442 15200 3450 15264
rect 3514 15200 3530 15264
rect 3594 15200 3610 15264
rect 3674 15200 3690 15264
rect 3754 15200 3763 15264
rect 3442 14176 3763 15200
rect 3442 14112 3450 14176
rect 3514 14112 3530 14176
rect 3594 14112 3610 14176
rect 3674 14112 3690 14176
rect 3754 14112 3763 14176
rect 3442 13088 3763 14112
rect 5941 16896 6261 17456
rect 5941 16832 5949 16896
rect 6013 16832 6029 16896
rect 6093 16832 6109 16896
rect 6173 16832 6189 16896
rect 6253 16832 6261 16896
rect 5941 15808 6261 16832
rect 8440 17440 8760 17456
rect 8440 17376 8448 17440
rect 8512 17376 8528 17440
rect 8592 17376 8608 17440
rect 8672 17376 8688 17440
rect 8752 17376 8760 17440
rect 6499 16420 6565 16421
rect 6499 16356 6500 16420
rect 6564 16356 6565 16420
rect 6499 16355 6565 16356
rect 5941 15744 5949 15808
rect 6013 15744 6029 15808
rect 6093 15744 6109 15808
rect 6173 15744 6189 15808
rect 6253 15744 6261 15808
rect 5941 14720 6261 15744
rect 5941 14656 5949 14720
rect 6013 14656 6029 14720
rect 6093 14656 6109 14720
rect 6173 14656 6189 14720
rect 6253 14656 6261 14720
rect 5763 13972 5829 13973
rect 5763 13908 5764 13972
rect 5828 13908 5829 13972
rect 5763 13907 5829 13908
rect 3442 13024 3450 13088
rect 3514 13024 3530 13088
rect 3594 13024 3610 13088
rect 3674 13024 3690 13088
rect 3754 13024 3763 13088
rect 3442 12000 3763 13024
rect 3442 11936 3450 12000
rect 3514 11936 3530 12000
rect 3594 11936 3610 12000
rect 3674 11936 3690 12000
rect 3754 11936 3763 12000
rect 3442 10912 3763 11936
rect 3442 10848 3450 10912
rect 3514 10848 3530 10912
rect 3594 10848 3610 10912
rect 3674 10848 3690 10912
rect 3754 10848 3763 10912
rect 3442 9824 3763 10848
rect 3442 9760 3450 9824
rect 3514 9760 3530 9824
rect 3594 9760 3610 9824
rect 3674 9760 3690 9824
rect 3754 9760 3763 9824
rect 3003 9620 3069 9621
rect 3003 9556 3004 9620
rect 3068 9556 3069 9620
rect 3003 9555 3069 9556
rect 3006 5269 3066 9555
rect 3442 8736 3763 9760
rect 3442 8672 3450 8736
rect 3514 8672 3530 8736
rect 3594 8672 3610 8736
rect 3674 8672 3690 8736
rect 3754 8672 3763 8736
rect 3442 7648 3763 8672
rect 4291 7988 4357 7989
rect 4291 7924 4292 7988
rect 4356 7924 4357 7988
rect 4291 7923 4357 7924
rect 3442 7584 3450 7648
rect 3514 7584 3530 7648
rect 3594 7584 3610 7648
rect 3674 7584 3690 7648
rect 3754 7584 3763 7648
rect 3442 6560 3763 7584
rect 3442 6496 3450 6560
rect 3514 6496 3530 6560
rect 3594 6496 3610 6560
rect 3674 6496 3690 6560
rect 3754 6496 3763 6560
rect 3442 5472 3763 6496
rect 3442 5408 3450 5472
rect 3514 5408 3530 5472
rect 3594 5408 3610 5472
rect 3674 5408 3690 5472
rect 3754 5408 3763 5472
rect 3003 5268 3069 5269
rect 3003 5204 3004 5268
rect 3068 5204 3069 5268
rect 3003 5203 3069 5204
rect 3187 4996 3253 4997
rect 3187 4932 3188 4996
rect 3252 4932 3253 4996
rect 3187 4931 3253 4932
rect 3190 2549 3250 4931
rect 3442 4384 3763 5408
rect 3442 4320 3450 4384
rect 3514 4320 3530 4384
rect 3594 4320 3610 4384
rect 3674 4320 3690 4384
rect 3754 4320 3763 4384
rect 3442 3296 3763 4320
rect 4294 3365 4354 7923
rect 5766 7717 5826 13907
rect 5941 13632 6261 14656
rect 5941 13568 5949 13632
rect 6013 13568 6029 13632
rect 6093 13568 6109 13632
rect 6173 13568 6189 13632
rect 6253 13568 6261 13632
rect 5941 12544 6261 13568
rect 5941 12480 5949 12544
rect 6013 12480 6029 12544
rect 6093 12480 6109 12544
rect 6173 12480 6189 12544
rect 6253 12480 6261 12544
rect 5941 11456 6261 12480
rect 5941 11392 5949 11456
rect 6013 11392 6029 11456
rect 6093 11392 6109 11456
rect 6173 11392 6189 11456
rect 6253 11392 6261 11456
rect 5941 10368 6261 11392
rect 5941 10304 5949 10368
rect 6013 10304 6029 10368
rect 6093 10304 6109 10368
rect 6173 10304 6189 10368
rect 6253 10304 6261 10368
rect 5941 9280 6261 10304
rect 5941 9216 5949 9280
rect 6013 9216 6029 9280
rect 6093 9216 6109 9280
rect 6173 9216 6189 9280
rect 6253 9216 6261 9280
rect 5941 8192 6261 9216
rect 5941 8128 5949 8192
rect 6013 8128 6029 8192
rect 6093 8128 6109 8192
rect 6173 8128 6189 8192
rect 6253 8128 6261 8192
rect 5763 7716 5829 7717
rect 5763 7652 5764 7716
rect 5828 7652 5829 7716
rect 5763 7651 5829 7652
rect 5941 7104 6261 8128
rect 5941 7040 5949 7104
rect 6013 7040 6029 7104
rect 6093 7040 6109 7104
rect 6173 7040 6189 7104
rect 6253 7040 6261 7104
rect 5941 6016 6261 7040
rect 5941 5952 5949 6016
rect 6013 5952 6029 6016
rect 6093 5952 6109 6016
rect 6173 5952 6189 6016
rect 6253 5952 6261 6016
rect 5941 4928 6261 5952
rect 6502 4997 6562 16355
rect 8440 16352 8760 17376
rect 10938 16896 11259 17456
rect 10938 16832 10946 16896
rect 11010 16832 11026 16896
rect 11090 16832 11106 16896
rect 11170 16832 11186 16896
rect 11250 16832 11259 16896
rect 9995 16556 10061 16557
rect 9995 16492 9996 16556
rect 10060 16492 10061 16556
rect 9995 16491 10061 16492
rect 8440 16288 8448 16352
rect 8512 16288 8528 16352
rect 8592 16288 8608 16352
rect 8672 16288 8688 16352
rect 8752 16288 8760 16352
rect 8440 15264 8760 16288
rect 9627 15876 9693 15877
rect 9627 15812 9628 15876
rect 9692 15812 9693 15876
rect 9627 15811 9693 15812
rect 8440 15200 8448 15264
rect 8512 15200 8528 15264
rect 8592 15200 8608 15264
rect 8672 15200 8688 15264
rect 8752 15200 8760 15264
rect 8440 14176 8760 15200
rect 8440 14112 8448 14176
rect 8512 14112 8528 14176
rect 8592 14112 8608 14176
rect 8672 14112 8688 14176
rect 8752 14112 8760 14176
rect 8155 13700 8221 13701
rect 8155 13636 8156 13700
rect 8220 13636 8221 13700
rect 8155 13635 8221 13636
rect 8158 10165 8218 13635
rect 8440 13088 8760 14112
rect 8440 13024 8448 13088
rect 8512 13024 8528 13088
rect 8592 13024 8608 13088
rect 8672 13024 8688 13088
rect 8752 13024 8760 13088
rect 8440 12000 8760 13024
rect 8440 11936 8448 12000
rect 8512 11936 8528 12000
rect 8592 11936 8608 12000
rect 8672 11936 8688 12000
rect 8752 11936 8760 12000
rect 8440 10912 8760 11936
rect 8440 10848 8448 10912
rect 8512 10848 8528 10912
rect 8592 10848 8608 10912
rect 8672 10848 8688 10912
rect 8752 10848 8760 10912
rect 8155 10164 8221 10165
rect 8155 10100 8156 10164
rect 8220 10100 8221 10164
rect 8155 10099 8221 10100
rect 8440 9824 8760 10848
rect 9630 10845 9690 15811
rect 9811 13972 9877 13973
rect 9811 13908 9812 13972
rect 9876 13908 9877 13972
rect 9811 13907 9877 13908
rect 9814 12613 9874 13907
rect 9811 12612 9877 12613
rect 9811 12548 9812 12612
rect 9876 12548 9877 12612
rect 9811 12547 9877 12548
rect 9998 12341 10058 16491
rect 10938 15808 11259 16832
rect 10938 15744 10946 15808
rect 11010 15744 11026 15808
rect 11090 15744 11106 15808
rect 11170 15744 11186 15808
rect 11250 15744 11259 15808
rect 10363 15060 10429 15061
rect 10363 14996 10364 15060
rect 10428 14996 10429 15060
rect 10363 14995 10429 14996
rect 9995 12340 10061 12341
rect 9995 12276 9996 12340
rect 10060 12276 10061 12340
rect 9995 12275 10061 12276
rect 10366 11525 10426 14995
rect 10938 14720 11259 15744
rect 10938 14656 10946 14720
rect 11010 14656 11026 14720
rect 11090 14656 11106 14720
rect 11170 14656 11186 14720
rect 11250 14656 11259 14720
rect 10938 13632 11259 14656
rect 10938 13568 10946 13632
rect 11010 13568 11026 13632
rect 11090 13568 11106 13632
rect 11170 13568 11186 13632
rect 11250 13568 11259 13632
rect 10547 12748 10613 12749
rect 10547 12684 10548 12748
rect 10612 12684 10613 12748
rect 10547 12683 10613 12684
rect 10363 11524 10429 11525
rect 10363 11460 10364 11524
rect 10428 11460 10429 11524
rect 10363 11459 10429 11460
rect 9627 10844 9693 10845
rect 9627 10780 9628 10844
rect 9692 10780 9693 10844
rect 9627 10779 9693 10780
rect 8440 9760 8448 9824
rect 8512 9760 8528 9824
rect 8592 9760 8608 9824
rect 8672 9760 8688 9824
rect 8752 9760 8760 9824
rect 8440 8736 8760 9760
rect 9811 9212 9877 9213
rect 9811 9148 9812 9212
rect 9876 9148 9877 9212
rect 9811 9147 9877 9148
rect 8440 8672 8448 8736
rect 8512 8672 8528 8736
rect 8592 8672 8608 8736
rect 8672 8672 8688 8736
rect 8752 8672 8760 8736
rect 8440 7648 8760 8672
rect 9627 8668 9693 8669
rect 9627 8604 9628 8668
rect 9692 8604 9693 8668
rect 9627 8603 9693 8604
rect 9630 8310 9690 8603
rect 8440 7584 8448 7648
rect 8512 7584 8528 7648
rect 8592 7584 8608 7648
rect 8672 7584 8688 7648
rect 8752 7584 8760 7648
rect 6683 7172 6749 7173
rect 6683 7108 6684 7172
rect 6748 7108 6749 7172
rect 6683 7107 6749 7108
rect 6499 4996 6565 4997
rect 6499 4932 6500 4996
rect 6564 4932 6565 4996
rect 6499 4931 6565 4932
rect 5941 4864 5949 4928
rect 6013 4864 6029 4928
rect 6093 4864 6109 4928
rect 6173 4864 6189 4928
rect 6253 4864 6261 4928
rect 4475 4316 4541 4317
rect 4475 4252 4476 4316
rect 4540 4252 4541 4316
rect 4475 4251 4541 4252
rect 4291 3364 4357 3365
rect 4291 3300 4292 3364
rect 4356 3300 4357 3364
rect 4291 3299 4357 3300
rect 3442 3232 3450 3296
rect 3514 3232 3530 3296
rect 3594 3232 3610 3296
rect 3674 3232 3690 3296
rect 3754 3232 3763 3296
rect 3187 2548 3253 2549
rect 3187 2484 3188 2548
rect 3252 2484 3253 2548
rect 3187 2483 3253 2484
rect 3442 2208 3763 3232
rect 4478 2277 4538 4251
rect 5941 3840 6261 4864
rect 6499 3908 6565 3909
rect 6499 3844 6500 3908
rect 6564 3844 6565 3908
rect 6499 3843 6565 3844
rect 5941 3776 5949 3840
rect 6013 3776 6029 3840
rect 6093 3776 6109 3840
rect 6173 3776 6189 3840
rect 6253 3776 6261 3840
rect 5941 2752 6261 3776
rect 6502 2821 6562 3843
rect 6686 2957 6746 7107
rect 8440 6560 8760 7584
rect 8440 6496 8448 6560
rect 8512 6496 8528 6560
rect 8592 6496 8608 6560
rect 8672 6496 8688 6560
rect 8752 6496 8760 6560
rect 8440 5472 8760 6496
rect 9446 8250 9690 8310
rect 8891 6220 8957 6221
rect 8891 6156 8892 6220
rect 8956 6156 8957 6220
rect 8891 6155 8957 6156
rect 8440 5408 8448 5472
rect 8512 5408 8528 5472
rect 8592 5408 8608 5472
rect 8672 5408 8688 5472
rect 8752 5408 8760 5472
rect 8440 4384 8760 5408
rect 8440 4320 8448 4384
rect 8512 4320 8528 4384
rect 8592 4320 8608 4384
rect 8672 4320 8688 4384
rect 8752 4320 8760 4384
rect 8440 3296 8760 4320
rect 8894 3365 8954 6155
rect 9075 5540 9141 5541
rect 9075 5476 9076 5540
rect 9140 5476 9141 5540
rect 9075 5475 9141 5476
rect 8891 3364 8957 3365
rect 8891 3300 8892 3364
rect 8956 3300 8957 3364
rect 8891 3299 8957 3300
rect 8440 3232 8448 3296
rect 8512 3232 8528 3296
rect 8592 3232 8608 3296
rect 8672 3232 8688 3296
rect 8752 3232 8760 3296
rect 6683 2956 6749 2957
rect 6683 2892 6684 2956
rect 6748 2892 6749 2956
rect 6683 2891 6749 2892
rect 6499 2820 6565 2821
rect 6499 2756 6500 2820
rect 6564 2756 6565 2820
rect 6499 2755 6565 2756
rect 5941 2688 5949 2752
rect 6013 2688 6029 2752
rect 6093 2688 6109 2752
rect 6173 2688 6189 2752
rect 6253 2688 6261 2752
rect 4475 2276 4541 2277
rect 4475 2212 4476 2276
rect 4540 2212 4541 2276
rect 4475 2211 4541 2212
rect 3442 2144 3450 2208
rect 3514 2144 3530 2208
rect 3594 2144 3610 2208
rect 3674 2144 3690 2208
rect 3754 2144 3763 2208
rect 3442 2128 3763 2144
rect 5941 2128 6261 2688
rect 8440 2208 8760 3232
rect 8440 2144 8448 2208
rect 8512 2144 8528 2208
rect 8592 2144 8608 2208
rect 8672 2144 8688 2208
rect 8752 2144 8760 2208
rect 8440 2128 8760 2144
rect 9078 2005 9138 5475
rect 9259 4452 9325 4453
rect 9259 4388 9260 4452
rect 9324 4388 9325 4452
rect 9259 4387 9325 4388
rect 9262 2549 9322 4387
rect 9446 3909 9506 8250
rect 9814 8122 9874 9147
rect 9630 8062 9874 8122
rect 9443 3908 9509 3909
rect 9443 3844 9444 3908
rect 9508 3844 9509 3908
rect 9443 3843 9509 3844
rect 9259 2548 9325 2549
rect 9259 2484 9260 2548
rect 9324 2484 9325 2548
rect 9259 2483 9325 2484
rect 9075 2004 9141 2005
rect 9075 1940 9076 2004
rect 9140 1940 9141 2004
rect 9075 1939 9141 1940
rect 9446 1869 9506 3843
rect 9630 2957 9690 8062
rect 9995 6628 10061 6629
rect 9995 6564 9996 6628
rect 10060 6564 10061 6628
rect 9995 6563 10061 6564
rect 10179 6628 10245 6629
rect 10179 6564 10180 6628
rect 10244 6564 10245 6628
rect 10179 6563 10245 6564
rect 9811 4452 9877 4453
rect 9811 4388 9812 4452
rect 9876 4388 9877 4452
rect 9811 4387 9877 4388
rect 9814 3365 9874 4387
rect 9811 3364 9877 3365
rect 9811 3300 9812 3364
rect 9876 3300 9877 3364
rect 9811 3299 9877 3300
rect 9627 2956 9693 2957
rect 9627 2892 9628 2956
rect 9692 2892 9693 2956
rect 9627 2891 9693 2892
rect 9998 2549 10058 6563
rect 10182 4453 10242 6563
rect 10366 5269 10426 11459
rect 10550 7173 10610 12683
rect 10938 12544 11259 13568
rect 13437 17440 13757 17456
rect 13437 17376 13445 17440
rect 13509 17376 13525 17440
rect 13589 17376 13605 17440
rect 13669 17376 13685 17440
rect 13749 17376 13757 17440
rect 13437 16352 13757 17376
rect 13437 16288 13445 16352
rect 13509 16288 13525 16352
rect 13589 16288 13605 16352
rect 13669 16288 13685 16352
rect 13749 16288 13757 16352
rect 13437 15264 13757 16288
rect 13437 15200 13445 15264
rect 13509 15200 13525 15264
rect 13589 15200 13605 15264
rect 13669 15200 13685 15264
rect 13749 15200 13757 15264
rect 13437 14176 13757 15200
rect 13437 14112 13445 14176
rect 13509 14112 13525 14176
rect 13589 14112 13605 14176
rect 13669 14112 13685 14176
rect 13749 14112 13757 14176
rect 11467 13156 11533 13157
rect 11467 13092 11468 13156
rect 11532 13092 11533 13156
rect 11467 13091 11533 13092
rect 10938 12480 10946 12544
rect 11010 12480 11026 12544
rect 11090 12480 11106 12544
rect 11170 12480 11186 12544
rect 11250 12480 11259 12544
rect 10938 11456 11259 12480
rect 10938 11392 10946 11456
rect 11010 11392 11026 11456
rect 11090 11392 11106 11456
rect 11170 11392 11186 11456
rect 11250 11392 11259 11456
rect 10731 11116 10797 11117
rect 10731 11052 10732 11116
rect 10796 11052 10797 11116
rect 10731 11051 10797 11052
rect 10734 9893 10794 11051
rect 10938 10368 11259 11392
rect 11470 10573 11530 13091
rect 13437 13088 13757 14112
rect 14043 13292 14109 13293
rect 14043 13228 14044 13292
rect 14108 13228 14109 13292
rect 14043 13227 14109 13228
rect 13437 13024 13445 13088
rect 13509 13024 13525 13088
rect 13589 13024 13605 13088
rect 13669 13024 13685 13088
rect 13749 13024 13757 13088
rect 11651 13020 11717 13021
rect 11651 12956 11652 13020
rect 11716 12956 11717 13020
rect 11651 12955 11717 12956
rect 11467 10572 11533 10573
rect 11467 10508 11468 10572
rect 11532 10508 11533 10572
rect 11467 10507 11533 10508
rect 10938 10304 10946 10368
rect 11010 10304 11026 10368
rect 11090 10304 11106 10368
rect 11170 10304 11186 10368
rect 11250 10304 11259 10368
rect 10731 9892 10797 9893
rect 10731 9828 10732 9892
rect 10796 9828 10797 9892
rect 10731 9827 10797 9828
rect 10938 9280 11259 10304
rect 10938 9216 10946 9280
rect 11010 9216 11026 9280
rect 11090 9216 11106 9280
rect 11170 9216 11186 9280
rect 11250 9216 11259 9280
rect 10938 8192 11259 9216
rect 10938 8128 10946 8192
rect 11010 8128 11026 8192
rect 11090 8128 11106 8192
rect 11170 8128 11186 8192
rect 11250 8128 11259 8192
rect 10731 8124 10797 8125
rect 10731 8060 10732 8124
rect 10796 8060 10797 8124
rect 10731 8059 10797 8060
rect 10547 7172 10613 7173
rect 10547 7108 10548 7172
rect 10612 7108 10613 7172
rect 10547 7107 10613 7108
rect 10734 6221 10794 8059
rect 10938 7104 11259 8128
rect 10938 7040 10946 7104
rect 11010 7040 11026 7104
rect 11090 7040 11106 7104
rect 11170 7040 11186 7104
rect 11250 7040 11259 7104
rect 10547 6220 10613 6221
rect 10547 6156 10548 6220
rect 10612 6156 10613 6220
rect 10547 6155 10613 6156
rect 10731 6220 10797 6221
rect 10731 6156 10732 6220
rect 10796 6156 10797 6220
rect 10731 6155 10797 6156
rect 10550 5813 10610 6155
rect 10938 6016 11259 7040
rect 11470 6354 11530 10507
rect 11654 8125 11714 12955
rect 12019 12884 12085 12885
rect 12019 12820 12020 12884
rect 12084 12820 12085 12884
rect 12019 12819 12085 12820
rect 11835 10980 11901 10981
rect 11835 10916 11836 10980
rect 11900 10916 11901 10980
rect 11835 10915 11901 10916
rect 11651 8124 11717 8125
rect 11651 8060 11652 8124
rect 11716 8060 11717 8124
rect 11651 8059 11717 8060
rect 11838 7853 11898 10915
rect 11835 7852 11901 7853
rect 11835 7788 11836 7852
rect 11900 7788 11901 7852
rect 11835 7787 11901 7788
rect 11470 6294 11714 6354
rect 11467 6220 11533 6221
rect 11467 6156 11468 6220
rect 11532 6156 11533 6220
rect 11467 6155 11533 6156
rect 10938 5952 10946 6016
rect 11010 5952 11026 6016
rect 11090 5952 11106 6016
rect 11170 5952 11186 6016
rect 11250 5952 11259 6016
rect 10547 5812 10613 5813
rect 10547 5748 10548 5812
rect 10612 5748 10613 5812
rect 10547 5747 10613 5748
rect 10363 5268 10429 5269
rect 10363 5204 10364 5268
rect 10428 5204 10429 5268
rect 10363 5203 10429 5204
rect 10938 4928 11259 5952
rect 10938 4864 10946 4928
rect 11010 4864 11026 4928
rect 11090 4864 11106 4928
rect 11170 4864 11186 4928
rect 11250 4864 11259 4928
rect 10179 4452 10245 4453
rect 10179 4388 10180 4452
rect 10244 4388 10245 4452
rect 10179 4387 10245 4388
rect 10731 4180 10797 4181
rect 10731 4116 10732 4180
rect 10796 4116 10797 4180
rect 10731 4115 10797 4116
rect 10734 3773 10794 4115
rect 10938 3840 11259 4864
rect 10938 3776 10946 3840
rect 11010 3776 11026 3840
rect 11090 3776 11106 3840
rect 11170 3776 11186 3840
rect 11250 3776 11259 3840
rect 10731 3772 10797 3773
rect 10731 3708 10732 3772
rect 10796 3708 10797 3772
rect 10731 3707 10797 3708
rect 10179 3364 10245 3365
rect 10179 3300 10180 3364
rect 10244 3300 10245 3364
rect 10179 3299 10245 3300
rect 10182 2821 10242 3299
rect 10179 2820 10245 2821
rect 10179 2756 10180 2820
rect 10244 2756 10245 2820
rect 10179 2755 10245 2756
rect 10938 2752 11259 3776
rect 10938 2688 10946 2752
rect 11010 2688 11026 2752
rect 11090 2688 11106 2752
rect 11170 2688 11186 2752
rect 11250 2688 11259 2752
rect 9995 2548 10061 2549
rect 9995 2484 9996 2548
rect 10060 2484 10061 2548
rect 9995 2483 10061 2484
rect 10938 2128 11259 2688
rect 11470 2277 11530 6155
rect 11654 6085 11714 6294
rect 11651 6084 11717 6085
rect 11651 6020 11652 6084
rect 11716 6020 11717 6084
rect 11651 6019 11717 6020
rect 11651 5132 11717 5133
rect 11651 5068 11652 5132
rect 11716 5068 11717 5132
rect 11651 5067 11717 5068
rect 11654 2549 11714 5067
rect 11838 2821 11898 7787
rect 12022 4725 12082 12819
rect 12939 12340 13005 12341
rect 12939 12276 12940 12340
rect 13004 12276 13005 12340
rect 12939 12275 13005 12276
rect 12203 11388 12269 11389
rect 12203 11324 12204 11388
rect 12268 11324 12269 11388
rect 12203 11323 12269 11324
rect 12206 9893 12266 11323
rect 12755 11116 12821 11117
rect 12755 11052 12756 11116
rect 12820 11052 12821 11116
rect 12755 11051 12821 11052
rect 12387 10164 12453 10165
rect 12387 10100 12388 10164
rect 12452 10100 12453 10164
rect 12387 10099 12453 10100
rect 12203 9892 12269 9893
rect 12203 9828 12204 9892
rect 12268 9828 12269 9892
rect 12203 9827 12269 9828
rect 12203 7852 12269 7853
rect 12203 7788 12204 7852
rect 12268 7788 12269 7852
rect 12203 7787 12269 7788
rect 12019 4724 12085 4725
rect 12019 4660 12020 4724
rect 12084 4660 12085 4724
rect 12019 4659 12085 4660
rect 12206 3909 12266 7787
rect 12390 6901 12450 10099
rect 12571 9484 12637 9485
rect 12571 9420 12572 9484
rect 12636 9420 12637 9484
rect 12571 9419 12637 9420
rect 12387 6900 12453 6901
rect 12387 6836 12388 6900
rect 12452 6836 12453 6900
rect 12387 6835 12453 6836
rect 12390 4997 12450 6835
rect 12574 6085 12634 9419
rect 12758 8261 12818 11051
rect 12942 10301 13002 12275
rect 13437 12000 13757 13024
rect 13437 11936 13445 12000
rect 13509 11936 13525 12000
rect 13589 11936 13605 12000
rect 13669 11936 13685 12000
rect 13749 11936 13757 12000
rect 13437 10912 13757 11936
rect 13437 10848 13445 10912
rect 13509 10848 13525 10912
rect 13589 10848 13605 10912
rect 13669 10848 13685 10912
rect 13749 10848 13757 10912
rect 13123 10844 13189 10845
rect 13123 10780 13124 10844
rect 13188 10780 13189 10844
rect 13123 10779 13189 10780
rect 12939 10300 13005 10301
rect 12939 10236 12940 10300
rect 13004 10236 13005 10300
rect 12939 10235 13005 10236
rect 12942 9213 13002 10235
rect 12939 9212 13005 9213
rect 12939 9148 12940 9212
rect 13004 9148 13005 9212
rect 12939 9147 13005 9148
rect 12755 8260 12821 8261
rect 12755 8196 12756 8260
rect 12820 8196 12821 8260
rect 12755 8195 12821 8196
rect 12571 6084 12637 6085
rect 12571 6020 12572 6084
rect 12636 6020 12637 6084
rect 12571 6019 12637 6020
rect 12571 5812 12637 5813
rect 12571 5748 12572 5812
rect 12636 5748 12637 5812
rect 12571 5747 12637 5748
rect 12387 4996 12453 4997
rect 12387 4932 12388 4996
rect 12452 4932 12453 4996
rect 12387 4931 12453 4932
rect 12019 3908 12085 3909
rect 12019 3844 12020 3908
rect 12084 3844 12085 3908
rect 12019 3843 12085 3844
rect 12203 3908 12269 3909
rect 12203 3844 12204 3908
rect 12268 3844 12269 3908
rect 12203 3843 12269 3844
rect 12022 3770 12082 3843
rect 12387 3772 12453 3773
rect 12022 3710 12266 3770
rect 12019 3500 12085 3501
rect 12019 3436 12020 3500
rect 12084 3436 12085 3500
rect 12019 3435 12085 3436
rect 11835 2820 11901 2821
rect 11835 2756 11836 2820
rect 11900 2756 11901 2820
rect 11835 2755 11901 2756
rect 11651 2548 11717 2549
rect 11651 2484 11652 2548
rect 11716 2484 11717 2548
rect 11651 2483 11717 2484
rect 11467 2276 11533 2277
rect 11467 2212 11468 2276
rect 11532 2212 11533 2276
rect 11467 2211 11533 2212
rect 9443 1868 9509 1869
rect 9443 1804 9444 1868
rect 9508 1804 9509 1868
rect 9443 1803 9509 1804
rect 12022 1733 12082 3435
rect 12206 2005 12266 3710
rect 12387 3708 12388 3772
rect 12452 3708 12453 3772
rect 12387 3707 12453 3708
rect 12390 2685 12450 3707
rect 12574 3093 12634 5747
rect 12758 4045 12818 8195
rect 12942 6357 13002 9147
rect 12939 6356 13005 6357
rect 12939 6292 12940 6356
rect 13004 6292 13005 6356
rect 12939 6291 13005 6292
rect 13126 4997 13186 10779
rect 13437 9824 13757 10848
rect 13437 9760 13445 9824
rect 13509 9760 13525 9824
rect 13589 9760 13605 9824
rect 13669 9760 13685 9824
rect 13749 9760 13757 9824
rect 13437 8736 13757 9760
rect 14046 9213 14106 13227
rect 14043 9212 14109 9213
rect 14043 9148 14044 9212
rect 14108 9148 14109 9212
rect 14043 9147 14109 9148
rect 13859 9076 13925 9077
rect 13859 9012 13860 9076
rect 13924 9012 13925 9076
rect 13859 9011 13925 9012
rect 13437 8672 13445 8736
rect 13509 8672 13525 8736
rect 13589 8672 13605 8736
rect 13669 8672 13685 8736
rect 13749 8672 13757 8736
rect 13307 8260 13373 8261
rect 13307 8196 13308 8260
rect 13372 8196 13373 8260
rect 13307 8195 13373 8196
rect 13123 4996 13189 4997
rect 13123 4932 13124 4996
rect 13188 4932 13189 4996
rect 13123 4931 13189 4932
rect 12755 4044 12821 4045
rect 12755 3980 12756 4044
rect 12820 3980 12821 4044
rect 12755 3979 12821 3980
rect 13310 3637 13370 8195
rect 13437 7648 13757 8672
rect 13437 7584 13445 7648
rect 13509 7584 13525 7648
rect 13589 7584 13605 7648
rect 13669 7584 13685 7648
rect 13749 7584 13757 7648
rect 13437 6560 13757 7584
rect 13437 6496 13445 6560
rect 13509 6496 13525 6560
rect 13589 6496 13605 6560
rect 13669 6496 13685 6560
rect 13749 6496 13757 6560
rect 13437 5472 13757 6496
rect 13862 5813 13922 9011
rect 13859 5812 13925 5813
rect 13859 5748 13860 5812
rect 13924 5748 13925 5812
rect 13859 5747 13925 5748
rect 13437 5408 13445 5472
rect 13509 5408 13525 5472
rect 13589 5408 13605 5472
rect 13669 5408 13685 5472
rect 13749 5408 13757 5472
rect 13437 4384 13757 5408
rect 13437 4320 13445 4384
rect 13509 4320 13525 4384
rect 13589 4320 13605 4384
rect 13669 4320 13685 4384
rect 13749 4320 13757 4384
rect 13307 3636 13373 3637
rect 13307 3572 13308 3636
rect 13372 3572 13373 3636
rect 13307 3571 13373 3572
rect 12755 3500 12821 3501
rect 12755 3436 12756 3500
rect 12820 3436 12821 3500
rect 12755 3435 12821 3436
rect 12571 3092 12637 3093
rect 12571 3028 12572 3092
rect 12636 3028 12637 3092
rect 12571 3027 12637 3028
rect 12387 2684 12453 2685
rect 12387 2620 12388 2684
rect 12452 2620 12453 2684
rect 12387 2619 12453 2620
rect 12758 2549 12818 3435
rect 13437 3296 13757 4320
rect 13437 3232 13445 3296
rect 13509 3232 13525 3296
rect 13589 3232 13605 3296
rect 13669 3232 13685 3296
rect 13749 3232 13757 3296
rect 12755 2548 12821 2549
rect 12755 2484 12756 2548
rect 12820 2484 12821 2548
rect 12755 2483 12821 2484
rect 13437 2208 13757 3232
rect 14046 2821 14106 9147
rect 14043 2820 14109 2821
rect 14043 2756 14044 2820
rect 14108 2756 14109 2820
rect 14043 2755 14109 2756
rect 13437 2144 13445 2208
rect 13509 2144 13525 2208
rect 13589 2144 13605 2208
rect 13669 2144 13685 2208
rect 13749 2144 13757 2208
rect 13437 2128 13757 2144
rect 12203 2004 12269 2005
rect 12203 1940 12204 2004
rect 12268 1940 12269 2004
rect 12203 1939 12269 1940
rect 12019 1732 12085 1733
rect 12019 1668 12020 1732
rect 12084 1668 12085 1732
rect 12019 1667 12085 1668
use sky130_fd_sc_hd__diode_2  ANTENNA__32__A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 1932 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output65 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 2116 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output64
timestamp 1624635492
transform -1 0 1748 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output58
timestamp 1624635492
transform 1 0 1932 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output53
timestamp 1624635492
transform -1 0 1748 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1624635492
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output69
timestamp 1624635492
transform -1 0 3220 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output68
timestamp 1624635492
transform -1 0 2852 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output67
timestamp 1624635492
transform -1 0 2484 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 2300 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l4_in_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 4692 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output54
timestamp 1624635492
transform -1 0 4232 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output55
timestamp 1624635492
transform -1 0 4600 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output56
timestamp 1624635492
transform -1 0 4968 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output59
timestamp 1624635492
transform 1 0 4324 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output70
timestamp 1624635492
transform -1 0 3588 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output71
timestamp 1624635492
transform -1 0 3956 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output72
timestamp 1624635492
transform -1 0 4324 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _36_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 5336 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_1_
timestamp 1624635492
transform 1 0 6440 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_0_
timestamp 1624635492
transform 1 0 5520 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_1_
timestamp 1624635492
transform 1 0 6532 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_1_
timestamp 1624635492
transform 1 0 5612 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1624635492
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1624635492
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output57
timestamp 1624635492
transform -1 0 5336 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_3_
timestamp 1624635492
transform 1 0 7268 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_1_
timestamp 1624635492
transform 1 0 7360 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_1_
timestamp 1624635492
transform 1 0 8096 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  input5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 8556 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input16
timestamp 1624635492
transform -1 0 8924 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1624635492
transform -1 0 9108 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1624635492
transform -1 0 9292 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input17
timestamp 1624635492
transform -1 0 9568 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1624635492
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1624635492
transform -1 0 9660 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input18
timestamp 1624635492
transform -1 0 9936 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _42_
timestamp 1624635492
transform 1 0 9660 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 9936 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1624635492
transform -1 0 10396 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _45_
timestamp 1624635492
transform 1 0 9936 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1624635492
transform -1 0 10764 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _48_
timestamp 1624635492
transform -1 0 10764 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _46_
timestamp 1624635492
transform 1 0 10212 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output61
timestamp 1624635492
transform -1 0 11500 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output60
timestamp 1624635492
transform -1 0 11132 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 11316 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _51_
timestamp 1624635492
transform 1 0 10764 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1624635492
transform -1 0 11592 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1624635492
transform -1 0 11776 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_118
timestamp 1624635492
transform 1 0 11960 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1624635492
transform -1 0 12236 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1624635492
transform 1 0 11684 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1624635492
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1624635492
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_122
timestamp 1624635492
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output62
timestamp 1624635492
transform -1 0 12604 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1624635492
transform -1 0 12696 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1624635492
transform -1 0 12328 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1624635492
transform -1 0 12788 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1624635492
transform -1 0 13064 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1624635492
transform -1 0 12880 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1624635492
transform -1 0 13156 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_134
timestamp 1624635492
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1624635492
transform -1 0 13432 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1624635492
transform -1 0 13248 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1624635492
transform -1 0 13524 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1624635492
transform -1 0 13892 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1624635492
transform -1 0 13708 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1624635492
transform -1 0 14076 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1624635492
transform -1 0 13800 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1624635492
transform 1 0 13800 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input45
timestamp 1624635492
transform -1 0 14352 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_3_S_FTB01
timestamp 1624635492
transform -1 0 14628 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_2_S_FTB01
timestamp 1624635492
transform -1 0 14444 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1624635492
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_146
timestamp 1624635492
transform 1 0 14536 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output116
timestamp 1624635492
transform 1 0 14628 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_3_S_FTB01
timestamp 1624635492
transform -1 0 14904 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_2_S_FTB01
timestamp 1624635492
transform 1 0 14904 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1624635492
transform -1 0 15364 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output118
timestamp 1624635492
transform 1 0 15364 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output96
timestamp 1624635492
transform 1 0 14996 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output94
timestamp 1624635492
transform 1 0 15364 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1624635492
transform -1 0 16008 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1624635492
transform -1 0 16008 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _32_
timestamp 1624635492
transform 1 0 2392 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _33_
timestamp 1624635492
transform 1 0 2668 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _34_
timestamp 1624635492
transform 1 0 2944 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 2116 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1624635492
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output66
timestamp 1624635492
transform -1 0 1748 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output97
timestamp 1624635492
transform -1 0 2116 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _35_
timestamp 1624635492
transform 1 0 3220 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _37_
timestamp 1624635492
transform 1 0 3496 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l4_in_0_
timestamp 1624635492
transform 1 0 4692 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l4_in_0_
timestamp 1624635492
transform 1 0 3864 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1624635492
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _38_
timestamp 1624635492
transform 1 0 5520 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_1_
timestamp 1624635492
transform 1 0 5796 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_2_
timestamp 1624635492
transform -1 0 7452 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _21_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 8648 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_2_
timestamp 1624635492
transform 1 0 7452 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  output63
timestamp 1624635492
transform -1 0 8648 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _47_
timestamp 1624635492
transform 1 0 9936 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _49_
timestamp 1624635492
transform -1 0 10488 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _50_
timestamp 1624635492
transform -1 0 10764 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_2_
timestamp 1624635492
transform 1 0 9108 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1624635492
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_85
timestamp 1624635492
transform 1 0 8924 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_S_FTB01 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 11868 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1624635492
transform 1 0 10764 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 1624635492
transform -1 0 11316 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1624635492
transform -1 0 11500 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1624635492
transform -1 0 11684 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1624635492
transform -1 0 11868 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1624635492
transform -1 0 12604 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1624635492
transform -1 0 12788 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1624635492
transform -1 0 12972 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 12972 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1624635492
transform 1 0 13340 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 13156 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 13524 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1624635492
transform 1 0 13892 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1624635492
transform 1 0 13708 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1624635492
transform 1 0 14076 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1624635492
transform -1 0 14536 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1624635492
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1624635492
transform -1 0 16008 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input46
timestamp 1624635492
transform -1 0 14812 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input47
timestamp 1624635492
transform 1 0 14812 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input48
timestamp 1624635492
transform -1 0 15364 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output52
timestamp 1624635492
transform 1 0 15364 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _40_
timestamp 1624635492
transform -1 0 3036 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _41_
timestamp 1624635492
transform -1 0 2760 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _43_
timestamp 1624635492
transform -1 0 2484 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1624635492
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output98
timestamp 1624635492
transform -1 0 1748 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output99
timestamp 1624635492
transform -1 0 2116 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_11
timestamp 1624635492
transform 1 0 2116 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_0_
timestamp 1624635492
transform 1 0 4692 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_1_
timestamp 1624635492
transform 1 0 3864 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l4_in_0_
timestamp 1624635492
transform 1 0 3036 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 6440 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_0_
timestamp 1624635492
transform 1 0 5520 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1624635492
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_1_
timestamp 1624635492
transform 1 0 7912 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_1_
timestamp 1624635492
transform 1 0 8740 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _44_
timestamp 1624635492
transform 1 0 10396 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_1_
timestamp 1624635492
transform 1 0 9568 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_right_ipin_0.prog_clk
timestamp 1624635492
transform 1 0 10672 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_right_ipin_0.prog_clk
timestamp 1624635492
transform 1 0 10948 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1624635492
transform -1 0 11408 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1624635492
transform -1 0 11868 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1624635492
transform -1 0 11592 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1624635492
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1624635492
transform -1 0 12236 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1624635492
transform -1 0 12052 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 12420 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_S_FTB01_A
timestamp 1624635492
transform -1 0 12420 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 12604 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 12788 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1624635492
transform 1 0 12972 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 13340 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 13156 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__33__A
timestamp 1624635492
transform 1 0 13524 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 13892 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__34__A
timestamp 1624635492
transform 1 0 13708 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 14076 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A0
timestamp 1624635492
transform -1 0 14444 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1624635492
transform 1 0 14444 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1624635492
transform -1 0 16008 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output114
timestamp 1624635492
transform 1 0 15456 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1624635492
transform -1 0 15272 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1624635492
transform -1 0 15456 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1624635492
transform 1 0 14628 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_149
timestamp 1624635492
transform 1 0 14812 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l4_in_0_
timestamp 1624635492
transform 1 0 2944 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 2392 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 2668 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 2116 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1624635492
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1624635492
transform -1 0 2024 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output100
timestamp 1624635492
transform -1 0 1748 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_10
timestamp 1624635492
transform 1 0 2024 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1624635492
transform -1 0 4508 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _39_
timestamp 1624635492
transform 1 0 3956 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_0_
timestamp 1624635492
transform -1 0 5336 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1624635492
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_30
timestamp 1624635492
transform 1 0 3864 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 6808 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 8280 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _16_
timestamp 1624635492
transform -1 0 8556 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1624635492
transform -1 0 8832 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_3_
timestamp 1624635492
transform 1 0 9108 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_3_
timestamp 1624635492
transform 1 0 9936 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1624635492
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1624635492
transform -1 0 9016 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  clk_3_N_FTB01
timestamp 1624635492
transform -1 0 11960 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_2_
timestamp 1624635492
transform -1 0 11592 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  prog_clk_2_N_FTB01
timestamp 1624635492
transform -1 0 12328 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  prog_clk_3_N_FTB01
timestamp 1624635492
transform -1 0 12696 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__35__A
timestamp 1624635492
transform 1 0 13432 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 13248 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 13064 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 12880 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__A1
timestamp 1624635492
transform -1 0 12880 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_142
timestamp 1624635492
transform 1 0 14168 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1624635492
transform 1 0 13984 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 13800 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1624635492
transform 1 0 13616 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1624635492
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_144 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 14352 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1624635492
transform -1 0 16008 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_156
timestamp 1624635492
transform 1 0 15456 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l1_in_0_
timestamp 1624635492
transform -1 0 3404 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l4_in_0_
timestamp 1624635492
transform -1 0 2576 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1624635492
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output101
timestamp 1624635492
transform -1 0 1748 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 6348 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 4876 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 6440 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1624635492
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 9384 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_1_
timestamp 1624635492
transform 1 0 9384 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_2_
timestamp 1624635492
transform 1 0 10212 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clk_2_N_FTB01
timestamp 1624635492
transform -1 0 11408 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_3_
timestamp 1624635492
transform 1 0 11684 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1624635492
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 11408 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 12512 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 12696 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 12880 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 13064 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 13248 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 13432 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1624635492
transform 1 0 13616 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_138
timestamp 1624635492
transform 1 0 13800 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1624635492
transform -1 0 16008 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_150 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 14904 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_158
timestamp 1624635492
transform 1 0 15640 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7
timestamp 1624635492
transform 1 0 1748 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 1564 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1624635492
transform -1 0 1748 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output102
timestamp 1624635492
transform -1 0 1748 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1624635492
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1624635492
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 1840 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_0_
timestamp 1624635492
transform -1 0 2576 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_0_
timestamp 1624635492
transform 1 0 2576 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_0_
timestamp 1624635492
transform -1 0 2944 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_0_
timestamp 1624635492
transform -1 0 3772 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1624635492
transform -1 0 4416 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 6348 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 4876 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l1_in_0_
timestamp 1624635492
transform -1 0 5244 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1624635492
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_right_ipin_0.prog_clk
timestamp 1624635492
transform -1 0 4140 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 5244 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 8188 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 6440 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1624635492
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 9384 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_0_
timestamp 1624635492
transform 1 0 8188 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 9108 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 10856 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_0_
timestamp 1624635492
transform 1 0 10580 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1624635492
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1624635492
transform -1 0 11132 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1624635492
transform -1 0 11408 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_2_
timestamp 1624635492
transform 1 0 11408 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_3_
timestamp 1624635492
transform 1 0 12236 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_1_
timestamp 1624635492
transform 1 0 11684 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l1_in_0_
timestamp 1624635492
transform 1 0 12512 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1624635492
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1624635492
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 13432 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0__A0
timestamp 1624635492
transform 1 0 13248 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 13064 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_3_
timestamp 1624635492
transform 1 0 13340 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_6_142
timestamp 1624635492
transform 1 0 14168 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 14352 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 13984 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 13800 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 13616 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 14168 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1624635492
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_144
timestamp 1624635492
transform 1 0 14352 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1624635492
transform -1 0 16008 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1624635492
transform -1 0 16008 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_156
timestamp 1624635492
transform 1 0 15456 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_146
timestamp 1624635492
transform 1 0 14536 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_158
timestamp 1624635492
transform 1 0 15640 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_0_
timestamp 1624635492
transform 1 0 2944 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_0_
timestamp 1624635492
transform -1 0 2944 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 1840 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1624635492
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0__A0
timestamp 1624635492
transform -1 0 1840 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0__A0
timestamp 1624635492
transform -1 0 1656 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3
timestamp 1624635492
transform 1 0 1380 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_0_
timestamp 1624635492
transform 1 0 4324 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1624635492
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_right_ipin_0.prog_clk
timestamp 1624635492
transform 1 0 4048 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 3864 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 6624 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 8096 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_2_
timestamp 1624635492
transform 1 0 8096 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_1_
timestamp 1624635492
transform 1 0 10212 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 10212 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1624635492
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_85
timestamp 1624635492
transform 1 0 8924 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_2_
timestamp 1624635492
transform 1 0 11040 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_1_
timestamp 1624635492
transform 1 0 11868 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_1_
timestamp 1624635492
transform 1 0 12696 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1624635492
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__A0
timestamp 1624635492
transform -1 0 13708 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 13708 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__A0
timestamp 1624635492
transform -1 0 14076 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 14076 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 14352 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1624635492
transform -1 0 16008 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 14536 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__A1
timestamp 1624635492
transform -1 0 14904 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_150
timestamp 1624635492
transform 1 0 14904 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_158
timestamp 1624635492
transform 1 0 15640 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_0_
timestamp 1624635492
transform -1 0 3404 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_1_
timestamp 1624635492
transform -1 0 2576 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1624635492
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output103
timestamp 1624635492
transform -1 0 1748 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 4876 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 3404 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 7912 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1624635492
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 7912 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 9384 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l1_in_0_
timestamp 1624635492
transform 1 0 11684 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_3_
timestamp 1624635492
transform 1 0 12512 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1624635492
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_right_ipin_0.prog_clk
timestamp 1624635492
transform -1 0 11132 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_right_ipin_0.prog_clk
timestamp 1624635492
transform -1 0 11408 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 11408 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_2_
timestamp 1624635492
transform 1 0 13340 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_2__A1
timestamp 1624635492
transform -1 0 14352 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 14352 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1624635492
transform -1 0 16008 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_2__A0
timestamp 1624635492
transform -1 0 14720 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_148
timestamp 1624635492
transform 1 0 14720 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_156
timestamp 1624635492
transform 1 0 15456 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_0_
timestamp 1624635492
transform -1 0 3772 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_0_
timestamp 1624635492
transform -1 0 2944 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 1840 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1624635492
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0__A0
timestamp 1624635492
transform -1 0 1840 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 1472 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3
timestamp 1624635492
transform 1 0 1380 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 4600 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 3864 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1624635492
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_right_ipin_0.prog_clk
timestamp 1624635492
transform -1 0 4600 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 4140 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 7544 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 9016 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 10580 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_2_
timestamp 1624635492
transform 1 0 10580 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1624635492
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_2_
timestamp 1624635492
transform 1 0 11408 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_1_
timestamp 1624635492
transform 1 0 12236 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_3_
timestamp 1624635492
transform 1 0 13064 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1624635492
transform 1 0 14260 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 13892 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 14076 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 14352 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1624635492
transform -1 0 16008 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_2__A1
timestamp 1624635492
transform -1 0 14720 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 14720 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1__A0
timestamp 1624635492
transform -1 0 15088 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__A1
timestamp 1624635492
transform -1 0 15272 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_154 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 15272 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_158
timestamp 1624635492
transform 1 0 15640 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_0_
timestamp 1624635492
transform 1 0 2576 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l4_in_0_
timestamp 1624635492
transform 1 0 1748 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1624635492
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output104
timestamp 1624635492
transform -1 0 1748 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 4876 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 3404 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1624635492
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_right_ipin_0.prog_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 8372 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_11_58
timestamp 1624635492
transform 1 0 6440 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 9844 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 11316 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_0_
timestamp 1624635492
transform 1 0 11684 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_2_
timestamp 1624635492
transform 1 0 12512 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1624635492
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 11316 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_113
timestamp 1624635492
transform 1 0 11500 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_1_
timestamp 1624635492
transform 1 0 13340 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_2_
timestamp 1624635492
transform -1 0 14996 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1624635492
transform -1 0 16008 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__A1
timestamp 1624635492
transform -1 0 15180 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 15180 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_155
timestamp 1624635492
transform 1 0 15364 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_1_
timestamp 1624635492
transform 1 0 2944 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_0_
timestamp 1624635492
transform -1 0 2944 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 1840 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1624635492
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_right_ipin_0.prog_clk
timestamp 1624635492
transform -1 0 1840 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 1564 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 5428 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1624635492
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_30
timestamp 1624635492
transform 1 0 3864 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 5428 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1624635492
transform -1 0 8648 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1624635492
transform -1 0 8924 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 8372 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 9108 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_0_
timestamp 1624635492
transform -1 0 11408 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1624635492
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_85
timestamp 1624635492
transform 1 0 8924 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_2_
timestamp 1624635492
transform -1 0 12236 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_1_
timestamp 1624635492
transform 1 0 12236 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_0_
timestamp 1624635492
transform 1 0 13064 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_1_
timestamp 1624635492
transform 1 0 14352 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1624635492
transform 1 0 14260 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 14076 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_1__A1
timestamp 1624635492
transform -1 0 14260 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1624635492
transform -1 0 16008 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 15364 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 15548 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_157 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 15548 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_3
timestamp 1624635492
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1624635492
transform -1 0 1840 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output105
timestamp 1624635492
transform -1 0 1748 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1624635492
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1624635492
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 1840 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l4_in_0_
timestamp 1624635492
transform -1 0 2576 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_0_
timestamp 1624635492
transform 1 0 2116 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_0_
timestamp 1624635492
transform 1 0 2576 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_1_
timestamp 1624635492
transform 1 0 2944 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 4876 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 3404 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_0_
timestamp 1624635492
transform 1 0 4324 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1624635492
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_right_ipin_0.prog_clk
timestamp 1624635492
transform -1 0 4324 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_0__A0
timestamp 1624635492
transform 1 0 3864 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 5152 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 6624 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l1_in_0_
timestamp 1624635492
transform 1 0 6440 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1624635492
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1624635492
transform -1 0 7544 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 7728 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_1_
timestamp 1624635492
transform 1 0 8096 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 7544 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 9384 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_0_
timestamp 1624635492
transform 1 0 9108 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_3_
timestamp 1624635492
transform -1 0 10764 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1624635492
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 9200 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_85
timestamp 1624635492
transform 1 0 8924 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1624635492
transform -1 0 11132 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_1_
timestamp 1624635492
transform 1 0 10764 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_1_
timestamp 1624635492
transform 1 0 11592 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_1_
timestamp 1624635492
transform 1 0 12420 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_0_
timestamp 1624635492
transform 1 0 11684 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_2_
timestamp 1624635492
transform -1 0 13340 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1624635492
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_right_ipin_0.prog_clk
timestamp 1624635492
transform 1 0 11132 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 11408 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_3_
timestamp 1624635492
transform 1 0 13248 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_1_
timestamp 1624635492
transform 1 0 13340 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_3_
timestamp 1624635492
transform -1 0 14996 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_0_
timestamp 1624635492
transform 1 0 14352 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1624635492
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_0__A0
timestamp 1624635492
transform 1 0 14076 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  Test_en_E_FTB01
timestamp 1624635492
transform -1 0 15272 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1624635492
transform -1 0 16008 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1624635492
transform -1 0 16008 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output49
timestamp 1624635492
transform 1 0 15364 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Test_en_E_FTB01_A
timestamp 1624635492
transform -1 0 15456 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__A1
timestamp 1624635492
transform -1 0 15640 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__A1
timestamp 1624635492
transform -1 0 15364 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_158
timestamp 1624635492
transform 1 0 15640 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_1_
timestamp 1624635492
transform -1 0 3404 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_0_
timestamp 1624635492
transform -1 0 2576 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1624635492
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output106
timestamp 1624635492
transform -1 0 1748 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 4876 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 3404 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 6440 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1624635492
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 7912 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_2_
timestamp 1624635492
transform 1 0 9384 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_1_
timestamp 1624635492
transform 1 0 10212 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_2_
timestamp 1624635492
transform -1 0 12512 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_1_
timestamp 1624635492
transform 1 0 12512 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1624635492
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 11040 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 11408 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 11224 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l1_in_0_
timestamp 1624635492
transform -1 0 14168 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_2_
timestamp 1624635492
transform 1 0 14168 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1624635492
transform -1 0 16008 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__A0
timestamp 1624635492
transform -1 0 15180 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_153 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 15180 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l4_in_0_
timestamp 1624635492
transform 1 0 2944 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 1840 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l4_in_0_
timestamp 1624635492
transform 1 0 2116 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1624635492
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output107
timestamp 1624635492
transform -1 0 1748 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_7
timestamp 1624635492
transform 1 0 1748 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 5428 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1624635492
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_30
timestamp 1624635492
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 6900 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1624635492
transform -1 0 8648 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1624635492
transform -1 0 8924 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 8372 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_3_
timestamp 1624635492
transform 1 0 9108 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_0_
timestamp 1624635492
transform 1 0 9936 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1624635492
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_85
timestamp 1624635492
transform 1 0 8924 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_2_
timestamp 1624635492
transform 1 0 10764 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_0_
timestamp 1624635492
transform -1 0 12420 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_1_
timestamp 1624635492
transform 1 0 12420 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_3_
timestamp 1624635492
transform 1 0 14352 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1624635492
transform 1 0 14260 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 13248 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 13432 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 13616 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 13800 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 13984 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_142
timestamp 1624635492
transform 1 0 14168 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1624635492
transform -1 0 16008 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 15180 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_155
timestamp 1624635492
transform 1 0 15364 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_0_
timestamp 1624635492
transform 1 0 2392 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_0_
timestamp 1624635492
transform -1 0 2392 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1624635492
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1624635492
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 4876 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_0_
timestamp 1624635492
transform 1 0 4048 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_0_
timestamp 1624635492
transform -1 0 4048 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 6440 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1624635492
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 9384 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_1_
timestamp 1624635492
transform 1 0 9384 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_2_
timestamp 1624635492
transform 1 0 10212 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l4_in_0_
timestamp 1624635492
transform 1 0 11684 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1624635492
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_right_ipin_0.prog_clk
timestamp 1624635492
transform -1 0 11316 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 11316 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 12512 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_113
timestamp 1624635492
transform 1 0 11500 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 12696 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 12880 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 13064 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_134
timestamp 1624635492
transform 1 0 13432 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1624635492
transform -1 0 16008 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_146
timestamp 1624635492
transform 1 0 14536 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_158
timestamp 1624635492
transform 1 0 15640 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 1840 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_0_
timestamp 1624635492
transform -1 0 3772 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_1_
timestamp 1624635492
transform -1 0 2944 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1624635492
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output108
timestamp 1624635492
transform -1 0 1748 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_7
timestamp 1624635492
transform 1 0 1748 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1624635492
transform -1 0 4600 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 4600 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1624635492
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_right_ipin_0.prog_clk
timestamp 1624635492
transform 1 0 4048 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_30
timestamp 1624635492
transform 1 0 3864 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 7544 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 9016 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 9108 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_3_
timestamp 1624635492
transform 1 0 10580 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1624635492
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_2_
timestamp 1624635492
transform 1 0 11408 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_3_
timestamp 1624635492
transform 1 0 12236 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1624635492
transform 1 0 14260 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 13064 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_132
timestamp 1624635492
transform 1 0 13248 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_140
timestamp 1624635492
transform 1 0 13984 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_144
timestamp 1624635492
transform 1 0 14352 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1624635492
transform -1 0 16008 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_156
timestamp 1624635492
transform 1 0 15456 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_7
timestamp 1624635492
transform 1 0 1748 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1624635492
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output109
timestamp 1624635492
transform -1 0 1748 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1624635492
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1624635492
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l4_in_0_
timestamp 1624635492
transform -1 0 2576 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_19
timestamp 1624635492
transform 1 0 2852 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_15
timestamp 1624635492
transform 1 0 2484 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 2576 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l4_in_0_
timestamp 1624635492
transform 1 0 2576 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_1_
timestamp 1624635492
transform 1 0 2944 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 4876 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 4876 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l4_in_0_
timestamp 1624635492
transform 1 0 4600 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 3864 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1624635492
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_right_ipin_0.prog_clk
timestamp 1624635492
transform -1 0 4600 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_33
timestamp 1624635492
transform 1 0 4140 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 6440 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 6900 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1624635492
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1624635492
transform -1 0 8648 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1624635492
transform -1 0 8924 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 6900 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 7912 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_2_
timestamp 1624635492
transform 1 0 9384 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_1_
timestamp 1624635492
transform 1 0 9108 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_2_
timestamp 1624635492
transform 1 0 10212 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_1_
timestamp 1624635492
transform 1 0 9936 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1624635492
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_85
timestamp 1624635492
transform 1 0 8924 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 11224 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 11224 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 11040 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 11040 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_right_ipin_0.prog_clk
timestamp 1624635492
transform 1 0 10764 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1624635492
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 11868 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 11684 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_124
timestamp 1624635492
transform 1 0 12512 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_112
timestamp 1624635492
transform 1 0 11408 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_119
timestamp 1624635492
transform 1 0 12052 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1624635492
transform 1 0 14260 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_131
timestamp 1624635492
transform 1 0 13156 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_143
timestamp 1624635492
transform 1 0 14260 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_136
timestamp 1624635492
transform 1 0 13616 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_142
timestamp 1624635492
transform 1 0 14168 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_144
timestamp 1624635492
transform 1 0 14352 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1624635492
transform -1 0 16008 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1624635492
transform -1 0 16008 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_155
timestamp 1624635492
transform 1 0 15364 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_156
timestamp 1624635492
transform 1 0 15456 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 2484 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 2760 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1624635492
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1624635492
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 4876 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l4_in_0_
timestamp 1624635492
transform 1 0 4048 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_21_21
timestamp 1624635492
transform 1 0 3036 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_29
timestamp 1624635492
transform 1 0 3772 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 7912 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1624635492
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_0_
timestamp 1624635492
transform 1 0 7912 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_0_
timestamp 1624635492
transform 1 0 8740 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_3_
timestamp 1624635492
transform 1 0 9568 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_0__A0
timestamp 1624635492
transform 1 0 10396 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 10580 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1624635492
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_105
timestamp 1624635492
transform 1 0 10764 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_113
timestamp 1624635492
transform 1 0 11500 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_115
timestamp 1624635492
transform 1 0 11684 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_127
timestamp 1624635492
transform 1 0 12788 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_139
timestamp 1624635492
transform 1 0 13892 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1624635492
transform -1 0 16008 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_151
timestamp 1624635492
transform 1 0 14996 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1624635492
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output110
timestamp 1624635492
transform -1 0 1748 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_7
timestamp 1624635492
transform 1 0 1748 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_19
timestamp 1624635492
transform 1 0 2852 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_1_
timestamp 1624635492
transform -1 0 5060 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1624635492
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1624635492
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_30
timestamp 1624635492
transform 1 0 3864 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 7360 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_0_
timestamp 1624635492
transform 1 0 5060 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_1_
timestamp 1624635492
transform 1 0 7360 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l1_in_0_
timestamp 1624635492
transform -1 0 9016 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1624635492
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 9108 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 9292 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 9476 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 9660 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 9844 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 10028 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_99
timestamp 1624635492
transform 1 0 10212 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_111
timestamp 1624635492
transform 1 0 11316 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_123
timestamp 1624635492
transform 1 0 12420 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1624635492
transform 1 0 14260 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_135
timestamp 1624635492
transform 1 0 13524 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_144
timestamp 1624635492
transform 1 0 14352 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1624635492
transform -1 0 16008 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_156
timestamp 1624635492
transform 1 0 15456 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1624635492
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1624635492
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1624635492
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l4_in_0_
timestamp 1624635492
transform 1 0 4692 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1624635492
transform 1 0 4416 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_27
timestamp 1624635492
transform 1 0 3588 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_35
timestamp 1624635492
transform 1 0 4324 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_38
timestamp 1624635492
transform 1 0 4600 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_0_
timestamp 1624635492
transform 1 0 6440 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_0_
timestamp 1624635492
transform 1 0 5520 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1624635492
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_1_
timestamp 1624635492
transform 1 0 7268 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_2_
timestamp 1624635492
transform 1 0 8096 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _65_
timestamp 1624635492
transform 1 0 8924 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 9200 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_2__A1
timestamp 1624635492
transform 1 0 9384 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_92
timestamp 1624635492
transform 1 0 9568 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_104
timestamp 1624635492
transform 1 0 10672 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1624635492
transform 1 0 11592 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_112
timestamp 1624635492
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_115
timestamp 1624635492
transform 1 0 11684 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_127
timestamp 1624635492
transform 1 0 12788 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_139
timestamp 1624635492
transform 1 0 13892 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1624635492
transform -1 0 16008 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_151
timestamp 1624635492
transform 1 0 14996 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1624635492
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output111
timestamp 1624635492
transform -1 0 1748 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_N_FTB01_A
timestamp 1624635492
transform 1 0 1748 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_9
timestamp 1624635492
transform 1 0 1932 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _52_
timestamp 1624635492
transform 1 0 3864 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _53_
timestamp 1624635492
transform 1 0 4140 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _54_
timestamp 1624635492
transform 1 0 4416 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _55_
timestamp 1624635492
transform 1 0 4692 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1624635492
transform 1 0 3772 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_21
timestamp 1624635492
transform 1 0 3036 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _57_
timestamp 1624635492
transform 1 0 5244 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _58_
timestamp 1624635492
transform 1 0 5520 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l1_in_0_
timestamp 1624635492
transform 1 0 6348 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1624635492
transform 1 0 4968 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_0__A0
timestamp 1624635492
transform 1 0 6164 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1624635492
transform 1 0 5796 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1624635492
transform 1 0 5980 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_44
timestamp 1624635492
transform 1 0 5152 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _63_
timestamp 1624635492
transform 1 0 8004 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _64_
timestamp 1624635492
transform 1 0 8280 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _66_
timestamp 1624635492
transform 1 0 8556 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_1_
timestamp 1624635492
transform 1 0 7176 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _67_
timestamp 1624635492
transform 1 0 9108 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _69_
timestamp 1624635492
transform 1 0 9384 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _70_
timestamp 1624635492
transform 1 0 9660 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _71_
timestamp 1624635492
transform 1 0 9936 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1624635492
transform 1 0 9016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1624635492
transform 1 0 10212 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_101
timestamp 1624635492
transform 1 0 10396 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_113
timestamp 1624635492
transform 1 0 11500 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_125
timestamp 1624635492
transform 1 0 12604 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1624635492
transform 1 0 14260 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_137
timestamp 1624635492
transform 1 0 13708 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_24_144
timestamp 1624635492
transform 1 0 14352 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1624635492
transform -1 0 16008 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1624635492
transform -1 0 15640 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1624635492
transform -1 0 15272 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1624635492
transform -1 0 15456 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1624635492
transform -1 0 15088 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_158
timestamp 1624635492
transform 1 0 15640 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1624635492
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1624635492
transform -1 0 2024 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output112
timestamp 1624635492
transform -1 0 1748 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  output113
timestamp 1624635492
transform -1 0 2300 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1624635492
transform -1 0 2484 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output93_A
timestamp 1624635492
transform 1 0 2484 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output95_A
timestamp 1624635492
transform 1 0 2668 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_19
timestamp 1624635492
transform 1 0 2852 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A
timestamp 1624635492
transform -1 0 4876 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_31
timestamp 1624635492
transform 1 0 3956 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_41
timestamp 1624635492
transform 1 0 4876 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _56_
timestamp 1624635492
transform 1 0 5152 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _59_
timestamp 1624635492
transform 1 0 6440 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _60_
timestamp 1624635492
transform 1 0 6716 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1624635492
transform 1 0 6348 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1624635492
transform -1 0 5612 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_49
timestamp 1624635492
transform 1 0 5612 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _61_
timestamp 1624635492
transform 1 0 6992 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _62_
timestamp 1624635492
transform 1 0 7268 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _68_
timestamp 1624635492
transform -1 0 8924 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 7728 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1624635492
transform -1 0 7912 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1624635492
transform -1 0 8096 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 8096 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 8280 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_80
timestamp 1624635492
transform 1 0 8464 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_85
timestamp 1624635492
transform 1 0 8924 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_97
timestamp 1624635492
transform 1 0 10028 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1624635492
transform 1 0 11592 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_109
timestamp 1624635492
transform 1 0 11132 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_113
timestamp 1624635492
transform 1 0 11500 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_115
timestamp 1624635492
transform 1 0 11684 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1624635492
transform -1 0 14628 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1624635492
transform -1 0 13984 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1624635492
transform -1 0 13800 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_127
timestamp 1624635492
transform 1 0 12788 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_135
timestamp 1624635492
transform 1 0 13524 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_140
timestamp 1624635492
transform 1 0 13984 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_144
timestamp 1624635492
transform 1 0 14352 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1624635492
transform -1 0 16008 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1624635492
transform -1 0 15732 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1624635492
transform -1 0 15364 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1624635492
transform -1 0 14996 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1624635492
transform -1 0 14812 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output93
timestamp 1624635492
transform -1 0 1748 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1624635492
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1624635492
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_N_FTB01
timestamp 1624635492
transform 1 0 1380 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_9
timestamp 1624635492
transform 1 0 1932 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output115
timestamp 1624635492
transform -1 0 2484 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output95
timestamp 1624635492
transform -1 0 2116 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output50
timestamp 1624635492
transform -1 0 2392 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output117
timestamp 1624635492
transform -1 0 2852 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output73
timestamp 1624635492
transform -1 0 3128 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output51
timestamp 1624635492
transform -1 0 2760 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Test_en_N_FTB01
timestamp 1624635492
transform 1 0 2852 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_28
timestamp 1624635492
transform 1 0 3680 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output117_A
timestamp 1624635492
transform 1 0 3496 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output115_A
timestamp 1624635492
transform 1 0 3312 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Test_en_N_FTB01_A
timestamp 1624635492
transform 1 0 3128 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output84
timestamp 1624635492
transform -1 0 3496 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1624635492
transform 1 0 3772 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1624635492
transform 1 0 3772 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  Test_en_W_FTB01
timestamp 1624635492
transform 1 0 3496 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_32
timestamp 1624635492
transform 1 0 4048 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Test_en_W_FTB01_A
timestamp 1624635492
transform 1 0 3864 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output87
timestamp 1624635492
transform -1 0 4968 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output86
timestamp 1624635492
transform -1 0 4600 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output85
timestamp 1624635492
transform -1 0 4232 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_40
timestamp 1624635492
transform 1 0 4784 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output91
timestamp 1624635492
transform -1 0 5704 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output90
timestamp 1624635492
transform -1 0 5336 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output89
timestamp 1624635492
transform -1 0 5704 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output88
timestamp 1624635492
transform -1 0 5336 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_54
timestamp 1624635492
transform 1 0 6072 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output92
timestamp 1624635492
transform -1 0 6072 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output83
timestamp 1624635492
transform 1 0 5704 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output82
timestamp 1624635492
transform 1 0 6072 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_60
timestamp 1624635492
transform 1 0 6624 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1624635492
transform -1 0 6900 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output74
timestamp 1624635492
transform -1 0 6900 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1624635492
transform 1 0 6440 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_63
timestamp 1624635492
transform 1 0 6900 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1624635492
transform -1 0 7176 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output77
timestamp 1624635492
transform -1 0 8004 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output76
timestamp 1624635492
transform -1 0 7636 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output75
timestamp 1624635492
transform -1 0 7268 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_78
timestamp 1624635492
transform 1 0 8280 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output80
timestamp 1624635492
transform -1 0 9108 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output79
timestamp 1624635492
transform -1 0 8740 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output78
timestamp 1624635492
transform -1 0 8372 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_66
timestamp 1624635492
transform 1 0 7176 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_92
timestamp 1624635492
transform 1 0 9568 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output81
timestamp 1624635492
transform -1 0 9568 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1624635492
transform 1 0 9108 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1624635492
transform 1 0 9016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_101
timestamp 1624635492
transform 1 0 10396 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1624635492
transform -1 0 10764 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1624635492
transform -1 0 10396 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  input37
timestamp 1624635492
transform -1 0 10948 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input36
timestamp 1624635492
transform -1 0 10580 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input25
timestamp 1624635492
transform -1 0 10212 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_87
timestamp 1624635492
transform 1 0 9108 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_109
timestamp 1624635492
transform 1 0 11132 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_105
timestamp 1624635492
transform 1 0 10764 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1624635492
transform -1 0 11132 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  input38
timestamp 1624635492
transform -1 0 11316 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_113
timestamp 1624635492
transform 1 0 11500 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1624635492
transform -1 0 11500 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1624635492
transform -1 0 11684 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_115
timestamp 1624635492
transform 1 0 11684 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_117
timestamp 1624635492
transform 1 0 11868 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1624635492
transform -1 0 11868 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1624635492
transform 1 0 11868 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1624635492
transform 1 0 11776 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_123
timestamp 1624635492
transform 1 0 12420 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1624635492
transform -1 0 12420 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1624635492
transform -1 0 12512 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1624635492
transform -1 0 12880 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1624635492
transform -1 0 12880 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1624635492
transform -1 0 13248 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1624635492
transform -1 0 13064 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1624635492
transform -1 0 13616 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1624635492
transform -1 0 14168 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1624635492
transform -1 0 14076 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1624635492
transform -1 0 13800 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_138
timestamp 1624635492
transform 1 0 13800 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1624635492
transform 1 0 14260 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1624635492
transform 1 0 14444 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1624635492
transform -1 0 14720 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1624635492
transform -1 0 14352 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1624635492
transform -1 0 14260 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_144
timestamp 1624635492
transform 1 0 14352 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input43 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 13800 0 1 16864
box -38 -48 958 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1624635492
transform -1 0 16008 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1624635492
transform -1 0 16008 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1624635492
transform -1 0 15732 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1624635492
transform 1 0 14536 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1624635492
transform -1 0 15272 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1624635492
transform -1 0 15640 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1624635492
transform -1 0 15456 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1624635492
transform -1 0 15088 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_158
timestamp 1624635492
transform 1 0 15640 0 1 16864
box -38 -48 130 592
<< labels >>
rlabel metal3 s 16400 16600 17200 16720 6 Test_en_E_in
port 0 nsew signal input
rlabel metal3 s 16400 9936 17200 10056 6 Test_en_E_out
port 1 nsew signal tristate
rlabel metal2 s 2042 19200 2098 20000 6 Test_en_N_out
port 2 nsew signal tristate
rlabel metal2 s 13818 0 13874 800 6 Test_en_S_in
port 3 nsew signal input
rlabel metal3 s 0 17280 800 17400 6 Test_en_W_in
port 4 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 Test_en_W_out
port 5 nsew signal tristate
rlabel metal3 s 0 416 800 536 6 ccff_head
port 6 nsew signal input
rlabel metal3 s 16400 3272 17200 3392 6 ccff_tail
port 7 nsew signal tristate
rlabel metal2 s 6918 0 6974 800 6 chany_bottom_in[0]
port 8 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 chany_bottom_in[10]
port 9 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 chany_bottom_in[11]
port 10 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 chany_bottom_in[12]
port 11 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 chany_bottom_in[13]
port 12 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 chany_bottom_in[14]
port 13 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 chany_bottom_in[15]
port 14 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 chany_bottom_in[16]
port 15 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 chany_bottom_in[17]
port 16 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 chany_bottom_in[18]
port 17 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 chany_bottom_in[19]
port 18 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 chany_bottom_in[1]
port 19 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 chany_bottom_in[2]
port 20 nsew signal input
rlabel metal2 s 8022 0 8078 800 6 chany_bottom_in[3]
port 21 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 chany_bottom_in[4]
port 22 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 chany_bottom_in[5]
port 23 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 chany_bottom_in[6]
port 24 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 chany_bottom_in[7]
port 25 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 chany_bottom_in[8]
port 26 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 chany_bottom_in[9]
port 27 nsew signal input
rlabel metal2 s 110 0 166 800 6 chany_bottom_out[0]
port 28 nsew signal tristate
rlabel metal2 s 3514 0 3570 800 6 chany_bottom_out[10]
port 29 nsew signal tristate
rlabel metal2 s 3882 0 3938 800 6 chany_bottom_out[11]
port 30 nsew signal tristate
rlabel metal2 s 4158 0 4214 800 6 chany_bottom_out[12]
port 31 nsew signal tristate
rlabel metal2 s 4526 0 4582 800 6 chany_bottom_out[13]
port 32 nsew signal tristate
rlabel metal2 s 4894 0 4950 800 6 chany_bottom_out[14]
port 33 nsew signal tristate
rlabel metal2 s 5262 0 5318 800 6 chany_bottom_out[15]
port 34 nsew signal tristate
rlabel metal2 s 5538 0 5594 800 6 chany_bottom_out[16]
port 35 nsew signal tristate
rlabel metal2 s 5906 0 5962 800 6 chany_bottom_out[17]
port 36 nsew signal tristate
rlabel metal2 s 6274 0 6330 800 6 chany_bottom_out[18]
port 37 nsew signal tristate
rlabel metal2 s 6642 0 6698 800 6 chany_bottom_out[19]
port 38 nsew signal tristate
rlabel metal2 s 386 0 442 800 6 chany_bottom_out[1]
port 39 nsew signal tristate
rlabel metal2 s 754 0 810 800 6 chany_bottom_out[2]
port 40 nsew signal tristate
rlabel metal2 s 1122 0 1178 800 6 chany_bottom_out[3]
port 41 nsew signal tristate
rlabel metal2 s 1398 0 1454 800 6 chany_bottom_out[4]
port 42 nsew signal tristate
rlabel metal2 s 1766 0 1822 800 6 chany_bottom_out[5]
port 43 nsew signal tristate
rlabel metal2 s 2134 0 2190 800 6 chany_bottom_out[6]
port 44 nsew signal tristate
rlabel metal2 s 2502 0 2558 800 6 chany_bottom_out[7]
port 45 nsew signal tristate
rlabel metal2 s 2778 0 2834 800 6 chany_bottom_out[8]
port 46 nsew signal tristate
rlabel metal2 s 3146 0 3202 800 6 chany_bottom_out[9]
port 47 nsew signal tristate
rlabel metal2 s 9862 19200 9918 20000 6 chany_top_in[0]
port 48 nsew signal input
rlabel metal2 s 13634 19200 13690 20000 6 chany_top_in[10]
port 49 nsew signal input
rlabel metal2 s 14002 19200 14058 20000 6 chany_top_in[11]
port 50 nsew signal input
rlabel metal2 s 14370 19200 14426 20000 6 chany_top_in[12]
port 51 nsew signal input
rlabel metal2 s 14738 19200 14794 20000 6 chany_top_in[13]
port 52 nsew signal input
rlabel metal2 s 15106 19200 15162 20000 6 chany_top_in[14]
port 53 nsew signal input
rlabel metal2 s 15474 19200 15530 20000 6 chany_top_in[15]
port 54 nsew signal input
rlabel metal2 s 15842 19200 15898 20000 6 chany_top_in[16]
port 55 nsew signal input
rlabel metal2 s 16210 19200 16266 20000 6 chany_top_in[17]
port 56 nsew signal input
rlabel metal2 s 16578 19200 16634 20000 6 chany_top_in[18]
port 57 nsew signal input
rlabel metal2 s 16946 19200 17002 20000 6 chany_top_in[19]
port 58 nsew signal input
rlabel metal2 s 10230 19200 10286 20000 6 chany_top_in[1]
port 59 nsew signal input
rlabel metal2 s 10598 19200 10654 20000 6 chany_top_in[2]
port 60 nsew signal input
rlabel metal2 s 10966 19200 11022 20000 6 chany_top_in[3]
port 61 nsew signal input
rlabel metal2 s 11334 19200 11390 20000 6 chany_top_in[4]
port 62 nsew signal input
rlabel metal2 s 11794 19200 11850 20000 6 chany_top_in[5]
port 63 nsew signal input
rlabel metal2 s 12162 19200 12218 20000 6 chany_top_in[6]
port 64 nsew signal input
rlabel metal2 s 12530 19200 12586 20000 6 chany_top_in[7]
port 65 nsew signal input
rlabel metal2 s 12898 19200 12954 20000 6 chany_top_in[8]
port 66 nsew signal input
rlabel metal2 s 13266 19200 13322 20000 6 chany_top_in[9]
port 67 nsew signal input
rlabel metal2 s 2410 19200 2466 20000 6 chany_top_out[0]
port 68 nsew signal tristate
rlabel metal2 s 6182 19200 6238 20000 6 chany_top_out[10]
port 69 nsew signal tristate
rlabel metal2 s 6550 19200 6606 20000 6 chany_top_out[11]
port 70 nsew signal tristate
rlabel metal2 s 6918 19200 6974 20000 6 chany_top_out[12]
port 71 nsew signal tristate
rlabel metal2 s 7286 19200 7342 20000 6 chany_top_out[13]
port 72 nsew signal tristate
rlabel metal2 s 7654 19200 7710 20000 6 chany_top_out[14]
port 73 nsew signal tristate
rlabel metal2 s 8022 19200 8078 20000 6 chany_top_out[15]
port 74 nsew signal tristate
rlabel metal2 s 8390 19200 8446 20000 6 chany_top_out[16]
port 75 nsew signal tristate
rlabel metal2 s 8758 19200 8814 20000 6 chany_top_out[17]
port 76 nsew signal tristate
rlabel metal2 s 9126 19200 9182 20000 6 chany_top_out[18]
port 77 nsew signal tristate
rlabel metal2 s 9494 19200 9550 20000 6 chany_top_out[19]
port 78 nsew signal tristate
rlabel metal2 s 2778 19200 2834 20000 6 chany_top_out[1]
port 79 nsew signal tristate
rlabel metal2 s 3146 19200 3202 20000 6 chany_top_out[2]
port 80 nsew signal tristate
rlabel metal2 s 3514 19200 3570 20000 6 chany_top_out[3]
port 81 nsew signal tristate
rlabel metal2 s 3882 19200 3938 20000 6 chany_top_out[4]
port 82 nsew signal tristate
rlabel metal2 s 4250 19200 4306 20000 6 chany_top_out[5]
port 83 nsew signal tristate
rlabel metal2 s 4618 19200 4674 20000 6 chany_top_out[6]
port 84 nsew signal tristate
rlabel metal2 s 4986 19200 5042 20000 6 chany_top_out[7]
port 85 nsew signal tristate
rlabel metal2 s 5354 19200 5410 20000 6 chany_top_out[8]
port 86 nsew signal tristate
rlabel metal2 s 5722 19200 5778 20000 6 chany_top_out[9]
port 87 nsew signal tristate
rlabel metal2 s 202 19200 258 20000 6 clk_2_N_out
port 88 nsew signal tristate
rlabel metal2 s 14186 0 14242 800 6 clk_2_S_in
port 89 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 clk_2_S_out
port 90 nsew signal tristate
rlabel metal2 s 570 19200 626 20000 6 clk_3_N_out
port 91 nsew signal tristate
rlabel metal2 s 14554 0 14610 800 6 clk_3_S_in
port 92 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 clk_3_S_out
port 93 nsew signal tristate
rlabel metal3 s 0 1368 800 1488 6 left_grid_pin_16_
port 94 nsew signal tristate
rlabel metal3 s 0 2320 800 2440 6 left_grid_pin_17_
port 95 nsew signal tristate
rlabel metal3 s 0 3408 800 3528 6 left_grid_pin_18_
port 96 nsew signal tristate
rlabel metal3 s 0 4360 800 4480 6 left_grid_pin_19_
port 97 nsew signal tristate
rlabel metal3 s 0 5312 800 5432 6 left_grid_pin_20_
port 98 nsew signal tristate
rlabel metal3 s 0 6400 800 6520 6 left_grid_pin_21_
port 99 nsew signal tristate
rlabel metal3 s 0 7352 800 7472 6 left_grid_pin_22_
port 100 nsew signal tristate
rlabel metal3 s 0 8304 800 8424 6 left_grid_pin_23_
port 101 nsew signal tristate
rlabel metal3 s 0 9392 800 9512 6 left_grid_pin_24_
port 102 nsew signal tristate
rlabel metal3 s 0 10344 800 10464 6 left_grid_pin_25_
port 103 nsew signal tristate
rlabel metal3 s 0 11296 800 11416 6 left_grid_pin_26_
port 104 nsew signal tristate
rlabel metal3 s 0 12384 800 12504 6 left_grid_pin_27_
port 105 nsew signal tristate
rlabel metal3 s 0 13336 800 13456 6 left_grid_pin_28_
port 106 nsew signal tristate
rlabel metal3 s 0 14288 800 14408 6 left_grid_pin_29_
port 107 nsew signal tristate
rlabel metal3 s 0 15376 800 15496 6 left_grid_pin_30_
port 108 nsew signal tristate
rlabel metal3 s 0 16328 800 16448 6 left_grid_pin_31_
port 109 nsew signal tristate
rlabel metal2 s 938 19200 994 20000 6 prog_clk_0_N_out
port 110 nsew signal tristate
rlabel metal2 s 16210 0 16266 800 6 prog_clk_0_S_out
port 111 nsew signal tristate
rlabel metal3 s 0 19320 800 19440 6 prog_clk_0_W_in
port 112 nsew signal input
rlabel metal2 s 1306 19200 1362 20000 6 prog_clk_2_N_out
port 113 nsew signal tristate
rlabel metal2 s 14830 0 14886 800 6 prog_clk_2_S_in
port 114 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 prog_clk_2_S_out
port 115 nsew signal tristate
rlabel metal2 s 1674 19200 1730 20000 6 prog_clk_3_N_out
port 116 nsew signal tristate
rlabel metal2 s 15198 0 15254 800 6 prog_clk_3_S_in
port 117 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 prog_clk_3_S_out
port 118 nsew signal tristate
rlabel metal4 s 13437 2128 13757 17456 6 VPWR
port 119 nsew power bidirectional
rlabel metal4 s 8440 2128 8760 17456 6 VPWR
port 120 nsew power bidirectional
rlabel metal4 s 3443 2128 3763 17456 6 VPWR
port 121 nsew power bidirectional
rlabel metal4 s 10939 2128 11259 17456 6 VGND
port 122 nsew ground bidirectional
rlabel metal4 s 5941 2128 6261 17456 6 VGND
port 123 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 17200 20000
<< end >>
