magic
tech sky130A
magscale 1 2
timestamp 1680088213
<< viali >>
rect 24593 24361 24627 24395
rect 25973 24361 26007 24395
rect 29745 24361 29779 24395
rect 32321 24361 32355 24395
rect 33609 24361 33643 24395
rect 45385 24361 45419 24395
rect 27905 24293 27939 24327
rect 31677 24293 31711 24327
rect 37473 24293 37507 24327
rect 44649 24293 44683 24327
rect 3249 24225 3283 24259
rect 5825 24225 5859 24259
rect 8217 24225 8251 24259
rect 10977 24225 11011 24259
rect 13553 24225 13587 24259
rect 16129 24225 16163 24259
rect 18705 24225 18739 24259
rect 20913 24225 20947 24259
rect 22477 24225 22511 24259
rect 25237 24225 25271 24259
rect 29193 24225 29227 24259
rect 34069 24225 34103 24259
rect 34253 24225 34287 24259
rect 35541 24225 35575 24259
rect 36553 24225 36587 24259
rect 36737 24225 36771 24259
rect 37933 24225 37967 24259
rect 38117 24225 38151 24259
rect 40693 24225 40727 24259
rect 40969 24225 41003 24259
rect 48513 24225 48547 24259
rect 2237 24157 2271 24191
rect 4169 24157 4203 24191
rect 4629 24157 4663 24191
rect 6745 24157 6779 24191
rect 7389 24157 7423 24191
rect 9321 24157 9355 24191
rect 9965 24157 9999 24191
rect 11897 24157 11931 24191
rect 12541 24157 12575 24191
rect 14473 24157 14507 24191
rect 15117 24157 15151 24191
rect 17601 24157 17635 24191
rect 19625 24157 19659 24191
rect 20269 24157 20303 24191
rect 22017 24157 22051 24191
rect 24041 24157 24075 24191
rect 25881 24157 25915 24191
rect 28089 24157 28123 24191
rect 28733 24157 28767 24191
rect 29929 24157 29963 24191
rect 30573 24157 30607 24191
rect 31217 24157 31251 24191
rect 32505 24157 32539 24191
rect 33149 24157 33183 24191
rect 33977 24157 34011 24191
rect 38669 24157 38703 24191
rect 38945 24157 38979 24191
rect 40233 24157 40267 24191
rect 42625 24157 42659 24191
rect 45293 24157 45327 24191
rect 45937 24157 45971 24191
rect 47225 24157 47259 24191
rect 47777 24157 47811 24191
rect 48789 24157 48823 24191
rect 27261 24089 27295 24123
rect 29009 24089 29043 24123
rect 31861 24089 31895 24123
rect 41889 24089 41923 24123
rect 46765 24089 46799 24123
rect 3985 24021 4019 24055
rect 6561 24021 6595 24055
rect 9137 24021 9171 24055
rect 11713 24021 11747 24055
rect 14289 24021 14323 24055
rect 16865 24021 16899 24055
rect 19441 24021 19475 24055
rect 23857 24021 23891 24055
rect 24961 24021 24995 24055
rect 25053 24021 25087 24055
rect 26341 24021 26375 24055
rect 26709 24021 26743 24055
rect 27353 24021 27387 24055
rect 28549 24021 28583 24055
rect 30389 24021 30423 24055
rect 31033 24021 31067 24055
rect 31493 24021 31527 24055
rect 32965 24021 32999 24055
rect 34897 24021 34931 24055
rect 35265 24021 35299 24055
rect 35357 24021 35391 24055
rect 36093 24021 36127 24055
rect 36461 24021 36495 24055
rect 37841 24021 37875 24055
rect 40049 24021 40083 24055
rect 41981 24021 42015 24055
rect 42165 24021 42199 24055
rect 43913 24021 43947 24055
rect 46121 24021 46155 24055
rect 46857 24021 46891 24055
rect 47961 24021 47995 24055
rect 2145 23817 2179 23851
rect 12035 23817 12069 23851
rect 21281 23817 21315 23851
rect 23305 23817 23339 23851
rect 23765 23817 23799 23851
rect 28457 23817 28491 23851
rect 36277 23817 36311 23851
rect 38853 23817 38887 23851
rect 39221 23817 39255 23851
rect 45661 23817 45695 23851
rect 48237 23817 48271 23851
rect 3985 23749 4019 23783
rect 9137 23749 9171 23783
rect 10701 23749 10735 23783
rect 14289 23749 14323 23783
rect 16129 23749 16163 23783
rect 18153 23749 18187 23783
rect 23673 23749 23707 23783
rect 24501 23749 24535 23783
rect 32781 23749 32815 23783
rect 37933 23749 37967 23783
rect 41981 23749 42015 23783
rect 46857 23749 46891 23783
rect 47317 23749 47351 23783
rect 2329 23681 2363 23715
rect 2973 23681 3007 23715
rect 4721 23681 4755 23715
rect 6837 23681 6871 23715
rect 7481 23681 7515 23715
rect 8125 23681 8159 23715
rect 9965 23681 9999 23715
rect 13093 23681 13127 23715
rect 15117 23681 15151 23715
rect 17141 23681 17175 23715
rect 21465 23681 21499 23715
rect 22017 23681 22051 23715
rect 27353 23681 27387 23715
rect 27997 23681 28031 23715
rect 28641 23681 28675 23715
rect 29285 23681 29319 23715
rect 29561 23681 29595 23715
rect 32689 23681 32723 23715
rect 36921 23681 36955 23715
rect 37841 23681 37875 23715
rect 40233 23681 40267 23715
rect 40693 23681 40727 23715
rect 42901 23681 42935 23715
rect 44189 23681 44223 23715
rect 45385 23681 45419 23715
rect 46305 23681 46339 23715
rect 47593 23681 47627 23715
rect 48053 23681 48087 23715
rect 48789 23681 48823 23715
rect 5457 23613 5491 23647
rect 11805 23613 11839 23647
rect 18797 23613 18831 23647
rect 19073 23613 19107 23647
rect 23857 23613 23891 23647
rect 24869 23613 24903 23647
rect 25145 23613 25179 23647
rect 30021 23613 30055 23647
rect 30297 23613 30331 23647
rect 32965 23613 32999 23647
rect 33609 23613 33643 23647
rect 33885 23613 33919 23647
rect 36369 23613 36403 23647
rect 36461 23613 36495 23647
rect 38025 23613 38059 23647
rect 39313 23613 39347 23647
rect 39405 23613 39439 23647
rect 40969 23613 41003 23647
rect 41797 23613 41831 23647
rect 42625 23613 42659 23647
rect 43913 23613 43947 23647
rect 24409 23545 24443 23579
rect 32321 23545 32355 23579
rect 37473 23545 37507 23579
rect 38485 23545 38519 23579
rect 45201 23545 45235 23579
rect 47041 23545 47075 23579
rect 6653 23477 6687 23511
rect 7297 23477 7331 23511
rect 20545 23477 20579 23511
rect 20913 23477 20947 23511
rect 22247 23477 22281 23511
rect 26617 23477 26651 23511
rect 27169 23477 27203 23511
rect 27813 23477 27847 23511
rect 29101 23477 29135 23511
rect 31769 23477 31803 23511
rect 35357 23477 35391 23511
rect 35909 23477 35943 23511
rect 40049 23477 40083 23511
rect 42165 23477 42199 23511
rect 46121 23477 46155 23511
rect 48973 23477 49007 23511
rect 49433 23477 49467 23511
rect 4721 23273 4755 23307
rect 14197 23273 14231 23307
rect 19809 23273 19843 23307
rect 24777 23273 24811 23307
rect 25237 23273 25271 23307
rect 27905 23273 27939 23307
rect 29009 23273 29043 23307
rect 29745 23273 29779 23307
rect 33149 23273 33183 23307
rect 39037 23273 39071 23307
rect 40049 23273 40083 23307
rect 44741 23273 44775 23307
rect 45661 23273 45695 23307
rect 46305 23273 46339 23307
rect 22109 23205 22143 23239
rect 31033 23205 31067 23239
rect 45201 23205 45235 23239
rect 47041 23205 47075 23239
rect 47685 23205 47719 23239
rect 6101 23137 6135 23171
rect 7849 23137 7883 23171
rect 9873 23137 9907 23171
rect 11253 23137 11287 23171
rect 13369 23137 13403 23171
rect 15761 23137 15795 23171
rect 19349 23137 19383 23171
rect 20361 23137 20395 23171
rect 22845 23137 22879 23171
rect 23949 23137 23983 23171
rect 25973 23137 26007 23171
rect 28457 23137 28491 23171
rect 30205 23137 30239 23171
rect 30389 23137 30423 23171
rect 31401 23137 31435 23171
rect 35081 23137 35115 23171
rect 35357 23137 35391 23171
rect 37289 23137 37323 23171
rect 40601 23137 40635 23171
rect 41153 23137 41187 23171
rect 41797 23137 41831 23171
rect 46489 23137 46523 23171
rect 46765 23137 46799 23171
rect 1777 23069 1811 23103
rect 4261 23069 4295 23103
rect 4905 23069 4939 23103
rect 5365 23069 5399 23103
rect 7205 23069 7239 23103
rect 9229 23069 9263 23103
rect 10701 23069 10735 23103
rect 12541 23069 12575 23103
rect 14841 23069 14875 23103
rect 15485 23069 15519 23103
rect 17141 23069 17175 23103
rect 23673 23069 23707 23103
rect 25697 23069 25731 23103
rect 33885 23069 33919 23103
rect 34345 23069 34379 23103
rect 41521 23069 41555 23103
rect 44281 23069 44315 23103
rect 45385 23069 45419 23103
rect 47225 23069 47259 23103
rect 47869 23069 47903 23103
rect 48329 23069 48363 23103
rect 49065 23069 49099 23103
rect 2789 23001 2823 23035
rect 17417 23001 17451 23035
rect 19717 23001 19751 23035
rect 20637 23001 20671 23035
rect 22661 23001 22695 23035
rect 24685 23001 24719 23035
rect 31677 23001 31711 23035
rect 34161 23001 34195 23035
rect 34713 23001 34747 23035
rect 37565 23001 37599 23035
rect 40509 23001 40543 23035
rect 43545 23001 43579 23035
rect 45017 23001 45051 23035
rect 46121 23001 46155 23035
rect 4077 22933 4111 22967
rect 9321 22933 9355 22967
rect 14657 22933 14691 22967
rect 18889 22933 18923 22967
rect 23305 22933 23339 22967
rect 23765 22933 23799 22967
rect 27445 22933 27479 22967
rect 28273 22933 28307 22967
rect 28365 22933 28399 22967
rect 29193 22933 29227 22967
rect 30113 22933 30147 22967
rect 33701 22933 33735 22967
rect 36829 22933 36863 22967
rect 39405 22933 39439 22967
rect 39589 22933 39623 22967
rect 40417 22933 40451 22967
rect 43821 22933 43855 22967
rect 44373 22933 44407 22967
rect 45937 22933 45971 22967
rect 48513 22933 48547 22967
rect 49249 22933 49283 22967
rect 12265 22729 12299 22763
rect 18613 22729 18647 22763
rect 23765 22729 23799 22763
rect 24409 22729 24443 22763
rect 30757 22729 30791 22763
rect 31493 22729 31527 22763
rect 36093 22729 36127 22763
rect 44557 22729 44591 22763
rect 46765 22729 46799 22763
rect 47961 22729 47995 22763
rect 48513 22729 48547 22763
rect 19717 22661 19751 22695
rect 21557 22661 21591 22695
rect 22293 22661 22327 22695
rect 25145 22661 25179 22695
rect 27629 22661 27663 22695
rect 32689 22661 32723 22695
rect 33977 22661 34011 22695
rect 47685 22661 47719 22695
rect 1777 22593 1811 22627
rect 3985 22593 4019 22627
rect 4813 22593 4847 22627
rect 6837 22593 6871 22627
rect 7481 22593 7515 22627
rect 9965 22593 9999 22627
rect 11805 22593 11839 22627
rect 12817 22593 12851 22627
rect 15025 22593 15059 22627
rect 16865 22593 16899 22627
rect 18981 22593 19015 22627
rect 22017 22593 22051 22627
rect 24869 22593 24903 22627
rect 27353 22593 27387 22627
rect 28089 22593 28123 22627
rect 30665 22593 30699 22627
rect 31677 22593 31711 22627
rect 32781 22593 32815 22627
rect 33701 22593 33735 22627
rect 36461 22593 36495 22627
rect 36553 22593 36587 22627
rect 37473 22593 37507 22627
rect 40049 22593 40083 22627
rect 41061 22593 41095 22627
rect 41705 22593 41739 22627
rect 41981 22593 42015 22627
rect 42809 22593 42843 22627
rect 43453 22593 43487 22627
rect 44097 22593 44131 22627
rect 44741 22593 44775 22627
rect 45017 22593 45051 22627
rect 47225 22593 47259 22627
rect 47869 22593 47903 22627
rect 48329 22593 48363 22627
rect 49065 22593 49099 22627
rect 2789 22525 2823 22559
rect 5089 22525 5123 22559
rect 7941 22525 7975 22559
rect 10241 22525 10275 22559
rect 13093 22525 13127 22559
rect 14381 22525 14415 22559
rect 15393 22525 15427 22559
rect 17141 22525 17175 22559
rect 19441 22525 19475 22559
rect 28365 22525 28399 22559
rect 30849 22525 30883 22559
rect 32873 22525 32907 22559
rect 36737 22525 36771 22559
rect 37749 22525 37783 22559
rect 40141 22525 40175 22559
rect 40233 22525 40267 22559
rect 4169 22457 4203 22491
rect 6653 22457 6687 22491
rect 21189 22457 21223 22491
rect 24225 22457 24259 22491
rect 27169 22457 27203 22491
rect 35449 22457 35483 22491
rect 39221 22457 39255 22491
rect 42625 22457 42659 22491
rect 47041 22457 47075 22491
rect 11897 22389 11931 22423
rect 26617 22389 26651 22423
rect 29837 22389 29871 22423
rect 30297 22389 30331 22423
rect 32321 22389 32355 22423
rect 33333 22389 33367 22423
rect 35725 22389 35759 22423
rect 39681 22389 39715 22423
rect 40877 22389 40911 22423
rect 41521 22389 41555 22423
rect 42165 22389 42199 22423
rect 43269 22389 43303 22423
rect 43913 22389 43947 22423
rect 49249 22389 49283 22423
rect 7849 22185 7883 22219
rect 8401 22185 8435 22219
rect 12357 22185 12391 22219
rect 13001 22185 13035 22219
rect 16957 22185 16991 22219
rect 23857 22185 23891 22219
rect 30205 22185 30239 22219
rect 32597 22185 32631 22219
rect 37552 22185 37586 22219
rect 41245 22185 41279 22219
rect 42625 22185 42659 22219
rect 42809 22185 42843 22219
rect 43177 22185 43211 22219
rect 43729 22185 43763 22219
rect 47501 22185 47535 22219
rect 29745 22117 29779 22151
rect 34437 22117 34471 22151
rect 42441 22117 42475 22151
rect 2053 22049 2087 22083
rect 4445 22049 4479 22083
rect 6285 22049 6319 22083
rect 10057 22049 10091 22083
rect 11069 22049 11103 22083
rect 13645 22049 13679 22083
rect 14749 22049 14783 22083
rect 15485 22049 15519 22083
rect 17969 22049 18003 22083
rect 19901 22049 19935 22083
rect 21097 22049 21131 22083
rect 22017 22049 22051 22083
rect 23213 22049 23247 22083
rect 25145 22049 25179 22083
rect 26525 22049 26559 22083
rect 27629 22049 27663 22083
rect 27721 22049 27755 22083
rect 28917 22049 28951 22083
rect 30849 22049 30883 22083
rect 33701 22049 33735 22083
rect 34161 22049 34195 22083
rect 35541 22049 35575 22083
rect 36737 22049 36771 22083
rect 37289 22049 37323 22083
rect 39037 22049 39071 22083
rect 40601 22049 40635 22083
rect 41705 22049 41739 22083
rect 41797 22049 41831 22083
rect 42349 22049 42383 22083
rect 1777 21981 1811 22015
rect 4077 21981 4111 22015
rect 6009 21981 6043 22015
rect 8585 21981 8619 22015
rect 9137 21981 9171 22015
rect 11345 21981 11379 22015
rect 12541 21981 12575 22015
rect 15209 21981 15243 22015
rect 17601 21981 17635 22015
rect 19441 21981 19475 22015
rect 23029 21981 23063 22015
rect 24041 21981 24075 22015
rect 28733 21981 28767 22015
rect 29929 21981 29963 22015
rect 35357 21981 35391 22015
rect 36553 21981 36587 22015
rect 40509 21981 40543 22015
rect 43269 21981 43303 22015
rect 47961 21981 47995 22015
rect 48605 21981 48639 22015
rect 7757 21913 7791 21947
rect 14565 21913 14599 21947
rect 21833 21913 21867 21947
rect 25697 21913 25731 21947
rect 26341 21913 26375 21947
rect 26433 21913 26467 21947
rect 31125 21913 31159 21947
rect 36461 21913 36495 21947
rect 39589 21913 39623 21947
rect 49157 21913 49191 21947
rect 13369 21845 13403 21879
rect 13461 21845 13495 21879
rect 21465 21845 21499 21879
rect 21925 21845 21959 21879
rect 22661 21845 22695 21879
rect 23121 21845 23155 21879
rect 24593 21845 24627 21879
rect 24961 21845 24995 21879
rect 25053 21845 25087 21879
rect 25973 21845 26007 21879
rect 27169 21845 27203 21879
rect 27537 21845 27571 21879
rect 28365 21845 28399 21879
rect 28825 21845 28859 21879
rect 33057 21845 33091 21879
rect 33425 21845 33459 21879
rect 33517 21845 33551 21879
rect 34897 21845 34931 21879
rect 35265 21845 35299 21879
rect 36093 21845 36127 21879
rect 40049 21845 40083 21879
rect 40417 21845 40451 21879
rect 41613 21845 41647 21879
rect 47777 21845 47811 21879
rect 48421 21845 48455 21879
rect 49249 21845 49283 21879
rect 10517 21641 10551 21675
rect 13277 21641 13311 21675
rect 13921 21641 13955 21675
rect 17141 21641 17175 21675
rect 17877 21641 17911 21675
rect 26433 21641 26467 21675
rect 28365 21641 28399 21675
rect 30021 21641 30055 21675
rect 32597 21641 32631 21675
rect 34437 21641 34471 21675
rect 34897 21641 34931 21675
rect 36093 21641 36127 21675
rect 40233 21641 40267 21675
rect 41981 21641 42015 21675
rect 42533 21641 42567 21675
rect 47869 21641 47903 21675
rect 48789 21641 48823 21675
rect 4353 21573 4387 21607
rect 14841 21573 14875 21607
rect 16773 21573 16807 21607
rect 16957 21573 16991 21607
rect 22753 21573 22787 21607
rect 27629 21573 27663 21607
rect 31217 21573 31251 21607
rect 36829 21573 36863 21607
rect 40601 21573 40635 21607
rect 48421 21573 48455 21607
rect 1777 21505 1811 21539
rect 3617 21505 3651 21539
rect 5917 21505 5951 21539
rect 6561 21505 6595 21539
rect 8585 21505 8619 21539
rect 10701 21505 10735 21539
rect 11897 21505 11931 21539
rect 12265 21505 12299 21539
rect 12817 21505 12851 21539
rect 13185 21505 13219 21539
rect 14105 21505 14139 21539
rect 14565 21505 14599 21539
rect 17785 21505 17819 21539
rect 21281 21505 21315 21539
rect 25145 21505 25179 21539
rect 26617 21505 26651 21539
rect 27537 21505 27571 21539
rect 28733 21505 28767 21539
rect 28825 21505 28859 21539
rect 29929 21505 29963 21539
rect 31125 21505 31159 21539
rect 33609 21505 33643 21539
rect 33701 21505 33735 21539
rect 34805 21505 34839 21539
rect 41613 21505 41647 21539
rect 42625 21505 42659 21539
rect 48053 21505 48087 21539
rect 48605 21505 48639 21539
rect 49065 21505 49099 21539
rect 2789 21437 2823 21471
rect 7021 21437 7055 21471
rect 8861 21437 8895 21471
rect 18061 21437 18095 21471
rect 18613 21437 18647 21471
rect 18889 21437 18923 21471
rect 22477 21437 22511 21471
rect 25237 21437 25271 21471
rect 25421 21437 25455 21471
rect 27721 21437 27755 21471
rect 28917 21437 28951 21471
rect 30113 21437 30147 21471
rect 31401 21437 31435 21471
rect 33793 21437 33827 21471
rect 35081 21437 35115 21471
rect 36185 21437 36219 21471
rect 36277 21437 36311 21471
rect 38025 21437 38059 21471
rect 38301 21437 38335 21471
rect 40693 21437 40727 21471
rect 40785 21437 40819 21471
rect 5733 21369 5767 21403
rect 12449 21369 12483 21403
rect 17417 21369 17451 21403
rect 21465 21369 21499 21403
rect 24777 21369 24811 21403
rect 27169 21369 27203 21403
rect 33241 21369 33275 21403
rect 41429 21369 41463 21403
rect 42165 21369 42199 21403
rect 16313 21301 16347 21335
rect 20361 21301 20395 21335
rect 20729 21301 20763 21335
rect 21925 21301 21959 21335
rect 22109 21301 22143 21335
rect 24225 21301 24259 21335
rect 25881 21301 25915 21335
rect 26065 21301 26099 21335
rect 29561 21301 29595 21335
rect 30757 21301 30791 21335
rect 35725 21301 35759 21335
rect 39773 21301 39807 21335
rect 49249 21301 49283 21335
rect 9229 21097 9263 21131
rect 11989 21097 12023 21131
rect 12909 21097 12943 21131
rect 17404 21097 17438 21131
rect 19349 21097 19383 21131
rect 21446 21097 21480 21131
rect 23581 21097 23615 21131
rect 24041 21097 24075 21131
rect 25329 21097 25363 21131
rect 26709 21097 26743 21131
rect 28365 21097 28399 21131
rect 40049 21097 40083 21131
rect 49249 21097 49283 21131
rect 19993 21029 20027 21063
rect 25697 21029 25731 21063
rect 30849 21029 30883 21063
rect 42257 21029 42291 21063
rect 4445 20961 4479 20995
rect 6285 20961 6319 20995
rect 20545 20961 20579 20995
rect 22937 20961 22971 20995
rect 26157 20961 26191 20995
rect 26249 20961 26283 20995
rect 27721 20961 27755 20995
rect 28917 20961 28951 20995
rect 30205 20961 30239 20995
rect 31309 20961 31343 20995
rect 31493 20961 31527 20995
rect 32781 20961 32815 20995
rect 34897 20961 34931 20995
rect 36921 20961 36955 20995
rect 37933 20961 37967 20995
rect 40509 20961 40543 20995
rect 40601 20961 40635 20995
rect 41797 20961 41831 20995
rect 1777 20893 1811 20927
rect 4169 20893 4203 20927
rect 5917 20893 5951 20927
rect 8033 20893 8067 20927
rect 9413 20893 9447 20927
rect 9873 20893 9907 20927
rect 11345 20893 11379 20927
rect 11897 20893 11931 20927
rect 13737 20893 13771 20927
rect 14289 20893 14323 20927
rect 17141 20893 17175 20927
rect 20361 20893 20395 20927
rect 21189 20893 21223 20927
rect 23489 20893 23523 20927
rect 24777 20893 24811 20927
rect 25053 20893 25087 20927
rect 29929 20893 29963 20927
rect 32505 20893 32539 20927
rect 37657 20893 37691 20927
rect 41613 20893 41647 20927
rect 48605 20893 48639 20927
rect 49065 20893 49099 20927
rect 2789 20825 2823 20859
rect 10517 20825 10551 20859
rect 12817 20825 12851 20859
rect 14565 20825 14599 20859
rect 26065 20825 26099 20859
rect 31217 20825 31251 20859
rect 35173 20825 35207 20859
rect 40417 20825 40451 20859
rect 41705 20825 41739 20859
rect 7849 20757 7883 20791
rect 11161 20757 11195 20791
rect 12449 20757 12483 20791
rect 13553 20757 13587 20791
rect 16037 20757 16071 20791
rect 16497 20757 16531 20791
rect 18889 20757 18923 20791
rect 20453 20757 20487 20791
rect 24133 20757 24167 20791
rect 24593 20757 24627 20791
rect 28733 20757 28767 20791
rect 28825 20757 28859 20791
rect 29745 20757 29779 20791
rect 34253 20757 34287 20791
rect 36645 20757 36679 20791
rect 39405 20757 39439 20791
rect 41245 20757 41279 20791
rect 48789 20757 48823 20791
rect 5273 20553 5307 20587
rect 9689 20553 9723 20587
rect 10333 20553 10367 20587
rect 13001 20553 13035 20587
rect 14105 20553 14139 20587
rect 14933 20553 14967 20587
rect 15577 20553 15611 20587
rect 15945 20553 15979 20587
rect 16037 20553 16071 20587
rect 18797 20553 18831 20587
rect 19165 20553 19199 20587
rect 23213 20553 23247 20587
rect 34069 20553 34103 20587
rect 34529 20553 34563 20587
rect 34897 20553 34931 20587
rect 40325 20553 40359 20587
rect 40417 20553 40451 20587
rect 12541 20485 12575 20519
rect 12725 20485 12759 20519
rect 13277 20485 13311 20519
rect 19993 20485 20027 20519
rect 29837 20485 29871 20519
rect 29929 20485 29963 20519
rect 31125 20485 31159 20519
rect 32597 20485 32631 20519
rect 38025 20485 38059 20519
rect 1777 20417 1811 20451
rect 3617 20417 3651 20451
rect 5457 20417 5491 20451
rect 6561 20417 6595 20451
rect 9229 20417 9263 20451
rect 9873 20417 9907 20451
rect 10517 20417 10551 20451
rect 11805 20417 11839 20451
rect 15117 20417 15151 20451
rect 19717 20417 19751 20451
rect 22385 20417 22419 20451
rect 23397 20417 23431 20451
rect 23857 20417 23891 20451
rect 26249 20417 26283 20451
rect 27261 20417 27295 20451
rect 31033 20417 31067 20451
rect 36461 20417 36495 20451
rect 41153 20417 41187 20451
rect 48605 20417 48639 20451
rect 49065 20417 49099 20451
rect 2789 20349 2823 20383
rect 3893 20349 3927 20383
rect 7021 20349 7055 20383
rect 10977 20349 11011 20383
rect 14197 20349 14231 20383
rect 14381 20349 14415 20383
rect 16221 20349 16255 20383
rect 16773 20349 16807 20383
rect 17049 20349 17083 20383
rect 17325 20349 17359 20383
rect 21465 20349 21499 20383
rect 22477 20349 22511 20383
rect 22569 20349 22603 20383
rect 24133 20349 24167 20383
rect 25605 20349 25639 20383
rect 27537 20349 27571 20383
rect 29009 20349 29043 20383
rect 30021 20349 30055 20383
rect 31217 20349 31251 20383
rect 32321 20349 32355 20383
rect 34989 20349 35023 20383
rect 35173 20349 35207 20383
rect 36553 20349 36587 20383
rect 36737 20349 36771 20383
rect 37749 20349 37783 20383
rect 40509 20349 40543 20383
rect 13737 20281 13771 20315
rect 31861 20281 31895 20315
rect 36093 20281 36127 20315
rect 41705 20281 41739 20315
rect 49249 20281 49283 20315
rect 9045 20213 9079 20247
rect 11897 20213 11931 20247
rect 13461 20213 13495 20247
rect 22017 20213 22051 20247
rect 26065 20213 26099 20247
rect 26617 20213 26651 20247
rect 29469 20213 29503 20247
rect 30665 20213 30699 20247
rect 35541 20213 35575 20247
rect 35817 20213 35851 20247
rect 39497 20213 39531 20247
rect 39957 20213 39991 20247
rect 48421 20213 48455 20247
rect 9965 20009 9999 20043
rect 14289 20009 14323 20043
rect 16865 20009 16899 20043
rect 18153 20009 18187 20043
rect 20269 20009 20303 20043
rect 20808 20009 20842 20043
rect 25605 20009 25639 20043
rect 26801 20009 26835 20043
rect 29193 20009 29227 20043
rect 30941 20009 30975 20043
rect 48789 20009 48823 20043
rect 11529 19941 11563 19975
rect 13737 19941 13771 19975
rect 15669 19941 15703 19975
rect 23305 19941 23339 19975
rect 25053 19941 25087 19975
rect 25237 19941 25271 19975
rect 36093 19941 36127 19975
rect 38853 19941 38887 19975
rect 41245 19941 41279 19975
rect 4905 19873 4939 19907
rect 6285 19873 6319 19907
rect 11989 19873 12023 19907
rect 16313 19873 16347 19907
rect 17509 19873 17543 19907
rect 18797 19873 18831 19907
rect 19349 19873 19383 19907
rect 20545 19873 20579 19907
rect 22293 19873 22327 19907
rect 23857 19873 23891 19907
rect 24593 19873 24627 19907
rect 26157 19873 26191 19907
rect 27353 19873 27387 19907
rect 28457 19873 28491 19907
rect 28641 19873 28675 19907
rect 29009 19873 29043 19907
rect 30297 19873 30331 19907
rect 31493 19873 31527 19907
rect 32689 19873 32723 19907
rect 33977 19873 34011 19907
rect 35541 19873 35575 19907
rect 36645 19873 36679 19907
rect 38393 19873 38427 19907
rect 39589 19873 39623 19907
rect 40509 19873 40543 19907
rect 40601 19873 40635 19907
rect 41061 19873 41095 19907
rect 1777 19805 1811 19839
rect 4077 19805 4111 19839
rect 6009 19805 6043 19839
rect 7941 19805 7975 19839
rect 10149 19805 10183 19839
rect 10793 19805 10827 19839
rect 14473 19805 14507 19839
rect 18521 19805 18555 19839
rect 18613 19805 18647 19839
rect 22569 19805 22603 19839
rect 30205 19805 30239 19839
rect 31401 19805 31435 19839
rect 32597 19805 32631 19839
rect 33885 19805 33919 19839
rect 35265 19805 35299 19839
rect 2789 19737 2823 19771
rect 11345 19737 11379 19771
rect 12265 19737 12299 19771
rect 15025 19737 15059 19771
rect 16037 19737 16071 19771
rect 17325 19737 17359 19771
rect 19717 19737 19751 19771
rect 22845 19737 22879 19771
rect 23673 19737 23707 19771
rect 23765 19737 23799 19771
rect 27169 19737 27203 19771
rect 30113 19737 30147 19771
rect 32505 19737 32539 19771
rect 33793 19737 33827 19771
rect 35357 19737 35391 19771
rect 36461 19737 36495 19771
rect 40417 19737 40451 19771
rect 48605 19737 48639 19771
rect 49157 19737 49191 19771
rect 7757 19669 7791 19703
rect 10609 19669 10643 19703
rect 15117 19669 15151 19703
rect 16129 19669 16163 19703
rect 17233 19669 17267 19703
rect 19809 19669 19843 19703
rect 22937 19669 22971 19703
rect 25973 19669 26007 19703
rect 26065 19669 26099 19703
rect 27261 19669 27295 19703
rect 27997 19669 28031 19703
rect 28365 19669 28399 19703
rect 29745 19669 29779 19703
rect 31309 19669 31343 19703
rect 32137 19669 32171 19703
rect 33425 19669 33459 19703
rect 34437 19669 34471 19703
rect 34897 19669 34931 19703
rect 36553 19669 36587 19703
rect 37841 19669 37875 19703
rect 38209 19669 38243 19703
rect 38301 19669 38335 19703
rect 39037 19669 39071 19703
rect 40049 19669 40083 19703
rect 49249 19669 49283 19703
rect 10977 19465 11011 19499
rect 14473 19465 14507 19499
rect 14841 19465 14875 19499
rect 16865 19465 16899 19499
rect 17325 19465 17359 19499
rect 20729 19465 20763 19499
rect 21189 19465 21223 19499
rect 28457 19465 28491 19499
rect 29745 19465 29779 19499
rect 30205 19465 30239 19499
rect 32321 19465 32355 19499
rect 33517 19465 33551 19499
rect 33977 19465 34011 19499
rect 34713 19465 34747 19499
rect 35909 19465 35943 19499
rect 40141 19465 40175 19499
rect 40601 19465 40635 19499
rect 41337 19465 41371 19499
rect 2789 19397 2823 19431
rect 4445 19397 4479 19431
rect 10333 19397 10367 19431
rect 16129 19397 16163 19431
rect 21097 19397 21131 19431
rect 22753 19397 22787 19431
rect 23765 19397 23799 19431
rect 28825 19397 28859 19431
rect 32689 19397 32723 19431
rect 32781 19397 32815 19431
rect 40509 19397 40543 19431
rect 1777 19329 1811 19363
rect 3617 19329 3651 19363
rect 5365 19329 5399 19363
rect 11161 19329 11195 19363
rect 11713 19329 11747 19363
rect 12081 19329 12115 19363
rect 12725 19329 12759 19363
rect 15393 19329 15427 19363
rect 17233 19329 17267 19363
rect 18061 19329 18095 19363
rect 20085 19329 20119 19363
rect 22017 19329 22051 19363
rect 23489 19329 23523 19363
rect 26157 19329 26191 19363
rect 27629 19329 27663 19363
rect 30757 19329 30791 19363
rect 31585 19329 31619 19363
rect 33885 19329 33919 19363
rect 35081 19329 35115 19363
rect 36277 19329 36311 19363
rect 36369 19329 36403 19363
rect 37933 19329 37967 19363
rect 48605 19329 48639 19363
rect 49157 19329 49191 19363
rect 9689 19261 9723 19295
rect 12265 19261 12299 19295
rect 13001 19261 13035 19295
rect 15025 19261 15059 19295
rect 15577 19261 15611 19295
rect 17417 19261 17451 19295
rect 18337 19261 18371 19295
rect 21373 19261 21407 19295
rect 26249 19261 26283 19295
rect 26433 19261 26467 19295
rect 27721 19261 27755 19295
rect 27905 19261 27939 19295
rect 28917 19261 28951 19295
rect 29101 19261 29135 19295
rect 32873 19261 32907 19295
rect 34161 19261 34195 19295
rect 35173 19261 35207 19295
rect 35357 19261 35391 19295
rect 36461 19261 36495 19295
rect 38209 19261 38243 19295
rect 40693 19261 40727 19295
rect 41153 19261 41187 19295
rect 36921 19193 36955 19227
rect 37381 19193 37415 19227
rect 49341 19193 49375 19227
rect 5457 19125 5491 19159
rect 16221 19125 16255 19159
rect 20361 19125 20395 19159
rect 25237 19125 25271 19159
rect 25789 19125 25823 19159
rect 27261 19125 27295 19159
rect 30389 19125 30423 19159
rect 39681 19125 39715 19159
rect 48789 19125 48823 19159
rect 12541 18921 12575 18955
rect 16037 18921 16071 18955
rect 16957 18921 16991 18955
rect 18153 18921 18187 18955
rect 19901 18921 19935 18955
rect 21097 18921 21131 18955
rect 24593 18921 24627 18955
rect 29009 18921 29043 18955
rect 33885 18921 33919 18955
rect 34161 18921 34195 18955
rect 34529 18921 34563 18955
rect 37381 18921 37415 18955
rect 10885 18853 10919 18887
rect 11897 18853 11931 18887
rect 13553 18853 13587 18887
rect 13829 18853 13863 18887
rect 24041 18853 24075 18887
rect 27905 18853 27939 18887
rect 31493 18853 31527 18887
rect 32689 18853 32723 18887
rect 37749 18853 37783 18887
rect 49249 18853 49283 18887
rect 4445 18785 4479 18819
rect 9137 18785 9171 18819
rect 13185 18785 13219 18819
rect 14289 18785 14323 18819
rect 14565 18785 14599 18819
rect 17509 18785 17543 18819
rect 18797 18785 18831 18819
rect 20545 18785 20579 18819
rect 21649 18785 21683 18819
rect 22293 18785 22327 18819
rect 25237 18785 25271 18819
rect 25789 18785 25823 18819
rect 27537 18785 27571 18819
rect 30205 18785 30239 18819
rect 30297 18785 30331 18819
rect 31953 18785 31987 18819
rect 32137 18785 32171 18819
rect 33333 18785 33367 18819
rect 34989 18785 35023 18819
rect 38577 18785 38611 18819
rect 1777 18717 1811 18751
rect 4077 18717 4111 18751
rect 8217 18717 8251 18751
rect 11253 18717 11287 18751
rect 11529 18717 11563 18751
rect 12081 18717 12115 18751
rect 12909 18717 12943 18751
rect 16405 18717 16439 18751
rect 17417 18717 17451 18751
rect 18521 18717 18555 18751
rect 18613 18717 18647 18751
rect 20269 18717 20303 18751
rect 28273 18717 28307 18751
rect 29193 18717 29227 18751
rect 30113 18717 30147 18751
rect 35633 18717 35667 18751
rect 40049 18717 40083 18751
rect 48605 18717 48639 18751
rect 49065 18717 49099 18751
rect 2789 18649 2823 18683
rect 9413 18649 9447 18683
rect 13001 18649 13035 18683
rect 17325 18649 17359 18683
rect 20361 18649 20395 18683
rect 22569 18649 22603 18683
rect 25053 18649 25087 18683
rect 26065 18649 26099 18683
rect 35909 18649 35943 18683
rect 40325 18649 40359 18683
rect 42073 18649 42107 18683
rect 8309 18581 8343 18615
rect 16681 18581 16715 18615
rect 19349 18581 19383 18615
rect 21465 18581 21499 18615
rect 21557 18581 21591 18615
rect 24961 18581 24995 18615
rect 27997 18581 28031 18615
rect 28457 18581 28491 18615
rect 29745 18581 29779 18615
rect 30757 18581 30791 18615
rect 31861 18581 31895 18615
rect 33057 18581 33091 18615
rect 33149 18581 33183 18615
rect 33793 18581 33827 18615
rect 34253 18581 34287 18615
rect 38025 18581 38059 18615
rect 38393 18581 38427 18615
rect 38485 18581 38519 18615
rect 41797 18581 41831 18615
rect 48421 18581 48455 18615
rect 3433 18377 3467 18411
rect 7849 18377 7883 18411
rect 10793 18377 10827 18411
rect 14289 18377 14323 18411
rect 15025 18377 15059 18411
rect 17969 18377 18003 18411
rect 18429 18377 18463 18411
rect 22109 18377 22143 18411
rect 22477 18377 22511 18411
rect 26249 18377 26283 18411
rect 27537 18377 27571 18411
rect 35909 18377 35943 18411
rect 39773 18377 39807 18411
rect 40877 18377 40911 18411
rect 48789 18377 48823 18411
rect 16681 18309 16715 18343
rect 17325 18309 17359 18343
rect 23305 18309 23339 18343
rect 24041 18309 24075 18343
rect 28825 18309 28859 18343
rect 40141 18309 40175 18343
rect 1777 18241 1811 18275
rect 3617 18241 3651 18275
rect 4445 18241 4479 18275
rect 7757 18241 7791 18275
rect 9965 18241 9999 18275
rect 10885 18241 10919 18275
rect 16313 18241 16347 18275
rect 17509 18241 17543 18275
rect 18337 18241 18371 18275
rect 19625 18241 19659 18275
rect 22569 18241 22603 18275
rect 25053 18241 25087 18275
rect 25145 18241 25179 18275
rect 26341 18241 26375 18275
rect 28733 18241 28767 18275
rect 30481 18241 30515 18275
rect 31309 18241 31343 18275
rect 32689 18241 32723 18275
rect 36277 18241 36311 18275
rect 36369 18241 36403 18275
rect 37657 18241 37691 18275
rect 38025 18241 38059 18275
rect 40785 18241 40819 18275
rect 48605 18241 48639 18275
rect 49065 18241 49099 18275
rect 2789 18173 2823 18207
rect 4169 18173 4203 18207
rect 10977 18173 11011 18207
rect 11713 18173 11747 18207
rect 11989 18173 12023 18207
rect 14381 18173 14415 18207
rect 14565 18173 14599 18207
rect 15485 18173 15519 18207
rect 18613 18173 18647 18207
rect 19901 18173 19935 18207
rect 22753 18173 22787 18207
rect 25329 18173 25363 18207
rect 26433 18173 26467 18207
rect 27629 18173 27663 18207
rect 27813 18173 27847 18207
rect 28917 18173 28951 18207
rect 30573 18173 30607 18207
rect 30757 18173 30791 18207
rect 32781 18173 32815 18207
rect 32965 18173 32999 18207
rect 33609 18173 33643 18207
rect 33885 18173 33919 18207
rect 35357 18173 35391 18207
rect 36553 18173 36587 18207
rect 38301 18173 38335 18207
rect 40969 18173 41003 18207
rect 9781 18105 9815 18139
rect 10425 18105 10459 18139
rect 13921 18105 13955 18139
rect 15209 18105 15243 18139
rect 16129 18105 16163 18139
rect 24685 18105 24719 18139
rect 28365 18105 28399 18139
rect 29745 18105 29779 18139
rect 30113 18105 30147 18139
rect 40417 18105 40451 18139
rect 13461 18037 13495 18071
rect 18981 18037 19015 18071
rect 21373 18037 21407 18071
rect 25881 18037 25915 18071
rect 27169 18037 27203 18071
rect 32321 18037 32355 18071
rect 49249 18037 49283 18071
rect 12357 17833 12391 17867
rect 12909 17833 12943 17867
rect 16037 17833 16071 17867
rect 16773 17833 16807 17867
rect 19441 17833 19475 17867
rect 23305 17833 23339 17867
rect 29285 17833 29319 17867
rect 34345 17833 34379 17867
rect 16497 17765 16531 17799
rect 24593 17765 24627 17799
rect 25789 17765 25823 17799
rect 26341 17765 26375 17799
rect 29101 17765 29135 17799
rect 34529 17765 34563 17799
rect 38025 17765 38059 17799
rect 40509 17765 40543 17799
rect 2053 17697 2087 17731
rect 10609 17697 10643 17731
rect 14289 17697 14323 17731
rect 17417 17697 17451 17731
rect 18797 17697 18831 17731
rect 20269 17697 20303 17731
rect 22017 17697 22051 17731
rect 23765 17697 23799 17731
rect 23857 17697 23891 17731
rect 25053 17697 25087 17731
rect 25145 17697 25179 17731
rect 27077 17697 27111 17731
rect 31953 17697 31987 17731
rect 33241 17697 33275 17731
rect 33425 17697 33459 17731
rect 35817 17697 35851 17731
rect 36093 17697 36127 17731
rect 37565 17697 37599 17731
rect 38485 17697 38519 17731
rect 38577 17697 38611 17731
rect 40969 17697 41003 17731
rect 41061 17697 41095 17731
rect 1777 17629 1811 17663
rect 13093 17629 13127 17663
rect 13737 17629 13771 17663
rect 17141 17629 17175 17663
rect 17969 17629 18003 17663
rect 19625 17629 19659 17663
rect 25973 17629 26007 17663
rect 29929 17629 29963 17663
rect 31677 17629 31711 17663
rect 48605 17629 48639 17663
rect 49065 17629 49099 17663
rect 10885 17561 10919 17595
rect 14565 17561 14599 17595
rect 20545 17561 20579 17595
rect 22661 17561 22695 17595
rect 23673 17561 23707 17595
rect 27353 17561 27387 17595
rect 30757 17561 30791 17595
rect 40877 17561 40911 17595
rect 13553 17493 13587 17527
rect 17233 17493 17267 17527
rect 22293 17493 22327 17527
rect 24961 17493 24995 17527
rect 26433 17493 26467 17527
rect 28825 17493 28859 17527
rect 29653 17493 29687 17527
rect 31309 17493 31343 17527
rect 31769 17493 31803 17527
rect 32413 17493 32447 17527
rect 32781 17493 32815 17527
rect 33149 17493 33183 17527
rect 33793 17493 33827 17527
rect 34897 17493 34931 17527
rect 35541 17493 35575 17527
rect 38393 17493 38427 17527
rect 48789 17493 48823 17527
rect 49249 17493 49283 17527
rect 10425 17289 10459 17323
rect 14933 17289 14967 17323
rect 15577 17289 15611 17323
rect 16037 17289 16071 17323
rect 20913 17289 20947 17323
rect 24409 17289 24443 17323
rect 24869 17289 24903 17323
rect 25329 17289 25363 17323
rect 27353 17289 27387 17323
rect 27813 17289 27847 17323
rect 28641 17289 28675 17323
rect 34069 17289 34103 17323
rect 37841 17289 37875 17323
rect 48421 17289 48455 17323
rect 49249 17289 49283 17323
rect 10149 17221 10183 17255
rect 11805 17221 11839 17255
rect 12449 17221 12483 17255
rect 13093 17221 13127 17255
rect 14197 17221 14231 17255
rect 17785 17221 17819 17255
rect 25973 17221 26007 17255
rect 29009 17221 29043 17255
rect 29101 17221 29135 17255
rect 30205 17221 30239 17255
rect 32597 17221 32631 17255
rect 34621 17221 34655 17255
rect 36461 17221 36495 17255
rect 41061 17221 41095 17255
rect 1777 17153 1811 17187
rect 10793 17153 10827 17187
rect 15117 17153 15151 17187
rect 15945 17153 15979 17187
rect 16957 17153 16991 17187
rect 19165 17153 19199 17187
rect 22661 17153 22695 17187
rect 25237 17153 25271 17187
rect 27721 17153 27755 17187
rect 30297 17153 30331 17187
rect 31401 17153 31435 17187
rect 32321 17153 32355 17187
rect 36369 17153 36403 17187
rect 37933 17153 37967 17187
rect 48605 17153 48639 17187
rect 49157 17153 49191 17187
rect 2053 17085 2087 17119
rect 10885 17085 10919 17119
rect 10977 17085 11011 17119
rect 13185 17085 13219 17119
rect 13277 17085 13311 17119
rect 13829 17085 13863 17119
rect 16129 17085 16163 17119
rect 17141 17085 17175 17119
rect 18613 17085 18647 17119
rect 19441 17085 19475 17119
rect 22937 17085 22971 17119
rect 25421 17085 25455 17119
rect 27997 17085 28031 17119
rect 29193 17085 29227 17119
rect 30389 17085 30423 17119
rect 31493 17085 31527 17119
rect 31585 17085 31619 17119
rect 35357 17085 35391 17119
rect 36645 17085 36679 17119
rect 38117 17085 38151 17119
rect 38485 17085 38519 17119
rect 38945 17085 38979 17119
rect 39221 17085 39255 17119
rect 14381 17017 14415 17051
rect 36001 17017 36035 17051
rect 37473 17017 37507 17051
rect 9873 16949 9907 16983
rect 11897 16949 11931 16983
rect 12725 16949 12759 16983
rect 17509 16949 17543 16983
rect 21281 16949 21315 16983
rect 21649 16949 21683 16983
rect 22201 16949 22235 16983
rect 29837 16949 29871 16983
rect 31033 16949 31067 16983
rect 37013 16949 37047 16983
rect 40693 16949 40727 16983
rect 14197 16745 14231 16779
rect 17404 16745 17438 16779
rect 27353 16745 27387 16779
rect 28641 16745 28675 16779
rect 34529 16745 34563 16779
rect 48789 16745 48823 16779
rect 22753 16677 22787 16711
rect 28181 16677 28215 16711
rect 34253 16677 34287 16711
rect 36277 16677 36311 16711
rect 37381 16677 37415 16711
rect 41245 16677 41279 16711
rect 41521 16677 41555 16711
rect 8217 16609 8251 16643
rect 8401 16609 8435 16643
rect 10609 16609 10643 16643
rect 11621 16609 11655 16643
rect 13645 16609 13679 16643
rect 15025 16609 15059 16643
rect 16129 16609 16163 16643
rect 16221 16609 16255 16643
rect 17141 16609 17175 16643
rect 21281 16609 21315 16643
rect 23765 16609 23799 16643
rect 23949 16609 23983 16643
rect 25605 16609 25639 16643
rect 25881 16609 25915 16643
rect 27997 16609 28031 16643
rect 29285 16609 29319 16643
rect 30297 16609 30331 16643
rect 31401 16609 31435 16643
rect 31585 16609 31619 16643
rect 32229 16609 32263 16643
rect 35725 16609 35759 16643
rect 36737 16609 36771 16643
rect 36829 16609 36863 16643
rect 40509 16609 40543 16643
rect 40601 16609 40635 16643
rect 41061 16609 41095 16643
rect 1777 16541 1811 16575
rect 12541 16541 12575 16575
rect 14841 16541 14875 16575
rect 16681 16541 16715 16575
rect 20269 16541 20303 16575
rect 21005 16541 21039 16575
rect 27629 16541 27663 16575
rect 34897 16541 34931 16575
rect 37749 16541 37783 16575
rect 40417 16541 40451 16575
rect 48605 16541 48639 16575
rect 49065 16541 49099 16575
rect 2513 16473 2547 16507
rect 10057 16473 10091 16507
rect 10425 16473 10459 16507
rect 11437 16473 11471 16507
rect 16037 16473 16071 16507
rect 24685 16473 24719 16507
rect 28365 16473 28399 16507
rect 30113 16473 30147 16507
rect 30205 16473 30239 16507
rect 32505 16473 32539 16507
rect 38025 16473 38059 16507
rect 7757 16405 7791 16439
rect 8125 16405 8159 16439
rect 11069 16405 11103 16439
rect 11529 16405 11563 16439
rect 12357 16405 12391 16439
rect 13001 16405 13035 16439
rect 13369 16405 13403 16439
rect 13461 16405 13495 16439
rect 14473 16405 14507 16439
rect 14933 16405 14967 16439
rect 15669 16405 15703 16439
rect 18889 16405 18923 16439
rect 19441 16405 19475 16439
rect 20085 16405 20119 16439
rect 20637 16405 20671 16439
rect 23305 16405 23339 16439
rect 23673 16405 23707 16439
rect 24593 16405 24627 16439
rect 29745 16405 29779 16439
rect 30941 16405 30975 16439
rect 31309 16405 31343 16439
rect 33977 16405 34011 16439
rect 36645 16405 36679 16439
rect 39497 16405 39531 16439
rect 40049 16405 40083 16439
rect 49249 16405 49283 16439
rect 8309 16201 8343 16235
rect 9321 16201 9355 16235
rect 11069 16201 11103 16235
rect 11989 16201 12023 16235
rect 12449 16201 12483 16235
rect 13185 16201 13219 16235
rect 13553 16201 13587 16235
rect 14381 16201 14415 16235
rect 14749 16201 14783 16235
rect 17417 16201 17451 16235
rect 18797 16201 18831 16235
rect 23121 16201 23155 16235
rect 26341 16201 26375 16235
rect 30113 16201 30147 16235
rect 30941 16201 30975 16235
rect 31033 16201 31067 16235
rect 33977 16201 34011 16235
rect 36829 16201 36863 16235
rect 40969 16201 41003 16235
rect 13645 16133 13679 16167
rect 15945 16133 15979 16167
rect 19441 16133 19475 16167
rect 21373 16133 21407 16167
rect 23489 16133 23523 16167
rect 27629 16133 27663 16167
rect 32781 16133 32815 16167
rect 34805 16133 34839 16167
rect 38485 16133 38519 16167
rect 1777 16065 1811 16099
rect 9229 16065 9263 16099
rect 10977 16065 11011 16099
rect 12357 16065 12391 16099
rect 17785 16065 17819 16099
rect 19165 16065 19199 16099
rect 24593 16065 24627 16099
rect 27537 16065 27571 16099
rect 28365 16065 28399 16099
rect 32689 16065 32723 16099
rect 33885 16065 33919 16099
rect 38209 16065 38243 16099
rect 40877 16065 40911 16099
rect 48789 16065 48823 16099
rect 49065 16065 49099 16099
rect 2053 15997 2087 16031
rect 8401 15997 8435 16031
rect 8493 15997 8527 16031
rect 10425 15997 10459 16031
rect 12541 15997 12575 16031
rect 13737 15997 13771 16031
rect 14841 15997 14875 16031
rect 15025 15997 15059 16031
rect 15761 15997 15795 16031
rect 15853 15997 15887 16031
rect 17877 15997 17911 16031
rect 18061 15997 18095 16031
rect 23581 15997 23615 16031
rect 23765 15997 23799 16031
rect 24869 15997 24903 16031
rect 27721 15997 27755 16031
rect 28641 15997 28675 16031
rect 31125 15997 31159 16031
rect 32873 15997 32907 16031
rect 34069 15997 34103 16031
rect 34621 15997 34655 16031
rect 35081 15997 35115 16031
rect 35357 15997 35391 16031
rect 37473 15997 37507 16031
rect 39957 15997 39991 16031
rect 41061 15997 41095 16031
rect 16773 15929 16807 15963
rect 20913 15929 20947 15963
rect 22845 15929 22879 15963
rect 49249 15929 49283 15963
rect 7941 15861 7975 15895
rect 10609 15861 10643 15895
rect 11713 15861 11747 15895
rect 15393 15861 15427 15895
rect 16313 15861 16347 15895
rect 16865 15861 16899 15895
rect 17141 15861 17175 15895
rect 26617 15861 26651 15895
rect 27169 15861 27203 15895
rect 30573 15861 30607 15895
rect 31585 15861 31619 15895
rect 31769 15861 31803 15895
rect 32321 15861 32355 15895
rect 33517 15861 33551 15895
rect 40509 15861 40543 15895
rect 41613 15861 41647 15895
rect 16773 15657 16807 15691
rect 18981 15657 19015 15691
rect 19349 15657 19383 15691
rect 19901 15657 19935 15691
rect 21189 15657 21223 15691
rect 22477 15657 22511 15691
rect 25881 15657 25915 15691
rect 27169 15657 27203 15691
rect 32229 15657 32263 15691
rect 34345 15657 34379 15691
rect 36645 15657 36679 15691
rect 39497 15657 39531 15691
rect 42073 15657 42107 15691
rect 49157 15657 49191 15691
rect 14289 15589 14323 15623
rect 15577 15589 15611 15623
rect 2053 15521 2087 15555
rect 10793 15521 10827 15555
rect 11069 15521 11103 15555
rect 13461 15521 13495 15555
rect 13645 15521 13679 15555
rect 14841 15521 14875 15555
rect 16037 15521 16071 15555
rect 16221 15521 16255 15555
rect 17233 15521 17267 15555
rect 17325 15521 17359 15555
rect 20545 15521 20579 15555
rect 21649 15521 21683 15555
rect 21833 15521 21867 15555
rect 23765 15521 23799 15555
rect 25145 15521 25179 15555
rect 25329 15521 25363 15555
rect 26525 15521 26559 15555
rect 27997 15521 28031 15555
rect 30757 15521 30791 15555
rect 33149 15521 33183 15555
rect 33333 15521 33367 15555
rect 35173 15521 35207 15555
rect 40049 15521 40083 15555
rect 40325 15521 40359 15555
rect 1777 15453 1811 15487
rect 13369 15453 13403 15487
rect 15945 15453 15979 15487
rect 17141 15453 17175 15487
rect 17785 15453 17819 15487
rect 18613 15453 18647 15487
rect 21557 15453 21591 15487
rect 22201 15453 22235 15487
rect 23581 15453 23615 15487
rect 27813 15453 27847 15487
rect 28457 15453 28491 15487
rect 30481 15453 30515 15487
rect 33057 15453 33091 15487
rect 34897 15453 34931 15487
rect 37749 15453 37783 15487
rect 48881 15453 48915 15487
rect 49341 15453 49375 15487
rect 6469 15385 6503 15419
rect 14749 15385 14783 15419
rect 20361 15385 20395 15419
rect 23489 15385 23523 15419
rect 25053 15385 25087 15419
rect 26341 15385 26375 15419
rect 27905 15385 27939 15419
rect 28641 15385 28675 15419
rect 29193 15385 29227 15419
rect 38025 15385 38059 15419
rect 6561 15317 6595 15351
rect 12541 15317 12575 15351
rect 13001 15317 13035 15351
rect 14657 15317 14691 15351
rect 18429 15317 18463 15351
rect 20269 15317 20303 15351
rect 23121 15317 23155 15351
rect 24685 15317 24719 15351
rect 26249 15317 26283 15351
rect 26985 15317 27019 15351
rect 27445 15317 27479 15351
rect 29285 15317 29319 15351
rect 29837 15317 29871 15351
rect 32689 15317 32723 15351
rect 33885 15317 33919 15351
rect 37105 15317 37139 15351
rect 41797 15317 41831 15351
rect 9781 15113 9815 15147
rect 15025 15113 15059 15147
rect 15577 15113 15611 15147
rect 15945 15113 15979 15147
rect 18337 15113 18371 15147
rect 18705 15113 18739 15147
rect 19533 15113 19567 15147
rect 21833 15113 21867 15147
rect 22937 15113 22971 15147
rect 23397 15113 23431 15147
rect 24133 15113 24167 15147
rect 29745 15113 29779 15147
rect 30665 15113 30699 15147
rect 31401 15113 31435 15147
rect 32689 15113 32723 15147
rect 33885 15113 33919 15147
rect 34713 15113 34747 15147
rect 35081 15113 35115 15147
rect 39681 15113 39715 15147
rect 40141 15113 40175 15147
rect 49249 15113 49283 15147
rect 9873 15045 9907 15079
rect 10609 15045 10643 15079
rect 10977 15045 11011 15079
rect 11161 15045 11195 15079
rect 16037 15045 16071 15079
rect 19901 15045 19935 15079
rect 21097 15045 21131 15079
rect 25329 15045 25363 15079
rect 26341 15045 26375 15079
rect 27629 15045 27663 15079
rect 30573 15045 30607 15079
rect 31861 15045 31895 15079
rect 32781 15045 32815 15079
rect 40049 15045 40083 15079
rect 1777 14977 1811 15011
rect 12265 14977 12299 15011
rect 13277 14977 13311 15011
rect 17233 14977 17267 15011
rect 18797 14977 18831 15011
rect 19993 14977 20027 15011
rect 23305 14977 23339 15011
rect 24501 14977 24535 15011
rect 25237 14977 25271 15011
rect 26249 14977 26283 15011
rect 26985 14977 27019 15011
rect 27997 14977 28031 15011
rect 36277 14977 36311 15011
rect 36921 14977 36955 15011
rect 37473 14977 37507 15011
rect 41061 14977 41095 15011
rect 48789 14977 48823 15011
rect 49065 14977 49099 15011
rect 2053 14909 2087 14943
rect 10057 14909 10091 14943
rect 11621 14909 11655 14943
rect 12357 14909 12391 14943
rect 12449 14909 12483 14943
rect 13553 14909 13587 14943
rect 16129 14909 16163 14943
rect 17325 14909 17359 14943
rect 17417 14909 17451 14943
rect 18061 14909 18095 14943
rect 18889 14909 18923 14943
rect 20085 14909 20119 14943
rect 21189 14909 21223 14943
rect 21281 14909 21315 14943
rect 23581 14909 23615 14943
rect 24593 14909 24627 14943
rect 24685 14909 24719 14943
rect 26433 14909 26467 14943
rect 28273 14909 28307 14943
rect 30757 14909 30791 14943
rect 32965 14909 32999 14943
rect 33977 14909 34011 14943
rect 34069 14909 34103 14943
rect 35173 14909 35207 14943
rect 35357 14909 35391 14943
rect 36369 14909 36403 14943
rect 36553 14909 36587 14943
rect 37749 14909 37783 14943
rect 40233 14909 40267 14943
rect 11897 14841 11931 14875
rect 20729 14841 20763 14875
rect 25881 14841 25915 14875
rect 27261 14841 27295 14875
rect 32321 14841 32355 14875
rect 35909 14841 35943 14875
rect 9413 14773 9447 14807
rect 12909 14773 12943 14807
rect 16865 14773 16899 14807
rect 22017 14773 22051 14807
rect 25605 14773 25639 14807
rect 27445 14773 27479 14807
rect 30205 14773 30239 14807
rect 33517 14773 33551 14807
rect 39221 14773 39255 14807
rect 40877 14773 40911 14807
rect 10425 14569 10459 14603
rect 11805 14569 11839 14603
rect 13001 14569 13035 14603
rect 17693 14569 17727 14603
rect 18153 14569 18187 14603
rect 22845 14569 22879 14603
rect 23305 14569 23339 14603
rect 23581 14569 23615 14603
rect 27353 14569 27387 14603
rect 29745 14569 29779 14603
rect 36645 14569 36679 14603
rect 38853 14569 38887 14603
rect 39865 14569 39899 14603
rect 40049 14569 40083 14603
rect 14473 14501 14507 14535
rect 27813 14501 27847 14535
rect 2053 14433 2087 14467
rect 12357 14433 12391 14467
rect 13553 14433 13587 14467
rect 15025 14433 15059 14467
rect 16957 14433 16991 14467
rect 18705 14433 18739 14467
rect 20085 14433 20119 14467
rect 21097 14433 21131 14467
rect 21373 14433 21407 14467
rect 25605 14433 25639 14467
rect 28273 14433 28307 14467
rect 28457 14433 28491 14467
rect 30389 14433 30423 14467
rect 31493 14433 31527 14467
rect 32597 14433 32631 14467
rect 32689 14433 32723 14467
rect 33885 14433 33919 14467
rect 34897 14433 34931 14467
rect 37105 14433 37139 14467
rect 49341 14433 49375 14467
rect 1777 14365 1811 14399
rect 9781 14365 9815 14399
rect 10333 14365 10367 14399
rect 11161 14365 11195 14399
rect 14197 14365 14231 14399
rect 14933 14365 14967 14399
rect 30113 14365 30147 14399
rect 31401 14365 31435 14399
rect 33701 14365 33735 14399
rect 33793 14365 33827 14399
rect 39497 14365 39531 14399
rect 48605 14365 48639 14399
rect 49157 14365 49191 14399
rect 9597 14297 9631 14331
rect 12173 14297 12207 14331
rect 13369 14297 13403 14331
rect 15761 14297 15795 14331
rect 16773 14297 16807 14331
rect 18613 14297 18647 14331
rect 19901 14297 19935 14331
rect 25888 14297 25922 14331
rect 28181 14297 28215 14331
rect 32505 14297 32539 14331
rect 35173 14297 35207 14331
rect 37381 14297 37415 14331
rect 11253 14229 11287 14263
rect 12265 14229 12299 14263
rect 13461 14229 13495 14263
rect 14841 14229 14875 14263
rect 16405 14229 16439 14263
rect 16865 14229 16899 14263
rect 17509 14229 17543 14263
rect 18521 14229 18555 14263
rect 19533 14229 19567 14263
rect 19993 14229 20027 14263
rect 20545 14229 20579 14263
rect 20729 14229 20763 14263
rect 23857 14229 23891 14263
rect 24409 14229 24443 14263
rect 24593 14229 24627 14263
rect 24961 14229 24995 14263
rect 29009 14229 29043 14263
rect 30205 14229 30239 14263
rect 30941 14229 30975 14263
rect 31309 14229 31343 14263
rect 32137 14229 32171 14263
rect 33333 14229 33367 14263
rect 34529 14229 34563 14263
rect 39313 14229 39347 14263
rect 48697 14229 48731 14263
rect 3617 14025 3651 14059
rect 10425 14025 10459 14059
rect 10701 14025 10735 14059
rect 11713 14025 11747 14059
rect 14749 14025 14783 14059
rect 15577 14025 15611 14059
rect 17141 14025 17175 14059
rect 17509 14025 17543 14059
rect 18337 14025 18371 14059
rect 18705 14025 18739 14059
rect 23765 14025 23799 14059
rect 26617 14025 26651 14059
rect 31125 14025 31159 14059
rect 31585 14025 31619 14059
rect 36093 14025 36127 14059
rect 36737 14025 36771 14059
rect 37473 14025 37507 14059
rect 45661 14025 45695 14059
rect 48421 14025 48455 14059
rect 49249 14025 49283 14059
rect 25145 13957 25179 13991
rect 28917 13957 28951 13991
rect 37933 13957 37967 13991
rect 45017 13957 45051 13991
rect 48145 13957 48179 13991
rect 49157 13957 49191 13991
rect 1777 13889 1811 13923
rect 3525 13889 3559 13923
rect 3985 13889 4019 13923
rect 10977 13889 11011 13923
rect 12081 13889 12115 13923
rect 12173 13889 12207 13923
rect 15945 13889 15979 13923
rect 17601 13889 17635 13923
rect 18797 13889 18831 13923
rect 24869 13889 24903 13923
rect 27169 13889 27203 13923
rect 29377 13889 29411 13923
rect 34897 13889 34931 13923
rect 34989 13889 35023 13923
rect 37841 13889 37875 13923
rect 39037 13889 39071 13923
rect 45845 13889 45879 13923
rect 48605 13889 48639 13923
rect 2053 13821 2087 13855
rect 9873 13821 9907 13855
rect 12265 13821 12299 13855
rect 13001 13821 13035 13855
rect 13277 13821 13311 13855
rect 15025 13821 15059 13855
rect 15209 13821 15243 13855
rect 16037 13821 16071 13855
rect 16221 13821 16255 13855
rect 16773 13821 16807 13855
rect 17693 13821 17727 13855
rect 18889 13821 18923 13855
rect 19717 13821 19751 13855
rect 21465 13821 21499 13855
rect 22017 13821 22051 13855
rect 22293 13821 22327 13855
rect 24225 13821 24259 13855
rect 32321 13821 32355 13855
rect 32597 13821 32631 13855
rect 35173 13821 35207 13855
rect 36185 13821 36219 13855
rect 36369 13821 36403 13855
rect 38025 13821 38059 13855
rect 45201 13821 45235 13855
rect 34069 13753 34103 13787
rect 34529 13753 34563 13787
rect 35725 13753 35759 13787
rect 19349 13685 19383 13719
rect 19980 13685 20014 13719
rect 29640 13685 29674 13719
rect 14473 13481 14507 13515
rect 14933 13481 14967 13515
rect 18153 13481 18187 13515
rect 19717 13481 19751 13515
rect 22109 13481 22143 13515
rect 23305 13481 23339 13515
rect 24869 13481 24903 13515
rect 28089 13481 28123 13515
rect 28457 13481 28491 13515
rect 32781 13481 32815 13515
rect 33333 13481 33367 13515
rect 34897 13481 34931 13515
rect 38485 13481 38519 13515
rect 12541 13413 12575 13447
rect 15209 13413 15243 13447
rect 19441 13413 19475 13447
rect 29745 13413 29779 13447
rect 10793 13345 10827 13379
rect 15669 13345 15703 13379
rect 15853 13345 15887 13379
rect 16405 13345 16439 13379
rect 20177 13345 20211 13379
rect 20269 13345 20303 13379
rect 21465 13345 21499 13379
rect 22569 13345 22603 13379
rect 22753 13345 22787 13379
rect 23949 13345 23983 13379
rect 25513 13345 25547 13379
rect 29101 13345 29135 13379
rect 30297 13345 30331 13379
rect 31033 13345 31067 13379
rect 33885 13345 33919 13379
rect 35541 13345 35575 13379
rect 1777 13277 1811 13311
rect 2789 13277 2823 13311
rect 23673 13277 23707 13311
rect 25237 13277 25271 13311
rect 28917 13277 28951 13311
rect 30113 13277 30147 13311
rect 33701 13277 33735 13311
rect 35265 13277 35299 13311
rect 36461 13277 36495 13311
rect 41521 13277 41555 13311
rect 47961 13277 47995 13311
rect 11069 13209 11103 13243
rect 13737 13209 13771 13243
rect 14381 13209 14415 13243
rect 15577 13209 15611 13243
rect 16681 13209 16715 13243
rect 18705 13209 18739 13243
rect 20085 13209 20119 13243
rect 22477 13209 22511 13243
rect 23765 13209 23799 13243
rect 31309 13209 31343 13243
rect 34345 13209 34379 13243
rect 35357 13209 35391 13243
rect 36093 13209 36127 13243
rect 36737 13209 36771 13243
rect 49157 13209 49191 13243
rect 13093 13141 13127 13175
rect 13921 13141 13955 13175
rect 20913 13141 20947 13175
rect 21281 13141 21315 13175
rect 21373 13141 21407 13175
rect 24501 13141 24535 13175
rect 25329 13141 25363 13175
rect 26065 13141 26099 13175
rect 26801 13141 26835 13175
rect 27721 13141 27755 13175
rect 28825 13141 28859 13175
rect 30205 13141 30239 13175
rect 33793 13141 33827 13175
rect 36001 13141 36035 13175
rect 38209 13141 38243 13175
rect 41337 13141 41371 13175
rect 2881 12937 2915 12971
rect 12173 12937 12207 12971
rect 14841 12937 14875 12971
rect 15945 12937 15979 12971
rect 16865 12937 16899 12971
rect 20729 12937 20763 12971
rect 22661 12937 22695 12971
rect 23121 12937 23155 12971
rect 25605 12937 25639 12971
rect 26709 12937 26743 12971
rect 31769 12937 31803 12971
rect 32689 12937 32723 12971
rect 32781 12937 32815 12971
rect 33793 12937 33827 12971
rect 35817 12937 35851 12971
rect 35909 12937 35943 12971
rect 36645 12937 36679 12971
rect 36921 12937 36955 12971
rect 37013 12937 37047 12971
rect 1685 12869 1719 12903
rect 2145 12869 2179 12903
rect 11345 12869 11379 12903
rect 12081 12869 12115 12903
rect 12817 12869 12851 12903
rect 17877 12869 17911 12903
rect 21189 12869 21223 12903
rect 26157 12869 26191 12903
rect 27445 12869 27479 12903
rect 29561 12869 29595 12903
rect 34897 12869 34931 12903
rect 37749 12869 37783 12903
rect 40049 12869 40083 12903
rect 40509 12869 40543 12903
rect 3065 12801 3099 12835
rect 3341 12801 3375 12835
rect 13093 12801 13127 12835
rect 16037 12801 16071 12835
rect 18705 12801 18739 12835
rect 19625 12801 19659 12835
rect 21097 12801 21131 12835
rect 23029 12801 23063 12835
rect 26341 12801 26375 12835
rect 27169 12801 27203 12835
rect 30021 12801 30055 12835
rect 34069 12801 34103 12835
rect 37473 12801 37507 12835
rect 46121 12801 46155 12835
rect 47961 12801 47995 12835
rect 49157 12801 49191 12835
rect 1869 12733 1903 12767
rect 12265 12733 12299 12767
rect 13369 12733 13403 12767
rect 16129 12733 16163 12767
rect 17233 12733 17267 12767
rect 19717 12733 19751 12767
rect 19901 12733 19935 12767
rect 21281 12733 21315 12767
rect 22017 12733 22051 12767
rect 23213 12733 23247 12767
rect 23857 12733 23891 12767
rect 24133 12733 24167 12767
rect 29193 12733 29227 12767
rect 30297 12733 30331 12767
rect 32873 12733 32907 12767
rect 36093 12733 36127 12767
rect 39497 12733 39531 12767
rect 15301 12665 15335 12699
rect 16773 12665 16807 12699
rect 20453 12665 20487 12699
rect 25881 12665 25915 12699
rect 35449 12665 35483 12699
rect 40233 12665 40267 12699
rect 11713 12597 11747 12631
rect 15577 12597 15611 12631
rect 19257 12597 19291 12631
rect 32321 12597 32355 12631
rect 33425 12597 33459 12631
rect 33609 12597 33643 12631
rect 36553 12597 36587 12631
rect 45937 12597 45971 12631
rect 16037 12393 16071 12427
rect 19441 12393 19475 12427
rect 20913 12393 20947 12427
rect 23305 12393 23339 12427
rect 26985 12393 27019 12427
rect 38301 12393 38335 12427
rect 33885 12325 33919 12359
rect 37105 12325 37139 12359
rect 1869 12257 1903 12291
rect 9505 12257 9539 12291
rect 11713 12257 11747 12291
rect 14289 12257 14323 12291
rect 14565 12257 14599 12291
rect 17325 12257 17359 12291
rect 19993 12257 20027 12291
rect 20637 12257 20671 12291
rect 21373 12257 21407 12291
rect 21557 12257 21591 12291
rect 22661 12257 22695 12291
rect 23949 12257 23983 12291
rect 24869 12257 24903 12291
rect 27537 12257 27571 12291
rect 29101 12257 29135 12291
rect 29745 12257 29779 12291
rect 32137 12257 32171 12291
rect 35173 12257 35207 12291
rect 37565 12257 37599 12291
rect 37657 12257 37691 12291
rect 38853 12257 38887 12291
rect 49157 12257 49191 12291
rect 1593 12189 1627 12223
rect 16497 12189 16531 12223
rect 17141 12189 17175 12223
rect 17969 12189 18003 12223
rect 19809 12189 19843 12223
rect 21281 12189 21315 12223
rect 24593 12189 24627 12223
rect 26617 12189 26651 12223
rect 28273 12189 28307 12223
rect 34897 12189 34931 12223
rect 38761 12189 38795 12223
rect 39405 12189 39439 12223
rect 40141 12189 40175 12223
rect 40969 12189 41003 12223
rect 41613 12189 41647 12223
rect 46121 12189 46155 12223
rect 47961 12189 47995 12223
rect 2697 12121 2731 12155
rect 9781 12121 9815 12155
rect 11989 12121 12023 12155
rect 13737 12121 13771 12155
rect 18705 12121 18739 12155
rect 23673 12121 23707 12155
rect 27445 12121 27479 12155
rect 30021 12121 30055 12155
rect 32413 12121 32447 12155
rect 39589 12121 39623 12155
rect 40325 12121 40359 12155
rect 11253 12053 11287 12087
rect 16773 12053 16807 12087
rect 17233 12053 17267 12087
rect 19901 12053 19935 12087
rect 22109 12053 22143 12087
rect 22477 12053 22511 12087
rect 22569 12053 22603 12087
rect 23765 12053 23799 12087
rect 26341 12053 26375 12087
rect 27353 12053 27387 12087
rect 31493 12053 31527 12087
rect 31861 12053 31895 12087
rect 34253 12053 34287 12087
rect 34437 12053 34471 12087
rect 36645 12053 36679 12087
rect 37473 12053 37507 12087
rect 38669 12053 38703 12087
rect 40785 12053 40819 12087
rect 41429 12053 41463 12087
rect 45937 12053 45971 12087
rect 2329 11849 2363 11883
rect 11621 11849 11655 11883
rect 12725 11849 12759 11883
rect 13553 11849 13587 11883
rect 14381 11849 14415 11883
rect 15577 11849 15611 11883
rect 16405 11849 16439 11883
rect 25697 11849 25731 11883
rect 26433 11849 26467 11883
rect 27629 11849 27663 11883
rect 30757 11849 30791 11883
rect 31769 11849 31803 11883
rect 32689 11849 32723 11883
rect 33885 11849 33919 11883
rect 36921 11849 36955 11883
rect 37933 11849 37967 11883
rect 38669 11849 38703 11883
rect 12817 11781 12851 11815
rect 14289 11781 14323 11815
rect 19165 11781 19199 11815
rect 19901 11781 19935 11815
rect 19993 11781 20027 11815
rect 24225 11781 24259 11815
rect 39129 11781 39163 11815
rect 45109 11781 45143 11815
rect 49157 11781 49191 11815
rect 1593 11713 1627 11747
rect 2513 11713 2547 11747
rect 15485 11713 15519 11747
rect 19073 11713 19107 11747
rect 21097 11713 21131 11747
rect 21833 11713 21867 11747
rect 22109 11713 22143 11747
rect 22293 11713 22327 11747
rect 22569 11713 22603 11747
rect 26157 11713 26191 11747
rect 27537 11713 27571 11747
rect 31125 11713 31159 11747
rect 37841 11713 37875 11747
rect 39037 11713 39071 11747
rect 39957 11713 39991 11747
rect 40417 11713 40451 11747
rect 47961 11713 47995 11747
rect 2789 11645 2823 11679
rect 12909 11645 12943 11679
rect 13461 11645 13495 11679
rect 14565 11645 14599 11679
rect 15669 11645 15703 11679
rect 16865 11645 16899 11679
rect 17141 11645 17175 11679
rect 20177 11645 20211 11679
rect 21189 11645 21223 11679
rect 21281 11645 21315 11679
rect 23397 11645 23431 11679
rect 23949 11645 23983 11679
rect 27721 11645 27755 11679
rect 28457 11645 28491 11679
rect 28733 11645 28767 11679
rect 31217 11645 31251 11679
rect 31309 11645 31343 11679
rect 32781 11645 32815 11679
rect 32873 11645 32907 11679
rect 33977 11645 34011 11679
rect 34069 11645 34103 11679
rect 35173 11645 35207 11679
rect 35449 11645 35483 11679
rect 38025 11645 38059 11679
rect 39221 11645 39255 11679
rect 1777 11577 1811 11611
rect 16313 11577 16347 11611
rect 19533 11577 19567 11611
rect 20729 11577 20763 11611
rect 27169 11577 27203 11611
rect 40141 11577 40175 11611
rect 45293 11577 45327 11611
rect 12357 11509 12391 11543
rect 13921 11509 13955 11543
rect 15117 11509 15151 11543
rect 18613 11509 18647 11543
rect 30205 11509 30239 11543
rect 32321 11509 32355 11543
rect 33517 11509 33551 11543
rect 37473 11509 37507 11543
rect 2145 11305 2179 11339
rect 13185 11305 13219 11339
rect 14381 11305 14415 11339
rect 16773 11305 16807 11339
rect 19073 11305 19107 11339
rect 19257 11305 19291 11339
rect 19533 11305 19567 11339
rect 20716 11305 20750 11339
rect 28917 11305 28951 11339
rect 29745 11305 29779 11339
rect 38761 11305 38795 11339
rect 39589 11305 39623 11339
rect 1777 11237 1811 11271
rect 12725 11237 12759 11271
rect 15577 11237 15611 11271
rect 22201 11237 22235 11271
rect 23305 11237 23339 11271
rect 26341 11237 26375 11271
rect 28641 11237 28675 11271
rect 29101 11237 29135 11271
rect 29377 11237 29411 11271
rect 38209 11237 38243 11271
rect 40785 11237 40819 11271
rect 10977 11169 11011 11203
rect 14841 11169 14875 11203
rect 14933 11169 14967 11203
rect 16037 11169 16071 11203
rect 16221 11169 16255 11203
rect 17417 11169 17451 11203
rect 18613 11169 18647 11203
rect 20453 11169 20487 11203
rect 23765 11169 23799 11203
rect 23949 11169 23983 11203
rect 24869 11169 24903 11203
rect 27169 11169 27203 11203
rect 30297 11169 30331 11203
rect 31401 11169 31435 11203
rect 32873 11169 32907 11203
rect 34069 11169 34103 11203
rect 35725 11169 35759 11203
rect 49157 11169 49191 11203
rect 1593 11101 1627 11135
rect 2329 11101 2363 11135
rect 13001 11101 13035 11135
rect 14749 11101 14783 11135
rect 17233 11101 17267 11135
rect 18429 11101 18463 11135
rect 24593 11101 24627 11135
rect 26893 11101 26927 11135
rect 31125 11101 31159 11135
rect 33333 11101 33367 11135
rect 34713 11101 34747 11135
rect 37749 11101 37783 11135
rect 38393 11101 38427 11135
rect 40141 11101 40175 11135
rect 40969 11101 41003 11135
rect 45661 11101 45695 11135
rect 47961 11101 47995 11135
rect 11253 11033 11287 11067
rect 13553 11033 13587 11067
rect 15945 11033 15979 11067
rect 17141 11033 17175 11067
rect 19809 11033 19843 11067
rect 23673 11033 23707 11067
rect 30205 11033 30239 11067
rect 30757 11033 30791 11067
rect 36001 11033 36035 11067
rect 40325 11033 40359 11067
rect 45845 11033 45879 11067
rect 17969 10965 18003 10999
rect 18337 10965 18371 10999
rect 22661 10965 22695 10999
rect 30113 10965 30147 10999
rect 1777 10761 1811 10795
rect 12633 10761 12667 10795
rect 13185 10761 13219 10795
rect 14381 10761 14415 10795
rect 15945 10761 15979 10795
rect 17141 10761 17175 10795
rect 18797 10761 18831 10795
rect 19533 10761 19567 10795
rect 19901 10761 19935 10795
rect 21097 10761 21131 10795
rect 24225 10761 24259 10795
rect 27629 10761 27663 10795
rect 28549 10761 28583 10795
rect 31401 10761 31435 10795
rect 32321 10761 32355 10795
rect 33333 10761 33367 10795
rect 36093 10761 36127 10795
rect 14749 10693 14783 10727
rect 17509 10693 17543 10727
rect 21189 10693 21223 10727
rect 28825 10693 28859 10727
rect 29561 10693 29595 10727
rect 37289 10693 37323 10727
rect 49157 10693 49191 10727
rect 1593 10625 1627 10659
rect 2329 10625 2363 10659
rect 2881 10625 2915 10659
rect 13553 10625 13587 10659
rect 13645 10625 13679 10659
rect 14841 10625 14875 10659
rect 16865 10625 16899 10659
rect 18705 10625 18739 10659
rect 24593 10625 24627 10659
rect 25421 10625 25455 10659
rect 26341 10625 26375 10659
rect 27537 10625 27571 10659
rect 30573 10625 30607 10659
rect 32689 10625 32723 10659
rect 33793 10625 33827 10659
rect 36461 10625 36495 10659
rect 39773 10625 39807 10659
rect 40233 10625 40267 10659
rect 47961 10625 47995 10659
rect 3065 10557 3099 10591
rect 12909 10557 12943 10591
rect 13829 10557 13863 10591
rect 14933 10557 14967 10591
rect 16037 10557 16071 10591
rect 16129 10557 16163 10591
rect 17601 10557 17635 10591
rect 17693 10557 17727 10591
rect 18889 10557 18923 10591
rect 19993 10557 20027 10591
rect 20177 10557 20211 10591
rect 21373 10557 21407 10591
rect 22017 10557 22051 10591
rect 22293 10557 22327 10591
rect 24685 10557 24719 10591
rect 24869 10557 24903 10591
rect 27813 10557 27847 10591
rect 30665 10557 30699 10591
rect 30757 10557 30791 10591
rect 32781 10557 32815 10591
rect 32873 10557 32907 10591
rect 34069 10557 34103 10591
rect 36553 10557 36587 10591
rect 36645 10557 36679 10591
rect 2513 10489 2547 10523
rect 27169 10489 27203 10523
rect 35541 10489 35575 10523
rect 39957 10489 39991 10523
rect 15577 10421 15611 10455
rect 18337 10421 18371 10455
rect 20729 10421 20763 10455
rect 23765 10421 23799 10455
rect 25973 10421 26007 10455
rect 26157 10421 26191 10455
rect 26525 10421 26559 10455
rect 26801 10421 26835 10455
rect 30205 10421 30239 10455
rect 31953 10421 31987 10455
rect 12725 10217 12759 10251
rect 16405 10217 16439 10251
rect 18153 10217 18187 10251
rect 26341 10217 26375 10251
rect 32137 10217 32171 10251
rect 32597 10217 32631 10251
rect 36645 10217 36679 10251
rect 36921 10217 36955 10251
rect 13921 10149 13955 10183
rect 23857 10149 23891 10183
rect 26709 10149 26743 10183
rect 28733 10149 28767 10183
rect 1869 10081 1903 10115
rect 13277 10081 13311 10115
rect 16589 10081 16623 10115
rect 17417 10081 17451 10115
rect 17509 10081 17543 10115
rect 18613 10081 18647 10115
rect 18797 10081 18831 10115
rect 19533 10081 19567 10115
rect 20269 10081 20303 10115
rect 23213 10081 23247 10115
rect 23765 10081 23799 10115
rect 24593 10081 24627 10115
rect 29009 10081 29043 10115
rect 29377 10081 29411 10115
rect 29745 10081 29779 10115
rect 33241 10081 33275 10115
rect 34897 10081 34931 10115
rect 35173 10081 35207 10115
rect 49157 10081 49191 10115
rect 1593 10013 1627 10047
rect 13185 10013 13219 10047
rect 14289 10013 14323 10047
rect 22477 10013 22511 10047
rect 26985 10013 27019 10047
rect 30389 10013 30423 10047
rect 38301 10013 38335 10047
rect 38761 10013 38795 10047
rect 40601 10013 40635 10047
rect 44373 10013 44407 10047
rect 46121 10013 46155 10047
rect 47961 10013 47995 10047
rect 14565 9945 14599 9979
rect 20545 9945 20579 9979
rect 24869 9945 24903 9979
rect 27261 9945 27295 9979
rect 30665 9945 30699 9979
rect 32965 9945 32999 9979
rect 33793 9945 33827 9979
rect 40141 9945 40175 9979
rect 40325 9945 40359 9979
rect 44557 9945 44591 9979
rect 47317 9945 47351 9979
rect 12449 9877 12483 9911
rect 13093 9877 13127 9911
rect 16037 9877 16071 9911
rect 16957 9877 16991 9911
rect 17325 9877 17359 9911
rect 18521 9877 18555 9911
rect 22017 9877 22051 9911
rect 24041 9877 24075 9911
rect 33057 9877 33091 9911
rect 38393 9877 38427 9911
rect 2145 9673 2179 9707
rect 21097 9673 21131 9707
rect 22293 9673 22327 9707
rect 31493 9673 31527 9707
rect 31861 9673 31895 9707
rect 32321 9673 32355 9707
rect 35909 9673 35943 9707
rect 12541 9605 12575 9639
rect 12633 9605 12667 9639
rect 15393 9605 15427 9639
rect 18889 9605 18923 9639
rect 19625 9605 19659 9639
rect 21557 9605 21591 9639
rect 22753 9605 22787 9639
rect 23765 9605 23799 9639
rect 27813 9605 27847 9639
rect 32965 9605 32999 9639
rect 34161 9605 34195 9639
rect 49157 9605 49191 9639
rect 1593 9537 1627 9571
rect 2329 9537 2363 9571
rect 16129 9537 16163 9571
rect 16497 9537 16531 9571
rect 22661 9537 22695 9571
rect 23489 9537 23523 9571
rect 26065 9537 26099 9571
rect 26157 9537 26191 9571
rect 33885 9537 33919 9571
rect 47961 9537 47995 9571
rect 12725 9469 12759 9503
rect 13369 9469 13403 9503
rect 13645 9469 13679 9503
rect 16865 9469 16899 9503
rect 17141 9469 17175 9503
rect 19349 9469 19383 9503
rect 22937 9469 22971 9503
rect 26341 9469 26375 9503
rect 27537 9469 27571 9503
rect 29745 9469 29779 9503
rect 30021 9469 30055 9503
rect 33057 9469 33091 9503
rect 33149 9469 33183 9503
rect 1777 9401 1811 9435
rect 15853 9401 15887 9435
rect 29285 9401 29319 9435
rect 35633 9401 35667 9435
rect 12173 9333 12207 9367
rect 15669 9333 15703 9367
rect 16221 9333 16255 9367
rect 21373 9333 21407 9367
rect 21925 9333 21959 9367
rect 25237 9333 25271 9367
rect 25697 9333 25731 9367
rect 32597 9333 32631 9367
rect 1777 9129 1811 9163
rect 14289 9129 14323 9163
rect 21189 9129 21223 9163
rect 24409 9129 24443 9163
rect 24685 9129 24719 9163
rect 25329 9129 25363 9163
rect 25605 9129 25639 9163
rect 28181 9129 28215 9163
rect 32505 9129 32539 9163
rect 32781 9129 32815 9163
rect 33333 9129 33367 9163
rect 36553 9129 36587 9163
rect 2881 8993 2915 9027
rect 15761 8993 15795 9027
rect 16405 8993 16439 9027
rect 18153 8993 18187 9027
rect 18705 8993 18739 9027
rect 19441 8993 19475 9027
rect 22293 8993 22327 9027
rect 22569 8993 22603 9027
rect 28825 8993 28859 9027
rect 30757 8993 30791 9027
rect 33977 8993 34011 9027
rect 35449 8993 35483 9027
rect 49157 8993 49191 9027
rect 2329 8925 2363 8959
rect 3065 8925 3099 8959
rect 14473 8925 14507 8959
rect 14933 8925 14967 8959
rect 15577 8925 15611 8959
rect 15669 8925 15703 8959
rect 33057 8925 33091 8959
rect 33701 8925 33735 8959
rect 36737 8925 36771 8959
rect 37841 8925 37875 8959
rect 39865 8925 39899 8959
rect 47961 8925 47995 8959
rect 1685 8857 1719 8891
rect 16681 8857 16715 8891
rect 19717 8857 19751 8891
rect 28549 8857 28583 8891
rect 29745 8857 29779 8891
rect 31033 8857 31067 8891
rect 35357 8857 35391 8891
rect 39313 8857 39347 8891
rect 39497 8857 39531 8891
rect 2513 8789 2547 8823
rect 15209 8789 15243 8823
rect 21649 8789 21683 8823
rect 24041 8789 24075 8823
rect 24869 8789 24903 8823
rect 25697 8789 25731 8823
rect 27813 8789 27847 8823
rect 28641 8789 28675 8823
rect 30297 8789 30331 8823
rect 33793 8789 33827 8823
rect 34897 8789 34931 8823
rect 35265 8789 35299 8823
rect 37657 8789 37691 8823
rect 15393 8585 15427 8619
rect 18613 8585 18647 8619
rect 21465 8585 21499 8619
rect 24041 8585 24075 8619
rect 30573 8585 30607 8619
rect 34069 8585 34103 8619
rect 34437 8585 34471 8619
rect 37473 8585 37507 8619
rect 40417 8585 40451 8619
rect 13921 8517 13955 8551
rect 17141 8517 17175 8551
rect 22293 8517 22327 8551
rect 29101 8517 29135 8551
rect 44189 8517 44223 8551
rect 49157 8517 49191 8551
rect 1869 8449 1903 8483
rect 13645 8449 13679 8483
rect 16865 8449 16899 8483
rect 19717 8449 19751 8483
rect 22017 8449 22051 8483
rect 31401 8449 31435 8483
rect 32321 8449 32355 8483
rect 37657 8449 37691 8483
rect 39129 8449 39163 8483
rect 40325 8449 40359 8483
rect 40785 8449 40819 8483
rect 45845 8449 45879 8483
rect 47961 8449 47995 8483
rect 1593 8381 1627 8415
rect 19073 8381 19107 8415
rect 19993 8381 20027 8415
rect 28825 8381 28859 8415
rect 31493 8381 31527 8415
rect 31585 8381 31619 8415
rect 32597 8381 32631 8415
rect 46857 8381 46891 8415
rect 15761 8313 15795 8347
rect 23765 8313 23799 8347
rect 31033 8313 31067 8347
rect 38945 8313 38979 8347
rect 44373 8313 44407 8347
rect 2145 8041 2179 8075
rect 15577 8041 15611 8075
rect 21189 8041 21223 8075
rect 22017 8041 22051 8075
rect 31033 8041 31067 8075
rect 37565 8041 37599 8075
rect 17877 7973 17911 8007
rect 17141 7905 17175 7939
rect 17233 7905 17267 7939
rect 18521 7905 18555 7939
rect 19441 7905 19475 7939
rect 22661 7905 22695 7939
rect 29745 7905 29779 7939
rect 30573 7905 30607 7939
rect 31677 7905 31711 7939
rect 32965 7905 32999 7939
rect 49157 7905 49191 7939
rect 1593 7837 1627 7871
rect 2329 7837 2363 7871
rect 15761 7837 15795 7871
rect 17049 7837 17083 7871
rect 22385 7837 22419 7871
rect 38025 7837 38059 7871
rect 47961 7837 47995 7871
rect 18245 7769 18279 7803
rect 18981 7769 19015 7803
rect 19717 7769 19751 7803
rect 30389 7769 30423 7803
rect 31493 7769 31527 7803
rect 32689 7769 32723 7803
rect 38761 7769 38795 7803
rect 38945 7769 38979 7803
rect 1777 7701 1811 7735
rect 16681 7701 16715 7735
rect 18337 7701 18371 7735
rect 21465 7701 21499 7735
rect 21649 7701 21683 7735
rect 22477 7701 22511 7735
rect 23029 7701 23063 7735
rect 30665 7701 30699 7735
rect 31401 7701 31435 7735
rect 32321 7701 32355 7735
rect 32781 7701 32815 7735
rect 38117 7701 38151 7735
rect 39221 7701 39255 7735
rect 18245 7497 18279 7531
rect 18705 7497 18739 7531
rect 22017 7497 22051 7531
rect 22477 7497 22511 7531
rect 23029 7497 23063 7531
rect 30941 7497 30975 7531
rect 32321 7497 32355 7531
rect 21373 7429 21407 7463
rect 22385 7429 22419 7463
rect 37381 7429 37415 7463
rect 37841 7429 37875 7463
rect 44925 7429 44959 7463
rect 49157 7429 49191 7463
rect 1593 7361 1627 7395
rect 2145 7361 2179 7395
rect 38577 7361 38611 7395
rect 39037 7361 39071 7395
rect 47961 7361 47995 7395
rect 22661 7293 22695 7327
rect 1777 7225 1811 7259
rect 38761 7225 38795 7259
rect 45109 7225 45143 7259
rect 21281 7157 21315 7191
rect 21649 7157 21683 7191
rect 32873 7157 32907 7191
rect 37933 7157 37967 7191
rect 49157 6817 49191 6851
rect 2513 6749 2547 6783
rect 2789 6749 2823 6783
rect 17877 6749 17911 6783
rect 19809 6749 19843 6783
rect 46121 6749 46155 6783
rect 47961 6749 47995 6783
rect 1685 6681 1719 6715
rect 1869 6681 1903 6715
rect 47317 6681 47351 6715
rect 2329 6613 2363 6647
rect 17693 6613 17727 6647
rect 19625 6613 19659 6647
rect 2145 6409 2179 6443
rect 44005 6341 44039 6375
rect 49157 6341 49191 6375
rect 1593 6273 1627 6307
rect 2329 6273 2363 6307
rect 18061 6273 18095 6307
rect 37565 6273 37599 6307
rect 47961 6273 47995 6307
rect 18245 6205 18279 6239
rect 1777 6137 1811 6171
rect 38025 6137 38059 6171
rect 44189 6137 44223 6171
rect 18705 6069 18739 6103
rect 37657 6069 37691 6103
rect 2513 5865 2547 5899
rect 3065 5729 3099 5763
rect 49157 5729 49191 5763
rect 1593 5661 1627 5695
rect 2329 5661 2363 5695
rect 2881 5661 2915 5695
rect 43729 5661 43763 5695
rect 47961 5661 47995 5695
rect 43913 5593 43947 5627
rect 1777 5525 1811 5559
rect 38485 5253 38519 5287
rect 38945 5253 38979 5287
rect 49157 5253 49191 5287
rect 18889 5185 18923 5219
rect 37381 5185 37415 5219
rect 37749 5185 37783 5219
rect 45845 5185 45879 5219
rect 47961 5185 47995 5219
rect 1593 5117 1627 5151
rect 1869 5117 1903 5151
rect 19073 5117 19107 5151
rect 46857 5117 46891 5151
rect 38669 5049 38703 5083
rect 19533 4981 19567 5015
rect 37841 4981 37875 5015
rect 2145 4777 2179 4811
rect 36829 4777 36863 4811
rect 46673 4777 46707 4811
rect 20453 4641 20487 4675
rect 21925 4641 21959 4675
rect 25329 4641 25363 4675
rect 25605 4641 25639 4675
rect 47501 4641 47535 4675
rect 49157 4641 49191 4675
rect 1593 4573 1627 4607
rect 2329 4573 2363 4607
rect 20637 4573 20671 4607
rect 22109 4573 22143 4607
rect 23096 4573 23130 4607
rect 25145 4573 25179 4607
rect 37289 4573 37323 4607
rect 38485 4573 38519 4607
rect 47961 4573 47995 4607
rect 22569 4505 22603 4539
rect 38025 4505 38059 4539
rect 38209 4505 38243 4539
rect 46581 4505 46615 4539
rect 47317 4505 47351 4539
rect 1777 4437 1811 4471
rect 21097 4437 21131 4471
rect 23167 4437 23201 4471
rect 37381 4437 37415 4471
rect 46213 4437 46247 4471
rect 1685 4165 1719 4199
rect 27353 4165 27387 4199
rect 2329 4097 2363 4131
rect 3065 4097 3099 4131
rect 22360 4096 22394 4130
rect 22972 4097 23006 4131
rect 23075 4097 23109 4131
rect 23616 4097 23650 4131
rect 45845 4097 45879 4131
rect 47961 4097 47995 4131
rect 49157 4097 49191 4131
rect 24225 4029 24259 4063
rect 24409 4029 24443 4063
rect 25421 4029 25455 4063
rect 27169 4029 27203 4063
rect 27629 4029 27663 4063
rect 46673 4029 46707 4063
rect 2513 3961 2547 3995
rect 23719 3961 23753 3995
rect 1777 3893 1811 3927
rect 2881 3893 2915 3927
rect 22431 3893 22465 3927
rect 47685 3893 47719 3927
rect 23857 3689 23891 3723
rect 23029 3621 23063 3655
rect 24041 3621 24075 3655
rect 1869 3553 1903 3587
rect 24777 3553 24811 3587
rect 25053 3553 25087 3587
rect 36645 3553 36679 3587
rect 49157 3553 49191 3587
rect 1593 3485 1627 3519
rect 16497 3485 16531 3519
rect 21005 3485 21039 3519
rect 23581 3485 23615 3519
rect 24593 3485 24627 3519
rect 36461 3485 36495 3519
rect 36921 3485 36955 3519
rect 46121 3485 46155 3519
rect 47961 3485 47995 3519
rect 21281 3417 21315 3451
rect 45109 3417 45143 3451
rect 45477 3417 45511 3451
rect 47317 3417 47351 3451
rect 16589 3349 16623 3383
rect 22753 3349 22787 3383
rect 45569 3349 45603 3383
rect 2145 3145 2179 3179
rect 16313 3145 16347 3179
rect 21281 3145 21315 3179
rect 16681 3077 16715 3111
rect 24501 3077 24535 3111
rect 49157 3077 49191 3111
rect 1593 3009 1627 3043
rect 2513 3009 2547 3043
rect 14565 3009 14599 3043
rect 17601 3009 17635 3043
rect 18337 3009 18371 3043
rect 20177 3009 20211 3043
rect 20821 3009 20855 3043
rect 21465 3009 21499 3043
rect 22201 3009 22235 3043
rect 23305 3009 23339 3043
rect 26617 3009 26651 3043
rect 27537 3009 27571 3043
rect 28917 3009 28951 3043
rect 44005 3009 44039 3043
rect 45845 3009 45879 3043
rect 47961 3009 47995 3043
rect 14841 2941 14875 2975
rect 18613 2941 18647 2975
rect 24225 2941 24259 2975
rect 25973 2941 26007 2975
rect 29193 2941 29227 2975
rect 31033 2941 31067 2975
rect 45201 2941 45235 2975
rect 46857 2941 46891 2975
rect 1777 2873 1811 2907
rect 17417 2873 17451 2907
rect 19993 2873 20027 2907
rect 20637 2873 20671 2907
rect 22661 2873 22695 2907
rect 2329 2805 2363 2839
rect 2789 2805 2823 2839
rect 22293 2805 22327 2839
rect 23397 2805 23431 2839
rect 23765 2805 23799 2839
rect 26433 2805 26467 2839
rect 27813 2805 27847 2839
rect 27997 2805 28031 2839
rect 30665 2805 30699 2839
rect 3065 2601 3099 2635
rect 9689 2601 9723 2635
rect 26341 2601 26375 2635
rect 29009 2601 29043 2635
rect 32965 2601 32999 2635
rect 35081 2601 35115 2635
rect 1777 2533 1811 2567
rect 18705 2533 18739 2567
rect 19441 2533 19475 2567
rect 30849 2533 30883 2567
rect 2605 2465 2639 2499
rect 12265 2465 12299 2499
rect 14749 2465 14783 2499
rect 17325 2465 17359 2499
rect 20545 2465 20579 2499
rect 22845 2465 22879 2499
rect 25053 2465 25087 2499
rect 27629 2465 27663 2499
rect 37749 2465 37783 2499
rect 41429 2465 41463 2499
rect 43821 2465 43855 2499
rect 49157 2465 49191 2499
rect 1593 2397 1627 2431
rect 3249 2397 3283 2431
rect 9873 2397 9907 2431
rect 10149 2397 10183 2431
rect 11989 2397 12023 2431
rect 14473 2397 14507 2431
rect 17049 2397 17083 2431
rect 18889 2397 18923 2431
rect 19625 2397 19659 2431
rect 20085 2397 20119 2431
rect 22385 2397 22419 2431
rect 24593 2397 24627 2431
rect 27169 2397 27203 2431
rect 29193 2397 29227 2431
rect 29561 2397 29595 2431
rect 31033 2397 31067 2431
rect 31309 2397 31343 2431
rect 33149 2397 33183 2431
rect 33425 2397 33459 2431
rect 35265 2397 35299 2431
rect 35541 2397 35575 2431
rect 37473 2397 37507 2431
rect 40693 2397 40727 2431
rect 43545 2397 43579 2431
rect 45845 2397 45879 2431
rect 47961 2397 47995 2431
rect 2421 2329 2455 2363
rect 47041 2329 47075 2363
rect 3525 2261 3559 2295
rect 37105 2261 37139 2295
rect 43269 2261 43303 2295
<< metal1 >>
rect 30650 26324 30656 26376
rect 30708 26364 30714 26376
rect 40126 26364 40132 26376
rect 30708 26336 40132 26364
rect 30708 26324 30714 26336
rect 40126 26324 40132 26336
rect 40184 26324 40190 26376
rect 3418 25032 3424 25084
rect 3476 25072 3482 25084
rect 10042 25072 10048 25084
rect 3476 25044 10048 25072
rect 3476 25032 3482 25044
rect 10042 25032 10048 25044
rect 10100 25032 10106 25084
rect 29362 25032 29368 25084
rect 29420 25072 29426 25084
rect 40402 25072 40408 25084
rect 29420 25044 40408 25072
rect 29420 25032 29426 25044
rect 40402 25032 40408 25044
rect 40460 25032 40466 25084
rect 31294 24964 31300 25016
rect 31352 25004 31358 25016
rect 42794 25004 42800 25016
rect 31352 24976 42800 25004
rect 31352 24964 31358 24976
rect 42794 24964 42800 24976
rect 42852 24964 42858 25016
rect 4062 24896 4068 24948
rect 4120 24936 4126 24948
rect 8846 24936 8852 24948
rect 4120 24908 8852 24936
rect 4120 24896 4126 24908
rect 8846 24896 8852 24908
rect 8904 24896 8910 24948
rect 29638 24896 29644 24948
rect 29696 24936 29702 24948
rect 44266 24936 44272 24948
rect 29696 24908 44272 24936
rect 29696 24896 29702 24908
rect 44266 24896 44272 24908
rect 44324 24896 44330 24948
rect 25590 24828 25596 24880
rect 25648 24868 25654 24880
rect 48314 24868 48320 24880
rect 25648 24840 48320 24868
rect 25648 24828 25654 24840
rect 48314 24828 48320 24840
rect 48372 24828 48378 24880
rect 25866 24760 25872 24812
rect 25924 24800 25930 24812
rect 35434 24800 35440 24812
rect 25924 24772 35440 24800
rect 25924 24760 25930 24772
rect 35434 24760 35440 24772
rect 35492 24800 35498 24812
rect 37918 24800 37924 24812
rect 35492 24772 37924 24800
rect 35492 24760 35498 24772
rect 37918 24760 37924 24772
rect 37976 24800 37982 24812
rect 40494 24800 40500 24812
rect 37976 24772 40500 24800
rect 37976 24760 37982 24772
rect 40494 24760 40500 24772
rect 40552 24760 40558 24812
rect 16022 24692 16028 24744
rect 16080 24732 16086 24744
rect 24578 24732 24584 24744
rect 16080 24704 24584 24732
rect 16080 24692 16086 24704
rect 24578 24692 24584 24704
rect 24636 24692 24642 24744
rect 27982 24692 27988 24744
rect 28040 24732 28046 24744
rect 29178 24732 29184 24744
rect 28040 24704 29184 24732
rect 28040 24692 28046 24704
rect 29178 24692 29184 24704
rect 29236 24692 29242 24744
rect 34790 24692 34796 24744
rect 34848 24732 34854 24744
rect 38654 24732 38660 24744
rect 34848 24704 38660 24732
rect 34848 24692 34854 24704
rect 38654 24692 38660 24704
rect 38712 24692 38718 24744
rect 17862 24624 17868 24676
rect 17920 24664 17926 24676
rect 23290 24664 23296 24676
rect 17920 24636 23296 24664
rect 17920 24624 17926 24636
rect 23290 24624 23296 24636
rect 23348 24624 23354 24676
rect 23382 24624 23388 24676
rect 23440 24664 23446 24676
rect 26694 24664 26700 24676
rect 23440 24636 26700 24664
rect 23440 24624 23446 24636
rect 26694 24624 26700 24636
rect 26752 24624 26758 24676
rect 29086 24624 29092 24676
rect 29144 24664 29150 24676
rect 29144 24636 31754 24664
rect 29144 24624 29150 24636
rect 3878 24556 3884 24608
rect 3936 24596 3942 24608
rect 6638 24596 6644 24608
rect 3936 24568 6644 24596
rect 3936 24556 3942 24568
rect 6638 24556 6644 24568
rect 6696 24556 6702 24608
rect 17034 24556 17040 24608
rect 17092 24596 17098 24608
rect 24302 24596 24308 24608
rect 17092 24568 24308 24596
rect 17092 24556 17098 24568
rect 24302 24556 24308 24568
rect 24360 24556 24366 24608
rect 24762 24556 24768 24608
rect 24820 24596 24826 24608
rect 30558 24596 30564 24608
rect 24820 24568 30564 24596
rect 24820 24556 24826 24568
rect 30558 24556 30564 24568
rect 30616 24556 30622 24608
rect 31726 24596 31754 24636
rect 31846 24624 31852 24676
rect 31904 24664 31910 24676
rect 40034 24664 40040 24676
rect 31904 24636 40040 24664
rect 31904 24624 31910 24636
rect 40034 24624 40040 24636
rect 40092 24624 40098 24676
rect 32306 24596 32312 24608
rect 31726 24568 32312 24596
rect 32306 24556 32312 24568
rect 32364 24556 32370 24608
rect 34054 24556 34060 24608
rect 34112 24596 34118 24608
rect 39666 24596 39672 24608
rect 34112 24568 39672 24596
rect 34112 24556 34118 24568
rect 39666 24556 39672 24568
rect 39724 24556 39730 24608
rect 1104 24506 49864 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 32950 24506
rect 33002 24454 33014 24506
rect 33066 24454 33078 24506
rect 33130 24454 33142 24506
rect 33194 24454 33206 24506
rect 33258 24454 42950 24506
rect 43002 24454 43014 24506
rect 43066 24454 43078 24506
rect 43130 24454 43142 24506
rect 43194 24454 43206 24506
rect 43258 24454 49864 24506
rect 1104 24432 49864 24454
rect 2774 24352 2780 24404
rect 2832 24392 2838 24404
rect 6178 24392 6184 24404
rect 2832 24364 6184 24392
rect 2832 24352 2838 24364
rect 6178 24352 6184 24364
rect 6236 24352 6242 24404
rect 7742 24352 7748 24404
rect 7800 24392 7806 24404
rect 20714 24392 20720 24404
rect 7800 24364 20720 24392
rect 7800 24352 7806 24364
rect 20714 24352 20720 24364
rect 20772 24352 20778 24404
rect 20824 24364 24532 24392
rect 6730 24324 6736 24336
rect 5828 24296 6736 24324
rect 3237 24259 3295 24265
rect 3237 24225 3249 24259
rect 3283 24256 3295 24259
rect 3510 24256 3516 24268
rect 3283 24228 3516 24256
rect 3283 24225 3295 24228
rect 3237 24219 3295 24225
rect 3510 24216 3516 24228
rect 3568 24216 3574 24268
rect 5828 24265 5856 24296
rect 6730 24284 6736 24296
rect 6788 24284 6794 24336
rect 10134 24324 10140 24336
rect 8128 24296 10140 24324
rect 5813 24259 5871 24265
rect 4172 24228 5764 24256
rect 2225 24191 2283 24197
rect 2225 24157 2237 24191
rect 2271 24188 2283 24191
rect 2314 24188 2320 24200
rect 2271 24160 2320 24188
rect 2271 24157 2283 24160
rect 2225 24151 2283 24157
rect 2314 24148 2320 24160
rect 2372 24148 2378 24200
rect 4172 24197 4200 24228
rect 4157 24191 4215 24197
rect 4157 24157 4169 24191
rect 4203 24157 4215 24191
rect 4157 24151 4215 24157
rect 4617 24191 4675 24197
rect 4617 24157 4629 24191
rect 4663 24157 4675 24191
rect 5736 24188 5764 24228
rect 5813 24225 5825 24259
rect 5859 24225 5871 24259
rect 8128 24256 8156 24296
rect 10134 24284 10140 24296
rect 10192 24284 10198 24336
rect 11882 24324 11888 24336
rect 10980 24296 11888 24324
rect 5813 24219 5871 24225
rect 6656 24228 8156 24256
rect 8205 24259 8263 24265
rect 6656 24188 6684 24228
rect 8205 24225 8217 24259
rect 8251 24256 8263 24259
rect 8662 24256 8668 24268
rect 8251 24228 8668 24256
rect 8251 24225 8263 24228
rect 8205 24219 8263 24225
rect 8662 24216 8668 24228
rect 8720 24216 8726 24268
rect 10980 24265 11008 24296
rect 11882 24284 11888 24296
rect 11940 24284 11946 24336
rect 14918 24324 14924 24336
rect 12406 24296 14924 24324
rect 10965 24259 11023 24265
rect 10965 24225 10977 24259
rect 11011 24225 11023 24259
rect 10965 24219 11023 24225
rect 5736 24160 6684 24188
rect 6733 24191 6791 24197
rect 4617 24151 4675 24157
rect 6733 24157 6745 24191
rect 6779 24157 6791 24191
rect 6733 24151 6791 24157
rect 2130 24080 2136 24132
rect 2188 24120 2194 24132
rect 4632 24120 4660 24151
rect 2188 24092 4660 24120
rect 6748 24120 6776 24151
rect 7374 24148 7380 24200
rect 7432 24148 7438 24200
rect 9309 24191 9367 24197
rect 9309 24157 9321 24191
rect 9355 24157 9367 24191
rect 9309 24151 9367 24157
rect 9953 24191 10011 24197
rect 9953 24157 9965 24191
rect 9999 24188 10011 24191
rect 11885 24191 11943 24197
rect 9999 24160 11100 24188
rect 9999 24157 10011 24160
rect 9953 24151 10011 24157
rect 9324 24120 9352 24151
rect 10870 24120 10876 24132
rect 6748 24092 9260 24120
rect 9324 24092 10876 24120
rect 2188 24080 2194 24092
rect 3973 24055 4031 24061
rect 3973 24021 3985 24055
rect 4019 24052 4031 24055
rect 5534 24052 5540 24064
rect 4019 24024 5540 24052
rect 4019 24021 4031 24024
rect 3973 24015 4031 24021
rect 5534 24012 5540 24024
rect 5592 24012 5598 24064
rect 6549 24055 6607 24061
rect 6549 24021 6561 24055
rect 6595 24052 6607 24055
rect 7466 24052 7472 24064
rect 6595 24024 7472 24052
rect 6595 24021 6607 24024
rect 6549 24015 6607 24021
rect 7466 24012 7472 24024
rect 7524 24012 7530 24064
rect 9122 24012 9128 24064
rect 9180 24012 9186 24064
rect 9232 24052 9260 24092
rect 10870 24080 10876 24092
rect 10928 24080 10934 24132
rect 11072 24120 11100 24160
rect 11885 24157 11897 24191
rect 11931 24188 11943 24191
rect 12406 24188 12434 24296
rect 14918 24284 14924 24296
rect 14976 24284 14982 24336
rect 19610 24324 19616 24336
rect 18708 24296 19616 24324
rect 13541 24259 13599 24265
rect 13541 24225 13553 24259
rect 13587 24256 13599 24259
rect 13814 24256 13820 24268
rect 13587 24228 13820 24256
rect 13587 24225 13599 24228
rect 13541 24219 13599 24225
rect 13814 24216 13820 24228
rect 13872 24216 13878 24268
rect 16117 24259 16175 24265
rect 16117 24225 16129 24259
rect 16163 24256 16175 24259
rect 17678 24256 17684 24268
rect 16163 24228 17684 24256
rect 16163 24225 16175 24228
rect 16117 24219 16175 24225
rect 17678 24216 17684 24228
rect 17736 24216 17742 24268
rect 18708 24265 18736 24296
rect 19610 24284 19616 24296
rect 19668 24284 19674 24336
rect 18693 24259 18751 24265
rect 18693 24225 18705 24259
rect 18739 24225 18751 24259
rect 20824 24256 20852 24364
rect 20990 24284 20996 24336
rect 21048 24324 21054 24336
rect 24026 24324 24032 24336
rect 21048 24296 24032 24324
rect 21048 24284 21054 24296
rect 24026 24284 24032 24296
rect 24084 24284 24090 24336
rect 24504 24324 24532 24364
rect 24578 24352 24584 24404
rect 24636 24352 24642 24404
rect 25958 24352 25964 24404
rect 26016 24352 26022 24404
rect 29733 24395 29791 24401
rect 29733 24392 29745 24395
rect 26068 24364 29745 24392
rect 26068 24324 26096 24364
rect 29733 24361 29745 24364
rect 29779 24361 29791 24395
rect 29733 24355 29791 24361
rect 29914 24352 29920 24404
rect 29972 24392 29978 24404
rect 29972 24364 31800 24392
rect 29972 24352 29978 24364
rect 24504 24296 26096 24324
rect 27246 24284 27252 24336
rect 27304 24324 27310 24336
rect 27893 24327 27951 24333
rect 27893 24324 27905 24327
rect 27304 24296 27905 24324
rect 27304 24284 27310 24296
rect 27893 24293 27905 24296
rect 27939 24293 27951 24327
rect 27893 24287 27951 24293
rect 28626 24284 28632 24336
rect 28684 24324 28690 24336
rect 31478 24324 31484 24336
rect 28684 24296 31484 24324
rect 28684 24284 28690 24296
rect 31478 24284 31484 24296
rect 31536 24324 31542 24336
rect 31665 24327 31723 24333
rect 31665 24324 31677 24327
rect 31536 24296 31677 24324
rect 31536 24284 31542 24296
rect 31665 24293 31677 24296
rect 31711 24293 31723 24327
rect 31772 24324 31800 24364
rect 32306 24352 32312 24404
rect 32364 24352 32370 24404
rect 32398 24352 32404 24404
rect 32456 24392 32462 24404
rect 33597 24395 33655 24401
rect 33597 24392 33609 24395
rect 32456 24364 33609 24392
rect 32456 24352 32462 24364
rect 33597 24361 33609 24364
rect 33643 24361 33655 24395
rect 40310 24392 40316 24404
rect 33597 24355 33655 24361
rect 36556 24364 40316 24392
rect 31772 24296 33180 24324
rect 31665 24287 31723 24293
rect 18693 24219 18751 24225
rect 19628 24228 20852 24256
rect 11931 24160 12434 24188
rect 12529 24191 12587 24197
rect 11931 24157 11943 24160
rect 11885 24151 11943 24157
rect 12529 24157 12541 24191
rect 12575 24188 12587 24191
rect 13722 24188 13728 24200
rect 12575 24160 13728 24188
rect 12575 24157 12587 24160
rect 12529 24151 12587 24157
rect 13722 24148 13728 24160
rect 13780 24148 13786 24200
rect 14366 24148 14372 24200
rect 14424 24188 14430 24200
rect 14461 24191 14519 24197
rect 14461 24188 14473 24191
rect 14424 24160 14473 24188
rect 14424 24148 14430 24160
rect 14461 24157 14473 24160
rect 14507 24157 14519 24191
rect 14461 24151 14519 24157
rect 15105 24191 15163 24197
rect 15105 24157 15117 24191
rect 15151 24157 15163 24191
rect 15105 24151 15163 24157
rect 17589 24191 17647 24197
rect 17589 24157 17601 24191
rect 17635 24188 17647 24191
rect 19334 24188 19340 24200
rect 17635 24160 19340 24188
rect 17635 24157 17647 24160
rect 17589 24151 17647 24157
rect 12618 24120 12624 24132
rect 11072 24092 12624 24120
rect 12618 24080 12624 24092
rect 12676 24080 12682 24132
rect 15120 24120 15148 24151
rect 19334 24148 19340 24160
rect 19392 24148 19398 24200
rect 19628 24197 19656 24228
rect 20898 24216 20904 24268
rect 20956 24216 20962 24268
rect 22465 24259 22523 24265
rect 22465 24256 22477 24259
rect 21100 24228 22477 24256
rect 19613 24191 19671 24197
rect 19613 24157 19625 24191
rect 19659 24157 19671 24191
rect 19613 24151 19671 24157
rect 20257 24191 20315 24197
rect 20257 24157 20269 24191
rect 20303 24157 20315 24191
rect 20257 24151 20315 24157
rect 18414 24120 18420 24132
rect 15120 24092 18420 24120
rect 18414 24080 18420 24092
rect 18472 24080 18478 24132
rect 9766 24052 9772 24064
rect 9232 24024 9772 24052
rect 9766 24012 9772 24024
rect 9824 24012 9830 24064
rect 11698 24012 11704 24064
rect 11756 24012 11762 24064
rect 11790 24012 11796 24064
rect 11848 24052 11854 24064
rect 14277 24055 14335 24061
rect 14277 24052 14289 24055
rect 11848 24024 14289 24052
rect 11848 24012 11854 24024
rect 14277 24021 14289 24024
rect 14323 24021 14335 24055
rect 14277 24015 14335 24021
rect 16853 24055 16911 24061
rect 16853 24021 16865 24055
rect 16899 24052 16911 24055
rect 18506 24052 18512 24064
rect 16899 24024 18512 24052
rect 16899 24021 16911 24024
rect 16853 24015 16911 24021
rect 18506 24012 18512 24024
rect 18564 24012 18570 24064
rect 19426 24012 19432 24064
rect 19484 24012 19490 24064
rect 20272 24052 20300 24151
rect 20530 24148 20536 24200
rect 20588 24188 20594 24200
rect 21100 24188 21128 24228
rect 22465 24225 22477 24228
rect 22511 24225 22523 24259
rect 22465 24219 22523 24225
rect 25225 24259 25283 24265
rect 25225 24225 25237 24259
rect 25271 24225 25283 24259
rect 25225 24219 25283 24225
rect 20588 24160 21128 24188
rect 20588 24148 20594 24160
rect 21266 24148 21272 24200
rect 21324 24188 21330 24200
rect 22005 24191 22063 24197
rect 22005 24188 22017 24191
rect 21324 24160 22017 24188
rect 21324 24148 21330 24160
rect 22005 24157 22017 24160
rect 22051 24157 22063 24191
rect 22005 24151 22063 24157
rect 24029 24191 24087 24197
rect 24029 24157 24041 24191
rect 24075 24188 24087 24191
rect 25038 24188 25044 24200
rect 24075 24160 25044 24188
rect 24075 24157 24087 24160
rect 24029 24151 24087 24157
rect 25038 24148 25044 24160
rect 25096 24148 25102 24200
rect 20438 24080 20444 24132
rect 20496 24120 20502 24132
rect 25240 24120 25268 24219
rect 27338 24216 27344 24268
rect 27396 24256 27402 24268
rect 29181 24259 29239 24265
rect 29181 24256 29193 24259
rect 27396 24228 29193 24256
rect 27396 24216 27402 24228
rect 25866 24148 25872 24200
rect 25924 24148 25930 24200
rect 26050 24148 26056 24200
rect 26108 24188 26114 24200
rect 28736 24197 28764 24228
rect 29181 24225 29193 24228
rect 29227 24225 29239 24259
rect 29181 24219 29239 24225
rect 28077 24191 28135 24197
rect 28077 24188 28089 24191
rect 26108 24160 28089 24188
rect 26108 24148 26114 24160
rect 28077 24157 28089 24160
rect 28123 24157 28135 24191
rect 28077 24151 28135 24157
rect 28721 24191 28779 24197
rect 28721 24157 28733 24191
rect 28767 24157 28779 24191
rect 28721 24151 28779 24157
rect 29917 24191 29975 24197
rect 29917 24157 29929 24191
rect 29963 24188 29975 24191
rect 30098 24188 30104 24200
rect 29963 24160 30104 24188
rect 29963 24157 29975 24160
rect 29917 24151 29975 24157
rect 20496 24092 25268 24120
rect 20496 24080 20502 24092
rect 27154 24080 27160 24132
rect 27212 24120 27218 24132
rect 27249 24123 27307 24129
rect 27249 24120 27261 24123
rect 27212 24092 27261 24120
rect 27212 24080 27218 24092
rect 27249 24089 27261 24092
rect 27295 24089 27307 24123
rect 28092 24120 28120 24151
rect 30098 24148 30104 24160
rect 30156 24148 30162 24200
rect 30558 24148 30564 24200
rect 30616 24188 30622 24200
rect 31110 24188 31116 24200
rect 30616 24160 31116 24188
rect 30616 24148 30622 24160
rect 31110 24148 31116 24160
rect 31168 24148 31174 24200
rect 31205 24191 31263 24197
rect 31205 24157 31217 24191
rect 31251 24188 31263 24191
rect 31478 24188 31484 24200
rect 31251 24160 31484 24188
rect 31251 24157 31263 24160
rect 31205 24151 31263 24157
rect 31478 24148 31484 24160
rect 31536 24148 31542 24200
rect 32122 24148 32128 24200
rect 32180 24188 32186 24200
rect 33152 24197 33180 24296
rect 34422 24284 34428 24336
rect 34480 24324 34486 24336
rect 34480 24296 36492 24324
rect 34480 24284 34486 24296
rect 34054 24216 34060 24268
rect 34112 24216 34118 24268
rect 34241 24259 34299 24265
rect 34241 24225 34253 24259
rect 34287 24256 34299 24259
rect 35342 24256 35348 24268
rect 34287 24228 35348 24256
rect 34287 24225 34299 24228
rect 34241 24219 34299 24225
rect 35342 24216 35348 24228
rect 35400 24216 35406 24268
rect 35526 24216 35532 24268
rect 35584 24216 35590 24268
rect 32493 24191 32551 24197
rect 32493 24188 32505 24191
rect 32180 24160 32505 24188
rect 32180 24148 32186 24160
rect 32493 24157 32505 24160
rect 32539 24157 32551 24191
rect 32493 24151 32551 24157
rect 33137 24191 33195 24197
rect 33137 24157 33149 24191
rect 33183 24188 33195 24191
rect 33965 24191 34023 24197
rect 33183 24160 33732 24188
rect 33183 24157 33195 24160
rect 33137 24151 33195 24157
rect 28997 24123 29055 24129
rect 28997 24120 29009 24123
rect 28092 24092 29009 24120
rect 27249 24083 27307 24089
rect 28997 24089 29009 24092
rect 29043 24089 29055 24123
rect 28997 24083 29055 24089
rect 30742 24080 30748 24132
rect 30800 24120 30806 24132
rect 31849 24123 31907 24129
rect 31849 24120 31861 24123
rect 30800 24092 31861 24120
rect 30800 24080 30806 24092
rect 31849 24089 31861 24092
rect 31895 24120 31907 24123
rect 31938 24120 31944 24132
rect 31895 24092 31944 24120
rect 31895 24089 31907 24092
rect 31849 24083 31907 24089
rect 31938 24080 31944 24092
rect 31996 24080 32002 24132
rect 33704 24120 33732 24160
rect 33965 24157 33977 24191
rect 34011 24188 34023 24191
rect 36078 24188 36084 24200
rect 34011 24160 36084 24188
rect 34011 24157 34023 24160
rect 33965 24151 34023 24157
rect 36078 24148 36084 24160
rect 36136 24148 36142 24200
rect 36464 24188 36492 24296
rect 36556 24265 36584 24364
rect 40310 24352 40316 24364
rect 40368 24352 40374 24404
rect 40494 24352 40500 24404
rect 40552 24392 40558 24404
rect 40862 24392 40868 24404
rect 40552 24364 40868 24392
rect 40552 24352 40558 24364
rect 40862 24352 40868 24364
rect 40920 24392 40926 24404
rect 45373 24395 45431 24401
rect 45373 24392 45385 24395
rect 40920 24364 45385 24392
rect 40920 24352 40926 24364
rect 45373 24361 45385 24364
rect 45419 24361 45431 24395
rect 45373 24355 45431 24361
rect 37461 24327 37519 24333
rect 37461 24293 37473 24327
rect 37507 24324 37519 24327
rect 39114 24324 39120 24336
rect 37507 24296 39120 24324
rect 37507 24293 37519 24296
rect 37461 24287 37519 24293
rect 39114 24284 39120 24296
rect 39172 24284 39178 24336
rect 44637 24327 44695 24333
rect 44637 24324 44649 24327
rect 40236 24296 44649 24324
rect 36541 24259 36599 24265
rect 36541 24225 36553 24259
rect 36587 24225 36599 24259
rect 36541 24219 36599 24225
rect 36725 24259 36783 24265
rect 36725 24225 36737 24259
rect 36771 24256 36783 24259
rect 37366 24256 37372 24268
rect 36771 24228 37372 24256
rect 36771 24225 36783 24228
rect 36725 24219 36783 24225
rect 37366 24216 37372 24228
rect 37424 24216 37430 24268
rect 37918 24216 37924 24268
rect 37976 24216 37982 24268
rect 38105 24259 38163 24265
rect 38105 24225 38117 24259
rect 38151 24256 38163 24259
rect 38286 24256 38292 24268
rect 38151 24228 38292 24256
rect 38151 24225 38163 24228
rect 38105 24219 38163 24225
rect 38286 24216 38292 24228
rect 38344 24216 38350 24268
rect 38657 24191 38715 24197
rect 38657 24188 38669 24191
rect 36464 24160 38669 24188
rect 38657 24157 38669 24160
rect 38703 24157 38715 24191
rect 38657 24151 38715 24157
rect 34146 24120 34152 24132
rect 33704 24092 34152 24120
rect 34146 24080 34152 24092
rect 34204 24080 34210 24132
rect 37734 24120 37740 24132
rect 34900 24092 37740 24120
rect 22554 24052 22560 24064
rect 20272 24024 22560 24052
rect 22554 24012 22560 24024
rect 22612 24012 22618 24064
rect 23845 24055 23903 24061
rect 23845 24021 23857 24055
rect 23891 24052 23903 24055
rect 24670 24052 24676 24064
rect 23891 24024 24676 24052
rect 23891 24021 23903 24024
rect 23845 24015 23903 24021
rect 24670 24012 24676 24024
rect 24728 24012 24734 24064
rect 24946 24012 24952 24064
rect 25004 24012 25010 24064
rect 25041 24055 25099 24061
rect 25041 24021 25053 24055
rect 25087 24052 25099 24055
rect 26142 24052 26148 24064
rect 25087 24024 26148 24052
rect 25087 24021 25099 24024
rect 25041 24015 25099 24021
rect 26142 24012 26148 24024
rect 26200 24012 26206 24064
rect 26234 24012 26240 24064
rect 26292 24052 26298 24064
rect 26329 24055 26387 24061
rect 26329 24052 26341 24055
rect 26292 24024 26341 24052
rect 26292 24012 26298 24024
rect 26329 24021 26341 24024
rect 26375 24021 26387 24055
rect 26329 24015 26387 24021
rect 26418 24012 26424 24064
rect 26476 24052 26482 24064
rect 26697 24055 26755 24061
rect 26697 24052 26709 24055
rect 26476 24024 26709 24052
rect 26476 24012 26482 24024
rect 26697 24021 26709 24024
rect 26743 24021 26755 24055
rect 26697 24015 26755 24021
rect 27338 24012 27344 24064
rect 27396 24012 27402 24064
rect 28537 24055 28595 24061
rect 28537 24021 28549 24055
rect 28583 24052 28595 24055
rect 28626 24052 28632 24064
rect 28583 24024 28632 24052
rect 28583 24021 28595 24024
rect 28537 24015 28595 24021
rect 28626 24012 28632 24024
rect 28684 24012 28690 24064
rect 30374 24012 30380 24064
rect 30432 24012 30438 24064
rect 30926 24012 30932 24064
rect 30984 24052 30990 24064
rect 31021 24055 31079 24061
rect 31021 24052 31033 24055
rect 30984 24024 31033 24052
rect 30984 24012 30990 24024
rect 31021 24021 31033 24024
rect 31067 24021 31079 24055
rect 31021 24015 31079 24021
rect 31110 24012 31116 24064
rect 31168 24052 31174 24064
rect 31481 24055 31539 24061
rect 31481 24052 31493 24055
rect 31168 24024 31493 24052
rect 31168 24012 31174 24024
rect 31481 24021 31493 24024
rect 31527 24021 31539 24055
rect 31481 24015 31539 24021
rect 32950 24012 32956 24064
rect 33008 24012 33014 24064
rect 34900 24061 34928 24092
rect 37734 24080 37740 24092
rect 37792 24080 37798 24132
rect 38672 24120 38700 24151
rect 38930 24148 38936 24200
rect 38988 24148 38994 24200
rect 40126 24148 40132 24200
rect 40184 24188 40190 24200
rect 40236 24197 40264 24296
rect 44637 24293 44649 24296
rect 44683 24293 44695 24327
rect 44637 24287 44695 24293
rect 40678 24216 40684 24268
rect 40736 24216 40742 24268
rect 40954 24216 40960 24268
rect 41012 24216 41018 24268
rect 47486 24216 47492 24268
rect 47544 24256 47550 24268
rect 48222 24256 48228 24268
rect 47544 24228 48228 24256
rect 47544 24216 47550 24228
rect 48222 24216 48228 24228
rect 48280 24256 48286 24268
rect 48501 24259 48559 24265
rect 48501 24256 48513 24259
rect 48280 24228 48513 24256
rect 48280 24216 48286 24228
rect 48501 24225 48513 24228
rect 48547 24225 48559 24259
rect 48501 24219 48559 24225
rect 40221 24191 40279 24197
rect 40221 24188 40233 24191
rect 40184 24160 40233 24188
rect 40184 24148 40190 24160
rect 40221 24157 40233 24160
rect 40267 24157 40279 24191
rect 40696 24188 40724 24216
rect 41322 24188 41328 24200
rect 40696 24160 41328 24188
rect 40221 24151 40279 24157
rect 41322 24148 41328 24160
rect 41380 24148 41386 24200
rect 42150 24148 42156 24200
rect 42208 24188 42214 24200
rect 42613 24191 42671 24197
rect 42613 24188 42625 24191
rect 42208 24160 42625 24188
rect 42208 24148 42214 24160
rect 42613 24157 42625 24160
rect 42659 24188 42671 24191
rect 44634 24188 44640 24200
rect 42659 24160 44640 24188
rect 42659 24157 42671 24160
rect 42613 24151 42671 24157
rect 44634 24148 44640 24160
rect 44692 24148 44698 24200
rect 44726 24148 44732 24200
rect 44784 24188 44790 24200
rect 45278 24188 45284 24200
rect 44784 24160 45284 24188
rect 44784 24148 44790 24160
rect 45278 24148 45284 24160
rect 45336 24148 45342 24200
rect 45554 24148 45560 24200
rect 45612 24188 45618 24200
rect 45925 24191 45983 24197
rect 45925 24188 45937 24191
rect 45612 24160 45937 24188
rect 45612 24148 45618 24160
rect 45925 24157 45937 24160
rect 45971 24188 45983 24191
rect 47213 24191 47271 24197
rect 47213 24188 47225 24191
rect 45971 24160 47225 24188
rect 45971 24157 45983 24160
rect 45925 24151 45983 24157
rect 47213 24157 47225 24160
rect 47259 24157 47271 24191
rect 47213 24151 47271 24157
rect 47302 24148 47308 24200
rect 47360 24188 47366 24200
rect 47765 24191 47823 24197
rect 47765 24188 47777 24191
rect 47360 24160 47777 24188
rect 47360 24148 47366 24160
rect 47765 24157 47777 24160
rect 47811 24157 47823 24191
rect 47765 24151 47823 24157
rect 48774 24148 48780 24200
rect 48832 24148 48838 24200
rect 41782 24120 41788 24132
rect 38672 24092 41788 24120
rect 41782 24080 41788 24092
rect 41840 24080 41846 24132
rect 41877 24123 41935 24129
rect 41877 24089 41889 24123
rect 41923 24120 41935 24123
rect 42242 24120 42248 24132
rect 41923 24092 42248 24120
rect 41923 24089 41935 24092
rect 41877 24083 41935 24089
rect 42242 24080 42248 24092
rect 42300 24080 42306 24132
rect 46014 24080 46020 24132
rect 46072 24120 46078 24132
rect 46750 24120 46756 24132
rect 46072 24092 46756 24120
rect 46072 24080 46078 24092
rect 46750 24080 46756 24092
rect 46808 24080 46814 24132
rect 34885 24055 34943 24061
rect 34885 24021 34897 24055
rect 34931 24021 34943 24055
rect 34885 24015 34943 24021
rect 35250 24012 35256 24064
rect 35308 24012 35314 24064
rect 35345 24055 35403 24061
rect 35345 24021 35357 24055
rect 35391 24052 35403 24055
rect 35434 24052 35440 24064
rect 35391 24024 35440 24052
rect 35391 24021 35403 24024
rect 35345 24015 35403 24021
rect 35434 24012 35440 24024
rect 35492 24012 35498 24064
rect 35986 24012 35992 24064
rect 36044 24052 36050 24064
rect 36081 24055 36139 24061
rect 36081 24052 36093 24055
rect 36044 24024 36093 24052
rect 36044 24012 36050 24024
rect 36081 24021 36093 24024
rect 36127 24021 36139 24055
rect 36081 24015 36139 24021
rect 36170 24012 36176 24064
rect 36228 24052 36234 24064
rect 36449 24055 36507 24061
rect 36449 24052 36461 24055
rect 36228 24024 36461 24052
rect 36228 24012 36234 24024
rect 36449 24021 36461 24024
rect 36495 24021 36507 24055
rect 36449 24015 36507 24021
rect 37642 24012 37648 24064
rect 37700 24052 37706 24064
rect 37829 24055 37887 24061
rect 37829 24052 37841 24055
rect 37700 24024 37841 24052
rect 37700 24012 37706 24024
rect 37829 24021 37841 24024
rect 37875 24021 37887 24055
rect 37829 24015 37887 24021
rect 40037 24055 40095 24061
rect 40037 24021 40049 24055
rect 40083 24052 40095 24055
rect 40494 24052 40500 24064
rect 40083 24024 40500 24052
rect 40083 24021 40095 24024
rect 40037 24015 40095 24021
rect 40494 24012 40500 24024
rect 40552 24012 40558 24064
rect 41966 24012 41972 24064
rect 42024 24012 42030 24064
rect 42150 24012 42156 24064
rect 42208 24012 42214 24064
rect 43901 24055 43959 24061
rect 43901 24021 43913 24055
rect 43947 24052 43959 24055
rect 43990 24052 43996 24064
rect 43947 24024 43996 24052
rect 43947 24021 43959 24024
rect 43901 24015 43959 24021
rect 43990 24012 43996 24024
rect 44048 24012 44054 24064
rect 46106 24012 46112 24064
rect 46164 24012 46170 24064
rect 46198 24012 46204 24064
rect 46256 24052 46262 24064
rect 46845 24055 46903 24061
rect 46845 24052 46857 24055
rect 46256 24024 46857 24052
rect 46256 24012 46262 24024
rect 46845 24021 46857 24024
rect 46891 24021 46903 24055
rect 46845 24015 46903 24021
rect 46934 24012 46940 24064
rect 46992 24052 46998 24064
rect 47949 24055 48007 24061
rect 47949 24052 47961 24055
rect 46992 24024 47961 24052
rect 46992 24012 46998 24024
rect 47949 24021 47961 24024
rect 47995 24021 48007 24055
rect 47949 24015 48007 24021
rect 1104 23962 49864 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 27950 23962
rect 28002 23910 28014 23962
rect 28066 23910 28078 23962
rect 28130 23910 28142 23962
rect 28194 23910 28206 23962
rect 28258 23910 37950 23962
rect 38002 23910 38014 23962
rect 38066 23910 38078 23962
rect 38130 23910 38142 23962
rect 38194 23910 38206 23962
rect 38258 23910 47950 23962
rect 48002 23910 48014 23962
rect 48066 23910 48078 23962
rect 48130 23910 48142 23962
rect 48194 23910 48206 23962
rect 48258 23910 49864 23962
rect 1104 23888 49864 23910
rect 2130 23808 2136 23860
rect 2188 23808 2194 23860
rect 11790 23848 11796 23860
rect 2332 23820 6592 23848
rect 2332 23721 2360 23820
rect 3973 23783 4031 23789
rect 3973 23749 3985 23783
rect 4019 23780 4031 23783
rect 4154 23780 4160 23792
rect 4019 23752 4160 23780
rect 4019 23749 4031 23752
rect 3973 23743 4031 23749
rect 4154 23740 4160 23752
rect 4212 23740 4218 23792
rect 2317 23715 2375 23721
rect 2317 23681 2329 23715
rect 2363 23681 2375 23715
rect 2317 23675 2375 23681
rect 2961 23715 3019 23721
rect 2961 23681 2973 23715
rect 3007 23712 3019 23715
rect 3694 23712 3700 23724
rect 3007 23684 3700 23712
rect 3007 23681 3019 23684
rect 2961 23675 3019 23681
rect 3694 23672 3700 23684
rect 3752 23672 3758 23724
rect 4706 23672 4712 23724
rect 4764 23672 4770 23724
rect 5442 23604 5448 23656
rect 5500 23604 5506 23656
rect 6564 23644 6592 23820
rect 8128 23820 11796 23848
rect 6825 23715 6883 23721
rect 6825 23681 6837 23715
rect 6871 23712 6883 23715
rect 7469 23715 7527 23721
rect 6871 23684 7420 23712
rect 6871 23681 6883 23684
rect 6825 23675 6883 23681
rect 7392 23644 7420 23684
rect 7469 23681 7481 23715
rect 7515 23712 7527 23715
rect 7742 23712 7748 23724
rect 7515 23684 7748 23712
rect 7515 23681 7527 23684
rect 7469 23675 7527 23681
rect 7742 23672 7748 23684
rect 7800 23672 7806 23724
rect 8128 23721 8156 23820
rect 11790 23808 11796 23820
rect 11848 23808 11854 23860
rect 12023 23851 12081 23857
rect 12023 23817 12035 23851
rect 12069 23848 12081 23851
rect 17034 23848 17040 23860
rect 12069 23820 17040 23848
rect 12069 23817 12081 23820
rect 12023 23811 12081 23817
rect 17034 23808 17040 23820
rect 17092 23808 17098 23860
rect 20990 23848 20996 23860
rect 17144 23820 20996 23848
rect 9125 23783 9183 23789
rect 9125 23749 9137 23783
rect 9171 23780 9183 23783
rect 9306 23780 9312 23792
rect 9171 23752 9312 23780
rect 9171 23749 9183 23752
rect 9125 23743 9183 23749
rect 9306 23740 9312 23752
rect 9364 23740 9370 23792
rect 10686 23740 10692 23792
rect 10744 23740 10750 23792
rect 10870 23740 10876 23792
rect 10928 23780 10934 23792
rect 12342 23780 12348 23792
rect 10928 23752 12348 23780
rect 10928 23740 10934 23752
rect 12342 23740 12348 23752
rect 12400 23740 12406 23792
rect 14182 23780 14188 23792
rect 13004 23752 14188 23780
rect 8113 23715 8171 23721
rect 8113 23681 8125 23715
rect 8159 23681 8171 23715
rect 8113 23675 8171 23681
rect 9953 23715 10011 23721
rect 9953 23681 9965 23715
rect 9999 23712 10011 23715
rect 12434 23712 12440 23724
rect 9999 23684 12440 23712
rect 9999 23681 10011 23684
rect 9953 23675 10011 23681
rect 12434 23672 12440 23684
rect 12492 23672 12498 23724
rect 8386 23644 8392 23656
rect 6564 23616 6868 23644
rect 7392 23616 8392 23644
rect 4062 23536 4068 23588
rect 4120 23576 4126 23588
rect 6730 23576 6736 23588
rect 4120 23548 6736 23576
rect 4120 23536 4126 23548
rect 6730 23536 6736 23548
rect 6788 23536 6794 23588
rect 6840 23576 6868 23616
rect 8386 23604 8392 23616
rect 8444 23604 8450 23656
rect 11793 23647 11851 23653
rect 11793 23613 11805 23647
rect 11839 23613 11851 23647
rect 13004 23644 13032 23752
rect 14182 23740 14188 23752
rect 14240 23740 14246 23792
rect 14277 23783 14335 23789
rect 14277 23749 14289 23783
rect 14323 23780 14335 23783
rect 14458 23780 14464 23792
rect 14323 23752 14464 23780
rect 14323 23749 14335 23752
rect 14277 23743 14335 23749
rect 14458 23740 14464 23752
rect 14516 23740 14522 23792
rect 16114 23740 16120 23792
rect 16172 23740 16178 23792
rect 17144 23721 17172 23820
rect 20990 23808 20996 23820
rect 21048 23808 21054 23860
rect 21266 23808 21272 23860
rect 21324 23808 21330 23860
rect 21468 23820 23244 23848
rect 18141 23783 18199 23789
rect 18141 23749 18153 23783
rect 18187 23780 18199 23783
rect 18322 23780 18328 23792
rect 18187 23752 18328 23780
rect 18187 23749 18199 23752
rect 18141 23743 18199 23749
rect 18322 23740 18328 23752
rect 18380 23740 18386 23792
rect 13081 23715 13139 23721
rect 13081 23681 13093 23715
rect 13127 23681 13139 23715
rect 13081 23675 13139 23681
rect 15105 23715 15163 23721
rect 15105 23681 15117 23715
rect 15151 23681 15163 23715
rect 15105 23675 15163 23681
rect 17129 23715 17187 23721
rect 17129 23681 17141 23715
rect 17175 23681 17187 23715
rect 17129 23675 17187 23681
rect 11793 23607 11851 23613
rect 12176 23616 13032 23644
rect 10318 23576 10324 23588
rect 6840 23548 10324 23576
rect 10318 23536 10324 23548
rect 10376 23536 10382 23588
rect 11808 23576 11836 23607
rect 12176 23576 12204 23616
rect 13096 23576 13124 23675
rect 15120 23644 15148 23675
rect 20162 23672 20168 23724
rect 20220 23672 20226 23724
rect 21468 23721 21496 23820
rect 22020 23752 23152 23780
rect 22020 23721 22048 23752
rect 21453 23715 21511 23721
rect 21453 23681 21465 23715
rect 21499 23681 21511 23715
rect 21453 23675 21511 23681
rect 22005 23715 22063 23721
rect 22005 23681 22017 23715
rect 22051 23681 22063 23715
rect 22005 23675 22063 23681
rect 17954 23644 17960 23656
rect 15120 23616 17960 23644
rect 17954 23604 17960 23616
rect 18012 23604 18018 23656
rect 18785 23647 18843 23653
rect 18785 23613 18797 23647
rect 18831 23613 18843 23647
rect 18785 23607 18843 23613
rect 11808 23548 12204 23576
rect 12268 23548 13124 23576
rect 4798 23468 4804 23520
rect 4856 23508 4862 23520
rect 6641 23511 6699 23517
rect 6641 23508 6653 23511
rect 4856 23480 6653 23508
rect 4856 23468 4862 23480
rect 6641 23477 6653 23480
rect 6687 23477 6699 23511
rect 6641 23471 6699 23477
rect 7285 23511 7343 23517
rect 7285 23477 7297 23511
rect 7331 23508 7343 23511
rect 12268 23508 12296 23548
rect 7331 23480 12296 23508
rect 7331 23477 7343 23480
rect 7285 23471 7343 23477
rect 12342 23468 12348 23520
rect 12400 23508 12406 23520
rect 15378 23508 15384 23520
rect 12400 23480 15384 23508
rect 12400 23468 12406 23480
rect 15378 23468 15384 23480
rect 15436 23468 15442 23520
rect 18800 23508 18828 23607
rect 19058 23604 19064 23656
rect 19116 23644 19122 23656
rect 22094 23644 22100 23656
rect 19116 23616 22100 23644
rect 19116 23604 19122 23616
rect 22094 23604 22100 23616
rect 22152 23644 22158 23656
rect 23124 23644 23152 23752
rect 23216 23712 23244 23820
rect 23290 23808 23296 23860
rect 23348 23808 23354 23860
rect 23753 23851 23811 23857
rect 23753 23817 23765 23851
rect 23799 23848 23811 23851
rect 23799 23820 24900 23848
rect 23799 23817 23811 23820
rect 23753 23811 23811 23817
rect 23661 23783 23719 23789
rect 23661 23749 23673 23783
rect 23707 23780 23719 23783
rect 23842 23780 23848 23792
rect 23707 23752 23848 23780
rect 23707 23749 23719 23752
rect 23661 23743 23719 23749
rect 23842 23740 23848 23752
rect 23900 23740 23906 23792
rect 23934 23740 23940 23792
rect 23992 23780 23998 23792
rect 24489 23783 24547 23789
rect 24489 23780 24501 23783
rect 23992 23752 24501 23780
rect 23992 23740 23998 23752
rect 24489 23749 24501 23752
rect 24535 23749 24547 23783
rect 24872 23780 24900 23820
rect 24946 23808 24952 23860
rect 25004 23848 25010 23860
rect 26142 23848 26148 23860
rect 25004 23820 26148 23848
rect 25004 23808 25010 23820
rect 26142 23808 26148 23820
rect 26200 23808 26206 23860
rect 26510 23808 26516 23860
rect 26568 23848 26574 23860
rect 28445 23851 28503 23857
rect 28445 23848 28457 23851
rect 26568 23820 28457 23848
rect 26568 23808 26574 23820
rect 28445 23817 28457 23820
rect 28491 23817 28503 23851
rect 31570 23848 31576 23860
rect 28445 23811 28503 23817
rect 28644 23820 31576 23848
rect 25406 23780 25412 23792
rect 24872 23752 25412 23780
rect 24489 23743 24547 23749
rect 25406 23740 25412 23752
rect 25464 23740 25470 23792
rect 26418 23780 26424 23792
rect 26358 23752 26424 23780
rect 26418 23740 26424 23752
rect 26476 23740 26482 23792
rect 26970 23740 26976 23792
rect 27028 23780 27034 23792
rect 27028 23752 28028 23780
rect 27028 23740 27034 23752
rect 28000 23724 28028 23752
rect 27341 23715 27399 23721
rect 23216 23684 24716 23712
rect 23750 23644 23756 23656
rect 22152 23616 22232 23644
rect 23124 23616 23756 23644
rect 22152 23604 22158 23616
rect 20162 23536 20168 23588
rect 20220 23576 20226 23588
rect 20220 23548 20668 23576
rect 20220 23536 20226 23548
rect 20346 23508 20352 23520
rect 18800 23480 20352 23508
rect 20346 23468 20352 23480
rect 20404 23468 20410 23520
rect 20530 23468 20536 23520
rect 20588 23468 20594 23520
rect 20640 23508 20668 23548
rect 20714 23536 20720 23588
rect 20772 23576 20778 23588
rect 22002 23576 22008 23588
rect 20772 23548 22008 23576
rect 20772 23536 20778 23548
rect 22002 23536 22008 23548
rect 22060 23536 22066 23588
rect 22204 23576 22232 23616
rect 23750 23604 23756 23616
rect 23808 23604 23814 23656
rect 23845 23647 23903 23653
rect 23845 23613 23857 23647
rect 23891 23613 23903 23647
rect 23845 23607 23903 23613
rect 23860 23576 23888 23607
rect 22204 23548 23888 23576
rect 24397 23579 24455 23585
rect 24397 23545 24409 23579
rect 24443 23576 24455 23579
rect 24486 23576 24492 23588
rect 24443 23548 24492 23576
rect 24443 23545 24455 23548
rect 24397 23539 24455 23545
rect 24486 23536 24492 23548
rect 24544 23536 24550 23588
rect 20901 23511 20959 23517
rect 20901 23508 20913 23511
rect 20640 23480 20913 23508
rect 20901 23477 20913 23480
rect 20947 23508 20959 23511
rect 21082 23508 21088 23520
rect 20947 23480 21088 23508
rect 20947 23477 20959 23480
rect 20901 23471 20959 23477
rect 21082 23468 21088 23480
rect 21140 23468 21146 23520
rect 22235 23511 22293 23517
rect 22235 23477 22247 23511
rect 22281 23508 22293 23511
rect 24578 23508 24584 23520
rect 22281 23480 24584 23508
rect 22281 23477 22293 23480
rect 22235 23471 22293 23477
rect 24578 23468 24584 23480
rect 24636 23468 24642 23520
rect 24688 23508 24716 23684
rect 27341 23681 27353 23715
rect 27387 23681 27399 23715
rect 27341 23675 27399 23681
rect 24854 23604 24860 23656
rect 24912 23604 24918 23656
rect 25133 23647 25191 23653
rect 25133 23613 25145 23647
rect 25179 23644 25191 23647
rect 25179 23616 27292 23644
rect 25179 23613 25191 23616
rect 25133 23607 25191 23613
rect 26510 23508 26516 23520
rect 24688 23480 26516 23508
rect 26510 23468 26516 23480
rect 26568 23468 26574 23520
rect 26602 23468 26608 23520
rect 26660 23468 26666 23520
rect 26694 23468 26700 23520
rect 26752 23508 26758 23520
rect 27157 23511 27215 23517
rect 27157 23508 27169 23511
rect 26752 23480 27169 23508
rect 26752 23468 26758 23480
rect 27157 23477 27169 23480
rect 27203 23477 27215 23511
rect 27264 23508 27292 23616
rect 27356 23576 27384 23675
rect 27982 23672 27988 23724
rect 28040 23672 28046 23724
rect 28644 23721 28672 23820
rect 31570 23808 31576 23820
rect 31628 23808 31634 23860
rect 31662 23808 31668 23860
rect 31720 23848 31726 23860
rect 32950 23848 32956 23860
rect 31720 23820 32956 23848
rect 31720 23808 31726 23820
rect 32950 23808 32956 23820
rect 33008 23808 33014 23860
rect 36265 23851 36323 23857
rect 34256 23820 35204 23848
rect 29454 23740 29460 23792
rect 29512 23780 29518 23792
rect 30742 23780 30748 23792
rect 29512 23752 30748 23780
rect 29512 23740 29518 23752
rect 30742 23740 30748 23752
rect 30800 23740 30806 23792
rect 32769 23783 32827 23789
rect 32769 23749 32781 23783
rect 32815 23780 32827 23783
rect 34256 23780 34284 23820
rect 32815 23752 34284 23780
rect 32815 23749 32827 23752
rect 32769 23743 32827 23749
rect 34422 23740 34428 23792
rect 34480 23740 34486 23792
rect 28629 23715 28687 23721
rect 28629 23681 28641 23715
rect 28675 23681 28687 23715
rect 28629 23675 28687 23681
rect 29178 23672 29184 23724
rect 29236 23712 29242 23724
rect 29273 23715 29331 23721
rect 29273 23712 29285 23715
rect 29236 23684 29285 23712
rect 29236 23672 29242 23684
rect 29273 23681 29285 23684
rect 29319 23712 29331 23715
rect 29549 23715 29607 23721
rect 29549 23712 29561 23715
rect 29319 23684 29561 23712
rect 29319 23681 29331 23684
rect 29273 23675 29331 23681
rect 29549 23681 29561 23684
rect 29595 23681 29607 23715
rect 29549 23675 29607 23681
rect 32674 23672 32680 23724
rect 32732 23672 32738 23724
rect 27798 23604 27804 23656
rect 27856 23644 27862 23656
rect 30009 23647 30067 23653
rect 30009 23644 30021 23647
rect 27856 23616 30021 23644
rect 27856 23604 27862 23616
rect 30009 23613 30021 23616
rect 30055 23613 30067 23647
rect 30009 23607 30067 23613
rect 30285 23647 30343 23653
rect 30285 23613 30297 23647
rect 30331 23644 30343 23647
rect 30650 23644 30656 23656
rect 30331 23616 30656 23644
rect 30331 23613 30343 23616
rect 30285 23607 30343 23613
rect 29730 23576 29736 23588
rect 27356 23548 29736 23576
rect 29730 23536 29736 23548
rect 29788 23536 29794 23588
rect 27614 23508 27620 23520
rect 27264 23480 27620 23508
rect 27157 23471 27215 23477
rect 27614 23468 27620 23480
rect 27672 23468 27678 23520
rect 27706 23468 27712 23520
rect 27764 23508 27770 23520
rect 27801 23511 27859 23517
rect 27801 23508 27813 23511
rect 27764 23480 27813 23508
rect 27764 23468 27770 23480
rect 27801 23477 27813 23480
rect 27847 23477 27859 23511
rect 27801 23471 27859 23477
rect 29089 23511 29147 23517
rect 29089 23477 29101 23511
rect 29135 23508 29147 23511
rect 29178 23508 29184 23520
rect 29135 23480 29184 23508
rect 29135 23477 29147 23480
rect 29089 23471 29147 23477
rect 29178 23468 29184 23480
rect 29236 23468 29242 23520
rect 30024 23508 30052 23607
rect 30650 23604 30656 23616
rect 30708 23644 30714 23656
rect 32582 23644 32588 23656
rect 30708 23616 32588 23644
rect 30708 23604 30714 23616
rect 32582 23604 32588 23616
rect 32640 23604 32646 23656
rect 32953 23647 33011 23653
rect 32953 23613 32965 23647
rect 32999 23613 33011 23647
rect 32953 23607 33011 23613
rect 31570 23536 31576 23588
rect 31628 23576 31634 23588
rect 32309 23579 32367 23585
rect 32309 23576 32321 23579
rect 31628 23548 32321 23576
rect 31628 23536 31634 23548
rect 32309 23545 32321 23548
rect 32355 23545 32367 23579
rect 32309 23539 32367 23545
rect 31386 23508 31392 23520
rect 30024 23480 31392 23508
rect 31386 23468 31392 23480
rect 31444 23468 31450 23520
rect 31754 23468 31760 23520
rect 31812 23468 31818 23520
rect 32968 23508 32996 23607
rect 33594 23604 33600 23656
rect 33652 23604 33658 23656
rect 33873 23647 33931 23653
rect 33873 23613 33885 23647
rect 33919 23644 33931 23647
rect 34330 23644 34336 23656
rect 33919 23616 34336 23644
rect 33919 23613 33931 23616
rect 33873 23607 33931 23613
rect 34330 23604 34336 23616
rect 34388 23604 34394 23656
rect 35176 23576 35204 23820
rect 36265 23817 36277 23851
rect 36311 23848 36323 23851
rect 38841 23851 38899 23857
rect 38841 23848 38853 23851
rect 36311 23820 38853 23848
rect 36311 23817 36323 23820
rect 36265 23811 36323 23817
rect 38841 23817 38853 23820
rect 38887 23817 38899 23851
rect 38841 23811 38899 23817
rect 39209 23851 39267 23857
rect 39209 23817 39221 23851
rect 39255 23848 39267 23851
rect 44174 23848 44180 23860
rect 39255 23820 44180 23848
rect 39255 23817 39267 23820
rect 39209 23811 39267 23817
rect 44174 23808 44180 23820
rect 44232 23808 44238 23860
rect 45278 23808 45284 23860
rect 45336 23848 45342 23860
rect 45649 23851 45707 23857
rect 45649 23848 45661 23851
rect 45336 23820 45661 23848
rect 45336 23808 45342 23820
rect 45649 23817 45661 23820
rect 45695 23817 45707 23851
rect 48225 23851 48283 23857
rect 48225 23848 48237 23851
rect 45649 23811 45707 23817
rect 46768 23820 48237 23848
rect 35342 23740 35348 23792
rect 35400 23780 35406 23792
rect 37550 23780 37556 23792
rect 35400 23752 37556 23780
rect 35400 23740 35406 23752
rect 37550 23740 37556 23752
rect 37608 23740 37614 23792
rect 37734 23740 37740 23792
rect 37792 23780 37798 23792
rect 37921 23783 37979 23789
rect 37921 23780 37933 23783
rect 37792 23752 37933 23780
rect 37792 23740 37798 23752
rect 37921 23749 37933 23752
rect 37967 23749 37979 23783
rect 37921 23743 37979 23749
rect 38378 23740 38384 23792
rect 38436 23780 38442 23792
rect 38436 23752 40724 23780
rect 38436 23740 38442 23752
rect 35802 23672 35808 23724
rect 35860 23712 35866 23724
rect 36909 23715 36967 23721
rect 36909 23712 36921 23715
rect 35860 23684 36921 23712
rect 35860 23672 35866 23684
rect 36909 23681 36921 23684
rect 36955 23681 36967 23715
rect 36909 23675 36967 23681
rect 37458 23672 37464 23724
rect 37516 23672 37522 23724
rect 37829 23715 37887 23721
rect 37829 23681 37841 23715
rect 37875 23712 37887 23715
rect 40034 23712 40040 23724
rect 37875 23684 40040 23712
rect 37875 23681 37887 23684
rect 37829 23675 37887 23681
rect 40034 23672 40040 23684
rect 40092 23672 40098 23724
rect 40126 23672 40132 23724
rect 40184 23712 40190 23724
rect 40221 23715 40279 23721
rect 40221 23712 40233 23715
rect 40184 23684 40233 23712
rect 40184 23672 40190 23684
rect 40221 23681 40233 23684
rect 40267 23712 40279 23715
rect 40586 23712 40592 23724
rect 40267 23684 40592 23712
rect 40267 23681 40279 23684
rect 40221 23675 40279 23681
rect 40586 23672 40592 23684
rect 40644 23672 40650 23724
rect 40696 23721 40724 23752
rect 40770 23740 40776 23792
rect 40828 23780 40834 23792
rect 41969 23783 42027 23789
rect 41969 23780 41981 23783
rect 40828 23752 41981 23780
rect 40828 23740 40834 23752
rect 41969 23749 41981 23752
rect 42015 23749 42027 23783
rect 41969 23743 42027 23749
rect 42426 23740 42432 23792
rect 42484 23780 42490 23792
rect 46768 23780 46796 23820
rect 48225 23817 48237 23820
rect 48271 23817 48283 23851
rect 48225 23811 48283 23817
rect 42484 23752 46796 23780
rect 42484 23740 42490 23752
rect 46842 23740 46848 23792
rect 46900 23780 46906 23792
rect 47305 23783 47363 23789
rect 47305 23780 47317 23783
rect 46900 23752 47317 23780
rect 46900 23740 46906 23752
rect 47305 23749 47317 23752
rect 47351 23749 47363 23783
rect 47305 23743 47363 23749
rect 40681 23715 40739 23721
rect 40681 23681 40693 23715
rect 40727 23712 40739 23715
rect 42150 23712 42156 23724
rect 40727 23684 42156 23712
rect 40727 23681 40739 23684
rect 40681 23675 40739 23681
rect 42150 23672 42156 23684
rect 42208 23672 42214 23724
rect 42794 23672 42800 23724
rect 42852 23712 42858 23724
rect 42889 23715 42947 23721
rect 42889 23712 42901 23715
rect 42852 23684 42901 23712
rect 42852 23672 42858 23684
rect 42889 23681 42901 23684
rect 42935 23681 42947 23715
rect 42889 23675 42947 23681
rect 44177 23715 44235 23721
rect 44177 23681 44189 23715
rect 44223 23712 44235 23715
rect 44266 23712 44272 23724
rect 44223 23684 44272 23712
rect 44223 23681 44235 23684
rect 44177 23675 44235 23681
rect 44266 23672 44272 23684
rect 44324 23672 44330 23724
rect 45370 23672 45376 23724
rect 45428 23672 45434 23724
rect 46293 23715 46351 23721
rect 46293 23681 46305 23715
rect 46339 23681 46351 23715
rect 46293 23675 46351 23681
rect 36354 23604 36360 23656
rect 36412 23604 36418 23656
rect 36446 23604 36452 23656
rect 36504 23604 36510 23656
rect 37476 23644 37504 23672
rect 38013 23647 38071 23653
rect 38013 23644 38025 23647
rect 37476 23616 38025 23644
rect 38013 23613 38025 23616
rect 38059 23613 38071 23647
rect 38013 23607 38071 23613
rect 39298 23604 39304 23656
rect 39356 23604 39362 23656
rect 39390 23604 39396 23656
rect 39448 23604 39454 23656
rect 40402 23604 40408 23656
rect 40460 23644 40466 23656
rect 40957 23647 41015 23653
rect 40957 23644 40969 23647
rect 40460 23616 40969 23644
rect 40460 23604 40466 23616
rect 40957 23613 40969 23616
rect 41003 23613 41015 23647
rect 40957 23607 41015 23613
rect 41782 23604 41788 23656
rect 41840 23604 41846 23656
rect 42610 23604 42616 23656
rect 42668 23604 42674 23656
rect 43898 23604 43904 23656
rect 43956 23604 43962 23656
rect 46308 23644 46336 23675
rect 46750 23672 46756 23724
rect 46808 23712 46814 23724
rect 47581 23715 47639 23721
rect 47581 23712 47593 23715
rect 46808 23684 47593 23712
rect 46808 23672 46814 23684
rect 47581 23681 47593 23684
rect 47627 23681 47639 23715
rect 47581 23675 47639 23681
rect 47854 23672 47860 23724
rect 47912 23712 47918 23724
rect 48041 23715 48099 23721
rect 48041 23712 48053 23715
rect 47912 23684 48053 23712
rect 47912 23672 47918 23684
rect 48041 23681 48053 23684
rect 48087 23681 48099 23715
rect 48041 23675 48099 23681
rect 48590 23672 48596 23724
rect 48648 23712 48654 23724
rect 48777 23715 48835 23721
rect 48777 23712 48789 23715
rect 48648 23684 48789 23712
rect 48648 23672 48654 23684
rect 48777 23681 48789 23684
rect 48823 23681 48835 23715
rect 48777 23675 48835 23681
rect 46474 23644 46480 23656
rect 46308 23616 46480 23644
rect 46474 23604 46480 23616
rect 46532 23644 46538 23656
rect 48406 23644 48412 23656
rect 46532 23616 48412 23644
rect 46532 23604 46538 23616
rect 48406 23604 48412 23616
rect 48464 23604 48470 23656
rect 37461 23579 37519 23585
rect 37461 23576 37473 23579
rect 35176 23548 37473 23576
rect 37461 23545 37473 23548
rect 37507 23545 37519 23579
rect 37461 23539 37519 23545
rect 37642 23536 37648 23588
rect 37700 23576 37706 23588
rect 38470 23576 38476 23588
rect 37700 23548 38476 23576
rect 37700 23536 37706 23548
rect 38470 23536 38476 23548
rect 38528 23536 38534 23588
rect 39316 23576 39344 23604
rect 42426 23576 42432 23588
rect 39316 23548 41414 23576
rect 34974 23508 34980 23520
rect 32968 23480 34980 23508
rect 34974 23468 34980 23480
rect 35032 23508 35038 23520
rect 35345 23511 35403 23517
rect 35345 23508 35357 23511
rect 35032 23480 35357 23508
rect 35032 23468 35038 23480
rect 35345 23477 35357 23480
rect 35391 23477 35403 23511
rect 35345 23471 35403 23477
rect 35894 23468 35900 23520
rect 35952 23468 35958 23520
rect 37274 23468 37280 23520
rect 37332 23508 37338 23520
rect 38378 23508 38384 23520
rect 37332 23480 38384 23508
rect 37332 23468 37338 23480
rect 38378 23468 38384 23480
rect 38436 23468 38442 23520
rect 38654 23468 38660 23520
rect 38712 23508 38718 23520
rect 40037 23511 40095 23517
rect 40037 23508 40049 23511
rect 38712 23480 40049 23508
rect 38712 23468 38718 23480
rect 40037 23477 40049 23480
rect 40083 23477 40095 23511
rect 41386 23508 41414 23548
rect 42168 23548 42432 23576
rect 41598 23508 41604 23520
rect 41386 23480 41604 23508
rect 40037 23471 40095 23477
rect 41598 23468 41604 23480
rect 41656 23508 41662 23520
rect 42168 23517 42196 23548
rect 42426 23536 42432 23548
rect 42484 23536 42490 23588
rect 45186 23536 45192 23588
rect 45244 23536 45250 23588
rect 47029 23579 47087 23585
rect 47029 23576 47041 23579
rect 45296 23548 47041 23576
rect 42153 23511 42211 23517
rect 42153 23508 42165 23511
rect 41656 23480 42165 23508
rect 41656 23468 41662 23480
rect 42153 23477 42165 23480
rect 42199 23477 42211 23511
rect 42153 23471 42211 23477
rect 42242 23468 42248 23520
rect 42300 23508 42306 23520
rect 45296 23508 45324 23548
rect 47029 23545 47041 23548
rect 47075 23545 47087 23579
rect 47029 23539 47087 23545
rect 42300 23480 45324 23508
rect 42300 23468 42306 23480
rect 45370 23468 45376 23520
rect 45428 23508 45434 23520
rect 46109 23511 46167 23517
rect 46109 23508 46121 23511
rect 45428 23480 46121 23508
rect 45428 23468 45434 23480
rect 46109 23477 46121 23480
rect 46155 23477 46167 23511
rect 46109 23471 46167 23477
rect 47118 23468 47124 23520
rect 47176 23508 47182 23520
rect 48961 23511 49019 23517
rect 48961 23508 48973 23511
rect 47176 23480 48973 23508
rect 47176 23468 47182 23480
rect 48961 23477 48973 23480
rect 49007 23477 49019 23511
rect 48961 23471 49019 23477
rect 49142 23468 49148 23520
rect 49200 23508 49206 23520
rect 49421 23511 49479 23517
rect 49421 23508 49433 23511
rect 49200 23480 49433 23508
rect 49200 23468 49206 23480
rect 49421 23477 49433 23480
rect 49467 23477 49479 23511
rect 49421 23471 49479 23477
rect 1104 23418 49864 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 32950 23418
rect 33002 23366 33014 23418
rect 33066 23366 33078 23418
rect 33130 23366 33142 23418
rect 33194 23366 33206 23418
rect 33258 23366 42950 23418
rect 43002 23366 43014 23418
rect 43066 23366 43078 23418
rect 43130 23366 43142 23418
rect 43194 23366 43206 23418
rect 43258 23366 49864 23418
rect 1104 23344 49864 23366
rect 2866 23264 2872 23316
rect 2924 23304 2930 23316
rect 4338 23304 4344 23316
rect 2924 23276 4344 23304
rect 2924 23264 2930 23276
rect 4338 23264 4344 23276
rect 4396 23264 4402 23316
rect 4706 23264 4712 23316
rect 4764 23264 4770 23316
rect 14182 23264 14188 23316
rect 14240 23304 14246 23316
rect 14240 23276 16252 23304
rect 14240 23264 14246 23276
rect 15838 23236 15844 23248
rect 9876 23208 15844 23236
rect 1578 23128 1584 23180
rect 1636 23168 1642 23180
rect 4430 23168 4436 23180
rect 1636 23140 4436 23168
rect 1636 23128 1642 23140
rect 4430 23128 4436 23140
rect 4488 23128 4494 23180
rect 6086 23128 6092 23180
rect 6144 23128 6150 23180
rect 7834 23128 7840 23180
rect 7892 23128 7898 23180
rect 9876 23177 9904 23208
rect 15838 23196 15844 23208
rect 15896 23196 15902 23248
rect 9861 23171 9919 23177
rect 9861 23137 9873 23171
rect 9907 23137 9919 23171
rect 9861 23131 9919 23137
rect 11238 23128 11244 23180
rect 11296 23128 11302 23180
rect 13354 23128 13360 23180
rect 13412 23128 13418 23180
rect 14844 23140 15700 23168
rect 1765 23103 1823 23109
rect 1765 23069 1777 23103
rect 1811 23100 1823 23103
rect 4249 23103 4307 23109
rect 1811 23072 4200 23100
rect 1811 23069 1823 23072
rect 1765 23063 1823 23069
rect 2774 22992 2780 23044
rect 2832 22992 2838 23044
rect 3602 22924 3608 22976
rect 3660 22964 3666 22976
rect 4065 22967 4123 22973
rect 4065 22964 4077 22967
rect 3660 22936 4077 22964
rect 3660 22924 3666 22936
rect 4065 22933 4077 22936
rect 4111 22933 4123 22967
rect 4172 22964 4200 23072
rect 4249 23069 4261 23103
rect 4295 23100 4307 23103
rect 4522 23100 4528 23112
rect 4295 23072 4528 23100
rect 4295 23069 4307 23072
rect 4249 23063 4307 23069
rect 4522 23060 4528 23072
rect 4580 23060 4586 23112
rect 4893 23103 4951 23109
rect 4893 23069 4905 23103
rect 4939 23069 4951 23103
rect 4893 23063 4951 23069
rect 4908 23032 4936 23063
rect 5074 23060 5080 23112
rect 5132 23100 5138 23112
rect 5353 23103 5411 23109
rect 5353 23100 5365 23103
rect 5132 23072 5365 23100
rect 5132 23060 5138 23072
rect 5353 23069 5365 23072
rect 5399 23069 5411 23103
rect 5353 23063 5411 23069
rect 5534 23060 5540 23112
rect 5592 23100 5598 23112
rect 7193 23103 7251 23109
rect 7193 23100 7205 23103
rect 5592 23072 7205 23100
rect 5592 23060 5598 23072
rect 7193 23069 7205 23072
rect 7239 23069 7251 23103
rect 7193 23063 7251 23069
rect 9122 23060 9128 23112
rect 9180 23100 9186 23112
rect 9217 23103 9275 23109
rect 9217 23100 9229 23103
rect 9180 23072 9229 23100
rect 9180 23060 9186 23072
rect 9217 23069 9229 23072
rect 9263 23069 9275 23103
rect 9217 23063 9275 23069
rect 10689 23103 10747 23109
rect 10689 23069 10701 23103
rect 10735 23100 10747 23103
rect 12342 23100 12348 23112
rect 10735 23072 12348 23100
rect 10735 23069 10747 23072
rect 10689 23063 10747 23069
rect 12342 23060 12348 23072
rect 12400 23060 12406 23112
rect 12529 23103 12587 23109
rect 12529 23069 12541 23103
rect 12575 23100 12587 23103
rect 13906 23100 13912 23112
rect 12575 23072 13912 23100
rect 12575 23069 12587 23072
rect 12529 23063 12587 23069
rect 13906 23060 13912 23072
rect 13964 23060 13970 23112
rect 14844 23109 14872 23140
rect 14829 23103 14887 23109
rect 14829 23069 14841 23103
rect 14875 23069 14887 23103
rect 14829 23063 14887 23069
rect 15473 23103 15531 23109
rect 15473 23069 15485 23103
rect 15519 23069 15531 23103
rect 15473 23063 15531 23069
rect 7742 23032 7748 23044
rect 4908 23004 7748 23032
rect 7742 22992 7748 23004
rect 7800 22992 7806 23044
rect 6914 22964 6920 22976
rect 4172 22936 6920 22964
rect 4065 22927 4123 22933
rect 6914 22924 6920 22936
rect 6972 22924 6978 22976
rect 7006 22924 7012 22976
rect 7064 22964 7070 22976
rect 9309 22967 9367 22973
rect 9309 22964 9321 22967
rect 7064 22936 9321 22964
rect 7064 22924 7070 22936
rect 9309 22933 9321 22936
rect 9355 22933 9367 22967
rect 9309 22927 9367 22933
rect 14642 22924 14648 22976
rect 14700 22924 14706 22976
rect 15488 22964 15516 23063
rect 15672 23032 15700 23140
rect 15746 23128 15752 23180
rect 15804 23128 15810 23180
rect 16224 23168 16252 23276
rect 17954 23264 17960 23316
rect 18012 23304 18018 23316
rect 19797 23307 19855 23313
rect 19797 23304 19809 23307
rect 18012 23276 19809 23304
rect 18012 23264 18018 23276
rect 19797 23273 19809 23276
rect 19843 23273 19855 23307
rect 22830 23304 22836 23316
rect 19797 23267 19855 23273
rect 19904 23276 22836 23304
rect 19904 23236 19932 23276
rect 22830 23264 22836 23276
rect 22888 23264 22894 23316
rect 23750 23304 23756 23316
rect 23216 23276 23756 23304
rect 18432 23208 19932 23236
rect 20272 23208 20484 23236
rect 18432 23168 18460 23208
rect 19334 23168 19340 23180
rect 16224 23140 18460 23168
rect 18524 23140 19340 23168
rect 17034 23060 17040 23112
rect 17092 23100 17098 23112
rect 17129 23103 17187 23109
rect 17129 23100 17141 23103
rect 17092 23072 17141 23100
rect 17092 23060 17098 23072
rect 17129 23069 17141 23072
rect 17175 23069 17187 23103
rect 18524 23086 18552 23140
rect 19334 23128 19340 23140
rect 19392 23168 19398 23180
rect 20162 23168 20168 23180
rect 19392 23140 20168 23168
rect 19392 23128 19398 23140
rect 20162 23128 20168 23140
rect 20220 23128 20226 23180
rect 17129 23063 17187 23069
rect 19242 23060 19248 23112
rect 19300 23100 19306 23112
rect 20272 23100 20300 23208
rect 20346 23128 20352 23180
rect 20404 23128 20410 23180
rect 20456 23168 20484 23208
rect 22002 23196 22008 23248
rect 22060 23196 22066 23248
rect 22094 23196 22100 23248
rect 22152 23196 22158 23248
rect 23216 23236 23244 23276
rect 23750 23264 23756 23276
rect 23808 23264 23814 23316
rect 24026 23264 24032 23316
rect 24084 23304 24090 23316
rect 24765 23307 24823 23313
rect 24765 23304 24777 23307
rect 24084 23276 24777 23304
rect 24084 23264 24090 23276
rect 24765 23273 24777 23276
rect 24811 23273 24823 23307
rect 24765 23267 24823 23273
rect 25222 23264 25228 23316
rect 25280 23264 25286 23316
rect 25406 23264 25412 23316
rect 25464 23304 25470 23316
rect 27893 23307 27951 23313
rect 27893 23304 27905 23307
rect 25464 23276 27905 23304
rect 25464 23264 25470 23276
rect 27893 23273 27905 23276
rect 27939 23273 27951 23307
rect 27893 23267 27951 23273
rect 27982 23264 27988 23316
rect 28040 23304 28046 23316
rect 28997 23307 29055 23313
rect 28997 23304 29009 23307
rect 28040 23276 29009 23304
rect 28040 23264 28046 23276
rect 28997 23273 29009 23276
rect 29043 23273 29055 23307
rect 28997 23267 29055 23273
rect 29730 23264 29736 23316
rect 29788 23264 29794 23316
rect 32122 23304 32128 23316
rect 31036 23276 32128 23304
rect 22296 23208 23244 23236
rect 22020 23168 22048 23196
rect 22296 23168 22324 23208
rect 24578 23196 24584 23248
rect 24636 23236 24642 23248
rect 25498 23236 25504 23248
rect 24636 23208 25504 23236
rect 24636 23196 24642 23208
rect 25498 23196 25504 23208
rect 25556 23196 25562 23248
rect 27522 23196 27528 23248
rect 27580 23236 27586 23248
rect 27580 23208 29224 23236
rect 27580 23196 27586 23208
rect 22833 23171 22891 23177
rect 22833 23168 22845 23171
rect 20456 23140 21956 23168
rect 22020 23140 22324 23168
rect 22388 23140 22845 23168
rect 19300 23072 20300 23100
rect 19300 23060 19306 23072
rect 17310 23032 17316 23044
rect 15672 23004 17316 23032
rect 17310 22992 17316 23004
rect 17368 22992 17374 23044
rect 17402 22992 17408 23044
rect 17460 22992 17466 23044
rect 19702 22992 19708 23044
rect 19760 22992 19766 23044
rect 20625 23035 20683 23041
rect 20625 23001 20637 23035
rect 20671 23032 20683 23035
rect 20714 23032 20720 23044
rect 20671 23004 20720 23032
rect 20671 23001 20683 23004
rect 20625 22995 20683 23001
rect 20714 22992 20720 23004
rect 20772 22992 20778 23044
rect 21082 22992 21088 23044
rect 21140 22992 21146 23044
rect 21928 23032 21956 23140
rect 22002 23060 22008 23112
rect 22060 23100 22066 23112
rect 22388 23100 22416 23140
rect 22833 23137 22845 23140
rect 22879 23137 22891 23171
rect 22833 23131 22891 23137
rect 23937 23171 23995 23177
rect 23937 23137 23949 23171
rect 23983 23168 23995 23171
rect 25961 23171 26019 23177
rect 25961 23168 25973 23171
rect 23983 23140 25973 23168
rect 23983 23137 23995 23140
rect 23937 23131 23995 23137
rect 25961 23137 25973 23140
rect 26007 23168 26019 23171
rect 26602 23168 26608 23180
rect 26007 23140 26608 23168
rect 26007 23137 26019 23140
rect 25961 23131 26019 23137
rect 26602 23128 26608 23140
rect 26660 23128 26666 23180
rect 26694 23128 26700 23180
rect 26752 23168 26758 23180
rect 28445 23171 28503 23177
rect 28445 23168 28457 23171
rect 26752 23140 28457 23168
rect 26752 23128 26758 23140
rect 28445 23137 28457 23140
rect 28491 23137 28503 23171
rect 29196 23168 29224 23208
rect 29270 23196 29276 23248
rect 29328 23236 29334 23248
rect 31036 23245 31064 23276
rect 32122 23264 32128 23276
rect 32180 23264 32186 23316
rect 33137 23307 33195 23313
rect 33137 23273 33149 23307
rect 33183 23304 33195 23307
rect 33962 23304 33968 23316
rect 33183 23276 33968 23304
rect 33183 23273 33195 23276
rect 33137 23267 33195 23273
rect 33962 23264 33968 23276
rect 34020 23264 34026 23316
rect 35066 23264 35072 23316
rect 35124 23304 35130 23316
rect 37274 23304 37280 23316
rect 35124 23276 37280 23304
rect 35124 23264 35130 23276
rect 37274 23264 37280 23276
rect 37332 23264 37338 23316
rect 37550 23264 37556 23316
rect 37608 23304 37614 23316
rect 39025 23307 39083 23313
rect 39025 23304 39037 23307
rect 37608 23276 39037 23304
rect 37608 23264 37614 23276
rect 39025 23273 39037 23276
rect 39071 23273 39083 23307
rect 39025 23267 39083 23273
rect 40034 23264 40040 23316
rect 40092 23264 40098 23316
rect 40218 23264 40224 23316
rect 40276 23304 40282 23316
rect 40862 23304 40868 23316
rect 40276 23276 40868 23304
rect 40276 23264 40282 23276
rect 40862 23264 40868 23276
rect 40920 23264 40926 23316
rect 42794 23304 42800 23316
rect 41616 23276 42800 23304
rect 31021 23239 31079 23245
rect 31021 23236 31033 23239
rect 29328 23208 31033 23236
rect 29328 23196 29334 23208
rect 31021 23205 31033 23208
rect 31067 23205 31079 23239
rect 31021 23199 31079 23205
rect 31312 23208 31524 23236
rect 29454 23168 29460 23180
rect 29196 23140 29460 23168
rect 28445 23131 28503 23137
rect 29454 23128 29460 23140
rect 29512 23128 29518 23180
rect 30190 23128 30196 23180
rect 30248 23128 30254 23180
rect 30377 23171 30435 23177
rect 30377 23137 30389 23171
rect 30423 23137 30435 23171
rect 30377 23131 30435 23137
rect 22060 23072 22416 23100
rect 23661 23103 23719 23109
rect 22060 23060 22066 23072
rect 23661 23069 23673 23103
rect 23707 23100 23719 23103
rect 24394 23100 24400 23112
rect 23707 23072 24400 23100
rect 23707 23069 23719 23072
rect 23661 23063 23719 23069
rect 24394 23060 24400 23072
rect 24452 23060 24458 23112
rect 25314 23100 25320 23112
rect 24596 23072 25320 23100
rect 22649 23035 22707 23041
rect 21928 23004 22416 23032
rect 17494 22964 17500 22976
rect 15488 22936 17500 22964
rect 17494 22924 17500 22936
rect 17552 22924 17558 22976
rect 18874 22924 18880 22976
rect 18932 22924 18938 22976
rect 20530 22924 20536 22976
rect 20588 22964 20594 22976
rect 22278 22964 22284 22976
rect 20588 22936 22284 22964
rect 20588 22924 20594 22936
rect 22278 22924 22284 22936
rect 22336 22924 22342 22976
rect 22388 22964 22416 23004
rect 22649 23001 22661 23035
rect 22695 23032 22707 23035
rect 24596 23032 24624 23072
rect 25314 23060 25320 23072
rect 25372 23060 25378 23112
rect 25682 23060 25688 23112
rect 25740 23060 25746 23112
rect 27614 23060 27620 23112
rect 27672 23100 27678 23112
rect 28534 23100 28540 23112
rect 27672 23072 28540 23100
rect 27672 23060 27678 23072
rect 28534 23060 28540 23072
rect 28592 23060 28598 23112
rect 22695 23004 24624 23032
rect 22695 23001 22707 23004
rect 22649 22995 22707 23001
rect 24670 22992 24676 23044
rect 24728 22992 24734 23044
rect 26418 22992 26424 23044
rect 26476 22992 26482 23044
rect 28442 23032 28448 23044
rect 27448 23004 28448 23032
rect 23293 22967 23351 22973
rect 23293 22964 23305 22967
rect 22388 22936 23305 22964
rect 23293 22933 23305 22936
rect 23339 22933 23351 22967
rect 23293 22927 23351 22933
rect 23753 22967 23811 22973
rect 23753 22933 23765 22967
rect 23799 22964 23811 22967
rect 24486 22964 24492 22976
rect 23799 22936 24492 22964
rect 23799 22933 23811 22936
rect 23753 22927 23811 22933
rect 24486 22924 24492 22936
rect 24544 22924 24550 22976
rect 25130 22924 25136 22976
rect 25188 22964 25194 22976
rect 27448 22973 27476 23004
rect 28442 22992 28448 23004
rect 28500 22992 28506 23044
rect 30392 23032 30420 23131
rect 31312 23032 31340 23208
rect 31386 23128 31392 23180
rect 31444 23128 31450 23180
rect 31496 23168 31524 23208
rect 34974 23196 34980 23248
rect 35032 23236 35038 23248
rect 35032 23208 35204 23236
rect 35032 23196 35038 23208
rect 31754 23168 31760 23180
rect 31496 23140 31760 23168
rect 31754 23128 31760 23140
rect 31812 23128 31818 23180
rect 33686 23128 33692 23180
rect 33744 23168 33750 23180
rect 35066 23168 35072 23180
rect 33744 23140 35072 23168
rect 33744 23128 33750 23140
rect 35066 23128 35072 23140
rect 35124 23128 35130 23180
rect 35176 23168 35204 23208
rect 39206 23196 39212 23248
rect 39264 23236 39270 23248
rect 41616 23236 41644 23276
rect 42794 23264 42800 23276
rect 42852 23264 42858 23316
rect 44634 23264 44640 23316
rect 44692 23304 44698 23316
rect 44729 23307 44787 23313
rect 44729 23304 44741 23307
rect 44692 23276 44741 23304
rect 44692 23264 44698 23276
rect 44729 23273 44741 23276
rect 44775 23273 44787 23307
rect 44729 23267 44787 23273
rect 45462 23264 45468 23316
rect 45520 23304 45526 23316
rect 45649 23307 45707 23313
rect 45649 23304 45661 23307
rect 45520 23276 45661 23304
rect 45520 23264 45526 23276
rect 45649 23273 45661 23276
rect 45695 23273 45707 23307
rect 45649 23267 45707 23273
rect 46293 23307 46351 23313
rect 46293 23273 46305 23307
rect 46339 23304 46351 23307
rect 47762 23304 47768 23316
rect 46339 23276 47768 23304
rect 46339 23273 46351 23276
rect 46293 23267 46351 23273
rect 47762 23264 47768 23276
rect 47820 23264 47826 23316
rect 39264 23208 41644 23236
rect 39264 23196 39270 23208
rect 43898 23196 43904 23248
rect 43956 23236 43962 23248
rect 45189 23239 45247 23245
rect 45189 23236 45201 23239
rect 43956 23208 45201 23236
rect 43956 23196 43962 23208
rect 45189 23205 45201 23208
rect 45235 23205 45247 23239
rect 47029 23239 47087 23245
rect 47029 23236 47041 23239
rect 45189 23199 45247 23205
rect 45526 23208 47041 23236
rect 35345 23171 35403 23177
rect 35345 23168 35357 23171
rect 35176 23140 35357 23168
rect 35345 23137 35357 23140
rect 35391 23137 35403 23171
rect 35345 23131 35403 23137
rect 37274 23128 37280 23180
rect 37332 23168 37338 23180
rect 37332 23140 38792 23168
rect 37332 23128 37338 23140
rect 33873 23103 33931 23109
rect 33873 23100 33885 23103
rect 33060 23072 33885 23100
rect 31665 23035 31723 23041
rect 31665 23032 31677 23035
rect 29012 23004 30328 23032
rect 30392 23004 31677 23032
rect 27433 22967 27491 22973
rect 27433 22964 27445 22967
rect 25188 22936 27445 22964
rect 25188 22924 25194 22936
rect 27433 22933 27445 22936
rect 27479 22933 27491 22967
rect 27433 22927 27491 22933
rect 28258 22924 28264 22976
rect 28316 22924 28322 22976
rect 28353 22967 28411 22973
rect 28353 22933 28365 22967
rect 28399 22964 28411 22967
rect 29012 22964 29040 23004
rect 28399 22936 29040 22964
rect 29181 22967 29239 22973
rect 28399 22933 28411 22936
rect 28353 22927 28411 22933
rect 29181 22933 29193 22967
rect 29227 22964 29239 22967
rect 29454 22964 29460 22976
rect 29227 22936 29460 22964
rect 29227 22933 29239 22936
rect 29181 22927 29239 22933
rect 29454 22924 29460 22936
rect 29512 22924 29518 22976
rect 30098 22924 30104 22976
rect 30156 22924 30162 22976
rect 30300 22964 30328 23004
rect 31665 23001 31677 23004
rect 31711 23001 31723 23035
rect 31665 22995 31723 23001
rect 31938 22992 31944 23044
rect 31996 23032 32002 23044
rect 31996 23004 32154 23032
rect 31996 22992 32002 23004
rect 31018 22964 31024 22976
rect 30300 22936 31024 22964
rect 31018 22924 31024 22936
rect 31076 22924 31082 22976
rect 31110 22924 31116 22976
rect 31168 22964 31174 22976
rect 33060 22964 33088 23072
rect 33873 23069 33885 23072
rect 33919 23100 33931 23103
rect 34333 23103 34391 23109
rect 34333 23100 34345 23103
rect 33919 23072 34345 23100
rect 33919 23069 33931 23072
rect 33873 23063 33931 23069
rect 34333 23069 34345 23072
rect 34379 23069 34391 23103
rect 38764 23100 38792 23140
rect 38838 23128 38844 23180
rect 38896 23168 38902 23180
rect 40589 23171 40647 23177
rect 40589 23168 40601 23171
rect 38896 23140 40601 23168
rect 38896 23128 38902 23140
rect 40589 23137 40601 23140
rect 40635 23137 40647 23171
rect 40589 23131 40647 23137
rect 41141 23171 41199 23177
rect 41141 23137 41153 23171
rect 41187 23168 41199 23171
rect 41414 23168 41420 23180
rect 41187 23140 41420 23168
rect 41187 23137 41199 23140
rect 41141 23131 41199 23137
rect 41414 23128 41420 23140
rect 41472 23128 41478 23180
rect 41785 23171 41843 23177
rect 41785 23137 41797 23171
rect 41831 23168 41843 23171
rect 45526 23168 45554 23208
rect 47029 23205 47041 23208
rect 47075 23205 47087 23239
rect 47029 23199 47087 23205
rect 47670 23196 47676 23248
rect 47728 23196 47734 23248
rect 41831 23140 45554 23168
rect 41831 23137 41843 23140
rect 41785 23131 41843 23137
rect 46474 23128 46480 23180
rect 46532 23128 46538 23180
rect 46753 23171 46811 23177
rect 46753 23137 46765 23171
rect 46799 23168 46811 23171
rect 49234 23168 49240 23180
rect 46799 23140 49240 23168
rect 46799 23137 46811 23140
rect 46753 23131 46811 23137
rect 41509 23103 41567 23109
rect 41509 23100 41521 23103
rect 38764 23072 41521 23100
rect 34333 23063 34391 23069
rect 41509 23069 41521 23072
rect 41555 23069 41567 23103
rect 41509 23063 41567 23069
rect 42886 23060 42892 23112
rect 42944 23100 42950 23112
rect 43990 23100 43996 23112
rect 42944 23072 43996 23100
rect 42944 23060 42950 23072
rect 43990 23060 43996 23072
rect 44048 23060 44054 23112
rect 44082 23060 44088 23112
rect 44140 23100 44146 23112
rect 47228 23109 47256 23140
rect 49234 23128 49240 23140
rect 49292 23128 49298 23180
rect 44269 23103 44327 23109
rect 44269 23100 44281 23103
rect 44140 23072 44281 23100
rect 44140 23060 44146 23072
rect 44269 23069 44281 23072
rect 44315 23100 44327 23103
rect 45373 23103 45431 23109
rect 45373 23100 45385 23103
rect 44315 23072 45385 23100
rect 44315 23069 44327 23072
rect 44269 23063 44327 23069
rect 45373 23069 45385 23072
rect 45419 23069 45431 23103
rect 45373 23063 45431 23069
rect 47213 23103 47271 23109
rect 47213 23069 47225 23103
rect 47259 23069 47271 23103
rect 47213 23063 47271 23069
rect 47854 23060 47860 23112
rect 47912 23060 47918 23112
rect 48314 23060 48320 23112
rect 48372 23060 48378 23112
rect 49053 23103 49111 23109
rect 49053 23069 49065 23103
rect 49099 23100 49111 23103
rect 49326 23100 49332 23112
rect 49099 23072 49332 23100
rect 49099 23069 49111 23072
rect 49053 23063 49111 23069
rect 49326 23060 49332 23072
rect 49384 23060 49390 23112
rect 33594 22992 33600 23044
rect 33652 23032 33658 23044
rect 34149 23035 34207 23041
rect 34149 23032 34161 23035
rect 33652 23004 34161 23032
rect 33652 22992 33658 23004
rect 34149 23001 34161 23004
rect 34195 23032 34207 23035
rect 34422 23032 34428 23044
rect 34195 23004 34428 23032
rect 34195 23001 34207 23004
rect 34149 22995 34207 23001
rect 34422 22992 34428 23004
rect 34480 23032 34486 23044
rect 34701 23035 34759 23041
rect 34701 23032 34713 23035
rect 34480 23004 34713 23032
rect 34480 22992 34486 23004
rect 34701 23001 34713 23004
rect 34747 23032 34759 23035
rect 35802 23032 35808 23044
rect 34747 23004 35808 23032
rect 34747 23001 34759 23004
rect 34701 22995 34759 23001
rect 35802 22992 35808 23004
rect 35860 22992 35866 23044
rect 37553 23035 37611 23041
rect 37553 23001 37565 23035
rect 37599 23032 37611 23035
rect 37826 23032 37832 23044
rect 37599 23004 37832 23032
rect 37599 23001 37611 23004
rect 37553 22995 37611 23001
rect 37826 22992 37832 23004
rect 37884 22992 37890 23044
rect 40497 23035 40555 23041
rect 38778 23004 39436 23032
rect 31168 22936 33088 22964
rect 33689 22967 33747 22973
rect 31168 22924 31174 22936
rect 33689 22933 33701 22967
rect 33735 22964 33747 22967
rect 33778 22964 33784 22976
rect 33735 22936 33784 22964
rect 33735 22933 33747 22936
rect 33689 22927 33747 22933
rect 33778 22924 33784 22936
rect 33836 22924 33842 22976
rect 33870 22924 33876 22976
rect 33928 22964 33934 22976
rect 34790 22964 34796 22976
rect 33928 22936 34796 22964
rect 33928 22924 33934 22936
rect 34790 22924 34796 22936
rect 34848 22964 34854 22976
rect 34974 22964 34980 22976
rect 34848 22936 34980 22964
rect 34848 22924 34854 22936
rect 34974 22924 34980 22936
rect 35032 22924 35038 22976
rect 35250 22924 35256 22976
rect 35308 22964 35314 22976
rect 36817 22967 36875 22973
rect 36817 22964 36829 22967
rect 35308 22936 36829 22964
rect 35308 22924 35314 22936
rect 36817 22933 36829 22936
rect 36863 22964 36875 22967
rect 38838 22964 38844 22976
rect 36863 22936 38844 22964
rect 36863 22933 36875 22936
rect 36817 22927 36875 22933
rect 38838 22924 38844 22936
rect 38896 22924 38902 22976
rect 39408 22973 39436 23004
rect 40497 23001 40509 23035
rect 40543 23032 40555 23035
rect 40543 23004 41184 23032
rect 40543 23001 40555 23004
rect 40497 22995 40555 23001
rect 39393 22967 39451 22973
rect 39393 22933 39405 22967
rect 39439 22964 39451 22967
rect 39574 22964 39580 22976
rect 39439 22936 39580 22964
rect 39439 22933 39451 22936
rect 39393 22927 39451 22933
rect 39574 22924 39580 22936
rect 39632 22924 39638 22976
rect 40402 22924 40408 22976
rect 40460 22924 40466 22976
rect 41156 22964 41184 23004
rect 41230 22992 41236 23044
rect 41288 23032 41294 23044
rect 42058 23032 42064 23044
rect 41288 23004 42064 23032
rect 41288 22992 41294 23004
rect 42058 22992 42064 23004
rect 42116 22992 42122 23044
rect 43530 22992 43536 23044
rect 43588 22992 43594 23044
rect 44008 23032 44036 23060
rect 45005 23035 45063 23041
rect 45005 23032 45017 23035
rect 44008 23004 45017 23032
rect 45005 23001 45017 23004
rect 45051 23001 45063 23035
rect 45005 22995 45063 23001
rect 46109 23035 46167 23041
rect 46109 23001 46121 23035
rect 46155 23032 46167 23035
rect 48332 23032 48360 23060
rect 48590 23032 48596 23044
rect 46155 23004 48360 23032
rect 48424 23004 48596 23032
rect 46155 23001 46167 23004
rect 46109 22995 46167 23001
rect 42150 22964 42156 22976
rect 41156 22936 42156 22964
rect 42150 22924 42156 22936
rect 42208 22924 42214 22976
rect 42610 22924 42616 22976
rect 42668 22964 42674 22976
rect 43809 22967 43867 22973
rect 43809 22964 43821 22967
rect 42668 22936 43821 22964
rect 42668 22924 42674 22936
rect 43809 22933 43821 22936
rect 43855 22933 43867 22967
rect 43809 22927 43867 22933
rect 43990 22924 43996 22976
rect 44048 22964 44054 22976
rect 44361 22967 44419 22973
rect 44361 22964 44373 22967
rect 44048 22936 44373 22964
rect 44048 22924 44054 22936
rect 44361 22933 44373 22936
rect 44407 22933 44419 22967
rect 44361 22927 44419 22933
rect 45925 22967 45983 22973
rect 45925 22933 45937 22967
rect 45971 22964 45983 22967
rect 48424 22964 48452 23004
rect 48590 22992 48596 23004
rect 48648 22992 48654 23044
rect 45971 22936 48452 22964
rect 45971 22933 45983 22936
rect 45925 22927 45983 22933
rect 48498 22924 48504 22976
rect 48556 22924 48562 22976
rect 49234 22924 49240 22976
rect 49292 22924 49298 22976
rect 1104 22874 49864 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 27950 22874
rect 28002 22822 28014 22874
rect 28066 22822 28078 22874
rect 28130 22822 28142 22874
rect 28194 22822 28206 22874
rect 28258 22822 37950 22874
rect 38002 22822 38014 22874
rect 38066 22822 38078 22874
rect 38130 22822 38142 22874
rect 38194 22822 38206 22874
rect 38258 22822 47950 22874
rect 48002 22822 48014 22874
rect 48066 22822 48078 22874
rect 48130 22822 48142 22874
rect 48194 22822 48206 22874
rect 48258 22822 49864 22874
rect 1104 22800 49864 22822
rect 4062 22720 4068 22772
rect 4120 22760 4126 22772
rect 5534 22760 5540 22772
rect 4120 22732 5540 22760
rect 4120 22720 4126 22732
rect 5534 22720 5540 22732
rect 5592 22720 5598 22772
rect 11054 22720 11060 22772
rect 11112 22760 11118 22772
rect 12250 22760 12256 22772
rect 11112 22732 12256 22760
rect 11112 22720 11118 22732
rect 12250 22720 12256 22732
rect 12308 22720 12314 22772
rect 12710 22720 12716 22772
rect 12768 22760 12774 22772
rect 13538 22760 13544 22772
rect 12768 22732 13544 22760
rect 12768 22720 12774 22732
rect 13538 22720 13544 22732
rect 13596 22720 13602 22772
rect 17402 22720 17408 22772
rect 17460 22760 17466 22772
rect 18601 22763 18659 22769
rect 18601 22760 18613 22763
rect 17460 22732 18613 22760
rect 17460 22720 17466 22732
rect 18601 22729 18613 22732
rect 18647 22760 18659 22763
rect 20438 22760 20444 22772
rect 18647 22732 20444 22760
rect 18647 22729 18659 22732
rect 18601 22723 18659 22729
rect 20438 22720 20444 22732
rect 20496 22720 20502 22772
rect 23753 22763 23811 22769
rect 21560 22732 22416 22760
rect 15286 22692 15292 22704
rect 2746 22664 15292 22692
rect 1765 22627 1823 22633
rect 1765 22593 1777 22627
rect 1811 22624 1823 22627
rect 2746 22624 2774 22664
rect 15286 22652 15292 22664
rect 15344 22652 15350 22704
rect 17034 22692 17040 22704
rect 16868 22664 17040 22692
rect 1811 22596 2774 22624
rect 3973 22627 4031 22633
rect 1811 22593 1823 22596
rect 1765 22587 1823 22593
rect 3973 22593 3985 22627
rect 4019 22593 4031 22627
rect 3973 22587 4031 22593
rect 2777 22559 2835 22565
rect 2777 22525 2789 22559
rect 2823 22556 2835 22559
rect 2866 22556 2872 22568
rect 2823 22528 2872 22556
rect 2823 22525 2835 22528
rect 2777 22519 2835 22525
rect 2866 22516 2872 22528
rect 2924 22516 2930 22568
rect 3988 22420 4016 22587
rect 4798 22584 4804 22636
rect 4856 22584 4862 22636
rect 6825 22627 6883 22633
rect 6825 22593 6837 22627
rect 6871 22593 6883 22627
rect 6825 22587 6883 22593
rect 4982 22516 4988 22568
rect 5040 22556 5046 22568
rect 5077 22559 5135 22565
rect 5077 22556 5089 22559
rect 5040 22528 5089 22556
rect 5040 22516 5046 22528
rect 5077 22525 5089 22528
rect 5123 22525 5135 22559
rect 6840 22556 6868 22587
rect 7466 22584 7472 22636
rect 7524 22584 7530 22636
rect 9953 22627 10011 22633
rect 7576 22596 9904 22624
rect 7576 22556 7604 22596
rect 6840 22528 7604 22556
rect 5077 22519 5135 22525
rect 7650 22516 7656 22568
rect 7708 22556 7714 22568
rect 7929 22559 7987 22565
rect 7929 22556 7941 22559
rect 7708 22528 7941 22556
rect 7708 22516 7714 22528
rect 7929 22525 7941 22528
rect 7975 22525 7987 22559
rect 7929 22519 7987 22525
rect 4154 22448 4160 22500
rect 4212 22448 4218 22500
rect 6641 22491 6699 22497
rect 6641 22457 6653 22491
rect 6687 22488 6699 22491
rect 9122 22488 9128 22500
rect 6687 22460 9128 22488
rect 6687 22457 6699 22460
rect 6641 22451 6699 22457
rect 9122 22448 9128 22460
rect 9180 22448 9186 22500
rect 9876 22488 9904 22596
rect 9953 22593 9965 22627
rect 9999 22624 10011 22627
rect 11698 22624 11704 22636
rect 9999 22596 11704 22624
rect 9999 22593 10011 22596
rect 9953 22587 10011 22593
rect 11698 22584 11704 22596
rect 11756 22584 11762 22636
rect 11793 22627 11851 22633
rect 11793 22593 11805 22627
rect 11839 22624 11851 22627
rect 12710 22624 12716 22636
rect 11839 22596 12716 22624
rect 11839 22593 11851 22596
rect 11793 22587 11851 22593
rect 12710 22584 12716 22596
rect 12768 22584 12774 22636
rect 12805 22627 12863 22633
rect 12805 22593 12817 22627
rect 12851 22624 12863 22627
rect 14642 22624 14648 22636
rect 12851 22596 14648 22624
rect 12851 22593 12863 22596
rect 12805 22587 12863 22593
rect 14642 22584 14648 22596
rect 14700 22584 14706 22636
rect 15013 22627 15071 22633
rect 15013 22593 15025 22627
rect 15059 22624 15071 22627
rect 16666 22624 16672 22636
rect 15059 22596 16672 22624
rect 15059 22593 15071 22596
rect 15013 22587 15071 22593
rect 16666 22584 16672 22596
rect 16724 22584 16730 22636
rect 16868 22633 16896 22664
rect 17034 22652 17040 22664
rect 17092 22652 17098 22704
rect 18782 22652 18788 22704
rect 18840 22692 18846 22704
rect 19705 22695 19763 22701
rect 19705 22692 19717 22695
rect 18840 22664 19717 22692
rect 18840 22652 18846 22664
rect 19705 22661 19717 22664
rect 19751 22661 19763 22695
rect 21082 22692 21088 22704
rect 20930 22664 21088 22692
rect 19705 22655 19763 22661
rect 21082 22652 21088 22664
rect 21140 22692 21146 22704
rect 21560 22701 21588 22732
rect 21545 22695 21603 22701
rect 21545 22692 21557 22695
rect 21140 22664 21557 22692
rect 21140 22652 21146 22664
rect 21545 22661 21557 22664
rect 21591 22661 21603 22695
rect 21545 22655 21603 22661
rect 22278 22652 22284 22704
rect 22336 22652 22342 22704
rect 22388 22692 22416 22732
rect 23753 22729 23765 22763
rect 23799 22760 23811 22763
rect 24210 22760 24216 22772
rect 23799 22732 24216 22760
rect 23799 22729 23811 22732
rect 23753 22723 23811 22729
rect 24210 22720 24216 22732
rect 24268 22720 24274 22772
rect 24302 22720 24308 22772
rect 24360 22760 24366 22772
rect 24397 22763 24455 22769
rect 24397 22760 24409 22763
rect 24360 22732 24409 22760
rect 24360 22720 24366 22732
rect 24397 22729 24409 22732
rect 24443 22729 24455 22763
rect 24397 22723 24455 22729
rect 24412 22692 24440 22723
rect 24854 22720 24860 22772
rect 24912 22760 24918 22772
rect 27798 22760 27804 22772
rect 24912 22732 27804 22760
rect 24912 22720 24918 22732
rect 27798 22720 27804 22732
rect 27856 22720 27862 22772
rect 28736 22732 30696 22760
rect 25038 22692 25044 22704
rect 22388 22664 22770 22692
rect 24412 22664 25044 22692
rect 25038 22652 25044 22664
rect 25096 22652 25102 22704
rect 25130 22652 25136 22704
rect 25188 22652 25194 22704
rect 26418 22692 26424 22704
rect 26358 22664 26424 22692
rect 26418 22652 26424 22664
rect 26476 22692 26482 22704
rect 27522 22692 27528 22704
rect 26476 22664 27528 22692
rect 26476 22652 26482 22664
rect 27522 22652 27528 22664
rect 27580 22692 27586 22704
rect 27617 22695 27675 22701
rect 27617 22692 27629 22695
rect 27580 22664 27629 22692
rect 27580 22652 27586 22664
rect 27617 22661 27629 22664
rect 27663 22661 27675 22695
rect 27617 22655 27675 22661
rect 28350 22652 28356 22704
rect 28408 22692 28414 22704
rect 28736 22692 28764 22732
rect 28408 22664 28764 22692
rect 30668 22692 30696 22732
rect 30742 22720 30748 22772
rect 30800 22720 30806 22772
rect 31202 22720 31208 22772
rect 31260 22760 31266 22772
rect 31386 22760 31392 22772
rect 31260 22732 31392 22760
rect 31260 22720 31266 22732
rect 31386 22720 31392 22732
rect 31444 22720 31450 22772
rect 31478 22720 31484 22772
rect 31536 22720 31542 22772
rect 35986 22760 35992 22772
rect 31680 22732 35992 22760
rect 31570 22692 31576 22704
rect 30668 22664 31576 22692
rect 28408 22652 28414 22664
rect 31570 22652 31576 22664
rect 31628 22652 31634 22704
rect 16853 22627 16911 22633
rect 16853 22593 16865 22627
rect 16899 22593 16911 22627
rect 16853 22587 16911 22593
rect 18230 22584 18236 22636
rect 18288 22624 18294 22636
rect 18969 22627 19027 22633
rect 18969 22624 18981 22627
rect 18288 22596 18981 22624
rect 18288 22584 18294 22596
rect 18969 22593 18981 22596
rect 19015 22624 19027 22627
rect 19334 22624 19340 22636
rect 19015 22596 19340 22624
rect 19015 22593 19027 22596
rect 18969 22587 19027 22593
rect 19334 22584 19340 22596
rect 19392 22584 19398 22636
rect 22005 22627 22063 22633
rect 22005 22624 22017 22627
rect 21468 22596 22017 22624
rect 10226 22516 10232 22568
rect 10284 22516 10290 22568
rect 11900 22528 12112 22556
rect 11900 22488 11928 22528
rect 9876 22460 11928 22488
rect 7098 22420 7104 22432
rect 3988 22392 7104 22420
rect 7098 22380 7104 22392
rect 7156 22380 7162 22432
rect 8662 22380 8668 22432
rect 8720 22420 8726 22432
rect 11885 22423 11943 22429
rect 11885 22420 11897 22423
rect 8720 22392 11897 22420
rect 8720 22380 8726 22392
rect 11885 22389 11897 22392
rect 11931 22389 11943 22423
rect 12084 22420 12112 22528
rect 12250 22516 12256 22568
rect 12308 22556 12314 22568
rect 12308 22528 12434 22556
rect 12308 22516 12314 22528
rect 12406 22488 12434 22528
rect 12526 22516 12532 22568
rect 12584 22556 12590 22568
rect 13081 22559 13139 22565
rect 13081 22556 13093 22559
rect 12584 22528 13093 22556
rect 12584 22516 12590 22528
rect 13081 22525 13093 22528
rect 13127 22525 13139 22559
rect 13081 22519 13139 22525
rect 13538 22516 13544 22568
rect 13596 22556 13602 22568
rect 14369 22559 14427 22565
rect 14369 22556 14381 22559
rect 13596 22528 14381 22556
rect 13596 22516 13602 22528
rect 14369 22525 14381 22528
rect 14415 22556 14427 22559
rect 14458 22556 14464 22568
rect 14415 22528 14464 22556
rect 14415 22525 14427 22528
rect 14369 22519 14427 22525
rect 14458 22516 14464 22528
rect 14516 22516 14522 22568
rect 15102 22516 15108 22568
rect 15160 22556 15166 22568
rect 15381 22559 15439 22565
rect 15381 22556 15393 22559
rect 15160 22528 15393 22556
rect 15160 22516 15166 22528
rect 15381 22525 15393 22528
rect 15427 22525 15439 22559
rect 15381 22519 15439 22525
rect 16758 22516 16764 22568
rect 16816 22556 16822 22568
rect 17129 22559 17187 22565
rect 17129 22556 17141 22559
rect 16816 22528 17141 22556
rect 16816 22516 16822 22528
rect 17129 22525 17141 22528
rect 17175 22525 17187 22559
rect 17129 22519 17187 22525
rect 18598 22516 18604 22568
rect 18656 22556 18662 22568
rect 19429 22559 19487 22565
rect 19429 22556 19441 22559
rect 18656 22528 19441 22556
rect 18656 22516 18662 22528
rect 19429 22525 19441 22528
rect 19475 22525 19487 22559
rect 19429 22519 19487 22525
rect 18690 22488 18696 22500
rect 12406 22460 16988 22488
rect 14182 22420 14188 22432
rect 12084 22392 14188 22420
rect 11885 22383 11943 22389
rect 14182 22380 14188 22392
rect 14240 22380 14246 22432
rect 16960 22420 16988 22460
rect 18156 22460 18696 22488
rect 18156 22420 18184 22460
rect 18690 22448 18696 22460
rect 18748 22448 18754 22500
rect 20714 22448 20720 22500
rect 20772 22488 20778 22500
rect 21174 22488 21180 22500
rect 20772 22460 21180 22488
rect 20772 22448 20778 22460
rect 21174 22448 21180 22460
rect 21232 22448 21238 22500
rect 16960 22392 18184 22420
rect 20346 22380 20352 22432
rect 20404 22420 20410 22432
rect 21468 22420 21496 22596
rect 22005 22593 22017 22596
rect 22051 22593 22063 22627
rect 22005 22587 22063 22593
rect 24854 22584 24860 22636
rect 24912 22584 24918 22636
rect 27338 22584 27344 22636
rect 27396 22584 27402 22636
rect 27798 22584 27804 22636
rect 27856 22624 27862 22636
rect 28077 22627 28135 22633
rect 28077 22624 28089 22627
rect 27856 22596 28089 22624
rect 27856 22584 27862 22596
rect 28077 22593 28089 22596
rect 28123 22593 28135 22627
rect 28077 22587 28135 22593
rect 29454 22584 29460 22636
rect 29512 22584 29518 22636
rect 30650 22584 30656 22636
rect 30708 22584 30714 22636
rect 31680 22633 31708 22732
rect 35986 22720 35992 22732
rect 36044 22720 36050 22772
rect 36078 22720 36084 22772
rect 36136 22720 36142 22772
rect 38562 22720 38568 22772
rect 38620 22760 38626 22772
rect 41230 22760 41236 22772
rect 38620 22732 41236 22760
rect 38620 22720 38626 22732
rect 41230 22720 41236 22732
rect 41288 22720 41294 22772
rect 41966 22760 41972 22772
rect 41340 22732 41972 22760
rect 32677 22695 32735 22701
rect 32677 22661 32689 22695
rect 32723 22692 32735 22695
rect 33870 22692 33876 22704
rect 32723 22664 33876 22692
rect 32723 22661 32735 22664
rect 32677 22655 32735 22661
rect 33870 22652 33876 22664
rect 33928 22652 33934 22704
rect 33962 22652 33968 22704
rect 34020 22652 34026 22704
rect 34422 22652 34428 22704
rect 34480 22652 34486 22704
rect 37826 22692 37832 22704
rect 37200 22664 37832 22692
rect 31665 22627 31723 22633
rect 31665 22593 31677 22627
rect 31711 22593 31723 22627
rect 31665 22587 31723 22593
rect 32769 22627 32827 22633
rect 32769 22593 32781 22627
rect 32815 22624 32827 22627
rect 32815 22596 33640 22624
rect 32815 22593 32827 22596
rect 32769 22587 32827 22593
rect 21542 22516 21548 22568
rect 21600 22556 21606 22568
rect 23474 22556 23480 22568
rect 21600 22528 23480 22556
rect 21600 22516 21606 22528
rect 23474 22516 23480 22528
rect 23532 22516 23538 22568
rect 24486 22516 24492 22568
rect 24544 22556 24550 22568
rect 27522 22556 27528 22568
rect 24544 22528 27528 22556
rect 24544 22516 24550 22528
rect 27522 22516 27528 22528
rect 27580 22516 27586 22568
rect 28350 22516 28356 22568
rect 28408 22516 28414 22568
rect 28442 22516 28448 22568
rect 28500 22556 28506 22568
rect 30837 22559 30895 22565
rect 30837 22556 30849 22559
rect 28500 22528 30849 22556
rect 28500 22516 28506 22528
rect 30837 22525 30849 22528
rect 30883 22525 30895 22559
rect 30837 22519 30895 22525
rect 32861 22559 32919 22565
rect 32861 22525 32873 22559
rect 32907 22525 32919 22559
rect 33612 22556 33640 22596
rect 33686 22584 33692 22636
rect 33744 22584 33750 22636
rect 35986 22584 35992 22636
rect 36044 22624 36050 22636
rect 36449 22627 36507 22633
rect 36449 22624 36461 22627
rect 36044 22596 36461 22624
rect 36044 22584 36050 22596
rect 36449 22593 36461 22596
rect 36495 22593 36507 22627
rect 36449 22587 36507 22593
rect 36541 22627 36599 22633
rect 36541 22593 36553 22627
rect 36587 22624 36599 22627
rect 36814 22624 36820 22636
rect 36587 22596 36820 22624
rect 36587 22593 36599 22596
rect 36541 22587 36599 22593
rect 36814 22584 36820 22596
rect 36872 22584 36878 22636
rect 33612 22528 33824 22556
rect 32861 22519 32919 22525
rect 24213 22491 24271 22497
rect 24213 22457 24225 22491
rect 24259 22488 24271 22491
rect 24578 22488 24584 22500
rect 24259 22460 24584 22488
rect 24259 22457 24271 22460
rect 24213 22451 24271 22457
rect 24578 22448 24584 22460
rect 24636 22448 24642 22500
rect 27154 22448 27160 22500
rect 27212 22448 27218 22500
rect 29362 22448 29368 22500
rect 29420 22488 29426 22500
rect 32876 22488 32904 22519
rect 29420 22460 32904 22488
rect 29420 22448 29426 22460
rect 22462 22420 22468 22432
rect 20404 22392 22468 22420
rect 20404 22380 20410 22392
rect 22462 22380 22468 22392
rect 22520 22380 22526 22432
rect 26602 22380 26608 22432
rect 26660 22380 26666 22432
rect 28902 22380 28908 22432
rect 28960 22420 28966 22432
rect 29825 22423 29883 22429
rect 29825 22420 29837 22423
rect 28960 22392 29837 22420
rect 28960 22380 28966 22392
rect 29825 22389 29837 22392
rect 29871 22389 29883 22423
rect 29825 22383 29883 22389
rect 29914 22380 29920 22432
rect 29972 22420 29978 22432
rect 30285 22423 30343 22429
rect 30285 22420 30297 22423
rect 29972 22392 30297 22420
rect 29972 22380 29978 22392
rect 30285 22389 30297 22392
rect 30331 22389 30343 22423
rect 30285 22383 30343 22389
rect 31846 22380 31852 22432
rect 31904 22420 31910 22432
rect 32309 22423 32367 22429
rect 32309 22420 32321 22423
rect 31904 22392 32321 22420
rect 31904 22380 31910 22392
rect 32309 22389 32321 22392
rect 32355 22389 32367 22423
rect 32309 22383 32367 22389
rect 32858 22380 32864 22432
rect 32916 22420 32922 22432
rect 33321 22423 33379 22429
rect 33321 22420 33333 22423
rect 32916 22392 33333 22420
rect 32916 22380 32922 22392
rect 33321 22389 33333 22392
rect 33367 22420 33379 22423
rect 33594 22420 33600 22432
rect 33367 22392 33600 22420
rect 33367 22389 33379 22392
rect 33321 22383 33379 22389
rect 33594 22380 33600 22392
rect 33652 22380 33658 22432
rect 33796 22420 33824 22528
rect 34330 22516 34336 22568
rect 34388 22556 34394 22568
rect 36725 22559 36783 22565
rect 34388 22528 35480 22556
rect 34388 22516 34394 22528
rect 35452 22497 35480 22528
rect 36725 22525 36737 22559
rect 36771 22556 36783 22559
rect 37200 22556 37228 22664
rect 37826 22652 37832 22664
rect 37884 22652 37890 22704
rect 39574 22692 39580 22704
rect 38962 22664 39580 22692
rect 39574 22652 39580 22664
rect 39632 22652 39638 22704
rect 41340 22692 41368 22732
rect 41966 22720 41972 22732
rect 42024 22720 42030 22772
rect 42242 22720 42248 22772
rect 42300 22760 42306 22772
rect 42886 22760 42892 22772
rect 42300 22732 42892 22760
rect 42300 22720 42306 22732
rect 42886 22720 42892 22732
rect 42944 22720 42950 22772
rect 44542 22720 44548 22772
rect 44600 22720 44606 22772
rect 46753 22763 46811 22769
rect 46753 22729 46765 22763
rect 46799 22760 46811 22763
rect 47302 22760 47308 22772
rect 46799 22732 47308 22760
rect 46799 22729 46811 22732
rect 46753 22723 46811 22729
rect 47302 22720 47308 22732
rect 47360 22720 47366 22772
rect 47854 22720 47860 22772
rect 47912 22760 47918 22772
rect 47949 22763 48007 22769
rect 47949 22760 47961 22763
rect 47912 22732 47961 22760
rect 47912 22720 47918 22732
rect 47949 22729 47961 22732
rect 47995 22729 48007 22763
rect 47949 22723 48007 22729
rect 48406 22720 48412 22772
rect 48464 22760 48470 22772
rect 48501 22763 48559 22769
rect 48501 22760 48513 22763
rect 48464 22732 48513 22760
rect 48464 22720 48470 22732
rect 48501 22729 48513 22732
rect 48547 22729 48559 22763
rect 48501 22723 48559 22729
rect 39960 22664 41368 22692
rect 37274 22584 37280 22636
rect 37332 22624 37338 22636
rect 37461 22627 37519 22633
rect 37461 22624 37473 22627
rect 37332 22596 37473 22624
rect 37332 22584 37338 22596
rect 37461 22593 37473 22596
rect 37507 22593 37519 22627
rect 37461 22587 37519 22593
rect 39482 22584 39488 22636
rect 39540 22624 39546 22636
rect 39960 22624 39988 22664
rect 39540 22596 39988 22624
rect 39540 22584 39546 22596
rect 40034 22584 40040 22636
rect 40092 22584 40098 22636
rect 41064 22633 41092 22664
rect 41414 22652 41420 22704
rect 41472 22692 41478 22704
rect 41472 22664 42012 22692
rect 41472 22652 41478 22664
rect 41049 22627 41107 22633
rect 41049 22593 41061 22627
rect 41095 22624 41107 22627
rect 41095 22596 41129 22624
rect 41095 22593 41107 22596
rect 41049 22587 41107 22593
rect 41690 22584 41696 22636
rect 41748 22584 41754 22636
rect 41984 22633 42012 22664
rect 42058 22652 42064 22704
rect 42116 22692 42122 22704
rect 43714 22692 43720 22704
rect 42116 22664 43720 22692
rect 42116 22652 42122 22664
rect 43714 22652 43720 22664
rect 43772 22692 43778 22704
rect 47673 22695 47731 22701
rect 47673 22692 47685 22695
rect 43772 22664 44128 22692
rect 43772 22652 43778 22664
rect 41969 22627 42027 22633
rect 41969 22593 41981 22627
rect 42015 22624 42027 22627
rect 42242 22624 42248 22636
rect 42015 22596 42248 22624
rect 42015 22593 42027 22596
rect 41969 22587 42027 22593
rect 42242 22584 42248 22596
rect 42300 22584 42306 22636
rect 42794 22584 42800 22636
rect 42852 22584 42858 22636
rect 44100 22633 44128 22664
rect 47228 22664 47685 22692
rect 43441 22627 43499 22633
rect 43441 22593 43453 22627
rect 43487 22593 43499 22627
rect 43441 22587 43499 22593
rect 44085 22627 44143 22633
rect 44085 22593 44097 22627
rect 44131 22593 44143 22627
rect 44085 22587 44143 22593
rect 44729 22627 44787 22633
rect 44729 22593 44741 22627
rect 44775 22624 44787 22627
rect 45005 22627 45063 22633
rect 45005 22624 45017 22627
rect 44775 22596 45017 22624
rect 44775 22593 44787 22596
rect 44729 22587 44787 22593
rect 45005 22593 45017 22596
rect 45051 22593 45063 22627
rect 45005 22587 45063 22593
rect 36771 22528 37228 22556
rect 36771 22525 36783 22528
rect 36725 22519 36783 22525
rect 37734 22516 37740 22568
rect 37792 22516 37798 22568
rect 37826 22516 37832 22568
rect 37884 22556 37890 22568
rect 37884 22528 39712 22556
rect 37884 22516 37890 22528
rect 35437 22491 35495 22497
rect 35437 22457 35449 22491
rect 35483 22488 35495 22491
rect 37458 22488 37464 22500
rect 35483 22460 37464 22488
rect 35483 22457 35495 22460
rect 35437 22451 35495 22457
rect 37458 22448 37464 22460
rect 37516 22448 37522 22500
rect 39224 22497 39252 22528
rect 39209 22491 39267 22497
rect 39209 22457 39221 22491
rect 39255 22457 39267 22491
rect 39684 22488 39712 22528
rect 40126 22516 40132 22568
rect 40184 22516 40190 22568
rect 40221 22559 40279 22565
rect 40221 22525 40233 22559
rect 40267 22525 40279 22559
rect 40221 22519 40279 22525
rect 40236 22488 40264 22519
rect 40862 22516 40868 22568
rect 40920 22556 40926 22568
rect 43346 22556 43352 22568
rect 40920 22528 43352 22556
rect 40920 22516 40926 22528
rect 43346 22516 43352 22528
rect 43404 22556 43410 22568
rect 43456 22556 43484 22587
rect 44744 22556 44772 22587
rect 46658 22584 46664 22636
rect 46716 22624 46722 22636
rect 47228 22633 47256 22664
rect 47673 22661 47685 22664
rect 47719 22661 47731 22695
rect 47673 22655 47731 22661
rect 47213 22627 47271 22633
rect 47213 22624 47225 22627
rect 46716 22596 47225 22624
rect 46716 22584 46722 22596
rect 47213 22593 47225 22596
rect 47259 22593 47271 22627
rect 47213 22587 47271 22593
rect 47578 22584 47584 22636
rect 47636 22624 47642 22636
rect 47857 22627 47915 22633
rect 47857 22624 47869 22627
rect 47636 22596 47869 22624
rect 47636 22584 47642 22596
rect 47857 22593 47869 22596
rect 47903 22624 47915 22627
rect 48317 22627 48375 22633
rect 48317 22624 48329 22627
rect 47903 22596 48329 22624
rect 47903 22593 47915 22596
rect 47857 22587 47915 22593
rect 48317 22593 48329 22596
rect 48363 22593 48375 22627
rect 48317 22587 48375 22593
rect 49050 22584 49056 22636
rect 49108 22584 49114 22636
rect 43404 22528 43484 22556
rect 44100 22528 44772 22556
rect 43404 22516 43410 22528
rect 39684 22460 40264 22488
rect 40512 22460 42564 22488
rect 39209 22451 39267 22457
rect 35342 22420 35348 22432
rect 33796 22392 35348 22420
rect 35342 22380 35348 22392
rect 35400 22380 35406 22432
rect 35526 22380 35532 22432
rect 35584 22420 35590 22432
rect 35713 22423 35771 22429
rect 35713 22420 35725 22423
rect 35584 22392 35725 22420
rect 35584 22380 35590 22392
rect 35713 22389 35725 22392
rect 35759 22389 35771 22423
rect 35713 22383 35771 22389
rect 37734 22380 37740 22432
rect 37792 22420 37798 22432
rect 39482 22420 39488 22432
rect 37792 22392 39488 22420
rect 37792 22380 37798 22392
rect 39482 22380 39488 22392
rect 39540 22380 39546 22432
rect 39666 22380 39672 22432
rect 39724 22380 39730 22432
rect 39850 22380 39856 22432
rect 39908 22420 39914 22432
rect 40512 22420 40540 22460
rect 39908 22392 40540 22420
rect 40865 22423 40923 22429
rect 39908 22380 39914 22392
rect 40865 22389 40877 22423
rect 40911 22420 40923 22423
rect 40954 22420 40960 22432
rect 40911 22392 40960 22420
rect 40911 22389 40923 22392
rect 40865 22383 40923 22389
rect 40954 22380 40960 22392
rect 41012 22380 41018 22432
rect 41506 22380 41512 22432
rect 41564 22380 41570 22432
rect 42150 22380 42156 22432
rect 42208 22380 42214 22432
rect 42536 22420 42564 22460
rect 42610 22448 42616 22500
rect 42668 22448 42674 22500
rect 44100 22488 44128 22528
rect 42720 22460 44128 22488
rect 42720 22420 42748 22460
rect 44174 22448 44180 22500
rect 44232 22488 44238 22500
rect 47029 22491 47087 22497
rect 47029 22488 47041 22491
rect 44232 22460 47041 22488
rect 44232 22448 44238 22460
rect 47029 22457 47041 22460
rect 47075 22457 47087 22491
rect 47029 22451 47087 22457
rect 42536 22392 42748 22420
rect 42794 22380 42800 22432
rect 42852 22420 42858 22432
rect 43257 22423 43315 22429
rect 43257 22420 43269 22423
rect 42852 22392 43269 22420
rect 42852 22380 42858 22392
rect 43257 22389 43269 22392
rect 43303 22389 43315 22423
rect 43257 22383 43315 22389
rect 43898 22380 43904 22432
rect 43956 22380 43962 22432
rect 48590 22380 48596 22432
rect 48648 22420 48654 22432
rect 49237 22423 49295 22429
rect 49237 22420 49249 22423
rect 48648 22392 49249 22420
rect 48648 22380 48654 22392
rect 49237 22389 49249 22392
rect 49283 22389 49295 22423
rect 49237 22383 49295 22389
rect 1104 22330 49864 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 32950 22330
rect 33002 22278 33014 22330
rect 33066 22278 33078 22330
rect 33130 22278 33142 22330
rect 33194 22278 33206 22330
rect 33258 22278 42950 22330
rect 43002 22278 43014 22330
rect 43066 22278 43078 22330
rect 43130 22278 43142 22330
rect 43194 22278 43206 22330
rect 43258 22278 49864 22330
rect 1104 22256 49864 22278
rect 2222 22176 2228 22228
rect 2280 22216 2286 22228
rect 4890 22216 4896 22228
rect 2280 22188 4896 22216
rect 2280 22176 2286 22188
rect 4890 22176 4896 22188
rect 4948 22176 4954 22228
rect 6914 22176 6920 22228
rect 6972 22216 6978 22228
rect 7837 22219 7895 22225
rect 7837 22216 7849 22219
rect 6972 22188 7849 22216
rect 6972 22176 6978 22188
rect 7837 22185 7849 22188
rect 7883 22185 7895 22219
rect 7837 22179 7895 22185
rect 8386 22176 8392 22228
rect 8444 22176 8450 22228
rect 12342 22176 12348 22228
rect 12400 22176 12406 22228
rect 12989 22219 13047 22225
rect 12989 22216 13001 22219
rect 12452 22188 13001 22216
rect 3970 22108 3976 22160
rect 4028 22148 4034 22160
rect 4028 22120 6316 22148
rect 4028 22108 4034 22120
rect 1302 22040 1308 22092
rect 1360 22080 1366 22092
rect 2041 22083 2099 22089
rect 2041 22080 2053 22083
rect 1360 22052 2053 22080
rect 1360 22040 1366 22052
rect 2041 22049 2053 22052
rect 2087 22049 2099 22083
rect 2041 22043 2099 22049
rect 3878 22040 3884 22092
rect 3936 22080 3942 22092
rect 6288 22089 6316 22120
rect 11146 22108 11152 22160
rect 11204 22148 11210 22160
rect 12452 22148 12480 22188
rect 12989 22185 13001 22188
rect 13035 22185 13047 22219
rect 16758 22216 16764 22228
rect 12989 22179 13047 22185
rect 13648 22188 16764 22216
rect 11204 22120 12480 22148
rect 11204 22108 11210 22120
rect 4433 22083 4491 22089
rect 4433 22080 4445 22083
rect 3936 22052 4445 22080
rect 3936 22040 3942 22052
rect 4433 22049 4445 22052
rect 4479 22049 4491 22083
rect 4433 22043 4491 22049
rect 6273 22083 6331 22089
rect 6273 22049 6285 22083
rect 6319 22049 6331 22083
rect 6273 22043 6331 22049
rect 7576 22052 9260 22080
rect 1765 22015 1823 22021
rect 1765 21981 1777 22015
rect 1811 22012 1823 22015
rect 1811 21984 2774 22012
rect 1811 21981 1823 21984
rect 1765 21975 1823 21981
rect 2746 21944 2774 21984
rect 4062 21972 4068 22024
rect 4120 21972 4126 22024
rect 5997 22015 6055 22021
rect 5997 21981 6009 22015
rect 6043 22012 6055 22015
rect 6454 22012 6460 22024
rect 6043 21984 6460 22012
rect 6043 21981 6055 21984
rect 5997 21975 6055 21981
rect 6454 21972 6460 21984
rect 6512 21972 6518 22024
rect 7576 21944 7604 22052
rect 8573 22015 8631 22021
rect 8573 21981 8585 22015
rect 8619 21981 8631 22015
rect 8573 21975 8631 21981
rect 2746 21916 7604 21944
rect 7745 21947 7803 21953
rect 7745 21913 7757 21947
rect 7791 21913 7803 21947
rect 8588 21944 8616 21975
rect 9122 21972 9128 22024
rect 9180 21972 9186 22024
rect 9232 22012 9260 22052
rect 10042 22040 10048 22092
rect 10100 22040 10106 22092
rect 11054 22040 11060 22092
rect 11112 22040 11118 22092
rect 13648 22089 13676 22188
rect 16758 22176 16764 22188
rect 16816 22216 16822 22228
rect 16945 22219 17003 22225
rect 16945 22216 16957 22219
rect 16816 22188 16957 22216
rect 16816 22176 16822 22188
rect 16945 22185 16957 22188
rect 16991 22185 17003 22219
rect 16945 22179 17003 22185
rect 17034 22176 17040 22228
rect 17092 22216 17098 22228
rect 18598 22216 18604 22228
rect 17092 22188 18604 22216
rect 17092 22176 17098 22188
rect 18598 22176 18604 22188
rect 18656 22176 18662 22228
rect 18690 22176 18696 22228
rect 18748 22216 18754 22228
rect 22186 22216 22192 22228
rect 18748 22188 22192 22216
rect 18748 22176 18754 22188
rect 22186 22176 22192 22188
rect 22244 22176 22250 22228
rect 23750 22176 23756 22228
rect 23808 22216 23814 22228
rect 23845 22219 23903 22225
rect 23845 22216 23857 22219
rect 23808 22188 23857 22216
rect 23808 22176 23814 22188
rect 23845 22185 23857 22188
rect 23891 22185 23903 22219
rect 23845 22179 23903 22185
rect 24394 22176 24400 22228
rect 24452 22216 24458 22228
rect 27798 22216 27804 22228
rect 24452 22188 27804 22216
rect 24452 22176 24458 22188
rect 27798 22176 27804 22188
rect 27856 22176 27862 22228
rect 28350 22176 28356 22228
rect 28408 22216 28414 22228
rect 28994 22216 29000 22228
rect 28408 22188 29000 22216
rect 28408 22176 28414 22188
rect 28994 22176 29000 22188
rect 29052 22216 29058 22228
rect 29362 22216 29368 22228
rect 29052 22188 29368 22216
rect 29052 22176 29058 22188
rect 29362 22176 29368 22188
rect 29420 22176 29426 22228
rect 29454 22176 29460 22228
rect 29512 22216 29518 22228
rect 30193 22219 30251 22225
rect 30193 22216 30205 22219
rect 29512 22188 30205 22216
rect 29512 22176 29518 22188
rect 30193 22185 30205 22188
rect 30239 22216 30251 22219
rect 31570 22216 31576 22228
rect 30239 22188 31576 22216
rect 30239 22185 30251 22188
rect 30193 22179 30251 22185
rect 31570 22176 31576 22188
rect 31628 22176 31634 22228
rect 32582 22176 32588 22228
rect 32640 22176 32646 22228
rect 33318 22176 33324 22228
rect 33376 22216 33382 22228
rect 37182 22216 37188 22228
rect 33376 22188 37188 22216
rect 33376 22176 33382 22188
rect 37182 22176 37188 22188
rect 37240 22176 37246 22228
rect 37550 22225 37556 22228
rect 37540 22219 37556 22225
rect 37540 22185 37552 22219
rect 37540 22179 37556 22185
rect 37550 22176 37556 22179
rect 37608 22176 37614 22228
rect 40034 22176 40040 22228
rect 40092 22216 40098 22228
rect 41233 22219 41291 22225
rect 41233 22216 41245 22219
rect 40092 22188 41245 22216
rect 40092 22176 40098 22188
rect 41233 22185 41245 22188
rect 41279 22185 41291 22219
rect 41233 22179 41291 22185
rect 41690 22176 41696 22228
rect 41748 22216 41754 22228
rect 42613 22219 42671 22225
rect 42613 22216 42625 22219
rect 41748 22188 42625 22216
rect 41748 22176 41754 22188
rect 42613 22185 42625 22188
rect 42659 22185 42671 22219
rect 42613 22179 42671 22185
rect 42702 22176 42708 22228
rect 42760 22216 42766 22228
rect 42797 22219 42855 22225
rect 42797 22216 42809 22219
rect 42760 22188 42809 22216
rect 42760 22176 42766 22188
rect 42797 22185 42809 22188
rect 42843 22185 42855 22219
rect 42797 22179 42855 22185
rect 43165 22219 43223 22225
rect 43165 22185 43177 22219
rect 43211 22216 43223 22219
rect 43346 22216 43352 22228
rect 43211 22188 43352 22216
rect 43211 22185 43223 22188
rect 43165 22179 43223 22185
rect 43346 22176 43352 22188
rect 43404 22176 43410 22228
rect 43714 22176 43720 22228
rect 43772 22176 43778 22228
rect 47489 22219 47547 22225
rect 47489 22185 47501 22219
rect 47535 22216 47547 22219
rect 49326 22216 49332 22228
rect 47535 22188 49332 22216
rect 47535 22185 47547 22188
rect 47489 22179 47547 22185
rect 49326 22176 49332 22188
rect 49384 22176 49390 22228
rect 17218 22108 17224 22160
rect 17276 22148 17282 22160
rect 17276 22120 18000 22148
rect 17276 22108 17282 22120
rect 13633 22083 13691 22089
rect 13633 22049 13645 22083
rect 13679 22049 13691 22083
rect 13633 22043 13691 22049
rect 13722 22040 13728 22092
rect 13780 22080 13786 22092
rect 14737 22083 14795 22089
rect 14737 22080 14749 22083
rect 13780 22052 14749 22080
rect 13780 22040 13786 22052
rect 14737 22049 14749 22052
rect 14783 22049 14795 22083
rect 14737 22043 14795 22049
rect 15473 22083 15531 22089
rect 15473 22049 15485 22083
rect 15519 22080 15531 22083
rect 16114 22080 16120 22092
rect 15519 22052 16120 22080
rect 15519 22049 15531 22052
rect 15473 22043 15531 22049
rect 16114 22040 16120 22052
rect 16172 22040 16178 22092
rect 16482 22040 16488 22092
rect 16540 22080 16546 22092
rect 17972 22089 18000 22120
rect 18966 22108 18972 22160
rect 19024 22148 19030 22160
rect 19024 22120 19932 22148
rect 19024 22108 19030 22120
rect 19904 22089 19932 22120
rect 21450 22108 21456 22160
rect 21508 22148 21514 22160
rect 26602 22148 26608 22160
rect 21508 22120 22048 22148
rect 21508 22108 21514 22120
rect 17957 22083 18015 22089
rect 16540 22052 17540 22080
rect 16540 22040 16546 22052
rect 9232 21984 11284 22012
rect 11146 21944 11152 21956
rect 8588 21916 11152 21944
rect 7745 21907 7803 21913
rect 7760 21876 7788 21907
rect 11146 21904 11152 21916
rect 11204 21904 11210 21956
rect 11256 21944 11284 21984
rect 11330 21972 11336 22024
rect 11388 21972 11394 22024
rect 12526 21972 12532 22024
rect 12584 21972 12590 22024
rect 15194 21972 15200 22024
rect 15252 21972 15258 22024
rect 12710 21944 12716 21956
rect 11256 21916 12716 21944
rect 12710 21904 12716 21916
rect 12768 21904 12774 21956
rect 14553 21947 14611 21953
rect 14553 21913 14565 21947
rect 14599 21944 14611 21947
rect 14734 21944 14740 21956
rect 14599 21916 14740 21944
rect 14599 21913 14611 21916
rect 14553 21907 14611 21913
rect 14734 21904 14740 21916
rect 14792 21904 14798 21956
rect 16758 21944 16764 21956
rect 16698 21916 16764 21944
rect 16758 21904 16764 21916
rect 16816 21904 16822 21956
rect 9674 21876 9680 21888
rect 7760 21848 9680 21876
rect 9674 21836 9680 21848
rect 9732 21836 9738 21888
rect 9858 21836 9864 21888
rect 9916 21876 9922 21888
rect 13357 21879 13415 21885
rect 13357 21876 13369 21879
rect 9916 21848 13369 21876
rect 9916 21836 9922 21848
rect 13357 21845 13369 21848
rect 13403 21845 13415 21879
rect 13357 21839 13415 21845
rect 13449 21879 13507 21885
rect 13449 21845 13461 21879
rect 13495 21876 13507 21879
rect 16482 21876 16488 21888
rect 13495 21848 16488 21876
rect 13495 21845 13507 21848
rect 13449 21839 13507 21845
rect 16482 21836 16488 21848
rect 16540 21836 16546 21888
rect 17512 21876 17540 22052
rect 17957 22049 17969 22083
rect 18003 22049 18015 22083
rect 17957 22043 18015 22049
rect 19889 22083 19947 22089
rect 19889 22049 19901 22083
rect 19935 22049 19947 22083
rect 19889 22043 19947 22049
rect 20714 22040 20720 22092
rect 20772 22080 20778 22092
rect 21082 22080 21088 22092
rect 20772 22052 21088 22080
rect 20772 22040 20778 22052
rect 21082 22040 21088 22052
rect 21140 22040 21146 22092
rect 22020 22089 22048 22120
rect 23216 22120 26608 22148
rect 23216 22092 23244 22120
rect 22005 22083 22063 22089
rect 22005 22049 22017 22083
rect 22051 22049 22063 22083
rect 22005 22043 22063 22049
rect 23198 22040 23204 22092
rect 23256 22040 23262 22092
rect 23566 22040 23572 22092
rect 23624 22080 23630 22092
rect 24578 22080 24584 22092
rect 23624 22052 24584 22080
rect 23624 22040 23630 22052
rect 24578 22040 24584 22052
rect 24636 22040 24642 22092
rect 25130 22040 25136 22092
rect 25188 22080 25194 22092
rect 26418 22080 26424 22092
rect 25188 22052 26424 22080
rect 25188 22040 25194 22052
rect 26418 22040 26424 22052
rect 26476 22040 26482 22092
rect 26528 22089 26556 22120
rect 26602 22108 26608 22120
rect 26660 22108 26666 22160
rect 27062 22108 27068 22160
rect 27120 22148 27126 22160
rect 29733 22151 29791 22157
rect 29733 22148 29745 22151
rect 27120 22120 27752 22148
rect 27120 22108 27126 22120
rect 26513 22083 26571 22089
rect 26513 22049 26525 22083
rect 26559 22049 26571 22083
rect 26513 22043 26571 22049
rect 27246 22040 27252 22092
rect 27304 22080 27310 22092
rect 27724 22089 27752 22120
rect 28460 22120 29040 22148
rect 27617 22083 27675 22089
rect 27617 22080 27629 22083
rect 27304 22052 27629 22080
rect 27304 22040 27310 22052
rect 27617 22049 27629 22052
rect 27663 22049 27675 22083
rect 27617 22043 27675 22049
rect 27709 22083 27767 22089
rect 27709 22049 27721 22083
rect 27755 22080 27767 22083
rect 27755 22052 27789 22080
rect 27755 22049 27767 22052
rect 27709 22043 27767 22049
rect 17589 22015 17647 22021
rect 17589 21981 17601 22015
rect 17635 21981 17647 22015
rect 17589 21975 17647 21981
rect 17604 21944 17632 21975
rect 17678 21972 17684 22024
rect 17736 22012 17742 22024
rect 18230 22012 18236 22024
rect 17736 21984 18236 22012
rect 17736 21972 17742 21984
rect 18230 21972 18236 21984
rect 18288 21972 18294 22024
rect 19426 21972 19432 22024
rect 19484 21972 19490 22024
rect 21910 22012 21916 22024
rect 19628 21984 21916 22012
rect 19628 21944 19656 21984
rect 21910 21972 21916 21984
rect 21968 21972 21974 22024
rect 23017 22015 23075 22021
rect 23017 21981 23029 22015
rect 23063 22012 23075 22015
rect 23750 22012 23756 22024
rect 23063 21984 23756 22012
rect 23063 21981 23075 21984
rect 23017 21975 23075 21981
rect 23750 21972 23756 21984
rect 23808 21972 23814 22024
rect 24029 22015 24087 22021
rect 24029 21981 24041 22015
rect 24075 22012 24087 22015
rect 24946 22012 24952 22024
rect 24075 21984 24952 22012
rect 24075 21981 24087 21984
rect 24029 21975 24087 21981
rect 24946 21972 24952 21984
rect 25004 21972 25010 22024
rect 25314 21972 25320 22024
rect 25372 22012 25378 22024
rect 28460 22012 28488 22120
rect 28534 22040 28540 22092
rect 28592 22080 28598 22092
rect 28902 22080 28908 22092
rect 28592 22052 28908 22080
rect 28592 22040 28598 22052
rect 28902 22040 28908 22052
rect 28960 22040 28966 22092
rect 29012 22080 29040 22120
rect 29656 22120 29745 22148
rect 29656 22080 29684 22120
rect 29733 22117 29745 22120
rect 29779 22117 29791 22151
rect 34330 22148 34336 22160
rect 29733 22111 29791 22117
rect 33704 22120 34336 22148
rect 30374 22080 30380 22092
rect 29012 22052 29684 22080
rect 29840 22052 30380 22080
rect 25372 21984 28488 22012
rect 28721 22015 28779 22021
rect 25372 21972 25378 21984
rect 28721 21981 28733 22015
rect 28767 22012 28779 22015
rect 29840 22012 29868 22052
rect 30374 22040 30380 22052
rect 30432 22040 30438 22092
rect 30837 22083 30895 22089
rect 30837 22049 30849 22083
rect 30883 22080 30895 22083
rect 31202 22080 31208 22092
rect 30883 22052 31208 22080
rect 30883 22049 30895 22052
rect 30837 22043 30895 22049
rect 31202 22040 31208 22052
rect 31260 22080 31266 22092
rect 32306 22080 32312 22092
rect 31260 22052 32312 22080
rect 31260 22040 31266 22052
rect 32306 22040 32312 22052
rect 32364 22040 32370 22092
rect 33704 22089 33732 22120
rect 34330 22108 34336 22120
rect 34388 22108 34394 22160
rect 34422 22108 34428 22160
rect 34480 22108 34486 22160
rect 35710 22108 35716 22160
rect 35768 22148 35774 22160
rect 35768 22120 37320 22148
rect 35768 22108 35774 22120
rect 37292 22092 37320 22120
rect 38838 22108 38844 22160
rect 38896 22148 38902 22160
rect 38896 22120 40632 22148
rect 38896 22108 38902 22120
rect 33689 22083 33747 22089
rect 33689 22049 33701 22083
rect 33735 22080 33747 22083
rect 33735 22052 33769 22080
rect 33735 22049 33747 22052
rect 33689 22043 33747 22049
rect 34146 22040 34152 22092
rect 34204 22040 34210 22092
rect 35066 22080 35072 22092
rect 34348 22052 35072 22080
rect 28767 21984 29868 22012
rect 29917 22015 29975 22021
rect 28767 21981 28779 21984
rect 28721 21975 28779 21981
rect 29917 21981 29929 22015
rect 29963 22012 29975 22015
rect 30558 22012 30564 22024
rect 29963 21984 30564 22012
rect 29963 21981 29975 21984
rect 29917 21975 29975 21981
rect 30558 21972 30564 21984
rect 30616 21972 30622 22024
rect 33042 21972 33048 22024
rect 33100 22012 33106 22024
rect 34348 22012 34376 22052
rect 35066 22040 35072 22052
rect 35124 22040 35130 22092
rect 35529 22083 35587 22089
rect 35529 22049 35541 22083
rect 35575 22080 35587 22083
rect 35618 22080 35624 22092
rect 35575 22052 35624 22080
rect 35575 22049 35587 22052
rect 35529 22043 35587 22049
rect 35618 22040 35624 22052
rect 35676 22040 35682 22092
rect 36725 22083 36783 22089
rect 36004 22052 36676 22080
rect 33100 21984 34376 22012
rect 33100 21972 33106 21984
rect 34422 21972 34428 22024
rect 34480 22012 34486 22024
rect 35345 22015 35403 22021
rect 35345 22012 35357 22015
rect 34480 21984 35357 22012
rect 34480 21972 34486 21984
rect 35345 21981 35357 21984
rect 35391 22012 35403 22015
rect 36004 22012 36032 22052
rect 36648 22024 36676 22052
rect 36725 22049 36737 22083
rect 36771 22049 36783 22083
rect 36725 22043 36783 22049
rect 35391 21984 36032 22012
rect 35391 21981 35403 21984
rect 35345 21975 35403 21981
rect 36078 21972 36084 22024
rect 36136 22012 36142 22024
rect 36541 22015 36599 22021
rect 36541 22012 36553 22015
rect 36136 21984 36553 22012
rect 36136 21972 36142 21984
rect 36541 21981 36553 21984
rect 36587 21981 36599 22015
rect 36541 21975 36599 21981
rect 36630 21972 36636 22024
rect 36688 21972 36694 22024
rect 36740 22012 36768 22043
rect 37274 22040 37280 22092
rect 37332 22080 37338 22092
rect 37642 22080 37648 22092
rect 37332 22052 37648 22080
rect 37332 22040 37338 22052
rect 37642 22040 37648 22052
rect 37700 22040 37706 22092
rect 38286 22040 38292 22092
rect 38344 22080 38350 22092
rect 40604 22089 40632 22120
rect 40770 22108 40776 22160
rect 40828 22148 40834 22160
rect 40828 22120 41828 22148
rect 40828 22108 40834 22120
rect 41800 22094 41828 22120
rect 42426 22108 42432 22160
rect 42484 22108 42490 22160
rect 39025 22083 39083 22089
rect 39025 22080 39037 22083
rect 38344 22052 39037 22080
rect 38344 22040 38350 22052
rect 39025 22049 39037 22052
rect 39071 22049 39083 22083
rect 39025 22043 39083 22049
rect 40589 22083 40647 22089
rect 40589 22049 40601 22083
rect 40635 22049 40647 22083
rect 40589 22043 40647 22049
rect 41598 22040 41604 22092
rect 41656 22080 41662 22092
rect 41800 22089 41865 22094
rect 41693 22083 41751 22089
rect 41693 22080 41705 22083
rect 41656 22052 41705 22080
rect 41656 22040 41662 22052
rect 41693 22049 41705 22052
rect 41739 22049 41751 22083
rect 41693 22043 41751 22049
rect 41785 22083 41865 22089
rect 41785 22049 41797 22083
rect 41831 22066 41865 22083
rect 41831 22049 41843 22066
rect 41785 22043 41843 22049
rect 42058 22040 42064 22092
rect 42116 22080 42122 22092
rect 42337 22083 42395 22089
rect 42337 22080 42349 22083
rect 42116 22052 42349 22080
rect 42116 22040 42122 22052
rect 42337 22049 42349 22052
rect 42383 22080 42395 22083
rect 49234 22080 49240 22092
rect 42383 22052 49240 22080
rect 42383 22049 42395 22052
rect 42337 22043 42395 22049
rect 49234 22040 49240 22052
rect 49292 22040 49298 22092
rect 40497 22015 40555 22021
rect 36740 21984 37320 22012
rect 37292 21956 37320 21984
rect 40497 21981 40509 22015
rect 40543 22012 40555 22015
rect 40543 21984 41920 22012
rect 40543 21981 40555 21984
rect 40497 21975 40555 21981
rect 21821 21947 21879 21953
rect 17604 21916 19656 21944
rect 21008 21916 21496 21944
rect 21008 21876 21036 21916
rect 21468 21885 21496 21916
rect 21821 21913 21833 21947
rect 21867 21944 21879 21947
rect 24762 21944 24768 21956
rect 21867 21916 24768 21944
rect 21867 21913 21879 21916
rect 21821 21907 21879 21913
rect 24762 21904 24768 21916
rect 24820 21904 24826 21956
rect 25685 21947 25743 21953
rect 25685 21944 25697 21947
rect 24964 21916 25697 21944
rect 17512 21848 21036 21876
rect 21453 21879 21511 21885
rect 21453 21845 21465 21879
rect 21499 21845 21511 21879
rect 21453 21839 21511 21845
rect 21910 21836 21916 21888
rect 21968 21836 21974 21888
rect 22646 21836 22652 21888
rect 22704 21836 22710 21888
rect 23109 21879 23167 21885
rect 23109 21845 23121 21879
rect 23155 21876 23167 21879
rect 23566 21876 23572 21888
rect 23155 21848 23572 21876
rect 23155 21845 23167 21848
rect 23109 21839 23167 21845
rect 23566 21836 23572 21848
rect 23624 21836 23630 21888
rect 23842 21836 23848 21888
rect 23900 21876 23906 21888
rect 24581 21879 24639 21885
rect 24581 21876 24593 21879
rect 23900 21848 24593 21876
rect 23900 21836 23906 21848
rect 24581 21845 24593 21848
rect 24627 21845 24639 21879
rect 24581 21839 24639 21845
rect 24854 21836 24860 21888
rect 24912 21876 24918 21888
rect 24964 21885 24992 21916
rect 25685 21913 25697 21916
rect 25731 21944 25743 21947
rect 25774 21944 25780 21956
rect 25731 21916 25780 21944
rect 25731 21913 25743 21916
rect 25685 21907 25743 21913
rect 25774 21904 25780 21916
rect 25832 21904 25838 21956
rect 26142 21904 26148 21956
rect 26200 21944 26206 21956
rect 26329 21947 26387 21953
rect 26329 21944 26341 21947
rect 26200 21916 26341 21944
rect 26200 21904 26206 21916
rect 26329 21913 26341 21916
rect 26375 21913 26387 21947
rect 26329 21907 26387 21913
rect 26421 21947 26479 21953
rect 26421 21913 26433 21947
rect 26467 21944 26479 21947
rect 29822 21944 29828 21956
rect 26467 21916 29828 21944
rect 26467 21913 26479 21916
rect 26421 21907 26479 21913
rect 29822 21904 29828 21916
rect 29880 21904 29886 21956
rect 30742 21904 30748 21956
rect 30800 21944 30806 21956
rect 31113 21947 31171 21953
rect 31113 21944 31125 21947
rect 30800 21916 31125 21944
rect 30800 21904 30806 21916
rect 31113 21913 31125 21916
rect 31159 21944 31171 21947
rect 31386 21944 31392 21956
rect 31159 21916 31392 21944
rect 31159 21913 31171 21916
rect 31113 21907 31171 21913
rect 31386 21904 31392 21916
rect 31444 21904 31450 21956
rect 31570 21904 31576 21956
rect 31628 21904 31634 21956
rect 36354 21944 36360 21956
rect 34900 21916 36360 21944
rect 24949 21879 25007 21885
rect 24949 21876 24961 21879
rect 24912 21848 24961 21876
rect 24912 21836 24918 21848
rect 24949 21845 24961 21848
rect 24995 21845 25007 21879
rect 24949 21839 25007 21845
rect 25038 21836 25044 21888
rect 25096 21836 25102 21888
rect 25958 21836 25964 21888
rect 26016 21836 26022 21888
rect 26510 21836 26516 21888
rect 26568 21876 26574 21888
rect 27157 21879 27215 21885
rect 27157 21876 27169 21879
rect 26568 21848 27169 21876
rect 26568 21836 26574 21848
rect 27157 21845 27169 21848
rect 27203 21845 27215 21879
rect 27157 21839 27215 21845
rect 27430 21836 27436 21888
rect 27488 21876 27494 21888
rect 27525 21879 27583 21885
rect 27525 21876 27537 21879
rect 27488 21848 27537 21876
rect 27488 21836 27494 21848
rect 27525 21845 27537 21848
rect 27571 21845 27583 21879
rect 27525 21839 27583 21845
rect 27614 21836 27620 21888
rect 27672 21876 27678 21888
rect 28353 21879 28411 21885
rect 28353 21876 28365 21879
rect 27672 21848 28365 21876
rect 27672 21836 27678 21848
rect 28353 21845 28365 21848
rect 28399 21845 28411 21879
rect 28353 21839 28411 21845
rect 28813 21879 28871 21885
rect 28813 21845 28825 21879
rect 28859 21876 28871 21879
rect 31846 21876 31852 21888
rect 28859 21848 31852 21876
rect 28859 21845 28871 21848
rect 28813 21839 28871 21845
rect 31846 21836 31852 21848
rect 31904 21836 31910 21888
rect 32674 21836 32680 21888
rect 32732 21876 32738 21888
rect 33045 21879 33103 21885
rect 33045 21876 33057 21879
rect 32732 21848 33057 21876
rect 32732 21836 32738 21848
rect 33045 21845 33057 21848
rect 33091 21845 33103 21879
rect 33045 21839 33103 21845
rect 33410 21836 33416 21888
rect 33468 21836 33474 21888
rect 33502 21836 33508 21888
rect 33560 21836 33566 21888
rect 34900 21885 34928 21916
rect 36354 21904 36360 21916
rect 36412 21904 36418 21956
rect 36449 21947 36507 21953
rect 36449 21913 36461 21947
rect 36495 21944 36507 21947
rect 36495 21916 37228 21944
rect 36495 21913 36507 21916
rect 36449 21907 36507 21913
rect 34885 21879 34943 21885
rect 34885 21845 34897 21879
rect 34931 21845 34943 21879
rect 34885 21839 34943 21845
rect 35158 21836 35164 21888
rect 35216 21876 35222 21888
rect 35253 21879 35311 21885
rect 35253 21876 35265 21879
rect 35216 21848 35265 21876
rect 35216 21836 35222 21848
rect 35253 21845 35265 21848
rect 35299 21876 35311 21879
rect 35526 21876 35532 21888
rect 35299 21848 35532 21876
rect 35299 21845 35311 21848
rect 35253 21839 35311 21845
rect 35526 21836 35532 21848
rect 35584 21836 35590 21888
rect 36081 21879 36139 21885
rect 36081 21845 36093 21879
rect 36127 21876 36139 21879
rect 36170 21876 36176 21888
rect 36127 21848 36176 21876
rect 36127 21845 36139 21848
rect 36081 21839 36139 21845
rect 36170 21836 36176 21848
rect 36228 21836 36234 21888
rect 37200 21876 37228 21916
rect 37274 21904 37280 21956
rect 37332 21904 37338 21956
rect 38838 21944 38844 21956
rect 38778 21916 38844 21944
rect 38838 21904 38844 21916
rect 38896 21944 38902 21956
rect 39574 21944 39580 21956
rect 38896 21916 39580 21944
rect 38896 21904 38902 21916
rect 39574 21904 39580 21916
rect 39632 21944 39638 21956
rect 41414 21944 41420 21956
rect 39632 21916 41420 21944
rect 39632 21904 39638 21916
rect 41414 21904 41420 21916
rect 41472 21904 41478 21956
rect 41782 21944 41788 21956
rect 41524 21916 41788 21944
rect 38562 21876 38568 21888
rect 37200 21848 38568 21876
rect 38562 21836 38568 21848
rect 38620 21836 38626 21888
rect 40034 21836 40040 21888
rect 40092 21836 40098 21888
rect 40405 21879 40463 21885
rect 40405 21845 40417 21879
rect 40451 21876 40463 21879
rect 40678 21876 40684 21888
rect 40451 21848 40684 21876
rect 40451 21845 40463 21848
rect 40405 21839 40463 21845
rect 40678 21836 40684 21848
rect 40736 21876 40742 21888
rect 41524 21876 41552 21916
rect 41782 21904 41788 21916
rect 41840 21904 41846 21956
rect 41892 21944 41920 21984
rect 41966 21972 41972 22024
rect 42024 22008 42030 22024
rect 43257 22015 43315 22021
rect 43257 22012 43269 22015
rect 42076 22008 43269 22012
rect 42024 21984 43269 22008
rect 42024 21980 42104 21984
rect 43257 21981 43269 21984
rect 43303 21981 43315 22015
rect 42024 21972 42030 21980
rect 43257 21975 43315 21981
rect 46566 21972 46572 22024
rect 46624 22012 46630 22024
rect 47854 22012 47860 22024
rect 46624 21984 47860 22012
rect 46624 21972 46630 21984
rect 47854 21972 47860 21984
rect 47912 22012 47918 22024
rect 47949 22015 48007 22021
rect 47949 22012 47961 22015
rect 47912 21984 47961 22012
rect 47912 21972 47918 21984
rect 47949 21981 47961 21984
rect 47995 21981 48007 22015
rect 47949 21975 48007 21981
rect 48593 22015 48651 22021
rect 48593 21981 48605 22015
rect 48639 22012 48651 22015
rect 48774 22012 48780 22024
rect 48639 21984 48780 22012
rect 48639 21981 48651 21984
rect 48593 21975 48651 21981
rect 48774 21972 48780 21984
rect 48832 21972 48838 22024
rect 45370 21944 45376 21956
rect 41892 21916 45376 21944
rect 45370 21904 45376 21916
rect 45428 21904 45434 21956
rect 49142 21904 49148 21956
rect 49200 21904 49206 21956
rect 40736 21848 41552 21876
rect 41601 21879 41659 21885
rect 40736 21836 40742 21848
rect 41601 21845 41613 21879
rect 41647 21876 41659 21879
rect 47670 21876 47676 21888
rect 41647 21848 47676 21876
rect 41647 21845 41659 21848
rect 41601 21839 41659 21845
rect 47670 21836 47676 21848
rect 47728 21836 47734 21888
rect 47762 21836 47768 21888
rect 47820 21836 47826 21888
rect 48406 21836 48412 21888
rect 48464 21836 48470 21888
rect 48498 21836 48504 21888
rect 48556 21876 48562 21888
rect 49237 21879 49295 21885
rect 49237 21876 49249 21879
rect 48556 21848 49249 21876
rect 48556 21836 48562 21848
rect 49237 21845 49249 21848
rect 49283 21845 49295 21879
rect 49237 21839 49295 21845
rect 1104 21786 49864 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 27950 21786
rect 28002 21734 28014 21786
rect 28066 21734 28078 21786
rect 28130 21734 28142 21786
rect 28194 21734 28206 21786
rect 28258 21734 37950 21786
rect 38002 21734 38014 21786
rect 38066 21734 38078 21786
rect 38130 21734 38142 21786
rect 38194 21734 38206 21786
rect 38258 21734 47950 21786
rect 48002 21734 48014 21786
rect 48066 21734 48078 21786
rect 48130 21734 48142 21786
rect 48194 21734 48206 21786
rect 48258 21734 49864 21786
rect 1104 21712 49864 21734
rect 4062 21632 4068 21684
rect 4120 21672 4126 21684
rect 4120 21644 8708 21672
rect 4120 21632 4126 21644
rect 4338 21564 4344 21616
rect 4396 21564 4402 21616
rect 8680 21604 8708 21644
rect 9766 21632 9772 21684
rect 9824 21672 9830 21684
rect 10505 21675 10563 21681
rect 10505 21672 10517 21675
rect 9824 21644 10517 21672
rect 9824 21632 9830 21644
rect 10505 21641 10517 21644
rect 10551 21641 10563 21675
rect 10505 21635 10563 21641
rect 12618 21632 12624 21684
rect 12676 21672 12682 21684
rect 13265 21675 13323 21681
rect 13265 21672 13277 21675
rect 12676 21644 13277 21672
rect 12676 21632 12682 21644
rect 13265 21641 13277 21644
rect 13311 21641 13323 21675
rect 13265 21635 13323 21641
rect 13906 21632 13912 21684
rect 13964 21632 13970 21684
rect 17034 21672 17040 21684
rect 14568 21644 17040 21672
rect 10042 21604 10048 21616
rect 8680 21576 10048 21604
rect 10042 21564 10048 21576
rect 10100 21564 10106 21616
rect 1765 21539 1823 21545
rect 1765 21505 1777 21539
rect 1811 21536 1823 21539
rect 1811 21508 3556 21536
rect 1811 21505 1823 21508
rect 1765 21499 1823 21505
rect 2777 21471 2835 21477
rect 2777 21437 2789 21471
rect 2823 21468 2835 21471
rect 3326 21468 3332 21480
rect 2823 21440 3332 21468
rect 2823 21437 2835 21440
rect 2777 21431 2835 21437
rect 3326 21428 3332 21440
rect 3384 21428 3390 21480
rect 3528 21400 3556 21508
rect 3602 21496 3608 21548
rect 3660 21496 3666 21548
rect 5902 21496 5908 21548
rect 5960 21496 5966 21548
rect 6549 21539 6607 21545
rect 6549 21505 6561 21539
rect 6595 21505 6607 21539
rect 6549 21499 6607 21505
rect 5258 21428 5264 21480
rect 5316 21468 5322 21480
rect 6564 21468 6592 21499
rect 8570 21496 8576 21548
rect 8628 21496 8634 21548
rect 10689 21539 10747 21545
rect 10689 21505 10701 21539
rect 10735 21505 10747 21539
rect 10689 21499 10747 21505
rect 11885 21539 11943 21545
rect 11885 21505 11897 21539
rect 11931 21536 11943 21539
rect 11974 21536 11980 21548
rect 11931 21508 11980 21536
rect 11931 21505 11943 21508
rect 11885 21499 11943 21505
rect 5316 21440 6592 21468
rect 5316 21428 5322 21440
rect 6730 21428 6736 21480
rect 6788 21468 6794 21480
rect 7009 21471 7067 21477
rect 7009 21468 7021 21471
rect 6788 21440 7021 21468
rect 6788 21428 6794 21440
rect 7009 21437 7021 21440
rect 7055 21437 7067 21471
rect 7009 21431 7067 21437
rect 8846 21428 8852 21480
rect 8904 21428 8910 21480
rect 10704 21468 10732 21499
rect 11974 21496 11980 21508
rect 12032 21536 12038 21548
rect 12253 21539 12311 21545
rect 12253 21536 12265 21539
rect 12032 21508 12265 21536
rect 12032 21496 12038 21508
rect 12253 21505 12265 21508
rect 12299 21505 12311 21539
rect 12253 21499 12311 21505
rect 12802 21496 12808 21548
rect 12860 21496 12866 21548
rect 13173 21539 13231 21545
rect 13173 21505 13185 21539
rect 13219 21536 13231 21539
rect 13998 21536 14004 21548
rect 13219 21508 14004 21536
rect 13219 21505 13231 21508
rect 13173 21499 13231 21505
rect 13998 21496 14004 21508
rect 14056 21496 14062 21548
rect 14093 21539 14151 21545
rect 14093 21505 14105 21539
rect 14139 21505 14151 21539
rect 14093 21499 14151 21505
rect 13446 21468 13452 21480
rect 10704 21440 13452 21468
rect 13446 21428 13452 21440
rect 13504 21428 13510 21480
rect 14108 21468 14136 21499
rect 14274 21496 14280 21548
rect 14332 21536 14338 21548
rect 14568 21545 14596 21644
rect 17034 21632 17040 21644
rect 17092 21632 17098 21684
rect 17129 21675 17187 21681
rect 17129 21641 17141 21675
rect 17175 21672 17187 21675
rect 17678 21672 17684 21684
rect 17175 21644 17684 21672
rect 17175 21641 17187 21644
rect 17129 21635 17187 21641
rect 14826 21564 14832 21616
rect 14884 21564 14890 21616
rect 16758 21604 16764 21616
rect 16054 21576 16764 21604
rect 16758 21564 16764 21576
rect 16816 21604 16822 21616
rect 16945 21607 17003 21613
rect 16945 21604 16957 21607
rect 16816 21576 16957 21604
rect 16816 21564 16822 21576
rect 16945 21573 16957 21576
rect 16991 21604 17003 21607
rect 17144 21604 17172 21635
rect 17678 21632 17684 21644
rect 17736 21632 17742 21684
rect 17862 21632 17868 21684
rect 17920 21632 17926 21684
rect 20530 21672 20536 21684
rect 18432 21644 20536 21672
rect 16991 21576 17172 21604
rect 16991 21573 17003 21576
rect 16945 21567 17003 21573
rect 14553 21539 14611 21545
rect 14553 21536 14565 21539
rect 14332 21508 14565 21536
rect 14332 21496 14338 21508
rect 14553 21505 14565 21508
rect 14599 21505 14611 21539
rect 14553 21499 14611 21505
rect 17773 21539 17831 21545
rect 17773 21505 17785 21539
rect 17819 21536 17831 21539
rect 18322 21536 18328 21548
rect 17819 21508 18328 21536
rect 17819 21505 17831 21508
rect 17773 21499 17831 21505
rect 18322 21496 18328 21508
rect 18380 21496 18386 21548
rect 16114 21468 16120 21480
rect 14108 21440 16120 21468
rect 16114 21428 16120 21440
rect 16172 21428 16178 21480
rect 18049 21471 18107 21477
rect 18049 21437 18061 21471
rect 18095 21468 18107 21471
rect 18432 21468 18460 21644
rect 20530 21632 20536 21644
rect 20588 21632 20594 21684
rect 21910 21632 21916 21684
rect 21968 21672 21974 21684
rect 22278 21672 22284 21684
rect 21968 21644 22284 21672
rect 21968 21632 21974 21644
rect 22278 21632 22284 21644
rect 22336 21632 22342 21684
rect 26421 21675 26479 21681
rect 26421 21672 26433 21675
rect 22388 21644 26433 21672
rect 20714 21604 20720 21616
rect 20102 21576 20720 21604
rect 20714 21564 20720 21576
rect 20772 21564 20778 21616
rect 21269 21539 21327 21545
rect 21269 21505 21281 21539
rect 21315 21536 21327 21539
rect 21315 21508 22094 21536
rect 21315 21505 21327 21508
rect 21269 21499 21327 21505
rect 18095 21440 18460 21468
rect 18095 21437 18107 21440
rect 18049 21431 18107 21437
rect 18598 21428 18604 21480
rect 18656 21428 18662 21480
rect 18874 21428 18880 21480
rect 18932 21428 18938 21480
rect 22066 21468 22094 21508
rect 22388 21468 22416 21644
rect 26421 21641 26433 21644
rect 26467 21641 26479 21675
rect 26421 21635 26479 21641
rect 27798 21632 27804 21684
rect 27856 21672 27862 21684
rect 28353 21675 28411 21681
rect 28353 21672 28365 21675
rect 27856 21644 28365 21672
rect 27856 21632 27862 21644
rect 28353 21641 28365 21644
rect 28399 21641 28411 21675
rect 28353 21635 28411 21641
rect 30009 21675 30067 21681
rect 30009 21641 30021 21675
rect 30055 21672 30067 21675
rect 32398 21672 32404 21684
rect 30055 21644 32404 21672
rect 30055 21641 30067 21644
rect 30009 21635 30067 21641
rect 32398 21632 32404 21644
rect 32456 21632 32462 21684
rect 32585 21675 32643 21681
rect 32585 21641 32597 21675
rect 32631 21672 32643 21675
rect 33410 21672 33416 21684
rect 32631 21644 33416 21672
rect 32631 21641 32643 21644
rect 32585 21635 32643 21641
rect 33410 21632 33416 21644
rect 33468 21632 33474 21684
rect 34425 21675 34483 21681
rect 34425 21641 34437 21675
rect 34471 21641 34483 21675
rect 34425 21635 34483 21641
rect 22738 21564 22744 21616
rect 22796 21564 22802 21616
rect 23198 21564 23204 21616
rect 23256 21564 23262 21616
rect 25038 21564 25044 21616
rect 25096 21604 25102 21616
rect 26970 21604 26976 21616
rect 25096 21576 26976 21604
rect 25096 21564 25102 21576
rect 26970 21564 26976 21576
rect 27028 21564 27034 21616
rect 27080 21576 27384 21604
rect 25133 21539 25191 21545
rect 25133 21505 25145 21539
rect 25179 21536 25191 21539
rect 25866 21536 25872 21548
rect 25179 21508 25872 21536
rect 25179 21505 25191 21508
rect 25133 21499 25191 21505
rect 25866 21496 25872 21508
rect 25924 21496 25930 21548
rect 26605 21539 26663 21545
rect 26605 21505 26617 21539
rect 26651 21536 26663 21539
rect 26878 21536 26884 21548
rect 26651 21508 26884 21536
rect 26651 21505 26663 21508
rect 26605 21499 26663 21505
rect 26878 21496 26884 21508
rect 26936 21496 26942 21548
rect 22066 21440 22416 21468
rect 22462 21428 22468 21480
rect 22520 21428 22526 21480
rect 22572 21440 24900 21468
rect 5626 21400 5632 21412
rect 3528 21372 5632 21400
rect 5626 21360 5632 21372
rect 5684 21360 5690 21412
rect 5721 21403 5779 21409
rect 5721 21369 5733 21403
rect 5767 21400 5779 21403
rect 8570 21400 8576 21412
rect 5767 21372 8576 21400
rect 5767 21369 5779 21372
rect 5721 21363 5779 21369
rect 8570 21360 8576 21372
rect 8628 21360 8634 21412
rect 12437 21403 12495 21409
rect 12437 21400 12449 21403
rect 8680 21372 12449 21400
rect 4338 21292 4344 21344
rect 4396 21332 4402 21344
rect 8680 21332 8708 21372
rect 12437 21369 12449 21372
rect 12483 21369 12495 21403
rect 17405 21403 17463 21409
rect 17405 21400 17417 21403
rect 12437 21363 12495 21369
rect 12636 21372 12848 21400
rect 4396 21304 8708 21332
rect 4396 21292 4402 21304
rect 8754 21292 8760 21344
rect 8812 21332 8818 21344
rect 9950 21332 9956 21344
rect 8812 21304 9956 21332
rect 8812 21292 8818 21304
rect 9950 21292 9956 21304
rect 10008 21292 10014 21344
rect 11882 21292 11888 21344
rect 11940 21332 11946 21344
rect 12636 21332 12664 21372
rect 11940 21304 12664 21332
rect 12820 21332 12848 21372
rect 15856 21372 17417 21400
rect 15856 21332 15884 21372
rect 17405 21369 17417 21372
rect 17451 21369 17463 21403
rect 21453 21403 21511 21409
rect 21453 21400 21465 21403
rect 17405 21363 17463 21369
rect 19904 21372 21465 21400
rect 12820 21304 15884 21332
rect 11940 21292 11946 21304
rect 16298 21292 16304 21344
rect 16356 21292 16362 21344
rect 18690 21292 18696 21344
rect 18748 21332 18754 21344
rect 19904 21332 19932 21372
rect 21453 21369 21465 21372
rect 21499 21369 21511 21403
rect 21453 21363 21511 21369
rect 22278 21360 22284 21412
rect 22336 21400 22342 21412
rect 22572 21400 22600 21440
rect 22336 21372 22600 21400
rect 22336 21360 22342 21372
rect 24762 21360 24768 21412
rect 24820 21360 24826 21412
rect 24872 21400 24900 21440
rect 25222 21428 25228 21480
rect 25280 21428 25286 21480
rect 25314 21428 25320 21480
rect 25372 21468 25378 21480
rect 25409 21471 25467 21477
rect 25409 21468 25421 21471
rect 25372 21440 25421 21468
rect 25372 21428 25378 21440
rect 25409 21437 25421 21440
rect 25455 21468 25467 21471
rect 27080 21468 27108 21576
rect 25455 21440 27108 21468
rect 27356 21468 27384 21576
rect 27430 21564 27436 21616
rect 27488 21604 27494 21616
rect 27617 21607 27675 21613
rect 27617 21604 27629 21607
rect 27488 21576 27629 21604
rect 27488 21564 27494 21576
rect 27617 21573 27629 21576
rect 27663 21573 27675 21607
rect 27617 21567 27675 21573
rect 27706 21564 27712 21616
rect 27764 21604 27770 21616
rect 29822 21604 29828 21616
rect 27764 21576 29828 21604
rect 27764 21564 27770 21576
rect 29822 21564 29828 21576
rect 29880 21564 29886 21616
rect 31202 21564 31208 21616
rect 31260 21564 31266 21616
rect 31570 21564 31576 21616
rect 31628 21604 31634 21616
rect 32858 21604 32864 21616
rect 31628 21576 32864 21604
rect 31628 21564 31634 21576
rect 32858 21564 32864 21576
rect 32916 21564 32922 21616
rect 34440 21604 34468 21635
rect 34882 21632 34888 21684
rect 34940 21632 34946 21684
rect 35066 21632 35072 21684
rect 35124 21672 35130 21684
rect 35894 21672 35900 21684
rect 35124 21644 35900 21672
rect 35124 21632 35130 21644
rect 35894 21632 35900 21644
rect 35952 21632 35958 21684
rect 36081 21675 36139 21681
rect 36081 21641 36093 21675
rect 36127 21672 36139 21675
rect 40034 21672 40040 21684
rect 36127 21644 40040 21672
rect 36127 21641 36139 21644
rect 36081 21635 36139 21641
rect 40034 21632 40040 21644
rect 40092 21632 40098 21684
rect 40126 21632 40132 21684
rect 40184 21672 40190 21684
rect 40221 21675 40279 21681
rect 40221 21672 40233 21675
rect 40184 21644 40233 21672
rect 40184 21632 40190 21644
rect 40221 21641 40233 21644
rect 40267 21641 40279 21675
rect 40221 21635 40279 21641
rect 40402 21632 40408 21684
rect 40460 21672 40466 21684
rect 41969 21675 42027 21681
rect 40460 21644 41920 21672
rect 40460 21632 40466 21644
rect 36446 21604 36452 21616
rect 34440 21576 36452 21604
rect 36446 21564 36452 21576
rect 36504 21564 36510 21616
rect 36630 21564 36636 21616
rect 36688 21604 36694 21616
rect 36817 21607 36875 21613
rect 36817 21604 36829 21607
rect 36688 21576 36829 21604
rect 36688 21564 36694 21576
rect 36817 21573 36829 21576
rect 36863 21604 36875 21607
rect 38378 21604 38384 21616
rect 36863 21576 38384 21604
rect 36863 21573 36875 21576
rect 36817 21567 36875 21573
rect 38378 21564 38384 21576
rect 38436 21564 38442 21616
rect 38838 21564 38844 21616
rect 38896 21564 38902 21616
rect 39850 21564 39856 21616
rect 39908 21604 39914 21616
rect 40589 21607 40647 21613
rect 40589 21604 40601 21607
rect 39908 21576 40601 21604
rect 39908 21564 39914 21576
rect 40589 21573 40601 21576
rect 40635 21573 40647 21607
rect 41230 21604 41236 21616
rect 40589 21567 40647 21573
rect 40696 21576 41236 21604
rect 27525 21539 27583 21545
rect 27525 21505 27537 21539
rect 27571 21536 27583 21539
rect 27571 21508 28672 21536
rect 27571 21505 27583 21508
rect 27525 21499 27583 21505
rect 27709 21471 27767 21477
rect 27709 21468 27721 21471
rect 27356 21440 27721 21468
rect 25455 21437 25467 21440
rect 25409 21431 25467 21437
rect 27709 21437 27721 21440
rect 27755 21437 27767 21471
rect 27709 21431 27767 21437
rect 27157 21403 27215 21409
rect 27157 21400 27169 21403
rect 24872 21372 27169 21400
rect 27157 21369 27169 21372
rect 27203 21369 27215 21403
rect 28644 21400 28672 21508
rect 28718 21496 28724 21548
rect 28776 21496 28782 21548
rect 28810 21496 28816 21548
rect 28868 21496 28874 21548
rect 29917 21539 29975 21545
rect 29917 21505 29929 21539
rect 29963 21536 29975 21539
rect 31113 21539 31171 21545
rect 29963 21508 30880 21536
rect 29963 21505 29975 21508
rect 29917 21499 29975 21505
rect 28902 21428 28908 21480
rect 28960 21428 28966 21480
rect 29270 21428 29276 21480
rect 29328 21468 29334 21480
rect 30101 21471 30159 21477
rect 30101 21468 30113 21471
rect 29328 21440 30113 21468
rect 29328 21428 29334 21440
rect 30101 21437 30113 21440
rect 30147 21437 30159 21471
rect 30101 21431 30159 21437
rect 29086 21400 29092 21412
rect 28644 21372 29092 21400
rect 27157 21363 27215 21369
rect 29086 21360 29092 21372
rect 29144 21400 29150 21412
rect 29914 21400 29920 21412
rect 29144 21372 29920 21400
rect 29144 21360 29150 21372
rect 29914 21360 29920 21372
rect 29972 21360 29978 21412
rect 18748 21304 19932 21332
rect 18748 21292 18754 21304
rect 20346 21292 20352 21344
rect 20404 21292 20410 21344
rect 20714 21292 20720 21344
rect 20772 21332 20778 21344
rect 21910 21332 21916 21344
rect 20772 21304 21916 21332
rect 20772 21292 20778 21304
rect 21910 21292 21916 21304
rect 21968 21332 21974 21344
rect 22097 21335 22155 21341
rect 22097 21332 22109 21335
rect 21968 21304 22109 21332
rect 21968 21292 21974 21304
rect 22097 21301 22109 21304
rect 22143 21332 22155 21335
rect 23198 21332 23204 21344
rect 22143 21304 23204 21332
rect 22143 21301 22155 21304
rect 22097 21295 22155 21301
rect 23198 21292 23204 21304
rect 23256 21292 23262 21344
rect 24213 21335 24271 21341
rect 24213 21301 24225 21335
rect 24259 21332 24271 21335
rect 25406 21332 25412 21344
rect 24259 21304 25412 21332
rect 24259 21301 24271 21304
rect 24213 21295 24271 21301
rect 25406 21292 25412 21304
rect 25464 21292 25470 21344
rect 25866 21292 25872 21344
rect 25924 21292 25930 21344
rect 26053 21335 26111 21341
rect 26053 21301 26065 21335
rect 26099 21332 26111 21335
rect 26142 21332 26148 21344
rect 26099 21304 26148 21332
rect 26099 21301 26111 21304
rect 26053 21295 26111 21301
rect 26142 21292 26148 21304
rect 26200 21332 26206 21344
rect 26326 21332 26332 21344
rect 26200 21304 26332 21332
rect 26200 21292 26206 21304
rect 26326 21292 26332 21304
rect 26384 21292 26390 21344
rect 29546 21292 29552 21344
rect 29604 21292 29610 21344
rect 30650 21292 30656 21344
rect 30708 21332 30714 21344
rect 30745 21335 30803 21341
rect 30745 21332 30757 21335
rect 30708 21304 30757 21332
rect 30708 21292 30714 21304
rect 30745 21301 30757 21304
rect 30791 21301 30803 21335
rect 30852 21332 30880 21508
rect 31113 21505 31125 21539
rect 31159 21536 31171 21539
rect 33594 21536 33600 21548
rect 31159 21508 33600 21536
rect 31159 21505 31171 21508
rect 31113 21499 31171 21505
rect 33594 21496 33600 21508
rect 33652 21496 33658 21548
rect 33686 21496 33692 21548
rect 33744 21496 33750 21548
rect 34790 21496 34796 21548
rect 34848 21496 34854 21548
rect 36722 21536 36728 21548
rect 35084 21508 36728 21536
rect 31389 21471 31447 21477
rect 31389 21437 31401 21471
rect 31435 21468 31447 21471
rect 31570 21468 31576 21480
rect 31435 21440 31576 21468
rect 31435 21437 31447 21440
rect 31389 21431 31447 21437
rect 31570 21428 31576 21440
rect 31628 21428 31634 21480
rect 33410 21428 33416 21480
rect 33468 21468 33474 21480
rect 35084 21477 35112 21508
rect 36722 21496 36728 21508
rect 36780 21496 36786 21548
rect 33781 21471 33839 21477
rect 33781 21468 33793 21471
rect 33468 21440 33793 21468
rect 33468 21428 33474 21440
rect 33781 21437 33793 21440
rect 33827 21437 33839 21471
rect 33781 21431 33839 21437
rect 35069 21471 35127 21477
rect 35069 21437 35081 21471
rect 35115 21437 35127 21471
rect 35069 21431 35127 21437
rect 36170 21428 36176 21480
rect 36228 21428 36234 21480
rect 36265 21471 36323 21477
rect 36265 21437 36277 21471
rect 36311 21468 36323 21471
rect 36630 21468 36636 21480
rect 36311 21440 36636 21468
rect 36311 21437 36323 21440
rect 36265 21431 36323 21437
rect 36630 21428 36636 21440
rect 36688 21428 36694 21480
rect 37734 21428 37740 21480
rect 37792 21468 37798 21480
rect 38013 21471 38071 21477
rect 38013 21468 38025 21471
rect 37792 21440 38025 21468
rect 37792 21428 37798 21440
rect 38013 21437 38025 21440
rect 38059 21437 38071 21471
rect 38286 21468 38292 21480
rect 38013 21431 38071 21437
rect 38120 21440 38292 21468
rect 33229 21403 33287 21409
rect 33229 21369 33241 21403
rect 33275 21400 33287 21403
rect 36354 21400 36360 21412
rect 33275 21372 36360 21400
rect 33275 21369 33287 21372
rect 33229 21363 33287 21369
rect 36354 21360 36360 21372
rect 36412 21360 36418 21412
rect 37458 21360 37464 21412
rect 37516 21400 37522 21412
rect 38120 21400 38148 21440
rect 38286 21428 38292 21440
rect 38344 21428 38350 21480
rect 38378 21428 38384 21480
rect 38436 21468 38442 21480
rect 40696 21477 40724 21576
rect 41230 21564 41236 21576
rect 41288 21604 41294 21616
rect 41782 21604 41788 21616
rect 41288 21576 41788 21604
rect 41288 21564 41294 21576
rect 41782 21564 41788 21576
rect 41840 21564 41846 21616
rect 41892 21604 41920 21644
rect 41969 21641 41981 21675
rect 42015 21672 42027 21675
rect 42242 21672 42248 21684
rect 42015 21644 42248 21672
rect 42015 21641 42027 21644
rect 41969 21635 42027 21641
rect 42242 21632 42248 21644
rect 42300 21632 42306 21684
rect 42521 21675 42579 21681
rect 42521 21641 42533 21675
rect 42567 21672 42579 21675
rect 42886 21672 42892 21684
rect 42567 21644 42892 21672
rect 42567 21641 42579 21644
rect 42521 21635 42579 21641
rect 42886 21632 42892 21644
rect 42944 21672 42950 21684
rect 43990 21672 43996 21684
rect 42944 21644 43996 21672
rect 42944 21632 42950 21644
rect 43990 21632 43996 21644
rect 44048 21632 44054 21684
rect 47486 21632 47492 21684
rect 47544 21672 47550 21684
rect 47857 21675 47915 21681
rect 47857 21672 47869 21675
rect 47544 21644 47869 21672
rect 47544 21632 47550 21644
rect 47857 21641 47869 21644
rect 47903 21641 47915 21675
rect 47857 21635 47915 21641
rect 48774 21632 48780 21684
rect 48832 21632 48838 21684
rect 49050 21632 49056 21684
rect 49108 21632 49114 21684
rect 47762 21604 47768 21616
rect 41892 21576 47768 21604
rect 47762 21564 47768 21576
rect 47820 21564 47826 21616
rect 48409 21607 48467 21613
rect 48409 21573 48421 21607
rect 48455 21604 48467 21607
rect 49068 21604 49096 21632
rect 48455 21576 49096 21604
rect 48455 21573 48467 21576
rect 48409 21567 48467 21573
rect 40862 21496 40868 21548
rect 40920 21536 40926 21548
rect 41601 21539 41659 21545
rect 41601 21536 41613 21539
rect 40920 21508 41613 21536
rect 40920 21496 40926 21508
rect 41601 21505 41613 21508
rect 41647 21536 41659 21539
rect 42613 21539 42671 21545
rect 42613 21536 42625 21539
rect 41647 21508 42625 21536
rect 41647 21505 41659 21508
rect 41601 21499 41659 21505
rect 42613 21505 42625 21508
rect 42659 21505 42671 21539
rect 42613 21499 42671 21505
rect 47854 21496 47860 21548
rect 47912 21536 47918 21548
rect 48041 21539 48099 21545
rect 48041 21536 48053 21539
rect 47912 21508 48053 21536
rect 47912 21496 47918 21508
rect 48041 21505 48053 21508
rect 48087 21505 48099 21539
rect 48041 21499 48099 21505
rect 48593 21539 48651 21545
rect 48593 21505 48605 21539
rect 48639 21536 48651 21539
rect 49050 21536 49056 21548
rect 48639 21508 49056 21536
rect 48639 21505 48651 21508
rect 48593 21499 48651 21505
rect 49050 21496 49056 21508
rect 49108 21496 49114 21548
rect 40681 21471 40739 21477
rect 40681 21468 40693 21471
rect 38436 21440 40693 21468
rect 38436 21428 38442 21440
rect 40681 21437 40693 21440
rect 40727 21437 40739 21471
rect 40681 21431 40739 21437
rect 40770 21428 40776 21480
rect 40828 21428 40834 21480
rect 40880 21440 41736 21468
rect 37516 21372 38148 21400
rect 37516 21360 37522 21372
rect 40034 21360 40040 21412
rect 40092 21400 40098 21412
rect 40494 21400 40500 21412
rect 40092 21372 40500 21400
rect 40092 21360 40098 21372
rect 40494 21360 40500 21372
rect 40552 21360 40558 21412
rect 32674 21332 32680 21344
rect 30852 21304 32680 21332
rect 30745 21295 30803 21301
rect 32674 21292 32680 21304
rect 32732 21332 32738 21344
rect 34330 21332 34336 21344
rect 32732 21304 34336 21332
rect 32732 21292 32738 21304
rect 34330 21292 34336 21304
rect 34388 21292 34394 21344
rect 34514 21292 34520 21344
rect 34572 21332 34578 21344
rect 35713 21335 35771 21341
rect 35713 21332 35725 21335
rect 34572 21304 35725 21332
rect 34572 21292 34578 21304
rect 35713 21301 35725 21304
rect 35759 21301 35771 21335
rect 35713 21295 35771 21301
rect 37274 21292 37280 21344
rect 37332 21332 37338 21344
rect 39758 21332 39764 21344
rect 37332 21304 39764 21332
rect 37332 21292 37338 21304
rect 39758 21292 39764 21304
rect 39816 21292 39822 21344
rect 39850 21292 39856 21344
rect 39908 21332 39914 21344
rect 40880 21332 40908 21440
rect 41414 21360 41420 21412
rect 41472 21360 41478 21412
rect 41708 21400 41736 21440
rect 41782 21428 41788 21480
rect 41840 21468 41846 21480
rect 42886 21468 42892 21480
rect 41840 21440 42892 21468
rect 41840 21428 41846 21440
rect 42886 21428 42892 21440
rect 42944 21428 42950 21480
rect 42153 21403 42211 21409
rect 42153 21400 42165 21403
rect 41708 21372 42165 21400
rect 42153 21369 42165 21372
rect 42199 21400 42211 21403
rect 46198 21400 46204 21412
rect 42199 21372 46204 21400
rect 42199 21369 42211 21372
rect 42153 21363 42211 21369
rect 46198 21360 46204 21372
rect 46256 21360 46262 21412
rect 39908 21304 40908 21332
rect 39908 21292 39914 21304
rect 49234 21292 49240 21344
rect 49292 21292 49298 21344
rect 1104 21242 49864 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 32950 21242
rect 33002 21190 33014 21242
rect 33066 21190 33078 21242
rect 33130 21190 33142 21242
rect 33194 21190 33206 21242
rect 33258 21190 42950 21242
rect 43002 21190 43014 21242
rect 43066 21190 43078 21242
rect 43130 21190 43142 21242
rect 43194 21190 43206 21242
rect 43258 21190 49864 21242
rect 1104 21168 49864 21190
rect 2746 21100 6408 21128
rect 2746 20992 2774 21100
rect 1780 20964 2774 20992
rect 1780 20933 1808 20964
rect 4246 20952 4252 21004
rect 4304 20992 4310 21004
rect 4433 20995 4491 21001
rect 4433 20992 4445 20995
rect 4304 20964 4445 20992
rect 4304 20952 4310 20964
rect 4433 20961 4445 20964
rect 4479 20961 4491 20995
rect 4433 20955 4491 20961
rect 5534 20952 5540 21004
rect 5592 20992 5598 21004
rect 6273 20995 6331 21001
rect 6273 20992 6285 20995
rect 5592 20964 6285 20992
rect 5592 20952 5598 20964
rect 6273 20961 6285 20964
rect 6319 20961 6331 20995
rect 6273 20955 6331 20961
rect 1765 20927 1823 20933
rect 1765 20893 1777 20927
rect 1811 20893 1823 20927
rect 1765 20887 1823 20893
rect 4157 20927 4215 20933
rect 4157 20893 4169 20927
rect 4203 20924 4215 20927
rect 4338 20924 4344 20936
rect 4203 20896 4344 20924
rect 4203 20893 4215 20896
rect 4157 20887 4215 20893
rect 4338 20884 4344 20896
rect 4396 20884 4402 20936
rect 5905 20927 5963 20933
rect 5905 20893 5917 20927
rect 5951 20893 5963 20927
rect 5905 20887 5963 20893
rect 2774 20816 2780 20868
rect 2832 20816 2838 20868
rect 5920 20788 5948 20887
rect 6380 20856 6408 21100
rect 7742 21088 7748 21140
rect 7800 21128 7806 21140
rect 9217 21131 9275 21137
rect 9217 21128 9229 21131
rect 7800 21100 9229 21128
rect 7800 21088 7806 21100
rect 9217 21097 9229 21100
rect 9263 21097 9275 21131
rect 11977 21131 12035 21137
rect 11977 21128 11989 21131
rect 9217 21091 9275 21097
rect 9324 21100 11989 21128
rect 6454 21020 6460 21072
rect 6512 21060 6518 21072
rect 9324 21060 9352 21100
rect 11977 21097 11989 21100
rect 12023 21097 12035 21131
rect 11977 21091 12035 21097
rect 12434 21088 12440 21140
rect 12492 21128 12498 21140
rect 12897 21131 12955 21137
rect 12897 21128 12909 21131
rect 12492 21100 12909 21128
rect 12492 21088 12498 21100
rect 12897 21097 12909 21100
rect 12943 21097 12955 21131
rect 12897 21091 12955 21097
rect 12986 21088 12992 21140
rect 13044 21128 13050 21140
rect 16574 21128 16580 21140
rect 13044 21100 16580 21128
rect 13044 21088 13050 21100
rect 16574 21088 16580 21100
rect 16632 21088 16638 21140
rect 17392 21131 17450 21137
rect 17392 21097 17404 21131
rect 17438 21128 17450 21131
rect 18966 21128 18972 21140
rect 17438 21100 18972 21128
rect 17438 21097 17450 21100
rect 17392 21091 17450 21097
rect 18966 21088 18972 21100
rect 19024 21088 19030 21140
rect 19150 21088 19156 21140
rect 19208 21128 19214 21140
rect 19337 21131 19395 21137
rect 19337 21128 19349 21131
rect 19208 21100 19349 21128
rect 19208 21088 19214 21100
rect 19337 21097 19349 21100
rect 19383 21128 19395 21131
rect 20714 21128 20720 21140
rect 19383 21100 20720 21128
rect 19383 21097 19395 21100
rect 19337 21091 19395 21097
rect 20714 21088 20720 21100
rect 20772 21088 20778 21140
rect 21266 21088 21272 21140
rect 21324 21128 21330 21140
rect 21434 21131 21492 21137
rect 21434 21128 21446 21131
rect 21324 21100 21446 21128
rect 21324 21088 21330 21100
rect 21434 21097 21446 21100
rect 21480 21097 21492 21131
rect 21434 21091 21492 21097
rect 21542 21088 21548 21140
rect 21600 21128 21606 21140
rect 22646 21128 22652 21140
rect 21600 21100 22652 21128
rect 21600 21088 21606 21100
rect 22646 21088 22652 21100
rect 22704 21088 22710 21140
rect 22830 21088 22836 21140
rect 22888 21128 22894 21140
rect 23569 21131 23627 21137
rect 23569 21128 23581 21131
rect 22888 21100 23581 21128
rect 22888 21088 22894 21100
rect 23569 21097 23581 21100
rect 23615 21097 23627 21131
rect 23569 21091 23627 21097
rect 24029 21131 24087 21137
rect 24029 21097 24041 21131
rect 24075 21128 24087 21131
rect 24670 21128 24676 21140
rect 24075 21100 24676 21128
rect 24075 21097 24087 21100
rect 24029 21091 24087 21097
rect 24670 21088 24676 21100
rect 24728 21128 24734 21140
rect 25317 21131 25375 21137
rect 25317 21128 25329 21131
rect 24728 21100 25329 21128
rect 24728 21088 24734 21100
rect 25317 21097 25329 21100
rect 25363 21097 25375 21131
rect 25317 21091 25375 21097
rect 26694 21088 26700 21140
rect 26752 21088 26758 21140
rect 27154 21088 27160 21140
rect 27212 21128 27218 21140
rect 27798 21128 27804 21140
rect 27212 21100 27804 21128
rect 27212 21088 27218 21100
rect 27798 21088 27804 21100
rect 27856 21088 27862 21140
rect 28353 21131 28411 21137
rect 28353 21097 28365 21131
rect 28399 21128 28411 21131
rect 30098 21128 30104 21140
rect 28399 21100 30104 21128
rect 28399 21097 28411 21100
rect 28353 21091 28411 21097
rect 30098 21088 30104 21100
rect 30156 21088 30162 21140
rect 30374 21088 30380 21140
rect 30432 21128 30438 21140
rect 31386 21128 31392 21140
rect 30432 21100 31392 21128
rect 30432 21088 30438 21100
rect 31386 21088 31392 21100
rect 31444 21088 31450 21140
rect 34514 21128 34520 21140
rect 31726 21100 34520 21128
rect 10502 21060 10508 21072
rect 6512 21032 9352 21060
rect 9416 21032 10508 21060
rect 6512 21020 6518 21032
rect 9416 20992 9444 21032
rect 10502 21020 10508 21032
rect 10560 21020 10566 21072
rect 12802 21060 12808 21072
rect 11900 21032 12808 21060
rect 11790 20992 11796 21004
rect 8036 20964 9444 20992
rect 9784 20964 11796 20992
rect 8036 20933 8064 20964
rect 8021 20927 8079 20933
rect 8021 20893 8033 20927
rect 8067 20893 8079 20927
rect 8021 20887 8079 20893
rect 9401 20927 9459 20933
rect 9401 20893 9413 20927
rect 9447 20924 9459 20927
rect 9784 20924 9812 20964
rect 11790 20952 11796 20964
rect 11848 20952 11854 21004
rect 9447 20896 9812 20924
rect 9447 20893 9459 20896
rect 9401 20887 9459 20893
rect 9858 20884 9864 20936
rect 9916 20884 9922 20936
rect 11238 20924 11244 20936
rect 9968 20896 11244 20924
rect 9968 20856 9996 20896
rect 11238 20884 11244 20896
rect 11296 20884 11302 20936
rect 11330 20884 11336 20936
rect 11388 20884 11394 20936
rect 11900 20933 11928 21032
rect 12802 21020 12808 21032
rect 12860 21060 12866 21072
rect 13722 21060 13728 21072
rect 12860 21032 13728 21060
rect 12860 21020 12866 21032
rect 13722 21020 13728 21032
rect 13780 21020 13786 21072
rect 19981 21063 20039 21069
rect 19981 21029 19993 21063
rect 20027 21029 20039 21063
rect 19981 21023 20039 21029
rect 13630 20992 13636 21004
rect 12406 20964 13636 20992
rect 11885 20927 11943 20933
rect 11885 20893 11897 20927
rect 11931 20893 11943 20927
rect 12406 20924 12434 20964
rect 13630 20952 13636 20964
rect 13688 20952 13694 21004
rect 19996 20992 20024 21023
rect 23842 21020 23848 21072
rect 23900 21060 23906 21072
rect 25685 21063 25743 21069
rect 25685 21060 25697 21063
rect 23900 21032 25697 21060
rect 23900 21020 23906 21032
rect 25685 21029 25697 21032
rect 25731 21029 25743 21063
rect 29546 21060 29552 21072
rect 25685 21023 25743 21029
rect 26160 21032 29552 21060
rect 13740 20964 20024 20992
rect 13740 20933 13768 20964
rect 20438 20952 20444 21004
rect 20496 20992 20502 21004
rect 20533 20995 20591 21001
rect 20533 20992 20545 20995
rect 20496 20964 20545 20992
rect 20496 20952 20502 20964
rect 20533 20961 20545 20964
rect 20579 20992 20591 20995
rect 22925 20995 22983 21001
rect 22925 20992 22937 20995
rect 20579 20964 22937 20992
rect 20579 20961 20591 20964
rect 20533 20955 20591 20961
rect 22925 20961 22937 20964
rect 22971 20961 22983 20995
rect 25590 20992 25596 21004
rect 22925 20955 22983 20961
rect 23492 20964 25596 20992
rect 13725 20927 13783 20933
rect 11885 20887 11943 20893
rect 11992 20896 12434 20924
rect 12728 20896 13584 20924
rect 6380 20828 9996 20856
rect 10505 20859 10563 20865
rect 10505 20825 10517 20859
rect 10551 20856 10563 20859
rect 11992 20856 12020 20896
rect 10551 20828 12020 20856
rect 10551 20825 10563 20828
rect 10505 20819 10563 20825
rect 12066 20816 12072 20868
rect 12124 20856 12130 20868
rect 12728 20856 12756 20896
rect 12124 20828 12756 20856
rect 12124 20816 12130 20828
rect 12802 20816 12808 20868
rect 12860 20816 12866 20868
rect 7837 20791 7895 20797
rect 7837 20788 7849 20791
rect 5920 20760 7849 20788
rect 7837 20757 7849 20760
rect 7883 20757 7895 20791
rect 7837 20751 7895 20757
rect 11054 20748 11060 20800
rect 11112 20788 11118 20800
rect 11149 20791 11207 20797
rect 11149 20788 11161 20791
rect 11112 20760 11161 20788
rect 11112 20748 11118 20760
rect 11149 20757 11161 20760
rect 11195 20757 11207 20791
rect 11149 20751 11207 20757
rect 12434 20748 12440 20800
rect 12492 20788 12498 20800
rect 12986 20788 12992 20800
rect 12492 20760 12992 20788
rect 12492 20748 12498 20760
rect 12986 20748 12992 20760
rect 13044 20748 13050 20800
rect 13556 20797 13584 20896
rect 13725 20893 13737 20927
rect 13771 20893 13783 20927
rect 13725 20887 13783 20893
rect 14274 20884 14280 20936
rect 14332 20884 14338 20936
rect 17034 20884 17040 20936
rect 17092 20924 17098 20936
rect 17129 20927 17187 20933
rect 17129 20924 17141 20927
rect 17092 20896 17141 20924
rect 17092 20884 17098 20896
rect 17129 20893 17141 20896
rect 17175 20893 17187 20927
rect 17129 20887 17187 20893
rect 20349 20927 20407 20933
rect 20349 20893 20361 20927
rect 20395 20924 20407 20927
rect 21082 20924 21088 20936
rect 20395 20896 21088 20924
rect 20395 20893 20407 20896
rect 20349 20887 20407 20893
rect 21082 20884 21088 20896
rect 21140 20884 21146 20936
rect 21174 20884 21180 20936
rect 21232 20884 21238 20936
rect 23492 20933 23520 20964
rect 25590 20952 25596 20964
rect 25648 20952 25654 21004
rect 26160 21001 26188 21032
rect 29546 21020 29552 21032
rect 29604 21020 29610 21072
rect 30466 21060 30472 21072
rect 29748 21032 30472 21060
rect 26145 20995 26203 21001
rect 26145 20961 26157 20995
rect 26191 20961 26203 20995
rect 26145 20955 26203 20961
rect 26237 20995 26295 21001
rect 26237 20961 26249 20995
rect 26283 20961 26295 20995
rect 26237 20955 26295 20961
rect 27709 20995 27767 21001
rect 27709 20961 27721 20995
rect 27755 20992 27767 20995
rect 28718 20992 28724 21004
rect 27755 20964 28724 20992
rect 27755 20961 27767 20964
rect 27709 20955 27767 20961
rect 23477 20927 23535 20933
rect 23477 20893 23489 20927
rect 23523 20893 23535 20927
rect 23477 20887 23535 20893
rect 24118 20884 24124 20936
rect 24176 20924 24182 20936
rect 24765 20927 24823 20933
rect 24765 20924 24777 20927
rect 24176 20896 24777 20924
rect 24176 20884 24182 20896
rect 24765 20893 24777 20896
rect 24811 20924 24823 20927
rect 25041 20927 25099 20933
rect 25041 20924 25053 20927
rect 24811 20896 25053 20924
rect 24811 20893 24823 20896
rect 24765 20887 24823 20893
rect 25041 20893 25053 20896
rect 25087 20893 25099 20927
rect 25041 20887 25099 20893
rect 25774 20884 25780 20936
rect 25832 20924 25838 20936
rect 26252 20924 26280 20955
rect 28718 20952 28724 20964
rect 28776 20952 28782 21004
rect 28905 20995 28963 21001
rect 28905 20961 28917 20995
rect 28951 20992 28963 20995
rect 29748 20992 29776 21032
rect 30466 21020 30472 21032
rect 30524 21020 30530 21072
rect 30834 21020 30840 21072
rect 30892 21020 30898 21072
rect 31726 21060 31754 21100
rect 34514 21088 34520 21100
rect 34572 21088 34578 21140
rect 39942 21128 39948 21140
rect 34624 21100 39948 21128
rect 31312 21032 31754 21060
rect 30190 20992 30196 21004
rect 28951 20964 29776 20992
rect 29840 20964 30196 20992
rect 28951 20961 28963 20964
rect 28905 20955 28963 20961
rect 25832 20896 26280 20924
rect 25832 20884 25838 20896
rect 27338 20884 27344 20936
rect 27396 20924 27402 20936
rect 28626 20924 28632 20936
rect 27396 20896 28632 20924
rect 27396 20884 27402 20896
rect 28626 20884 28632 20896
rect 28684 20884 28690 20936
rect 28810 20884 28816 20936
rect 28868 20924 28874 20936
rect 29840 20924 29868 20964
rect 30190 20952 30196 20964
rect 30248 20952 30254 21004
rect 31312 21001 31340 21032
rect 34330 21020 34336 21072
rect 34388 21060 34394 21072
rect 34624 21060 34652 21100
rect 39942 21088 39948 21100
rect 40000 21088 40006 21140
rect 40037 21131 40095 21137
rect 40037 21097 40049 21131
rect 40083 21128 40095 21131
rect 40218 21128 40224 21140
rect 40083 21100 40224 21128
rect 40083 21097 40095 21100
rect 40037 21091 40095 21097
rect 40218 21088 40224 21100
rect 40276 21088 40282 21140
rect 40310 21088 40316 21140
rect 40368 21128 40374 21140
rect 41046 21128 41052 21140
rect 40368 21100 41052 21128
rect 40368 21088 40374 21100
rect 41046 21088 41052 21100
rect 41104 21128 41110 21140
rect 49237 21131 49295 21137
rect 49237 21128 49249 21131
rect 41104 21100 49249 21128
rect 41104 21088 41110 21100
rect 49237 21097 49249 21100
rect 49283 21097 49295 21131
rect 49237 21091 49295 21097
rect 34388 21032 34652 21060
rect 34388 21020 34394 21032
rect 39114 21020 39120 21072
rect 39172 21060 39178 21072
rect 39172 21032 39712 21060
rect 39172 21020 39178 21032
rect 31297 20995 31355 21001
rect 31297 20961 31309 20995
rect 31343 20961 31355 20995
rect 31297 20955 31355 20961
rect 31481 20995 31539 21001
rect 31481 20961 31493 20995
rect 31527 20992 31539 20995
rect 32769 20995 32827 21001
rect 32769 20992 32781 20995
rect 31527 20964 32781 20992
rect 31527 20961 31539 20964
rect 31481 20955 31539 20961
rect 32769 20961 32781 20964
rect 32815 20992 32827 20995
rect 34054 20992 34060 21004
rect 32815 20964 34060 20992
rect 32815 20961 32827 20964
rect 32769 20955 32827 20961
rect 34054 20952 34060 20964
rect 34112 20952 34118 21004
rect 34885 20995 34943 21001
rect 34885 20961 34897 20995
rect 34931 20992 34943 20995
rect 35710 20992 35716 21004
rect 34931 20964 35716 20992
rect 34931 20961 34943 20964
rect 34885 20955 34943 20961
rect 35710 20952 35716 20964
rect 35768 20952 35774 21004
rect 35802 20952 35808 21004
rect 35860 20992 35866 21004
rect 36909 20995 36967 21001
rect 36909 20992 36921 20995
rect 35860 20964 36921 20992
rect 35860 20952 35866 20964
rect 36909 20961 36921 20964
rect 36955 20992 36967 20995
rect 36998 20992 37004 21004
rect 36955 20964 37004 20992
rect 36955 20961 36967 20964
rect 36909 20955 36967 20961
rect 36998 20952 37004 20964
rect 37056 20952 37062 21004
rect 37274 20952 37280 21004
rect 37332 20992 37338 21004
rect 37921 20995 37979 21001
rect 37921 20992 37933 20995
rect 37332 20964 37933 20992
rect 37332 20952 37338 20964
rect 37921 20961 37933 20964
rect 37967 20961 37979 20995
rect 37921 20955 37979 20961
rect 38286 20952 38292 21004
rect 38344 20992 38350 21004
rect 39684 20992 39712 21032
rect 39758 21020 39764 21072
rect 39816 21060 39822 21072
rect 39816 21032 40632 21060
rect 39816 21020 39822 21032
rect 40604 21001 40632 21032
rect 42150 21020 42156 21072
rect 42208 21060 42214 21072
rect 42245 21063 42303 21069
rect 42245 21060 42257 21063
rect 42208 21032 42257 21060
rect 42208 21020 42214 21032
rect 42245 21029 42257 21032
rect 42291 21029 42303 21063
rect 42245 21023 42303 21029
rect 40497 20995 40555 21001
rect 40497 20992 40509 20995
rect 38344 20964 39620 20992
rect 39684 20964 40509 20992
rect 38344 20952 38350 20964
rect 28868 20896 29868 20924
rect 29917 20927 29975 20933
rect 28868 20884 28874 20896
rect 29917 20893 29929 20927
rect 29963 20924 29975 20927
rect 30282 20924 30288 20936
rect 29963 20896 30288 20924
rect 29963 20893 29975 20896
rect 29917 20887 29975 20893
rect 30282 20884 30288 20896
rect 30340 20884 30346 20936
rect 30558 20884 30564 20936
rect 30616 20924 30622 20936
rect 30616 20896 31340 20924
rect 30616 20884 30622 20896
rect 14550 20816 14556 20868
rect 14608 20816 14614 20868
rect 16758 20856 16764 20868
rect 15778 20828 16764 20856
rect 16758 20816 16764 20828
rect 16816 20816 16822 20868
rect 19150 20856 19156 20868
rect 18630 20828 19156 20856
rect 19150 20816 19156 20828
rect 19208 20816 19214 20868
rect 21542 20816 21548 20868
rect 21600 20856 21606 20868
rect 21910 20856 21916 20868
rect 21600 20828 21916 20856
rect 21600 20816 21606 20828
rect 21910 20816 21916 20828
rect 21968 20816 21974 20868
rect 25958 20856 25964 20868
rect 23860 20828 25964 20856
rect 13541 20791 13599 20797
rect 13541 20757 13553 20791
rect 13587 20757 13599 20791
rect 13541 20751 13599 20757
rect 14826 20748 14832 20800
rect 14884 20788 14890 20800
rect 16025 20791 16083 20797
rect 16025 20788 16037 20791
rect 14884 20760 16037 20788
rect 14884 20748 14890 20760
rect 16025 20757 16037 20760
rect 16071 20757 16083 20791
rect 16025 20751 16083 20757
rect 16485 20791 16543 20797
rect 16485 20757 16497 20791
rect 16531 20788 16543 20791
rect 17770 20788 17776 20800
rect 16531 20760 17776 20788
rect 16531 20757 16543 20760
rect 16485 20751 16543 20757
rect 17770 20748 17776 20760
rect 17828 20748 17834 20800
rect 18782 20748 18788 20800
rect 18840 20788 18846 20800
rect 18877 20791 18935 20797
rect 18877 20788 18889 20791
rect 18840 20760 18889 20788
rect 18840 20748 18846 20760
rect 18877 20757 18889 20760
rect 18923 20757 18935 20791
rect 18877 20751 18935 20757
rect 20441 20791 20499 20797
rect 20441 20757 20453 20791
rect 20487 20788 20499 20791
rect 23860 20788 23888 20828
rect 25958 20816 25964 20828
rect 26016 20816 26022 20868
rect 26053 20859 26111 20865
rect 26053 20825 26065 20859
rect 26099 20856 26111 20859
rect 26786 20856 26792 20868
rect 26099 20828 26792 20856
rect 26099 20825 26111 20828
rect 26053 20819 26111 20825
rect 26786 20816 26792 20828
rect 26844 20816 26850 20868
rect 27154 20816 27160 20868
rect 27212 20856 27218 20868
rect 29270 20856 29276 20868
rect 27212 20828 29276 20856
rect 27212 20816 27218 20828
rect 29270 20816 29276 20828
rect 29328 20816 29334 20868
rect 30098 20816 30104 20868
rect 30156 20856 30162 20868
rect 31205 20859 31263 20865
rect 31205 20856 31217 20859
rect 30156 20828 31217 20856
rect 30156 20816 30162 20828
rect 31205 20825 31217 20828
rect 31251 20825 31263 20859
rect 31205 20819 31263 20825
rect 20487 20760 23888 20788
rect 20487 20757 20499 20760
rect 20441 20751 20499 20757
rect 24026 20748 24032 20800
rect 24084 20788 24090 20800
rect 24121 20791 24179 20797
rect 24121 20788 24133 20791
rect 24084 20760 24133 20788
rect 24084 20748 24090 20760
rect 24121 20757 24133 20760
rect 24167 20757 24179 20791
rect 24121 20751 24179 20757
rect 24581 20791 24639 20797
rect 24581 20757 24593 20791
rect 24627 20788 24639 20791
rect 28626 20788 28632 20800
rect 24627 20760 28632 20788
rect 24627 20757 24639 20760
rect 24581 20751 24639 20757
rect 28626 20748 28632 20760
rect 28684 20748 28690 20800
rect 28718 20748 28724 20800
rect 28776 20748 28782 20800
rect 28810 20748 28816 20800
rect 28868 20748 28874 20800
rect 29362 20748 29368 20800
rect 29420 20788 29426 20800
rect 29546 20788 29552 20800
rect 29420 20760 29552 20788
rect 29420 20748 29426 20760
rect 29546 20748 29552 20760
rect 29604 20748 29610 20800
rect 29730 20748 29736 20800
rect 29788 20748 29794 20800
rect 31312 20788 31340 20896
rect 32306 20884 32312 20936
rect 32364 20924 32370 20936
rect 32493 20927 32551 20933
rect 32493 20924 32505 20927
rect 32364 20896 32505 20924
rect 32364 20884 32370 20896
rect 32493 20893 32505 20896
rect 32539 20893 32551 20927
rect 32493 20887 32551 20893
rect 37642 20884 37648 20936
rect 37700 20884 37706 20936
rect 39592 20924 39620 20964
rect 40497 20961 40509 20964
rect 40543 20961 40555 20995
rect 40497 20955 40555 20961
rect 40589 20995 40647 21001
rect 40589 20961 40601 20995
rect 40635 20961 40647 20995
rect 41785 20995 41843 21001
rect 41785 20992 41797 20995
rect 40589 20955 40647 20961
rect 41386 20964 41797 20992
rect 41386 20924 41414 20964
rect 41785 20961 41797 20964
rect 41831 20961 41843 20995
rect 41785 20955 41843 20961
rect 39592 20896 41414 20924
rect 41601 20927 41659 20933
rect 41601 20893 41613 20927
rect 41647 20924 41659 20927
rect 48406 20924 48412 20936
rect 41647 20896 48412 20924
rect 41647 20893 41659 20896
rect 41601 20887 41659 20893
rect 48406 20884 48412 20896
rect 48464 20884 48470 20936
rect 48593 20927 48651 20933
rect 48593 20893 48605 20927
rect 48639 20924 48651 20927
rect 49050 20924 49056 20936
rect 48639 20896 49056 20924
rect 48639 20893 48651 20896
rect 48593 20887 48651 20893
rect 49050 20884 49056 20896
rect 49108 20884 49114 20936
rect 31386 20816 31392 20868
rect 31444 20856 31450 20868
rect 32766 20856 32772 20868
rect 31444 20828 32772 20856
rect 31444 20816 31450 20828
rect 32766 20816 32772 20828
rect 32824 20816 32830 20868
rect 32858 20816 32864 20868
rect 32916 20856 32922 20868
rect 33226 20856 33232 20868
rect 32916 20828 33232 20856
rect 32916 20816 32922 20828
rect 33226 20816 33232 20828
rect 33284 20816 33290 20868
rect 35066 20856 35072 20868
rect 34164 20828 35072 20856
rect 34164 20788 34192 20828
rect 35066 20816 35072 20828
rect 35124 20816 35130 20868
rect 35161 20859 35219 20865
rect 35161 20825 35173 20859
rect 35207 20856 35219 20859
rect 35250 20856 35256 20868
rect 35207 20828 35256 20856
rect 35207 20825 35219 20828
rect 35161 20819 35219 20825
rect 35250 20816 35256 20828
rect 35308 20816 35314 20868
rect 35802 20816 35808 20868
rect 35860 20816 35866 20868
rect 38654 20816 38660 20868
rect 38712 20816 38718 20868
rect 40405 20859 40463 20865
rect 40405 20825 40417 20859
rect 40451 20856 40463 20859
rect 40451 20828 41276 20856
rect 40451 20825 40463 20828
rect 40405 20819 40463 20825
rect 31312 20760 34192 20788
rect 34238 20748 34244 20800
rect 34296 20748 34302 20800
rect 34698 20748 34704 20800
rect 34756 20788 34762 20800
rect 36170 20788 36176 20800
rect 34756 20760 36176 20788
rect 34756 20748 34762 20760
rect 36170 20748 36176 20760
rect 36228 20748 36234 20800
rect 36630 20748 36636 20800
rect 36688 20748 36694 20800
rect 38286 20748 38292 20800
rect 38344 20788 38350 20800
rect 41248 20797 41276 20828
rect 41414 20816 41420 20868
rect 41472 20856 41478 20868
rect 41693 20859 41751 20865
rect 41693 20856 41705 20859
rect 41472 20828 41705 20856
rect 41472 20816 41478 20828
rect 41693 20825 41705 20828
rect 41739 20856 41751 20859
rect 42150 20856 42156 20868
rect 41739 20828 42156 20856
rect 41739 20825 41751 20828
rect 41693 20819 41751 20825
rect 42150 20816 42156 20828
rect 42208 20816 42214 20868
rect 39393 20791 39451 20797
rect 39393 20788 39405 20791
rect 38344 20760 39405 20788
rect 38344 20748 38350 20760
rect 39393 20757 39405 20760
rect 39439 20757 39451 20791
rect 39393 20751 39451 20757
rect 41233 20791 41291 20797
rect 41233 20757 41245 20791
rect 41279 20757 41291 20791
rect 41233 20751 41291 20757
rect 48777 20791 48835 20797
rect 48777 20757 48789 20791
rect 48823 20788 48835 20791
rect 48958 20788 48964 20800
rect 48823 20760 48964 20788
rect 48823 20757 48835 20760
rect 48777 20751 48835 20757
rect 48958 20748 48964 20760
rect 49016 20748 49022 20800
rect 1104 20698 49864 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 27950 20698
rect 28002 20646 28014 20698
rect 28066 20646 28078 20698
rect 28130 20646 28142 20698
rect 28194 20646 28206 20698
rect 28258 20646 37950 20698
rect 38002 20646 38014 20698
rect 38066 20646 38078 20698
rect 38130 20646 38142 20698
rect 38194 20646 38206 20698
rect 38258 20646 47950 20698
rect 48002 20646 48014 20698
rect 48066 20646 48078 20698
rect 48130 20646 48142 20698
rect 48194 20646 48206 20698
rect 48258 20646 49864 20698
rect 1104 20624 49864 20646
rect 5258 20544 5264 20596
rect 5316 20544 5322 20596
rect 9674 20544 9680 20596
rect 9732 20544 9738 20596
rect 10318 20544 10324 20596
rect 10376 20544 10382 20596
rect 11882 20584 11888 20596
rect 10428 20556 11888 20584
rect 8386 20516 8392 20528
rect 6472 20488 8392 20516
rect 1765 20451 1823 20457
rect 1765 20417 1777 20451
rect 1811 20448 1823 20451
rect 1946 20448 1952 20460
rect 1811 20420 1952 20448
rect 1811 20417 1823 20420
rect 1765 20411 1823 20417
rect 1946 20408 1952 20420
rect 2004 20408 2010 20460
rect 3605 20451 3663 20457
rect 3605 20417 3617 20451
rect 3651 20448 3663 20451
rect 5445 20451 5503 20457
rect 3651 20420 4108 20448
rect 3651 20417 3663 20420
rect 3605 20411 3663 20417
rect 2777 20383 2835 20389
rect 2777 20349 2789 20383
rect 2823 20380 2835 20383
rect 2866 20380 2872 20392
rect 2823 20352 2872 20380
rect 2823 20349 2835 20352
rect 2777 20343 2835 20349
rect 2866 20340 2872 20352
rect 2924 20340 2930 20392
rect 3878 20340 3884 20392
rect 3936 20340 3942 20392
rect 4080 20312 4108 20420
rect 5445 20417 5457 20451
rect 5491 20448 5503 20451
rect 6472 20448 6500 20488
rect 8386 20476 8392 20488
rect 8444 20476 8450 20528
rect 5491 20420 6500 20448
rect 6549 20451 6607 20457
rect 5491 20417 5503 20420
rect 5445 20411 5503 20417
rect 6549 20417 6561 20451
rect 6595 20417 6607 20451
rect 6549 20411 6607 20417
rect 9217 20451 9275 20457
rect 9217 20417 9229 20451
rect 9263 20417 9275 20451
rect 9217 20411 9275 20417
rect 9861 20451 9919 20457
rect 9861 20417 9873 20451
rect 9907 20448 9919 20451
rect 10428 20448 10456 20556
rect 11882 20544 11888 20556
rect 11940 20544 11946 20596
rect 12989 20587 13047 20593
rect 12989 20584 13001 20587
rect 12544 20556 13001 20584
rect 10594 20476 10600 20528
rect 10652 20516 10658 20528
rect 12544 20525 12572 20556
rect 12989 20553 13001 20556
rect 13035 20584 13047 20587
rect 13354 20584 13360 20596
rect 13035 20556 13360 20584
rect 13035 20553 13047 20556
rect 12989 20547 13047 20553
rect 13354 20544 13360 20556
rect 13412 20544 13418 20596
rect 13630 20544 13636 20596
rect 13688 20584 13694 20596
rect 14093 20587 14151 20593
rect 14093 20584 14105 20587
rect 13688 20556 14105 20584
rect 13688 20544 13694 20556
rect 14093 20553 14105 20556
rect 14139 20553 14151 20587
rect 14093 20547 14151 20553
rect 14918 20544 14924 20596
rect 14976 20544 14982 20596
rect 15102 20544 15108 20596
rect 15160 20544 15166 20596
rect 15378 20544 15384 20596
rect 15436 20584 15442 20596
rect 15565 20587 15623 20593
rect 15565 20584 15577 20587
rect 15436 20556 15577 20584
rect 15436 20544 15442 20556
rect 15565 20553 15577 20556
rect 15611 20553 15623 20587
rect 15565 20547 15623 20553
rect 15838 20544 15844 20596
rect 15896 20584 15902 20596
rect 15933 20587 15991 20593
rect 15933 20584 15945 20587
rect 15896 20556 15945 20584
rect 15896 20544 15902 20556
rect 15933 20553 15945 20556
rect 15979 20553 15991 20587
rect 15933 20547 15991 20553
rect 16022 20544 16028 20596
rect 16080 20544 16086 20596
rect 18785 20587 18843 20593
rect 16132 20556 18644 20584
rect 12529 20519 12587 20525
rect 10652 20488 12480 20516
rect 10652 20476 10658 20488
rect 9907 20420 10456 20448
rect 10505 20451 10563 20457
rect 9907 20417 9919 20420
rect 9861 20411 9919 20417
rect 10505 20417 10517 20451
rect 10551 20448 10563 20451
rect 11422 20448 11428 20460
rect 10551 20420 11428 20448
rect 10551 20417 10563 20420
rect 10505 20411 10563 20417
rect 4154 20340 4160 20392
rect 4212 20380 4218 20392
rect 6564 20380 6592 20411
rect 4212 20352 6592 20380
rect 4212 20340 4218 20352
rect 6638 20340 6644 20392
rect 6696 20380 6702 20392
rect 7009 20383 7067 20389
rect 7009 20380 7021 20383
rect 6696 20352 7021 20380
rect 6696 20340 6702 20352
rect 7009 20349 7021 20352
rect 7055 20349 7067 20383
rect 9232 20380 9260 20411
rect 11422 20408 11428 20420
rect 11480 20408 11486 20460
rect 11793 20451 11851 20457
rect 11793 20417 11805 20451
rect 11839 20417 11851 20451
rect 11793 20411 11851 20417
rect 10410 20380 10416 20392
rect 9232 20352 10416 20380
rect 7009 20343 7067 20349
rect 10410 20340 10416 20352
rect 10468 20340 10474 20392
rect 10962 20340 10968 20392
rect 11020 20340 11026 20392
rect 11808 20380 11836 20411
rect 11882 20408 11888 20460
rect 11940 20448 11946 20460
rect 12452 20448 12480 20488
rect 12529 20485 12541 20519
rect 12575 20485 12587 20519
rect 12529 20479 12587 20485
rect 12710 20476 12716 20528
rect 12768 20476 12774 20528
rect 13262 20476 13268 20528
rect 13320 20516 13326 20528
rect 15120 20516 15148 20544
rect 16132 20516 16160 20556
rect 13320 20488 15056 20516
rect 15120 20488 16160 20516
rect 18616 20516 18644 20556
rect 18785 20553 18797 20587
rect 18831 20584 18843 20587
rect 18874 20584 18880 20596
rect 18831 20556 18880 20584
rect 18831 20553 18843 20556
rect 18785 20547 18843 20553
rect 18874 20544 18880 20556
rect 18932 20544 18938 20596
rect 19150 20544 19156 20596
rect 19208 20544 19214 20596
rect 20254 20584 20260 20596
rect 19720 20556 20260 20584
rect 19334 20516 19340 20528
rect 18616 20488 19340 20516
rect 13320 20476 13326 20488
rect 14918 20448 14924 20460
rect 11940 20420 12204 20448
rect 12452 20420 14924 20448
rect 11940 20408 11946 20420
rect 12176 20380 12204 20420
rect 14918 20408 14924 20420
rect 14976 20408 14982 20460
rect 14185 20383 14243 20389
rect 11808 20352 12020 20380
rect 12176 20352 13768 20380
rect 10870 20312 10876 20324
rect 4080 20284 10876 20312
rect 10870 20272 10876 20284
rect 10928 20272 10934 20324
rect 1762 20204 1768 20256
rect 1820 20244 1826 20256
rect 4798 20244 4804 20256
rect 1820 20216 4804 20244
rect 1820 20204 1826 20216
rect 4798 20204 4804 20216
rect 4856 20204 4862 20256
rect 4982 20204 4988 20256
rect 5040 20244 5046 20256
rect 9033 20247 9091 20253
rect 9033 20244 9045 20247
rect 5040 20216 9045 20244
rect 5040 20204 5046 20216
rect 9033 20213 9045 20216
rect 9079 20213 9091 20247
rect 9033 20207 9091 20213
rect 10042 20204 10048 20256
rect 10100 20244 10106 20256
rect 11885 20247 11943 20253
rect 11885 20244 11897 20247
rect 10100 20216 11897 20244
rect 10100 20204 10106 20216
rect 11885 20213 11897 20216
rect 11931 20213 11943 20247
rect 11992 20244 12020 20352
rect 13740 20321 13768 20352
rect 14185 20349 14197 20383
rect 14231 20349 14243 20383
rect 14185 20343 14243 20349
rect 14369 20383 14427 20389
rect 14369 20349 14381 20383
rect 14415 20380 14427 20383
rect 14826 20380 14832 20392
rect 14415 20352 14832 20380
rect 14415 20349 14427 20352
rect 14369 20343 14427 20349
rect 13725 20315 13783 20321
rect 13725 20281 13737 20315
rect 13771 20281 13783 20315
rect 14200 20312 14228 20343
rect 14826 20340 14832 20352
rect 14884 20340 14890 20392
rect 15028 20380 15056 20488
rect 19334 20476 19340 20488
rect 19392 20476 19398 20528
rect 15105 20451 15163 20457
rect 15105 20417 15117 20451
rect 15151 20448 15163 20451
rect 15930 20448 15936 20460
rect 15151 20420 15936 20448
rect 15151 20417 15163 20420
rect 15105 20411 15163 20417
rect 15930 20408 15936 20420
rect 15988 20408 15994 20460
rect 19150 20448 19156 20460
rect 18446 20420 19156 20448
rect 19150 20408 19156 20420
rect 19208 20408 19214 20460
rect 19720 20457 19748 20556
rect 20254 20544 20260 20556
rect 20312 20584 20318 20596
rect 22462 20584 22468 20596
rect 20312 20556 22468 20584
rect 20312 20544 20318 20556
rect 22462 20544 22468 20556
rect 22520 20584 22526 20596
rect 22738 20584 22744 20596
rect 22520 20556 22744 20584
rect 22520 20544 22526 20556
rect 22738 20544 22744 20556
rect 22796 20544 22802 20596
rect 22830 20544 22836 20596
rect 22888 20584 22894 20596
rect 23201 20587 23259 20593
rect 23201 20584 23213 20587
rect 22888 20556 23213 20584
rect 22888 20544 22894 20556
rect 23201 20553 23213 20556
rect 23247 20553 23259 20587
rect 25682 20584 25688 20596
rect 23201 20547 23259 20553
rect 23860 20556 25688 20584
rect 19978 20476 19984 20528
rect 20036 20476 20042 20528
rect 21266 20476 21272 20528
rect 21324 20516 21330 20528
rect 21324 20488 23520 20516
rect 21324 20476 21330 20488
rect 23492 20460 23520 20488
rect 19705 20451 19763 20457
rect 19705 20417 19717 20451
rect 19751 20417 19763 20451
rect 21542 20448 21548 20460
rect 21114 20420 21548 20448
rect 19705 20411 19763 20417
rect 21542 20408 21548 20420
rect 21600 20408 21606 20460
rect 22373 20451 22431 20457
rect 22373 20417 22385 20451
rect 22419 20448 22431 20451
rect 22419 20420 23336 20448
rect 22419 20417 22431 20420
rect 22373 20411 22431 20417
rect 15470 20380 15476 20392
rect 15028 20352 15476 20380
rect 15470 20340 15476 20352
rect 15528 20340 15534 20392
rect 16206 20340 16212 20392
rect 16264 20340 16270 20392
rect 16758 20340 16764 20392
rect 16816 20340 16822 20392
rect 17034 20340 17040 20392
rect 17092 20340 17098 20392
rect 17313 20383 17371 20389
rect 17313 20349 17325 20383
rect 17359 20380 17371 20383
rect 17678 20380 17684 20392
rect 17359 20352 17684 20380
rect 17359 20349 17371 20352
rect 17313 20343 17371 20349
rect 17678 20340 17684 20352
rect 17736 20340 17742 20392
rect 18046 20340 18052 20392
rect 18104 20380 18110 20392
rect 18782 20380 18788 20392
rect 18104 20352 18788 20380
rect 18104 20340 18110 20352
rect 18782 20340 18788 20352
rect 18840 20340 18846 20392
rect 18966 20340 18972 20392
rect 19024 20380 19030 20392
rect 21450 20380 21456 20392
rect 19024 20352 21456 20380
rect 19024 20340 19030 20352
rect 21450 20340 21456 20352
rect 21508 20340 21514 20392
rect 22462 20340 22468 20392
rect 22520 20340 22526 20392
rect 22557 20383 22615 20389
rect 22557 20349 22569 20383
rect 22603 20349 22615 20383
rect 23308 20380 23336 20420
rect 23382 20408 23388 20460
rect 23440 20408 23446 20460
rect 23474 20408 23480 20460
rect 23532 20448 23538 20460
rect 23860 20457 23888 20556
rect 25682 20544 25688 20556
rect 25740 20544 25746 20596
rect 32306 20584 32312 20596
rect 27264 20556 32312 20584
rect 24670 20476 24676 20528
rect 24728 20476 24734 20528
rect 25498 20476 25504 20528
rect 25556 20516 25562 20528
rect 26878 20516 26884 20528
rect 25556 20488 26884 20516
rect 25556 20476 25562 20488
rect 26878 20476 26884 20488
rect 26936 20476 26942 20528
rect 23845 20451 23903 20457
rect 23845 20448 23857 20451
rect 23532 20420 23857 20448
rect 23532 20408 23538 20420
rect 23845 20417 23857 20420
rect 23891 20417 23903 20451
rect 26237 20451 26295 20457
rect 23845 20411 23903 20417
rect 25516 20420 26188 20448
rect 23750 20380 23756 20392
rect 23308 20352 23756 20380
rect 22557 20343 22615 20349
rect 16850 20312 16856 20324
rect 14200 20284 16856 20312
rect 13725 20275 13783 20281
rect 16850 20272 16856 20284
rect 16908 20272 16914 20324
rect 13262 20244 13268 20256
rect 11992 20216 13268 20244
rect 11885 20207 11943 20213
rect 13262 20204 13268 20216
rect 13320 20204 13326 20256
rect 13449 20247 13507 20253
rect 13449 20213 13461 20247
rect 13495 20244 13507 20247
rect 13538 20244 13544 20256
rect 13495 20216 13544 20244
rect 13495 20213 13507 20216
rect 13449 20207 13507 20213
rect 13538 20204 13544 20216
rect 13596 20204 13602 20256
rect 13814 20204 13820 20256
rect 13872 20244 13878 20256
rect 15746 20244 15752 20256
rect 13872 20216 15752 20244
rect 13872 20204 13878 20216
rect 15746 20204 15752 20216
rect 15804 20204 15810 20256
rect 17052 20244 17080 20340
rect 22186 20272 22192 20324
rect 22244 20312 22250 20324
rect 22572 20312 22600 20343
rect 23750 20340 23756 20352
rect 23808 20340 23814 20392
rect 24121 20383 24179 20389
rect 24121 20349 24133 20383
rect 24167 20380 24179 20383
rect 24486 20380 24492 20392
rect 24167 20352 24492 20380
rect 24167 20349 24179 20352
rect 24121 20343 24179 20349
rect 24486 20340 24492 20352
rect 24544 20380 24550 20392
rect 25516 20380 25544 20420
rect 24544 20352 25544 20380
rect 25593 20383 25651 20389
rect 24544 20340 24550 20352
rect 25593 20349 25605 20383
rect 25639 20380 25651 20383
rect 25774 20380 25780 20392
rect 25639 20352 25780 20380
rect 25639 20349 25651 20352
rect 25593 20343 25651 20349
rect 25774 20340 25780 20352
rect 25832 20340 25838 20392
rect 26160 20380 26188 20420
rect 26237 20417 26249 20451
rect 26283 20448 26295 20451
rect 26694 20448 26700 20460
rect 26283 20420 26700 20448
rect 26283 20417 26295 20420
rect 26237 20411 26295 20417
rect 26694 20408 26700 20420
rect 26752 20408 26758 20460
rect 27264 20457 27292 20556
rect 32306 20544 32312 20556
rect 32364 20544 32370 20596
rect 32600 20556 34008 20584
rect 28258 20476 28264 20528
rect 28316 20476 28322 20528
rect 29822 20476 29828 20528
rect 29880 20476 29886 20528
rect 29917 20519 29975 20525
rect 29917 20485 29929 20519
rect 29963 20516 29975 20519
rect 30006 20516 30012 20528
rect 29963 20488 30012 20516
rect 29963 20485 29975 20488
rect 29917 20479 29975 20485
rect 30006 20476 30012 20488
rect 30064 20476 30070 20528
rect 31110 20476 31116 20528
rect 31168 20476 31174 20528
rect 31662 20516 31668 20528
rect 31312 20488 31668 20516
rect 27249 20451 27307 20457
rect 27249 20417 27261 20451
rect 27295 20417 27307 20451
rect 30834 20448 30840 20460
rect 27249 20411 27307 20417
rect 28736 20420 30840 20448
rect 27154 20380 27160 20392
rect 26160 20352 27160 20380
rect 27154 20340 27160 20352
rect 27212 20340 27218 20392
rect 27522 20340 27528 20392
rect 27580 20340 27586 20392
rect 27614 20340 27620 20392
rect 27672 20380 27678 20392
rect 28736 20380 28764 20420
rect 30834 20408 30840 20420
rect 30892 20408 30898 20460
rect 31021 20451 31079 20457
rect 31021 20417 31033 20451
rect 31067 20448 31079 20451
rect 31312 20448 31340 20488
rect 31662 20476 31668 20488
rect 31720 20476 31726 20528
rect 32600 20525 32628 20556
rect 32585 20519 32643 20525
rect 32585 20516 32597 20519
rect 32324 20488 32597 20516
rect 31067 20420 31340 20448
rect 31067 20417 31079 20420
rect 31021 20411 31079 20417
rect 31386 20408 31392 20460
rect 31444 20448 31450 20460
rect 32324 20448 32352 20488
rect 32585 20485 32597 20488
rect 32631 20485 32643 20519
rect 32585 20479 32643 20485
rect 33226 20476 33232 20528
rect 33284 20476 33290 20528
rect 33980 20516 34008 20556
rect 34054 20544 34060 20596
rect 34112 20544 34118 20596
rect 34517 20587 34575 20593
rect 34517 20553 34529 20587
rect 34563 20584 34575 20587
rect 34698 20584 34704 20596
rect 34563 20556 34704 20584
rect 34563 20553 34575 20556
rect 34517 20547 34575 20553
rect 34698 20544 34704 20556
rect 34756 20544 34762 20596
rect 34885 20587 34943 20593
rect 34885 20584 34897 20587
rect 34808 20556 34897 20584
rect 34422 20516 34428 20528
rect 33980 20488 34428 20516
rect 34422 20476 34428 20488
rect 34480 20476 34486 20528
rect 34606 20476 34612 20528
rect 34664 20516 34670 20528
rect 34808 20516 34836 20556
rect 34885 20553 34897 20556
rect 34931 20553 34943 20587
rect 40313 20587 40371 20593
rect 40313 20584 40325 20587
rect 34885 20547 34943 20553
rect 37246 20556 40325 20584
rect 37246 20516 37274 20556
rect 40313 20553 40325 20556
rect 40359 20553 40371 20587
rect 40313 20547 40371 20553
rect 40405 20587 40463 20593
rect 40405 20553 40417 20587
rect 40451 20584 40463 20587
rect 40586 20584 40592 20596
rect 40451 20556 40592 20584
rect 40451 20553 40463 20556
rect 40405 20547 40463 20553
rect 34664 20488 34836 20516
rect 34900 20488 37274 20516
rect 34664 20476 34670 20488
rect 31444 20420 32352 20448
rect 31444 20408 31450 20420
rect 27672 20352 28764 20380
rect 27672 20340 27678 20352
rect 28994 20340 29000 20392
rect 29052 20340 29058 20392
rect 29270 20380 29276 20392
rect 29104 20352 29276 20380
rect 22244 20284 22600 20312
rect 22244 20272 22250 20284
rect 25406 20272 25412 20324
rect 25464 20312 25470 20324
rect 29104 20312 29132 20352
rect 29270 20340 29276 20352
rect 29328 20380 29334 20392
rect 30009 20383 30067 20389
rect 30009 20380 30021 20383
rect 29328 20352 30021 20380
rect 29328 20340 29334 20352
rect 30009 20349 30021 20352
rect 30055 20349 30067 20383
rect 30009 20343 30067 20349
rect 31202 20340 31208 20392
rect 31260 20340 31266 20392
rect 32306 20340 32312 20392
rect 32364 20340 32370 20392
rect 25464 20284 27384 20312
rect 25464 20272 25470 20284
rect 18782 20244 18788 20256
rect 17052 20216 18788 20244
rect 18782 20204 18788 20216
rect 18840 20204 18846 20256
rect 22002 20204 22008 20256
rect 22060 20204 22066 20256
rect 25498 20204 25504 20256
rect 25556 20244 25562 20256
rect 26053 20247 26111 20253
rect 26053 20244 26065 20247
rect 25556 20216 26065 20244
rect 25556 20204 25562 20216
rect 26053 20213 26065 20216
rect 26099 20213 26111 20247
rect 26053 20207 26111 20213
rect 26602 20204 26608 20256
rect 26660 20204 26666 20256
rect 27356 20244 27384 20284
rect 28552 20284 29132 20312
rect 29196 20284 31156 20312
rect 28552 20244 28580 20284
rect 27356 20216 28580 20244
rect 28994 20204 29000 20256
rect 29052 20244 29058 20256
rect 29196 20244 29224 20284
rect 29052 20216 29224 20244
rect 29457 20247 29515 20253
rect 29052 20204 29058 20216
rect 29457 20213 29469 20247
rect 29503 20244 29515 20247
rect 30558 20244 30564 20256
rect 29503 20216 30564 20244
rect 29503 20213 29515 20216
rect 29457 20207 29515 20213
rect 30558 20204 30564 20216
rect 30616 20204 30622 20256
rect 30653 20247 30711 20253
rect 30653 20213 30665 20247
rect 30699 20244 30711 20247
rect 31018 20244 31024 20256
rect 30699 20216 31024 20244
rect 30699 20213 30711 20216
rect 30653 20207 30711 20213
rect 31018 20204 31024 20216
rect 31076 20204 31082 20256
rect 31128 20244 31156 20284
rect 31846 20272 31852 20324
rect 31904 20272 31910 20324
rect 34900 20244 34928 20488
rect 37366 20476 37372 20528
rect 37424 20516 37430 20528
rect 38013 20519 38071 20525
rect 38013 20516 38025 20519
rect 37424 20488 38025 20516
rect 37424 20476 37430 20488
rect 38013 20485 38025 20488
rect 38059 20516 38071 20519
rect 38286 20516 38292 20528
rect 38059 20488 38292 20516
rect 38059 20485 38071 20488
rect 38013 20479 38071 20485
rect 38286 20476 38292 20488
rect 38344 20476 38350 20528
rect 38654 20476 38660 20528
rect 38712 20476 38718 20528
rect 40328 20516 40356 20547
rect 40586 20544 40592 20556
rect 40644 20544 40650 20596
rect 40328 20488 41736 20516
rect 36449 20451 36507 20457
rect 36449 20417 36461 20451
rect 36495 20448 36507 20451
rect 37182 20448 37188 20460
rect 36495 20420 37188 20448
rect 36495 20417 36507 20420
rect 36449 20411 36507 20417
rect 37182 20408 37188 20420
rect 37240 20408 37246 20460
rect 41141 20451 41199 20457
rect 41141 20448 41153 20451
rect 39224 20420 41153 20448
rect 34977 20383 35035 20389
rect 34977 20349 34989 20383
rect 35023 20349 35035 20383
rect 34977 20343 35035 20349
rect 35161 20383 35219 20389
rect 35161 20349 35173 20383
rect 35207 20380 35219 20383
rect 35250 20380 35256 20392
rect 35207 20352 35256 20380
rect 35207 20349 35219 20352
rect 35161 20343 35219 20349
rect 31128 20216 34928 20244
rect 34992 20244 35020 20343
rect 35250 20340 35256 20352
rect 35308 20340 35314 20392
rect 35526 20340 35532 20392
rect 35584 20380 35590 20392
rect 36541 20383 36599 20389
rect 35584 20352 36492 20380
rect 35584 20340 35590 20352
rect 35066 20272 35072 20324
rect 35124 20312 35130 20324
rect 36081 20315 36139 20321
rect 36081 20312 36093 20315
rect 35124 20284 36093 20312
rect 35124 20272 35130 20284
rect 36081 20281 36093 20284
rect 36127 20281 36139 20315
rect 36081 20275 36139 20281
rect 35250 20244 35256 20256
rect 34992 20216 35256 20244
rect 35250 20204 35256 20216
rect 35308 20244 35314 20256
rect 35529 20247 35587 20253
rect 35529 20244 35541 20247
rect 35308 20216 35541 20244
rect 35308 20204 35314 20216
rect 35529 20213 35541 20216
rect 35575 20213 35587 20247
rect 35529 20207 35587 20213
rect 35802 20204 35808 20256
rect 35860 20204 35866 20256
rect 36464 20244 36492 20352
rect 36541 20349 36553 20383
rect 36587 20380 36599 20383
rect 36630 20380 36636 20392
rect 36587 20352 36636 20380
rect 36587 20349 36599 20352
rect 36541 20343 36599 20349
rect 36630 20340 36636 20352
rect 36688 20340 36694 20392
rect 36725 20383 36783 20389
rect 36725 20349 36737 20383
rect 36771 20380 36783 20383
rect 37550 20380 37556 20392
rect 36771 20352 37556 20380
rect 36771 20349 36783 20352
rect 36725 20343 36783 20349
rect 37550 20340 37556 20352
rect 37608 20340 37614 20392
rect 37734 20340 37740 20392
rect 37792 20340 37798 20392
rect 38562 20340 38568 20392
rect 38620 20380 38626 20392
rect 39224 20380 39252 20420
rect 41141 20417 41153 20420
rect 41187 20417 41199 20451
rect 41141 20411 41199 20417
rect 38620 20352 39252 20380
rect 38620 20340 38626 20352
rect 40494 20340 40500 20392
rect 40552 20340 40558 20392
rect 39022 20272 39028 20324
rect 39080 20312 39086 20324
rect 41322 20312 41328 20324
rect 39080 20284 41328 20312
rect 39080 20272 39086 20284
rect 41322 20272 41328 20284
rect 41380 20272 41386 20324
rect 41708 20321 41736 20488
rect 48593 20451 48651 20457
rect 48593 20417 48605 20451
rect 48639 20448 48651 20451
rect 48774 20448 48780 20460
rect 48639 20420 48780 20448
rect 48639 20417 48651 20420
rect 48593 20411 48651 20417
rect 48774 20408 48780 20420
rect 48832 20408 48838 20460
rect 49050 20408 49056 20460
rect 49108 20408 49114 20460
rect 41693 20315 41751 20321
rect 41693 20281 41705 20315
rect 41739 20312 41751 20315
rect 49237 20315 49295 20321
rect 49237 20312 49249 20315
rect 41739 20284 49249 20312
rect 41739 20281 41751 20284
rect 41693 20275 41751 20281
rect 49237 20281 49249 20284
rect 49283 20281 49295 20315
rect 49237 20275 49295 20281
rect 38654 20244 38660 20256
rect 36464 20216 38660 20244
rect 38654 20204 38660 20216
rect 38712 20204 38718 20256
rect 39206 20204 39212 20256
rect 39264 20244 39270 20256
rect 39485 20247 39543 20253
rect 39485 20244 39497 20247
rect 39264 20216 39497 20244
rect 39264 20204 39270 20216
rect 39485 20213 39497 20216
rect 39531 20213 39543 20247
rect 39485 20207 39543 20213
rect 39942 20204 39948 20256
rect 40000 20204 40006 20256
rect 48406 20204 48412 20256
rect 48464 20204 48470 20256
rect 1104 20154 49864 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 32950 20154
rect 33002 20102 33014 20154
rect 33066 20102 33078 20154
rect 33130 20102 33142 20154
rect 33194 20102 33206 20154
rect 33258 20102 42950 20154
rect 43002 20102 43014 20154
rect 43066 20102 43078 20154
rect 43130 20102 43142 20154
rect 43194 20102 43206 20154
rect 43258 20102 49864 20154
rect 1104 20080 49864 20102
rect 7006 20040 7012 20052
rect 4080 20012 7012 20040
rect 1762 19796 1768 19848
rect 1820 19796 1826 19848
rect 4080 19845 4108 20012
rect 7006 20000 7012 20012
rect 7064 20000 7070 20052
rect 9950 20000 9956 20052
rect 10008 20000 10014 20052
rect 14277 20043 14335 20049
rect 10796 20012 14044 20040
rect 4798 19932 4804 19984
rect 4856 19972 4862 19984
rect 4856 19944 10732 19972
rect 4856 19932 4862 19944
rect 4890 19864 4896 19916
rect 4948 19864 4954 19916
rect 6178 19864 6184 19916
rect 6236 19904 6242 19916
rect 6273 19907 6331 19913
rect 6273 19904 6285 19907
rect 6236 19876 6285 19904
rect 6236 19864 6242 19876
rect 6273 19873 6285 19876
rect 6319 19873 6331 19907
rect 6273 19867 6331 19873
rect 4065 19839 4123 19845
rect 4065 19805 4077 19839
rect 4111 19805 4123 19839
rect 4065 19799 4123 19805
rect 5997 19839 6055 19845
rect 5997 19805 6009 19839
rect 6043 19805 6055 19839
rect 5997 19799 6055 19805
rect 7929 19839 7987 19845
rect 7929 19805 7941 19839
rect 7975 19836 7987 19839
rect 9766 19836 9772 19848
rect 7975 19808 9772 19836
rect 7975 19805 7987 19808
rect 7929 19799 7987 19805
rect 2774 19728 2780 19780
rect 2832 19728 2838 19780
rect 6012 19700 6040 19799
rect 9766 19796 9772 19808
rect 9824 19796 9830 19848
rect 10137 19839 10195 19845
rect 10137 19805 10149 19839
rect 10183 19836 10195 19839
rect 10594 19836 10600 19848
rect 10183 19808 10600 19836
rect 10183 19805 10195 19808
rect 10137 19799 10195 19805
rect 10594 19796 10600 19808
rect 10652 19796 10658 19848
rect 7098 19728 7104 19780
rect 7156 19768 7162 19780
rect 7834 19768 7840 19780
rect 7156 19740 7840 19768
rect 7156 19728 7162 19740
rect 7834 19728 7840 19740
rect 7892 19768 7898 19780
rect 10042 19768 10048 19780
rect 7892 19740 10048 19768
rect 7892 19728 7898 19740
rect 10042 19728 10048 19740
rect 10100 19728 10106 19780
rect 7745 19703 7803 19709
rect 7745 19700 7757 19703
rect 6012 19672 7757 19700
rect 7745 19669 7757 19672
rect 7791 19669 7803 19703
rect 7745 19663 7803 19669
rect 10502 19660 10508 19712
rect 10560 19700 10566 19712
rect 10597 19703 10655 19709
rect 10597 19700 10609 19703
rect 10560 19672 10609 19700
rect 10560 19660 10566 19672
rect 10597 19669 10609 19672
rect 10643 19669 10655 19703
rect 10704 19700 10732 19944
rect 10796 19845 10824 20012
rect 10870 19932 10876 19984
rect 10928 19972 10934 19984
rect 11517 19975 11575 19981
rect 11517 19972 11529 19975
rect 10928 19944 11529 19972
rect 10928 19932 10934 19944
rect 11517 19941 11529 19944
rect 11563 19941 11575 19975
rect 11517 19935 11575 19941
rect 13725 19975 13783 19981
rect 13725 19941 13737 19975
rect 13771 19972 13783 19975
rect 13906 19972 13912 19984
rect 13771 19944 13912 19972
rect 13771 19941 13783 19944
rect 13725 19935 13783 19941
rect 13906 19932 13912 19944
rect 13964 19932 13970 19984
rect 14016 19972 14044 20012
rect 14277 20009 14289 20043
rect 14323 20040 14335 20043
rect 14366 20040 14372 20052
rect 14323 20012 14372 20040
rect 14323 20009 14335 20012
rect 14277 20003 14335 20009
rect 14366 20000 14372 20012
rect 14424 20000 14430 20052
rect 14918 20000 14924 20052
rect 14976 20040 14982 20052
rect 16853 20043 16911 20049
rect 16853 20040 16865 20043
rect 14976 20012 16865 20040
rect 14976 20000 14982 20012
rect 16853 20009 16865 20012
rect 16899 20009 16911 20043
rect 18046 20040 18052 20052
rect 16853 20003 16911 20009
rect 17420 20012 18052 20040
rect 15657 19975 15715 19981
rect 15657 19972 15669 19975
rect 14016 19944 15669 19972
rect 15657 19941 15669 19944
rect 15703 19941 15715 19975
rect 17420 19972 17448 20012
rect 18046 20000 18052 20012
rect 18104 20000 18110 20052
rect 18141 20043 18199 20049
rect 18141 20009 18153 20043
rect 18187 20040 18199 20043
rect 18322 20040 18328 20052
rect 18187 20012 18328 20040
rect 18187 20009 18199 20012
rect 18141 20003 18199 20009
rect 18322 20000 18328 20012
rect 18380 20000 18386 20052
rect 20257 20043 20315 20049
rect 20257 20009 20269 20043
rect 20303 20040 20315 20043
rect 20530 20040 20536 20052
rect 20303 20012 20536 20040
rect 20303 20009 20315 20012
rect 20257 20003 20315 20009
rect 20530 20000 20536 20012
rect 20588 20000 20594 20052
rect 20796 20043 20854 20049
rect 20796 20009 20808 20043
rect 20842 20040 20854 20043
rect 20842 20012 22416 20040
rect 20842 20009 20854 20012
rect 20796 20003 20854 20009
rect 18874 19972 18880 19984
rect 15657 19935 15715 19941
rect 16316 19944 17448 19972
rect 17512 19944 18880 19972
rect 11977 19907 12035 19913
rect 11977 19873 11989 19907
rect 12023 19904 12035 19907
rect 14274 19904 14280 19916
rect 12023 19876 14280 19904
rect 12023 19873 12035 19876
rect 11977 19867 12035 19873
rect 14274 19864 14280 19876
rect 14332 19864 14338 19916
rect 15562 19904 15568 19916
rect 14476 19876 15568 19904
rect 10781 19839 10839 19845
rect 10781 19805 10793 19839
rect 10827 19805 10839 19839
rect 14090 19836 14096 19848
rect 10781 19799 10839 19805
rect 13556 19808 14096 19836
rect 13556 19780 13584 19808
rect 14090 19796 14096 19808
rect 14148 19796 14154 19848
rect 14476 19845 14504 19876
rect 15562 19864 15568 19876
rect 15620 19864 15626 19916
rect 16316 19913 16344 19944
rect 17512 19913 17540 19944
rect 18874 19932 18880 19944
rect 18932 19932 18938 19984
rect 16301 19907 16359 19913
rect 16301 19873 16313 19907
rect 16347 19873 16359 19907
rect 16301 19867 16359 19873
rect 17497 19907 17555 19913
rect 17497 19873 17509 19907
rect 17543 19873 17555 19907
rect 17497 19867 17555 19873
rect 18785 19907 18843 19913
rect 18785 19873 18797 19907
rect 18831 19904 18843 19907
rect 19058 19904 19064 19916
rect 18831 19876 19064 19904
rect 18831 19873 18843 19876
rect 18785 19867 18843 19873
rect 19058 19864 19064 19876
rect 19116 19864 19122 19916
rect 19334 19864 19340 19916
rect 19392 19864 19398 19916
rect 20533 19907 20591 19913
rect 20533 19873 20545 19907
rect 20579 19904 20591 19907
rect 21174 19904 21180 19916
rect 20579 19876 21180 19904
rect 20579 19873 20591 19876
rect 20533 19867 20591 19873
rect 21174 19864 21180 19876
rect 21232 19864 21238 19916
rect 21358 19864 21364 19916
rect 21416 19904 21422 19916
rect 22281 19907 22339 19913
rect 22281 19904 22293 19907
rect 21416 19876 22293 19904
rect 21416 19864 21422 19876
rect 22281 19873 22293 19876
rect 22327 19873 22339 19907
rect 22388 19904 22416 20012
rect 22462 20000 22468 20052
rect 22520 20040 22526 20052
rect 25593 20043 25651 20049
rect 25593 20040 25605 20043
rect 22520 20012 25605 20040
rect 22520 20000 22526 20012
rect 25593 20009 25605 20012
rect 25639 20009 25651 20043
rect 25593 20003 25651 20009
rect 26786 20000 26792 20052
rect 26844 20000 26850 20052
rect 28350 20000 28356 20052
rect 28408 20040 28414 20052
rect 29181 20043 29239 20049
rect 29181 20040 29193 20043
rect 28408 20012 29193 20040
rect 28408 20000 28414 20012
rect 29181 20009 29193 20012
rect 29227 20040 29239 20043
rect 29454 20040 29460 20052
rect 29227 20012 29460 20040
rect 29227 20009 29239 20012
rect 29181 20003 29239 20009
rect 29454 20000 29460 20012
rect 29512 20000 29518 20052
rect 30374 20040 30380 20052
rect 29564 20012 30380 20040
rect 23293 19975 23351 19981
rect 23293 19941 23305 19975
rect 23339 19972 23351 19975
rect 23382 19972 23388 19984
rect 23339 19944 23388 19972
rect 23339 19941 23351 19944
rect 23293 19935 23351 19941
rect 23382 19932 23388 19944
rect 23440 19932 23446 19984
rect 24118 19972 24124 19984
rect 23860 19944 24124 19972
rect 23658 19904 23664 19916
rect 22388 19876 23664 19904
rect 22281 19867 22339 19873
rect 23658 19864 23664 19876
rect 23716 19864 23722 19916
rect 23860 19913 23888 19944
rect 24118 19932 24124 19944
rect 24176 19932 24182 19984
rect 24670 19932 24676 19984
rect 24728 19972 24734 19984
rect 25041 19975 25099 19981
rect 25041 19972 25053 19975
rect 24728 19944 25053 19972
rect 24728 19932 24734 19944
rect 25041 19941 25053 19944
rect 25087 19972 25099 19975
rect 25225 19975 25283 19981
rect 25225 19972 25237 19975
rect 25087 19944 25237 19972
rect 25087 19941 25099 19944
rect 25041 19935 25099 19941
rect 25225 19941 25237 19944
rect 25271 19941 25283 19975
rect 25225 19935 25283 19941
rect 26418 19932 26424 19984
rect 26476 19972 26482 19984
rect 29564 19972 29592 20012
rect 30374 20000 30380 20012
rect 30432 20000 30438 20052
rect 30929 20043 30987 20049
rect 30929 20009 30941 20043
rect 30975 20040 30987 20043
rect 33502 20040 33508 20052
rect 30975 20012 33508 20040
rect 30975 20009 30987 20012
rect 30929 20003 30987 20009
rect 33502 20000 33508 20012
rect 33560 20000 33566 20052
rect 34606 20000 34612 20052
rect 34664 20040 34670 20052
rect 35802 20040 35808 20052
rect 34664 20012 35808 20040
rect 34664 20000 34670 20012
rect 35802 20000 35808 20012
rect 35860 20040 35866 20052
rect 35860 20012 36768 20040
rect 35860 20000 35866 20012
rect 26476 19944 27614 19972
rect 26476 19932 26482 19944
rect 23845 19907 23903 19913
rect 23845 19873 23857 19907
rect 23891 19873 23903 19907
rect 23845 19867 23903 19873
rect 23934 19864 23940 19916
rect 23992 19904 23998 19916
rect 24581 19907 24639 19913
rect 24581 19904 24593 19907
rect 23992 19876 24593 19904
rect 23992 19864 23998 19876
rect 24581 19873 24593 19876
rect 24627 19873 24639 19907
rect 24581 19867 24639 19873
rect 25406 19864 25412 19916
rect 25464 19904 25470 19916
rect 26050 19904 26056 19916
rect 25464 19876 26056 19904
rect 25464 19864 25470 19876
rect 26050 19864 26056 19876
rect 26108 19864 26114 19916
rect 26142 19864 26148 19916
rect 26200 19864 26206 19916
rect 27154 19864 27160 19916
rect 27212 19904 27218 19916
rect 27341 19907 27399 19913
rect 27341 19904 27353 19907
rect 27212 19876 27353 19904
rect 27212 19864 27218 19876
rect 27341 19873 27353 19876
rect 27387 19873 27399 19907
rect 27341 19867 27399 19873
rect 14461 19839 14519 19845
rect 14461 19805 14473 19839
rect 14507 19805 14519 19839
rect 17402 19836 17408 19848
rect 14461 19799 14519 19805
rect 14936 19808 17408 19836
rect 11333 19771 11391 19777
rect 11333 19737 11345 19771
rect 11379 19768 11391 19771
rect 12158 19768 12164 19780
rect 11379 19740 12164 19768
rect 11379 19737 11391 19740
rect 11333 19731 11391 19737
rect 12158 19728 12164 19740
rect 12216 19728 12222 19780
rect 12250 19728 12256 19780
rect 12308 19728 12314 19780
rect 13538 19768 13544 19780
rect 13478 19740 13544 19768
rect 13538 19728 13544 19740
rect 13596 19728 13602 19780
rect 13648 19740 13860 19768
rect 13648 19700 13676 19740
rect 10704 19672 13676 19700
rect 13832 19700 13860 19740
rect 13906 19728 13912 19780
rect 13964 19768 13970 19780
rect 14550 19768 14556 19780
rect 13964 19740 14556 19768
rect 13964 19728 13970 19740
rect 14550 19728 14556 19740
rect 14608 19768 14614 19780
rect 14936 19768 14964 19808
rect 17402 19796 17408 19808
rect 17460 19796 17466 19848
rect 18506 19796 18512 19848
rect 18564 19796 18570 19848
rect 18601 19839 18659 19845
rect 18601 19805 18613 19839
rect 18647 19836 18659 19839
rect 18647 19808 20392 19836
rect 18647 19805 18659 19808
rect 18601 19799 18659 19805
rect 14608 19740 14964 19768
rect 14608 19728 14614 19740
rect 15010 19728 15016 19780
rect 15068 19728 15074 19780
rect 16025 19771 16083 19777
rect 16025 19737 16037 19771
rect 16071 19768 16083 19771
rect 17034 19768 17040 19780
rect 16071 19740 17040 19768
rect 16071 19737 16083 19740
rect 16025 19731 16083 19737
rect 17034 19728 17040 19740
rect 17092 19728 17098 19780
rect 17313 19771 17371 19777
rect 17313 19737 17325 19771
rect 17359 19768 17371 19771
rect 19610 19768 19616 19780
rect 17359 19740 19616 19768
rect 17359 19737 17371 19740
rect 17313 19731 17371 19737
rect 19610 19728 19616 19740
rect 19668 19728 19674 19780
rect 19705 19771 19763 19777
rect 19705 19737 19717 19771
rect 19751 19768 19763 19771
rect 20162 19768 20168 19780
rect 19751 19740 20168 19768
rect 19751 19737 19763 19740
rect 19705 19731 19763 19737
rect 20162 19728 20168 19740
rect 20220 19728 20226 19780
rect 15105 19703 15163 19709
rect 15105 19700 15117 19703
rect 13832 19672 15117 19700
rect 10597 19663 10655 19669
rect 15105 19669 15117 19672
rect 15151 19669 15163 19703
rect 15105 19663 15163 19669
rect 16117 19703 16175 19709
rect 16117 19669 16129 19703
rect 16163 19700 16175 19703
rect 16390 19700 16396 19712
rect 16163 19672 16396 19700
rect 16163 19669 16175 19672
rect 16117 19663 16175 19669
rect 16390 19660 16396 19672
rect 16448 19660 16454 19712
rect 17218 19660 17224 19712
rect 17276 19660 17282 19712
rect 17494 19660 17500 19712
rect 17552 19700 17558 19712
rect 19797 19703 19855 19709
rect 19797 19700 19809 19703
rect 17552 19672 19809 19700
rect 17552 19660 17558 19672
rect 19797 19669 19809 19672
rect 19843 19669 19855 19703
rect 20364 19700 20392 19808
rect 22370 19796 22376 19848
rect 22428 19836 22434 19848
rect 22557 19839 22615 19845
rect 22557 19836 22569 19839
rect 22428 19808 22569 19836
rect 22428 19796 22434 19808
rect 22557 19805 22569 19808
rect 22603 19805 22615 19839
rect 27586 19836 27614 19944
rect 28460 19944 29592 19972
rect 30300 19944 31754 19972
rect 28460 19913 28488 19944
rect 28445 19907 28503 19913
rect 28445 19873 28457 19907
rect 28491 19873 28503 19907
rect 28445 19867 28503 19873
rect 28629 19907 28687 19913
rect 28629 19873 28641 19907
rect 28675 19873 28687 19907
rect 28994 19904 29000 19916
rect 28629 19867 28687 19873
rect 28828 19876 29000 19904
rect 28644 19836 28672 19867
rect 27586 19808 28672 19836
rect 22557 19799 22615 19805
rect 21542 19728 21548 19780
rect 21600 19728 21606 19780
rect 22833 19771 22891 19777
rect 22833 19768 22845 19771
rect 22480 19740 22845 19768
rect 21082 19700 21088 19712
rect 20364 19672 21088 19700
rect 19797 19663 19855 19669
rect 21082 19660 21088 19672
rect 21140 19660 21146 19712
rect 21174 19660 21180 19712
rect 21232 19700 21238 19712
rect 22480 19700 22508 19740
rect 22833 19737 22845 19740
rect 22879 19768 22891 19771
rect 23661 19771 23719 19777
rect 23661 19768 23673 19771
rect 22879 19740 23673 19768
rect 22879 19737 22891 19740
rect 22833 19731 22891 19737
rect 23661 19737 23673 19740
rect 23707 19737 23719 19771
rect 23661 19731 23719 19737
rect 23753 19771 23811 19777
rect 23753 19737 23765 19771
rect 23799 19768 23811 19771
rect 24026 19768 24032 19780
rect 23799 19740 24032 19768
rect 23799 19737 23811 19740
rect 23753 19731 23811 19737
rect 24026 19728 24032 19740
rect 24084 19768 24090 19780
rect 25222 19768 25228 19780
rect 24084 19740 25228 19768
rect 24084 19728 24090 19740
rect 25222 19728 25228 19740
rect 25280 19728 25286 19780
rect 25866 19728 25872 19780
rect 25924 19768 25930 19780
rect 27157 19771 27215 19777
rect 27157 19768 27169 19771
rect 25924 19740 27169 19768
rect 25924 19728 25930 19740
rect 27157 19737 27169 19740
rect 27203 19768 27215 19771
rect 28828 19768 28856 19876
rect 28994 19864 29000 19876
rect 29052 19864 29058 19916
rect 29454 19864 29460 19916
rect 29512 19904 29518 19916
rect 30300 19913 30328 19944
rect 30285 19907 30343 19913
rect 30285 19904 30297 19907
rect 29512 19876 30297 19904
rect 29512 19864 29518 19876
rect 30285 19873 30297 19876
rect 30331 19873 30343 19907
rect 30285 19867 30343 19873
rect 30374 19864 30380 19916
rect 30432 19904 30438 19916
rect 31294 19904 31300 19916
rect 30432 19876 31300 19904
rect 30432 19864 30438 19876
rect 31294 19864 31300 19876
rect 31352 19864 31358 19916
rect 31478 19864 31484 19916
rect 31536 19864 31542 19916
rect 31726 19904 31754 19944
rect 31938 19932 31944 19984
rect 31996 19972 32002 19984
rect 36081 19975 36139 19981
rect 36081 19972 36093 19975
rect 31996 19944 36093 19972
rect 31996 19932 32002 19944
rect 36081 19941 36093 19944
rect 36127 19941 36139 19975
rect 36081 19935 36139 19941
rect 32677 19907 32735 19913
rect 32677 19904 32689 19907
rect 31726 19876 32689 19904
rect 32677 19873 32689 19876
rect 32723 19873 32735 19907
rect 32677 19867 32735 19873
rect 33502 19864 33508 19916
rect 33560 19904 33566 19916
rect 33965 19907 34023 19913
rect 33965 19904 33977 19907
rect 33560 19876 33977 19904
rect 33560 19864 33566 19876
rect 33965 19873 33977 19876
rect 34011 19873 34023 19907
rect 33965 19867 34023 19873
rect 34900 19876 35388 19904
rect 28902 19796 28908 19848
rect 28960 19836 28966 19848
rect 30193 19839 30251 19845
rect 30193 19836 30205 19839
rect 28960 19808 30205 19836
rect 28960 19796 28966 19808
rect 30193 19805 30205 19808
rect 30239 19805 30251 19839
rect 30193 19799 30251 19805
rect 27203 19740 28856 19768
rect 29656 19740 29960 19768
rect 27203 19737 27215 19740
rect 27157 19731 27215 19737
rect 21232 19672 22508 19700
rect 21232 19660 21238 19672
rect 22922 19660 22928 19712
rect 22980 19660 22986 19712
rect 25958 19660 25964 19712
rect 26016 19660 26022 19712
rect 26050 19660 26056 19712
rect 26108 19660 26114 19712
rect 26878 19660 26884 19712
rect 26936 19700 26942 19712
rect 27249 19703 27307 19709
rect 27249 19700 27261 19703
rect 26936 19672 27261 19700
rect 26936 19660 26942 19672
rect 27249 19669 27261 19672
rect 27295 19669 27307 19703
rect 27249 19663 27307 19669
rect 27614 19660 27620 19712
rect 27672 19700 27678 19712
rect 27985 19703 28043 19709
rect 27985 19700 27997 19703
rect 27672 19672 27997 19700
rect 27672 19660 27678 19672
rect 27985 19669 27997 19672
rect 28031 19669 28043 19703
rect 27985 19663 28043 19669
rect 28353 19703 28411 19709
rect 28353 19669 28365 19703
rect 28399 19700 28411 19703
rect 28718 19700 28724 19712
rect 28399 19672 28724 19700
rect 28399 19669 28411 19672
rect 28353 19663 28411 19669
rect 28718 19660 28724 19672
rect 28776 19660 28782 19712
rect 28902 19660 28908 19712
rect 28960 19700 28966 19712
rect 29656 19700 29684 19740
rect 28960 19672 29684 19700
rect 28960 19660 28966 19672
rect 29730 19660 29736 19712
rect 29788 19660 29794 19712
rect 29932 19700 29960 19740
rect 30006 19728 30012 19780
rect 30064 19768 30070 19780
rect 30101 19771 30159 19777
rect 30101 19768 30113 19771
rect 30064 19740 30113 19768
rect 30064 19728 30070 19740
rect 30101 19737 30113 19740
rect 30147 19737 30159 19771
rect 30208 19768 30236 19799
rect 31110 19796 31116 19848
rect 31168 19836 31174 19848
rect 31389 19839 31447 19845
rect 31389 19836 31401 19839
rect 31168 19808 31401 19836
rect 31168 19796 31174 19808
rect 31389 19805 31401 19808
rect 31435 19836 31447 19839
rect 31846 19836 31852 19848
rect 31435 19808 31852 19836
rect 31435 19805 31447 19808
rect 31389 19799 31447 19805
rect 31846 19796 31852 19808
rect 31904 19796 31910 19848
rect 32585 19839 32643 19845
rect 32585 19805 32597 19839
rect 32631 19836 32643 19839
rect 33873 19839 33931 19845
rect 33873 19836 33885 19839
rect 32631 19808 33885 19836
rect 32631 19805 32643 19808
rect 32585 19799 32643 19805
rect 33873 19805 33885 19808
rect 33919 19836 33931 19839
rect 34900 19836 34928 19876
rect 33919 19808 34928 19836
rect 33919 19805 33931 19808
rect 33873 19799 33931 19805
rect 34974 19796 34980 19848
rect 35032 19836 35038 19848
rect 35253 19839 35311 19845
rect 35253 19836 35265 19839
rect 35032 19808 35265 19836
rect 35032 19796 35038 19808
rect 35253 19805 35265 19808
rect 35299 19805 35311 19839
rect 35360 19836 35388 19876
rect 35526 19864 35532 19916
rect 35584 19864 35590 19916
rect 36170 19864 36176 19916
rect 36228 19904 36234 19916
rect 36633 19907 36691 19913
rect 36633 19904 36645 19907
rect 36228 19876 36645 19904
rect 36228 19864 36234 19876
rect 36633 19873 36645 19876
rect 36679 19873 36691 19907
rect 36740 19904 36768 20012
rect 37274 20000 37280 20052
rect 37332 20040 37338 20052
rect 48590 20040 48596 20052
rect 37332 20012 48596 20040
rect 37332 20000 37338 20012
rect 48590 20000 48596 20012
rect 48648 20000 48654 20052
rect 48774 20000 48780 20052
rect 48832 20000 48838 20052
rect 37090 19932 37096 19984
rect 37148 19972 37154 19984
rect 38194 19972 38200 19984
rect 37148 19944 38200 19972
rect 37148 19932 37154 19944
rect 38194 19932 38200 19944
rect 38252 19972 38258 19984
rect 38841 19975 38899 19981
rect 38841 19972 38853 19975
rect 38252 19944 38853 19972
rect 38252 19932 38258 19944
rect 38841 19941 38853 19944
rect 38887 19972 38899 19975
rect 39758 19972 39764 19984
rect 38887 19944 39764 19972
rect 38887 19941 38899 19944
rect 38841 19935 38899 19941
rect 39758 19932 39764 19944
rect 39816 19932 39822 19984
rect 41230 19972 41236 19984
rect 40512 19944 41236 19972
rect 37366 19904 37372 19916
rect 36740 19876 37372 19904
rect 36633 19867 36691 19873
rect 37366 19864 37372 19876
rect 37424 19864 37430 19916
rect 37642 19864 37648 19916
rect 37700 19904 37706 19916
rect 38381 19907 38439 19913
rect 38381 19904 38393 19907
rect 37700 19876 38393 19904
rect 37700 19864 37706 19876
rect 38381 19873 38393 19876
rect 38427 19873 38439 19907
rect 38381 19867 38439 19873
rect 38746 19864 38752 19916
rect 38804 19904 38810 19916
rect 39482 19904 39488 19916
rect 38804 19876 39488 19904
rect 38804 19864 38810 19876
rect 39482 19864 39488 19876
rect 39540 19904 39546 19916
rect 40512 19913 40540 19944
rect 41230 19932 41236 19944
rect 41288 19932 41294 19984
rect 39577 19907 39635 19913
rect 39577 19904 39589 19907
rect 39540 19876 39589 19904
rect 39540 19864 39546 19876
rect 39577 19873 39589 19876
rect 39623 19873 39635 19907
rect 39577 19867 39635 19873
rect 40497 19907 40555 19913
rect 40497 19873 40509 19907
rect 40543 19873 40555 19907
rect 40497 19867 40555 19873
rect 40586 19864 40592 19916
rect 40644 19864 40650 19916
rect 41046 19864 41052 19916
rect 41104 19864 41110 19916
rect 43898 19836 43904 19848
rect 35360 19808 43904 19836
rect 35253 19799 35311 19805
rect 43898 19796 43904 19808
rect 43956 19796 43962 19848
rect 32214 19768 32220 19780
rect 30208 19740 32220 19768
rect 30101 19731 30159 19737
rect 32214 19728 32220 19740
rect 32272 19728 32278 19780
rect 32493 19771 32551 19777
rect 32493 19737 32505 19771
rect 32539 19768 32551 19771
rect 33778 19768 33784 19780
rect 32539 19740 33784 19768
rect 32539 19737 32551 19740
rect 32493 19731 32551 19737
rect 33778 19728 33784 19740
rect 33836 19728 33842 19780
rect 35066 19768 35072 19780
rect 34256 19740 35072 19768
rect 30834 19700 30840 19712
rect 29932 19672 30840 19700
rect 30834 19660 30840 19672
rect 30892 19660 30898 19712
rect 31297 19703 31355 19709
rect 31297 19669 31309 19703
rect 31343 19700 31355 19703
rect 31662 19700 31668 19712
rect 31343 19672 31668 19700
rect 31343 19669 31355 19672
rect 31297 19663 31355 19669
rect 31662 19660 31668 19672
rect 31720 19660 31726 19712
rect 32122 19660 32128 19712
rect 32180 19660 32186 19712
rect 32398 19660 32404 19712
rect 32456 19700 32462 19712
rect 32766 19700 32772 19712
rect 32456 19672 32772 19700
rect 32456 19660 32462 19672
rect 32766 19660 32772 19672
rect 32824 19660 32830 19712
rect 33413 19703 33471 19709
rect 33413 19669 33425 19703
rect 33459 19700 33471 19703
rect 34256 19700 34284 19740
rect 35066 19728 35072 19740
rect 35124 19728 35130 19780
rect 35345 19771 35403 19777
rect 35345 19737 35357 19771
rect 35391 19768 35403 19771
rect 35434 19768 35440 19780
rect 35391 19740 35440 19768
rect 35391 19737 35403 19740
rect 35345 19731 35403 19737
rect 35434 19728 35440 19740
rect 35492 19728 35498 19780
rect 35618 19728 35624 19780
rect 35676 19768 35682 19780
rect 36449 19771 36507 19777
rect 35676 19740 35940 19768
rect 35676 19728 35682 19740
rect 33459 19672 34284 19700
rect 33459 19669 33471 19672
rect 33413 19663 33471 19669
rect 34330 19660 34336 19712
rect 34388 19700 34394 19712
rect 34425 19703 34483 19709
rect 34425 19700 34437 19703
rect 34388 19672 34437 19700
rect 34388 19660 34394 19672
rect 34425 19669 34437 19672
rect 34471 19669 34483 19703
rect 34425 19663 34483 19669
rect 34885 19703 34943 19709
rect 34885 19669 34897 19703
rect 34931 19700 34943 19703
rect 35802 19700 35808 19712
rect 34931 19672 35808 19700
rect 34931 19669 34943 19672
rect 34885 19663 34943 19669
rect 35802 19660 35808 19672
rect 35860 19660 35866 19712
rect 35912 19700 35940 19740
rect 36449 19737 36461 19771
rect 36495 19768 36507 19771
rect 40126 19768 40132 19780
rect 36495 19740 40132 19768
rect 36495 19737 36507 19740
rect 36449 19731 36507 19737
rect 40126 19728 40132 19740
rect 40184 19728 40190 19780
rect 40405 19771 40463 19777
rect 40405 19737 40417 19771
rect 40451 19768 40463 19771
rect 41046 19768 41052 19780
rect 40451 19740 41052 19768
rect 40451 19737 40463 19740
rect 40405 19731 40463 19737
rect 41046 19728 41052 19740
rect 41104 19728 41110 19780
rect 48593 19771 48651 19777
rect 48593 19737 48605 19771
rect 48639 19768 48651 19771
rect 49145 19771 49203 19777
rect 49145 19768 49157 19771
rect 48639 19740 49157 19768
rect 48639 19737 48651 19740
rect 48593 19731 48651 19737
rect 49145 19737 49157 19740
rect 49191 19768 49203 19771
rect 49326 19768 49332 19780
rect 49191 19740 49332 19768
rect 49191 19737 49203 19740
rect 49145 19731 49203 19737
rect 49326 19728 49332 19740
rect 49384 19728 49390 19780
rect 36541 19703 36599 19709
rect 36541 19700 36553 19703
rect 35912 19672 36553 19700
rect 36541 19669 36553 19672
rect 36587 19669 36599 19703
rect 36541 19663 36599 19669
rect 37826 19660 37832 19712
rect 37884 19660 37890 19712
rect 38194 19660 38200 19712
rect 38252 19660 38258 19712
rect 38289 19703 38347 19709
rect 38289 19669 38301 19703
rect 38335 19700 38347 19703
rect 38654 19700 38660 19712
rect 38335 19672 38660 19700
rect 38335 19669 38347 19672
rect 38289 19663 38347 19669
rect 38654 19660 38660 19672
rect 38712 19700 38718 19712
rect 39025 19703 39083 19709
rect 39025 19700 39037 19703
rect 38712 19672 39037 19700
rect 38712 19660 38718 19672
rect 39025 19669 39037 19672
rect 39071 19700 39083 19703
rect 39850 19700 39856 19712
rect 39071 19672 39856 19700
rect 39071 19669 39083 19672
rect 39025 19663 39083 19669
rect 39850 19660 39856 19672
rect 39908 19660 39914 19712
rect 40034 19660 40040 19712
rect 40092 19660 40098 19712
rect 45278 19660 45284 19712
rect 45336 19700 45342 19712
rect 49237 19703 49295 19709
rect 49237 19700 49249 19703
rect 45336 19672 49249 19700
rect 45336 19660 45342 19672
rect 49237 19669 49249 19672
rect 49283 19669 49295 19703
rect 49237 19663 49295 19669
rect 1104 19610 49864 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 27950 19610
rect 28002 19558 28014 19610
rect 28066 19558 28078 19610
rect 28130 19558 28142 19610
rect 28194 19558 28206 19610
rect 28258 19558 37950 19610
rect 38002 19558 38014 19610
rect 38066 19558 38078 19610
rect 38130 19558 38142 19610
rect 38194 19558 38206 19610
rect 38258 19558 47950 19610
rect 48002 19558 48014 19610
rect 48066 19558 48078 19610
rect 48130 19558 48142 19610
rect 48194 19558 48206 19610
rect 48258 19558 49864 19610
rect 1104 19536 49864 19558
rect 9306 19496 9312 19508
rect 3528 19468 9312 19496
rect 2777 19431 2835 19437
rect 2777 19397 2789 19431
rect 2823 19428 2835 19431
rect 2866 19428 2872 19440
rect 2823 19400 2872 19428
rect 2823 19397 2835 19400
rect 2777 19391 2835 19397
rect 2866 19388 2872 19400
rect 2924 19388 2930 19440
rect 1765 19363 1823 19369
rect 1765 19329 1777 19363
rect 1811 19360 1823 19363
rect 3528 19360 3556 19468
rect 9306 19456 9312 19468
rect 9364 19456 9370 19508
rect 10042 19456 10048 19508
rect 10100 19496 10106 19508
rect 10965 19499 11023 19505
rect 10965 19496 10977 19499
rect 10100 19468 10977 19496
rect 10100 19456 10106 19468
rect 10965 19465 10977 19468
rect 11011 19465 11023 19499
rect 10965 19459 11023 19465
rect 13354 19456 13360 19508
rect 13412 19496 13418 19508
rect 14461 19499 14519 19505
rect 14461 19496 14473 19499
rect 13412 19468 14473 19496
rect 13412 19456 13418 19468
rect 14461 19465 14473 19468
rect 14507 19465 14519 19499
rect 14461 19459 14519 19465
rect 14829 19499 14887 19505
rect 14829 19465 14841 19499
rect 14875 19496 14887 19499
rect 15010 19496 15016 19508
rect 14875 19468 15016 19496
rect 14875 19465 14887 19468
rect 14829 19459 14887 19465
rect 15010 19456 15016 19468
rect 15068 19456 15074 19508
rect 16850 19456 16856 19508
rect 16908 19456 16914 19508
rect 17313 19499 17371 19505
rect 17313 19465 17325 19499
rect 17359 19496 17371 19499
rect 19334 19496 19340 19508
rect 17359 19468 19340 19496
rect 17359 19465 17371 19468
rect 17313 19459 17371 19465
rect 19334 19456 19340 19468
rect 19392 19456 19398 19508
rect 19702 19456 19708 19508
rect 19760 19496 19766 19508
rect 20717 19499 20775 19505
rect 20717 19496 20729 19499
rect 19760 19468 20729 19496
rect 19760 19456 19766 19468
rect 20717 19465 20729 19468
rect 20763 19465 20775 19499
rect 20717 19459 20775 19465
rect 21177 19499 21235 19505
rect 21177 19465 21189 19499
rect 21223 19496 21235 19499
rect 23842 19496 23848 19508
rect 21223 19468 23848 19496
rect 21223 19465 21235 19468
rect 21177 19459 21235 19465
rect 23842 19456 23848 19468
rect 23900 19456 23906 19508
rect 25774 19496 25780 19508
rect 24136 19468 25780 19496
rect 4430 19388 4436 19440
rect 4488 19388 4494 19440
rect 10321 19431 10379 19437
rect 5276 19400 9352 19428
rect 1811 19332 3556 19360
rect 3605 19363 3663 19369
rect 1811 19329 1823 19332
rect 1765 19323 1823 19329
rect 3605 19329 3617 19363
rect 3651 19360 3663 19363
rect 5276 19360 5304 19400
rect 3651 19332 5304 19360
rect 3651 19329 3663 19332
rect 3605 19323 3663 19329
rect 5350 19320 5356 19372
rect 5408 19320 5414 19372
rect 9324 19292 9352 19400
rect 10321 19397 10333 19431
rect 10367 19428 10379 19431
rect 12618 19428 12624 19440
rect 10367 19400 12624 19428
rect 10367 19397 10379 19400
rect 10321 19391 10379 19397
rect 12618 19388 12624 19400
rect 12676 19388 12682 19440
rect 13538 19388 13544 19440
rect 13596 19388 13602 19440
rect 16117 19431 16175 19437
rect 16117 19397 16129 19431
rect 16163 19428 16175 19431
rect 16758 19428 16764 19440
rect 16163 19400 16764 19428
rect 16163 19397 16175 19400
rect 16117 19391 16175 19397
rect 16758 19388 16764 19400
rect 16816 19388 16822 19440
rect 18598 19428 18604 19440
rect 18064 19400 18604 19428
rect 10870 19360 10876 19372
rect 9600 19332 10876 19360
rect 9600 19292 9628 19332
rect 10870 19320 10876 19332
rect 10928 19320 10934 19372
rect 11146 19320 11152 19372
rect 11204 19320 11210 19372
rect 11701 19363 11759 19369
rect 11701 19329 11713 19363
rect 11747 19360 11759 19363
rect 12066 19360 12072 19372
rect 11747 19332 12072 19360
rect 11747 19329 11759 19332
rect 11701 19323 11759 19329
rect 12066 19320 12072 19332
rect 12124 19320 12130 19372
rect 12710 19320 12716 19372
rect 12768 19320 12774 19372
rect 15378 19360 15384 19372
rect 15120 19332 15384 19360
rect 9324 19264 9628 19292
rect 9674 19252 9680 19304
rect 9732 19252 9738 19304
rect 11330 19252 11336 19304
rect 11388 19292 11394 19304
rect 12253 19295 12311 19301
rect 12253 19292 12265 19295
rect 11388 19264 12265 19292
rect 11388 19252 11394 19264
rect 12253 19261 12265 19264
rect 12299 19261 12311 19295
rect 12253 19255 12311 19261
rect 12989 19295 13047 19301
rect 12989 19261 13001 19295
rect 13035 19292 13047 19295
rect 15013 19295 15071 19301
rect 13035 19264 14964 19292
rect 13035 19261 13047 19264
rect 12989 19255 13047 19261
rect 9398 19184 9404 19236
rect 9456 19224 9462 19236
rect 11238 19224 11244 19236
rect 9456 19196 11244 19224
rect 9456 19184 9462 19196
rect 11238 19184 11244 19196
rect 11296 19184 11302 19236
rect 14936 19224 14964 19264
rect 15013 19261 15025 19295
rect 15059 19292 15071 19295
rect 15120 19292 15148 19332
rect 15378 19320 15384 19332
rect 15436 19320 15442 19372
rect 18064 19369 18092 19400
rect 18598 19388 18604 19400
rect 18656 19388 18662 19440
rect 20530 19428 20536 19440
rect 19550 19400 20536 19428
rect 20530 19388 20536 19400
rect 20588 19388 20594 19440
rect 21085 19431 21143 19437
rect 21085 19397 21097 19431
rect 21131 19428 21143 19431
rect 21726 19428 21732 19440
rect 21131 19400 21732 19428
rect 21131 19397 21143 19400
rect 21085 19391 21143 19397
rect 21726 19388 21732 19400
rect 21784 19388 21790 19440
rect 22738 19388 22744 19440
rect 22796 19388 22802 19440
rect 23753 19431 23811 19437
rect 23753 19397 23765 19431
rect 23799 19428 23811 19431
rect 24026 19428 24032 19440
rect 23799 19400 24032 19428
rect 23799 19397 23811 19400
rect 23753 19391 23811 19397
rect 24026 19388 24032 19400
rect 24084 19428 24090 19440
rect 24136 19428 24164 19468
rect 25774 19456 25780 19468
rect 25832 19456 25838 19508
rect 25958 19456 25964 19508
rect 26016 19496 26022 19508
rect 27338 19496 27344 19508
rect 26016 19468 27344 19496
rect 26016 19456 26022 19468
rect 27338 19456 27344 19468
rect 27396 19496 27402 19508
rect 27706 19496 27712 19508
rect 27396 19468 27712 19496
rect 27396 19456 27402 19468
rect 27706 19456 27712 19468
rect 27764 19456 27770 19508
rect 28442 19456 28448 19508
rect 28500 19456 28506 19508
rect 29733 19499 29791 19505
rect 29733 19496 29745 19499
rect 29012 19468 29745 19496
rect 24084 19400 24164 19428
rect 24084 19388 24090 19400
rect 24762 19388 24768 19440
rect 24820 19388 24826 19440
rect 25222 19388 25228 19440
rect 25280 19428 25286 19440
rect 25280 19400 26648 19428
rect 25280 19388 25286 19400
rect 17221 19363 17279 19369
rect 17221 19329 17233 19363
rect 17267 19329 17279 19363
rect 17221 19323 17279 19329
rect 18049 19363 18107 19369
rect 18049 19329 18061 19363
rect 18095 19329 18107 19363
rect 18049 19323 18107 19329
rect 15059 19264 15148 19292
rect 15059 19261 15071 19264
rect 15013 19255 15071 19261
rect 15286 19252 15292 19304
rect 15344 19292 15350 19304
rect 15565 19295 15623 19301
rect 15565 19292 15577 19295
rect 15344 19264 15577 19292
rect 15344 19252 15350 19264
rect 15565 19261 15577 19264
rect 15611 19261 15623 19295
rect 15565 19255 15623 19261
rect 15746 19252 15752 19304
rect 15804 19292 15810 19304
rect 15804 19264 16344 19292
rect 15804 19252 15810 19264
rect 16022 19224 16028 19236
rect 14936 19196 16028 19224
rect 16022 19184 16028 19196
rect 16080 19184 16086 19236
rect 2314 19116 2320 19168
rect 2372 19156 2378 19168
rect 5445 19159 5503 19165
rect 5445 19156 5457 19159
rect 2372 19128 5457 19156
rect 2372 19116 2378 19128
rect 5445 19125 5457 19128
rect 5491 19125 5503 19159
rect 5445 19119 5503 19125
rect 8386 19116 8392 19168
rect 8444 19156 8450 19168
rect 11882 19156 11888 19168
rect 8444 19128 11888 19156
rect 8444 19116 8450 19128
rect 11882 19116 11888 19128
rect 11940 19116 11946 19168
rect 16206 19116 16212 19168
rect 16264 19116 16270 19168
rect 16316 19156 16344 19264
rect 16758 19252 16764 19304
rect 16816 19292 16822 19304
rect 17236 19292 17264 19323
rect 20070 19320 20076 19372
rect 20128 19320 20134 19372
rect 22005 19363 22063 19369
rect 21284 19332 21496 19360
rect 16816 19264 17264 19292
rect 16816 19252 16822 19264
rect 17402 19252 17408 19304
rect 17460 19252 17466 19304
rect 18325 19295 18383 19301
rect 18325 19261 18337 19295
rect 18371 19292 18383 19295
rect 18371 19264 19932 19292
rect 18371 19261 18383 19264
rect 18325 19255 18383 19261
rect 19904 19224 19932 19264
rect 20162 19252 20168 19304
rect 20220 19292 20226 19304
rect 21284 19292 21312 19332
rect 20220 19264 21312 19292
rect 21361 19295 21419 19301
rect 20220 19252 20226 19264
rect 21361 19261 21373 19295
rect 21407 19261 21419 19295
rect 21468 19292 21496 19332
rect 22005 19329 22017 19363
rect 22051 19360 22063 19363
rect 22922 19360 22928 19372
rect 22051 19332 22928 19360
rect 22051 19329 22063 19332
rect 22005 19323 22063 19329
rect 22922 19320 22928 19332
rect 22980 19320 22986 19372
rect 23474 19320 23480 19372
rect 23532 19320 23538 19372
rect 25498 19320 25504 19372
rect 25556 19360 25562 19372
rect 25958 19360 25964 19372
rect 25556 19332 25964 19360
rect 25556 19320 25562 19332
rect 25958 19320 25964 19332
rect 26016 19360 26022 19372
rect 26145 19363 26203 19369
rect 26016 19332 26096 19360
rect 26016 19320 26022 19332
rect 25130 19292 25136 19304
rect 21468 19264 25136 19292
rect 21361 19255 21419 19261
rect 20438 19224 20444 19236
rect 19904 19196 20444 19224
rect 20438 19184 20444 19196
rect 20496 19184 20502 19236
rect 21376 19224 21404 19255
rect 25130 19252 25136 19264
rect 25188 19252 25194 19304
rect 26068 19224 26096 19332
rect 26145 19329 26157 19363
rect 26191 19360 26203 19363
rect 26620 19360 26648 19400
rect 28258 19388 28264 19440
rect 28316 19428 28322 19440
rect 28534 19428 28540 19440
rect 28316 19400 28540 19428
rect 28316 19388 28322 19400
rect 28534 19388 28540 19400
rect 28592 19388 28598 19440
rect 28813 19431 28871 19437
rect 28813 19397 28825 19431
rect 28859 19428 28871 19431
rect 29012 19428 29040 19468
rect 29733 19465 29745 19468
rect 29779 19465 29791 19499
rect 29733 19459 29791 19465
rect 30006 19456 30012 19508
rect 30064 19496 30070 19508
rect 30193 19499 30251 19505
rect 30193 19496 30205 19499
rect 30064 19468 30205 19496
rect 30064 19456 30070 19468
rect 30193 19465 30205 19468
rect 30239 19465 30251 19499
rect 30193 19459 30251 19465
rect 30742 19456 30748 19508
rect 30800 19456 30806 19508
rect 32309 19499 32367 19505
rect 32309 19465 32321 19499
rect 32355 19496 32367 19499
rect 32858 19496 32864 19508
rect 32355 19468 32864 19496
rect 32355 19465 32367 19468
rect 32309 19459 32367 19465
rect 32858 19456 32864 19468
rect 32916 19456 32922 19508
rect 33505 19499 33563 19505
rect 33505 19465 33517 19499
rect 33551 19465 33563 19499
rect 33505 19459 33563 19465
rect 30760 19428 30788 19456
rect 28859 19400 29040 19428
rect 29840 19400 30788 19428
rect 28859 19397 28871 19400
rect 28813 19391 28871 19397
rect 27617 19363 27675 19369
rect 26191 19332 26372 19360
rect 26191 19329 26203 19332
rect 26145 19323 26203 19329
rect 26237 19295 26295 19301
rect 26237 19261 26249 19295
rect 26283 19261 26295 19295
rect 26237 19255 26295 19261
rect 26252 19224 26280 19255
rect 21376 19196 22094 19224
rect 26068 19196 26280 19224
rect 26344 19224 26372 19332
rect 26418 19294 26424 19346
rect 26476 19294 26482 19346
rect 26620 19334 27476 19360
rect 27617 19334 27629 19363
rect 26620 19332 27629 19334
rect 27448 19329 27629 19332
rect 27663 19360 27675 19363
rect 28626 19360 28632 19372
rect 27663 19332 28632 19360
rect 27663 19329 27675 19332
rect 27448 19323 27675 19329
rect 27448 19306 27660 19323
rect 28626 19320 28632 19332
rect 28684 19320 28690 19372
rect 26421 19261 26433 19294
rect 26467 19261 26479 19294
rect 26602 19292 26608 19304
rect 26421 19255 26479 19261
rect 26528 19264 26608 19292
rect 26528 19224 26556 19264
rect 26602 19252 26608 19264
rect 26660 19252 26666 19304
rect 27709 19295 27767 19301
rect 27709 19261 27721 19295
rect 27755 19261 27767 19295
rect 27709 19255 27767 19261
rect 27893 19295 27951 19301
rect 27893 19261 27905 19295
rect 27939 19292 27951 19295
rect 27939 19264 28672 19292
rect 27939 19261 27951 19264
rect 27893 19255 27951 19261
rect 26344 19196 26556 19224
rect 27724 19224 27752 19255
rect 28644 19236 28672 19264
rect 28718 19252 28724 19304
rect 28776 19292 28782 19304
rect 28905 19295 28963 19301
rect 28905 19292 28917 19295
rect 28776 19264 28917 19292
rect 28776 19252 28782 19264
rect 28905 19261 28917 19264
rect 28951 19261 28963 19295
rect 28905 19255 28963 19261
rect 29089 19295 29147 19301
rect 29089 19261 29101 19295
rect 29135 19292 29147 19295
rect 29178 19292 29184 19304
rect 29135 19264 29184 19292
rect 29135 19261 29147 19264
rect 29089 19255 29147 19261
rect 29178 19252 29184 19264
rect 29236 19292 29242 19304
rect 29840 19292 29868 19400
rect 32674 19388 32680 19440
rect 32732 19388 32738 19440
rect 32766 19388 32772 19440
rect 32824 19388 32830 19440
rect 33520 19428 33548 19459
rect 33962 19456 33968 19508
rect 34020 19496 34026 19508
rect 34422 19496 34428 19508
rect 34020 19468 34428 19496
rect 34020 19456 34026 19468
rect 34422 19456 34428 19468
rect 34480 19456 34486 19508
rect 34701 19499 34759 19505
rect 34701 19465 34713 19499
rect 34747 19496 34759 19499
rect 35618 19496 35624 19508
rect 34747 19468 35624 19496
rect 34747 19465 34759 19468
rect 34701 19459 34759 19465
rect 35618 19456 35624 19468
rect 35676 19456 35682 19508
rect 35894 19456 35900 19508
rect 35952 19456 35958 19508
rect 37918 19456 37924 19508
rect 37976 19496 37982 19508
rect 38378 19496 38384 19508
rect 37976 19468 38384 19496
rect 37976 19456 37982 19468
rect 38378 19456 38384 19468
rect 38436 19456 38442 19508
rect 40126 19456 40132 19508
rect 40184 19456 40190 19508
rect 40402 19456 40408 19508
rect 40460 19496 40466 19508
rect 40589 19499 40647 19505
rect 40589 19496 40601 19499
rect 40460 19468 40601 19496
rect 40460 19456 40466 19468
rect 40589 19465 40601 19468
rect 40635 19496 40647 19499
rect 41325 19499 41383 19505
rect 41325 19496 41337 19499
rect 40635 19468 41337 19496
rect 40635 19465 40647 19468
rect 40589 19459 40647 19465
rect 41325 19465 41337 19468
rect 41371 19496 41383 19499
rect 49234 19496 49240 19508
rect 41371 19468 49240 19496
rect 41371 19465 41383 19468
rect 41325 19459 41383 19465
rect 49234 19456 49240 19468
rect 49292 19456 49298 19508
rect 33520 19400 35204 19428
rect 30374 19320 30380 19372
rect 30432 19360 30438 19372
rect 30745 19363 30803 19369
rect 30745 19360 30757 19363
rect 30432 19332 30757 19360
rect 30432 19320 30438 19332
rect 30745 19329 30757 19332
rect 30791 19329 30803 19363
rect 30745 19323 30803 19329
rect 31573 19363 31631 19369
rect 31573 19329 31585 19363
rect 31619 19360 31631 19363
rect 32306 19360 32312 19372
rect 31619 19332 32312 19360
rect 31619 19329 31631 19332
rect 31573 19323 31631 19329
rect 32306 19320 32312 19332
rect 32364 19360 32370 19372
rect 32582 19360 32588 19372
rect 32364 19332 32588 19360
rect 32364 19320 32370 19332
rect 32582 19320 32588 19332
rect 32640 19320 32646 19372
rect 33873 19363 33931 19369
rect 33873 19329 33885 19363
rect 33919 19360 33931 19363
rect 34238 19360 34244 19372
rect 33919 19332 34244 19360
rect 33919 19329 33931 19332
rect 33873 19323 33931 19329
rect 34238 19320 34244 19332
rect 34296 19320 34302 19372
rect 34606 19320 34612 19372
rect 34664 19360 34670 19372
rect 35069 19363 35127 19369
rect 35069 19360 35081 19363
rect 34664 19332 35081 19360
rect 34664 19320 34670 19332
rect 35069 19329 35081 19332
rect 35115 19329 35127 19363
rect 35176 19360 35204 19400
rect 36538 19388 36544 19440
rect 36596 19428 36602 19440
rect 38470 19428 38476 19440
rect 36596 19400 38476 19428
rect 36596 19388 36602 19400
rect 38470 19388 38476 19400
rect 38528 19388 38534 19440
rect 39482 19428 39488 19440
rect 39422 19400 39488 19428
rect 39482 19388 39488 19400
rect 39540 19388 39546 19440
rect 40497 19431 40555 19437
rect 40497 19397 40509 19431
rect 40543 19428 40555 19431
rect 48406 19428 48412 19440
rect 40543 19400 48412 19428
rect 40543 19397 40555 19400
rect 40497 19391 40555 19397
rect 48406 19388 48412 19400
rect 48464 19388 48470 19440
rect 36078 19360 36084 19372
rect 35176 19332 36084 19360
rect 35069 19323 35127 19329
rect 36078 19320 36084 19332
rect 36136 19320 36142 19372
rect 36262 19320 36268 19372
rect 36320 19320 36326 19372
rect 36354 19320 36360 19372
rect 36412 19320 36418 19372
rect 37734 19320 37740 19372
rect 37792 19360 37798 19372
rect 37921 19363 37979 19369
rect 37921 19360 37933 19363
rect 37792 19332 37933 19360
rect 37792 19320 37798 19332
rect 37921 19329 37933 19332
rect 37967 19329 37979 19363
rect 37921 19323 37979 19329
rect 40126 19320 40132 19372
rect 40184 19360 40190 19372
rect 41230 19360 41236 19372
rect 40184 19332 41236 19360
rect 40184 19320 40190 19332
rect 41230 19320 41236 19332
rect 41288 19360 41294 19372
rect 45278 19360 45284 19372
rect 41288 19332 45284 19360
rect 41288 19320 41294 19332
rect 45278 19320 45284 19332
rect 45336 19320 45342 19372
rect 48593 19363 48651 19369
rect 48593 19329 48605 19363
rect 48639 19360 48651 19363
rect 49142 19360 49148 19372
rect 48639 19332 49148 19360
rect 48639 19329 48651 19332
rect 48593 19323 48651 19329
rect 49142 19320 49148 19332
rect 49200 19320 49206 19372
rect 31478 19292 31484 19304
rect 29236 19264 29868 19292
rect 29932 19264 31484 19292
rect 29236 19252 29242 19264
rect 27798 19224 27804 19236
rect 27724 19196 27804 19224
rect 19794 19156 19800 19168
rect 16316 19128 19800 19156
rect 19794 19116 19800 19128
rect 19852 19116 19858 19168
rect 20349 19159 20407 19165
rect 20349 19125 20361 19159
rect 20395 19156 20407 19159
rect 20530 19156 20536 19168
rect 20395 19128 20536 19156
rect 20395 19125 20407 19128
rect 20349 19119 20407 19125
rect 20530 19116 20536 19128
rect 20588 19156 20594 19168
rect 21542 19156 21548 19168
rect 20588 19128 21548 19156
rect 20588 19116 20594 19128
rect 21542 19116 21548 19128
rect 21600 19116 21606 19168
rect 22066 19156 22094 19196
rect 27798 19184 27804 19196
rect 27856 19224 27862 19236
rect 28534 19224 28540 19236
rect 27856 19196 28540 19224
rect 27856 19184 27862 19196
rect 28534 19184 28540 19196
rect 28592 19184 28598 19236
rect 28626 19184 28632 19236
rect 28684 19224 28690 19236
rect 29932 19224 29960 19264
rect 31478 19252 31484 19264
rect 31536 19252 31542 19304
rect 32861 19295 32919 19301
rect 32861 19261 32873 19295
rect 32907 19261 32919 19295
rect 32861 19255 32919 19261
rect 34149 19295 34207 19301
rect 34149 19261 34161 19295
rect 34195 19261 34207 19295
rect 34149 19255 34207 19261
rect 35161 19295 35219 19301
rect 35161 19261 35173 19295
rect 35207 19292 35219 19295
rect 35250 19292 35256 19304
rect 35207 19264 35256 19292
rect 35207 19261 35219 19264
rect 35161 19255 35219 19261
rect 31110 19224 31116 19236
rect 28684 19196 29960 19224
rect 30024 19196 31116 19224
rect 28684 19184 28690 19196
rect 25222 19156 25228 19168
rect 22066 19128 25228 19156
rect 25222 19116 25228 19128
rect 25280 19116 25286 19168
rect 25774 19116 25780 19168
rect 25832 19116 25838 19168
rect 27246 19116 27252 19168
rect 27304 19116 27310 19168
rect 27982 19116 27988 19168
rect 28040 19156 28046 19168
rect 30024 19156 30052 19196
rect 31110 19184 31116 19196
rect 31168 19184 31174 19236
rect 32876 19224 32904 19255
rect 32784 19196 32904 19224
rect 34164 19224 34192 19255
rect 35250 19252 35256 19264
rect 35308 19252 35314 19304
rect 35345 19295 35403 19301
rect 35345 19261 35357 19295
rect 35391 19292 35403 19295
rect 35894 19292 35900 19304
rect 35391 19264 35900 19292
rect 35391 19261 35403 19264
rect 35345 19255 35403 19261
rect 35894 19252 35900 19264
rect 35952 19252 35958 19304
rect 36449 19295 36507 19301
rect 36449 19292 36461 19295
rect 36372 19264 36461 19292
rect 36372 19236 36400 19264
rect 36449 19261 36461 19264
rect 36495 19261 36507 19295
rect 36449 19255 36507 19261
rect 38194 19252 38200 19304
rect 38252 19252 38258 19304
rect 39206 19252 39212 19304
rect 39264 19292 39270 19304
rect 40681 19295 40739 19301
rect 40681 19292 40693 19295
rect 39264 19264 40693 19292
rect 39264 19252 39270 19264
rect 40681 19261 40693 19264
rect 40727 19261 40739 19295
rect 41138 19292 41144 19304
rect 40681 19255 40739 19261
rect 40788 19264 41144 19292
rect 34164 19196 36308 19224
rect 32784 19168 32812 19196
rect 28040 19128 30052 19156
rect 28040 19116 28046 19128
rect 30374 19116 30380 19168
rect 30432 19116 30438 19168
rect 32766 19116 32772 19168
rect 32824 19116 32830 19168
rect 35894 19116 35900 19168
rect 35952 19156 35958 19168
rect 36170 19156 36176 19168
rect 35952 19128 36176 19156
rect 35952 19116 35958 19128
rect 36170 19116 36176 19128
rect 36228 19116 36234 19168
rect 36280 19156 36308 19196
rect 36354 19184 36360 19236
rect 36412 19184 36418 19236
rect 36906 19184 36912 19236
rect 36964 19184 36970 19236
rect 37366 19184 37372 19236
rect 37424 19224 37430 19236
rect 37918 19224 37924 19236
rect 37424 19196 37924 19224
rect 37424 19184 37430 19196
rect 37918 19184 37924 19196
rect 37976 19184 37982 19236
rect 39482 19184 39488 19236
rect 39540 19224 39546 19236
rect 40218 19224 40224 19236
rect 39540 19196 40224 19224
rect 39540 19184 39546 19196
rect 40218 19184 40224 19196
rect 40276 19224 40282 19236
rect 40788 19224 40816 19264
rect 41138 19252 41144 19264
rect 41196 19252 41202 19304
rect 49329 19227 49387 19233
rect 49329 19224 49341 19227
rect 40276 19196 40816 19224
rect 40880 19196 49341 19224
rect 40276 19184 40282 19196
rect 37458 19156 37464 19168
rect 36280 19128 37464 19156
rect 37458 19116 37464 19128
rect 37516 19116 37522 19168
rect 38286 19116 38292 19168
rect 38344 19156 38350 19168
rect 39669 19159 39727 19165
rect 39669 19156 39681 19159
rect 38344 19128 39681 19156
rect 38344 19116 38350 19128
rect 39669 19125 39681 19128
rect 39715 19125 39727 19159
rect 39669 19119 39727 19125
rect 39758 19116 39764 19168
rect 39816 19156 39822 19168
rect 40880 19156 40908 19196
rect 49329 19193 49341 19196
rect 49375 19193 49387 19227
rect 49329 19187 49387 19193
rect 39816 19128 40908 19156
rect 39816 19116 39822 19128
rect 41138 19116 41144 19168
rect 41196 19156 41202 19168
rect 41598 19156 41604 19168
rect 41196 19128 41604 19156
rect 41196 19116 41202 19128
rect 41598 19116 41604 19128
rect 41656 19116 41662 19168
rect 48777 19159 48835 19165
rect 48777 19125 48789 19159
rect 48823 19156 48835 19159
rect 49050 19156 49056 19168
rect 48823 19128 49056 19156
rect 48823 19125 48835 19128
rect 48777 19119 48835 19125
rect 49050 19116 49056 19128
rect 49108 19116 49114 19168
rect 1104 19066 49864 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 32950 19066
rect 33002 19014 33014 19066
rect 33066 19014 33078 19066
rect 33130 19014 33142 19066
rect 33194 19014 33206 19066
rect 33258 19014 42950 19066
rect 43002 19014 43014 19066
rect 43066 19014 43078 19066
rect 43130 19014 43142 19066
rect 43194 19014 43206 19066
rect 43258 19014 49864 19066
rect 1104 18992 49864 19014
rect 11054 18952 11060 18964
rect 8956 18924 11060 18952
rect 3786 18776 3792 18828
rect 3844 18816 3850 18828
rect 4433 18819 4491 18825
rect 4433 18816 4445 18819
rect 3844 18788 4445 18816
rect 3844 18776 3850 18788
rect 4433 18785 4445 18788
rect 4479 18785 4491 18819
rect 8662 18816 8668 18828
rect 4433 18779 4491 18785
rect 5000 18788 8668 18816
rect 1765 18751 1823 18757
rect 1765 18717 1777 18751
rect 1811 18748 1823 18751
rect 4065 18751 4123 18757
rect 1811 18720 3924 18748
rect 1811 18717 1823 18720
rect 1765 18711 1823 18717
rect 2774 18640 2780 18692
rect 2832 18640 2838 18692
rect 3896 18680 3924 18720
rect 4065 18717 4077 18751
rect 4111 18748 4123 18751
rect 5000 18748 5028 18788
rect 8662 18776 8668 18788
rect 8720 18776 8726 18828
rect 4111 18720 5028 18748
rect 8205 18751 8263 18757
rect 4111 18717 4123 18720
rect 4065 18711 4123 18717
rect 8205 18717 8217 18751
rect 8251 18748 8263 18751
rect 8956 18748 8984 18924
rect 11054 18912 11060 18924
rect 11112 18912 11118 18964
rect 11422 18912 11428 18964
rect 11480 18952 11486 18964
rect 12529 18955 12587 18961
rect 12529 18952 12541 18955
rect 11480 18924 12541 18952
rect 11480 18912 11486 18924
rect 12529 18921 12541 18924
rect 12575 18921 12587 18955
rect 12529 18915 12587 18921
rect 15102 18912 15108 18964
rect 15160 18952 15166 18964
rect 15160 18924 15700 18952
rect 15160 18912 15166 18924
rect 10870 18844 10876 18896
rect 10928 18844 10934 18896
rect 11882 18844 11888 18896
rect 11940 18844 11946 18896
rect 13541 18887 13599 18893
rect 13541 18884 13553 18887
rect 13096 18856 13553 18884
rect 9125 18819 9183 18825
rect 9125 18785 9137 18819
rect 9171 18816 9183 18819
rect 10594 18816 10600 18828
rect 9171 18788 10600 18816
rect 9171 18785 9183 18788
rect 9125 18779 9183 18785
rect 10594 18776 10600 18788
rect 10652 18776 10658 18828
rect 13096 18816 13124 18856
rect 13541 18853 13553 18856
rect 13587 18884 13599 18887
rect 13817 18887 13875 18893
rect 13817 18884 13829 18887
rect 13587 18856 13829 18884
rect 13587 18853 13599 18856
rect 13541 18847 13599 18853
rect 13817 18853 13829 18856
rect 13863 18884 13875 18887
rect 14090 18884 14096 18896
rect 13863 18856 14096 18884
rect 13863 18853 13875 18856
rect 13817 18847 13875 18853
rect 14090 18844 14096 18856
rect 14148 18844 14154 18896
rect 11900 18788 13124 18816
rect 13173 18819 13231 18825
rect 11900 18760 11928 18788
rect 13173 18785 13185 18819
rect 13219 18816 13231 18819
rect 13354 18816 13360 18828
rect 13219 18788 13360 18816
rect 13219 18785 13231 18788
rect 13173 18779 13231 18785
rect 13354 18776 13360 18788
rect 13412 18776 13418 18828
rect 14274 18776 14280 18828
rect 14332 18776 14338 18828
rect 14553 18819 14611 18825
rect 14553 18785 14565 18819
rect 14599 18816 14611 18819
rect 15286 18816 15292 18828
rect 14599 18788 15292 18816
rect 14599 18785 14611 18788
rect 14553 18779 14611 18785
rect 15286 18776 15292 18788
rect 15344 18776 15350 18828
rect 11241 18751 11299 18757
rect 11241 18748 11253 18751
rect 8251 18720 8984 18748
rect 10534 18720 11253 18748
rect 8251 18717 8263 18720
rect 8205 18711 8263 18717
rect 11241 18717 11253 18720
rect 11287 18748 11299 18751
rect 11514 18748 11520 18760
rect 11287 18720 11520 18748
rect 11287 18717 11299 18720
rect 11241 18711 11299 18717
rect 11514 18708 11520 18720
rect 11572 18748 11578 18760
rect 11882 18748 11888 18760
rect 11572 18720 11888 18748
rect 11572 18708 11578 18720
rect 11882 18708 11888 18720
rect 11940 18708 11946 18760
rect 12069 18751 12127 18757
rect 12069 18717 12081 18751
rect 12115 18748 12127 18751
rect 12115 18720 12434 18748
rect 12115 18717 12127 18720
rect 12069 18711 12127 18717
rect 3896 18652 8432 18680
rect 8294 18572 8300 18624
rect 8352 18572 8358 18624
rect 8404 18612 8432 18652
rect 9398 18640 9404 18692
rect 9456 18640 9462 18692
rect 11698 18680 11704 18692
rect 10704 18652 11704 18680
rect 10704 18612 10732 18652
rect 11698 18640 11704 18652
rect 11756 18640 11762 18692
rect 8404 18584 10732 18612
rect 12406 18612 12434 18720
rect 12618 18708 12624 18760
rect 12676 18748 12682 18760
rect 12897 18751 12955 18757
rect 12897 18748 12909 18751
rect 12676 18720 12909 18748
rect 12676 18708 12682 18720
rect 12897 18717 12909 18720
rect 12943 18717 12955 18751
rect 12897 18711 12955 18717
rect 13262 18708 13268 18760
rect 13320 18748 13326 18760
rect 13446 18748 13452 18760
rect 13320 18720 13452 18748
rect 13320 18708 13326 18720
rect 13446 18708 13452 18720
rect 13504 18708 13510 18760
rect 15672 18748 15700 18924
rect 16022 18912 16028 18964
rect 16080 18912 16086 18964
rect 16482 18912 16488 18964
rect 16540 18952 16546 18964
rect 16945 18955 17003 18961
rect 16945 18952 16957 18955
rect 16540 18924 16957 18952
rect 16540 18912 16546 18924
rect 16945 18921 16957 18924
rect 16991 18921 17003 18955
rect 16945 18915 17003 18921
rect 17034 18912 17040 18964
rect 17092 18952 17098 18964
rect 18141 18955 18199 18961
rect 18141 18952 18153 18955
rect 17092 18924 18153 18952
rect 17092 18912 17098 18924
rect 18141 18921 18153 18924
rect 18187 18921 18199 18955
rect 18141 18915 18199 18921
rect 19610 18912 19616 18964
rect 19668 18952 19674 18964
rect 19889 18955 19947 18961
rect 19889 18952 19901 18955
rect 19668 18924 19901 18952
rect 19668 18912 19674 18924
rect 19889 18921 19901 18924
rect 19935 18921 19947 18955
rect 19889 18915 19947 18921
rect 21082 18912 21088 18964
rect 21140 18912 21146 18964
rect 24581 18955 24639 18961
rect 24581 18952 24593 18955
rect 22204 18924 24593 18952
rect 15930 18844 15936 18896
rect 15988 18884 15994 18896
rect 15988 18856 17632 18884
rect 15988 18844 15994 18856
rect 16298 18776 16304 18828
rect 16356 18816 16362 18828
rect 17497 18819 17555 18825
rect 17497 18816 17509 18819
rect 16356 18788 17509 18816
rect 16356 18776 16362 18788
rect 17497 18785 17509 18788
rect 17543 18785 17555 18819
rect 17604 18816 17632 18856
rect 17678 18844 17684 18896
rect 17736 18884 17742 18896
rect 17736 18856 20576 18884
rect 17736 18844 17742 18856
rect 18690 18816 18696 18828
rect 17604 18788 18696 18816
rect 17497 18779 17555 18785
rect 18690 18776 18696 18788
rect 18748 18776 18754 18828
rect 18785 18819 18843 18825
rect 18785 18785 18797 18819
rect 18831 18816 18843 18819
rect 18966 18816 18972 18828
rect 18831 18788 18972 18816
rect 18831 18785 18843 18788
rect 18785 18779 18843 18785
rect 18966 18776 18972 18788
rect 19024 18776 19030 18828
rect 20548 18825 20576 18856
rect 20533 18819 20591 18825
rect 20533 18785 20545 18819
rect 20579 18816 20591 18819
rect 21358 18816 21364 18828
rect 20579 18788 21364 18816
rect 20579 18785 20591 18788
rect 20533 18779 20591 18785
rect 21358 18776 21364 18788
rect 21416 18776 21422 18828
rect 21634 18776 21640 18828
rect 21692 18776 21698 18828
rect 16393 18751 16451 18757
rect 16393 18748 16405 18751
rect 15672 18734 16405 18748
rect 15686 18720 16405 18734
rect 16393 18717 16405 18720
rect 16439 18748 16451 18751
rect 16666 18748 16672 18760
rect 16439 18720 16672 18748
rect 16439 18717 16451 18720
rect 16393 18711 16451 18717
rect 16666 18708 16672 18720
rect 16724 18708 16730 18760
rect 17402 18708 17408 18760
rect 17460 18708 17466 18760
rect 17770 18708 17776 18760
rect 17828 18748 17834 18760
rect 18509 18751 18567 18757
rect 18509 18748 18521 18751
rect 17828 18720 18521 18748
rect 17828 18708 17834 18720
rect 18509 18717 18521 18720
rect 18555 18717 18567 18751
rect 18509 18711 18567 18717
rect 18601 18751 18659 18757
rect 18601 18717 18613 18751
rect 18647 18748 18659 18751
rect 18647 18720 18828 18748
rect 18647 18717 18659 18720
rect 18601 18711 18659 18717
rect 12989 18683 13047 18689
rect 12989 18649 13001 18683
rect 13035 18680 13047 18683
rect 13035 18652 14964 18680
rect 13035 18649 13047 18652
rect 12989 18643 13047 18649
rect 13446 18612 13452 18624
rect 12406 18584 13452 18612
rect 13446 18572 13452 18584
rect 13504 18572 13510 18624
rect 14936 18612 14964 18652
rect 16942 18640 16948 18692
rect 17000 18680 17006 18692
rect 17313 18683 17371 18689
rect 17313 18680 17325 18683
rect 17000 18652 17325 18680
rect 17000 18640 17006 18652
rect 17313 18649 17325 18652
rect 17359 18649 17371 18683
rect 17313 18643 17371 18649
rect 15562 18612 15568 18624
rect 14936 18584 15568 18612
rect 15562 18572 15568 18584
rect 15620 18572 15626 18624
rect 16669 18615 16727 18621
rect 16669 18581 16681 18615
rect 16715 18612 16727 18615
rect 16758 18612 16764 18624
rect 16715 18584 16764 18612
rect 16715 18581 16727 18584
rect 16669 18575 16727 18581
rect 16758 18572 16764 18584
rect 16816 18572 16822 18624
rect 18800 18612 18828 18720
rect 19058 18708 19064 18760
rect 19116 18748 19122 18760
rect 20257 18751 20315 18757
rect 19116 18720 19472 18748
rect 19116 18708 19122 18720
rect 18874 18640 18880 18692
rect 18932 18680 18938 18692
rect 18932 18652 19380 18680
rect 18932 18640 18938 18652
rect 19352 18624 19380 18652
rect 19150 18612 19156 18624
rect 18800 18584 19156 18612
rect 19150 18572 19156 18584
rect 19208 18572 19214 18624
rect 19334 18572 19340 18624
rect 19392 18572 19398 18624
rect 19444 18612 19472 18720
rect 20257 18717 20269 18751
rect 20303 18748 20315 18751
rect 22204 18748 22232 18924
rect 24581 18921 24593 18924
rect 24627 18921 24639 18955
rect 24581 18915 24639 18921
rect 25130 18912 25136 18964
rect 25188 18952 25194 18964
rect 28997 18955 29055 18961
rect 28997 18952 29009 18955
rect 25188 18924 29009 18952
rect 25188 18912 25194 18924
rect 28997 18921 29009 18924
rect 29043 18921 29055 18955
rect 28997 18915 29055 18921
rect 33042 18912 33048 18964
rect 33100 18952 33106 18964
rect 33873 18955 33931 18961
rect 33873 18952 33885 18955
rect 33100 18924 33885 18952
rect 33100 18912 33106 18924
rect 33873 18921 33885 18924
rect 33919 18921 33931 18955
rect 33873 18915 33931 18921
rect 33962 18912 33968 18964
rect 34020 18952 34026 18964
rect 34149 18955 34207 18961
rect 34149 18952 34161 18955
rect 34020 18924 34161 18952
rect 34020 18912 34026 18924
rect 34149 18921 34161 18924
rect 34195 18952 34207 18955
rect 34330 18952 34336 18964
rect 34195 18924 34336 18952
rect 34195 18921 34207 18924
rect 34149 18915 34207 18921
rect 34330 18912 34336 18924
rect 34388 18912 34394 18964
rect 34514 18912 34520 18964
rect 34572 18912 34578 18964
rect 36906 18952 36912 18964
rect 34624 18924 36912 18952
rect 23658 18844 23664 18896
rect 23716 18884 23722 18896
rect 24029 18887 24087 18893
rect 24029 18884 24041 18887
rect 23716 18856 24041 18884
rect 23716 18844 23722 18856
rect 24029 18853 24041 18856
rect 24075 18884 24087 18887
rect 27893 18887 27951 18893
rect 24075 18856 25912 18884
rect 24075 18853 24087 18856
rect 24029 18847 24087 18853
rect 22281 18819 22339 18825
rect 22281 18785 22293 18819
rect 22327 18816 22339 18819
rect 22646 18816 22652 18828
rect 22327 18788 22652 18816
rect 22327 18785 22339 18788
rect 22281 18779 22339 18785
rect 22646 18776 22652 18788
rect 22704 18816 22710 18828
rect 23290 18816 23296 18828
rect 22704 18788 23296 18816
rect 22704 18776 22710 18788
rect 23290 18776 23296 18788
rect 23348 18776 23354 18828
rect 25240 18825 25268 18856
rect 25225 18819 25283 18825
rect 25225 18785 25237 18819
rect 25271 18785 25283 18819
rect 25225 18779 25283 18785
rect 25682 18776 25688 18828
rect 25740 18816 25746 18828
rect 25777 18819 25835 18825
rect 25777 18816 25789 18819
rect 25740 18788 25789 18816
rect 25740 18776 25746 18788
rect 25777 18785 25789 18788
rect 25823 18785 25835 18819
rect 25884 18816 25912 18856
rect 27893 18853 27905 18887
rect 27939 18884 27951 18887
rect 28350 18884 28356 18896
rect 27939 18856 28356 18884
rect 27939 18853 27951 18856
rect 27893 18847 27951 18853
rect 28350 18844 28356 18856
rect 28408 18844 28414 18896
rect 28902 18844 28908 18896
rect 28960 18884 28966 18896
rect 31481 18887 31539 18893
rect 31481 18884 31493 18887
rect 28960 18856 31493 18884
rect 28960 18844 28966 18856
rect 31481 18853 31493 18856
rect 31527 18853 31539 18887
rect 31481 18847 31539 18853
rect 32677 18887 32735 18893
rect 32677 18853 32689 18887
rect 32723 18884 32735 18887
rect 34624 18884 34652 18924
rect 36906 18912 36912 18924
rect 36964 18912 36970 18964
rect 37369 18955 37427 18961
rect 37369 18921 37381 18955
rect 37415 18952 37427 18955
rect 38194 18952 38200 18964
rect 37415 18924 38200 18952
rect 37415 18921 37427 18924
rect 37369 18915 37427 18921
rect 38194 18912 38200 18924
rect 38252 18912 38258 18964
rect 32723 18856 34652 18884
rect 32723 18853 32735 18856
rect 32677 18847 32735 18853
rect 37458 18844 37464 18896
rect 37516 18884 37522 18896
rect 37737 18887 37795 18893
rect 37737 18884 37749 18887
rect 37516 18856 37749 18884
rect 37516 18844 37522 18856
rect 37737 18853 37749 18856
rect 37783 18884 37795 18887
rect 38746 18884 38752 18896
rect 37783 18856 38752 18884
rect 37783 18853 37795 18856
rect 37737 18847 37795 18853
rect 38746 18844 38752 18856
rect 38804 18844 38810 18896
rect 42702 18844 42708 18896
rect 42760 18884 42766 18896
rect 49237 18887 49295 18893
rect 49237 18884 49249 18887
rect 42760 18856 49249 18884
rect 42760 18844 42766 18856
rect 49237 18853 49249 18856
rect 49283 18853 49295 18887
rect 49237 18847 49295 18853
rect 27062 18816 27068 18828
rect 25884 18788 27068 18816
rect 25777 18779 25835 18785
rect 27062 18776 27068 18788
rect 27120 18776 27126 18828
rect 27338 18776 27344 18828
rect 27396 18816 27402 18828
rect 27525 18819 27583 18825
rect 27525 18816 27537 18819
rect 27396 18788 27537 18816
rect 27396 18776 27402 18788
rect 27525 18785 27537 18788
rect 27571 18816 27583 18819
rect 29454 18816 29460 18828
rect 27571 18788 29460 18816
rect 27571 18785 27583 18788
rect 27525 18779 27583 18785
rect 29454 18776 29460 18788
rect 29512 18776 29518 18828
rect 29638 18776 29644 18828
rect 29696 18816 29702 18828
rect 30193 18819 30251 18825
rect 30193 18816 30205 18819
rect 29696 18788 30205 18816
rect 29696 18776 29702 18788
rect 30193 18785 30205 18788
rect 30239 18785 30251 18819
rect 30193 18779 30251 18785
rect 30282 18776 30288 18828
rect 30340 18776 30346 18828
rect 31938 18776 31944 18828
rect 31996 18776 32002 18828
rect 32125 18819 32183 18825
rect 32125 18785 32137 18819
rect 32171 18785 32183 18819
rect 32125 18779 32183 18785
rect 33321 18819 33379 18825
rect 33321 18785 33333 18819
rect 33367 18816 33379 18819
rect 34146 18816 34152 18828
rect 33367 18788 34152 18816
rect 33367 18785 33379 18788
rect 33321 18779 33379 18785
rect 20303 18720 22232 18748
rect 20303 18717 20315 18720
rect 20257 18711 20315 18717
rect 27430 18708 27436 18760
rect 27488 18748 27494 18760
rect 28261 18751 28319 18757
rect 27488 18720 27936 18748
rect 27488 18708 27494 18720
rect 20349 18683 20407 18689
rect 20349 18649 20361 18683
rect 20395 18680 20407 18683
rect 22278 18680 22284 18692
rect 20395 18652 22284 18680
rect 20395 18649 20407 18652
rect 20349 18643 20407 18649
rect 22278 18640 22284 18652
rect 22336 18640 22342 18692
rect 22557 18683 22615 18689
rect 22557 18649 22569 18683
rect 22603 18649 22615 18683
rect 24118 18680 24124 18692
rect 23782 18652 24124 18680
rect 22557 18643 22615 18649
rect 21174 18612 21180 18624
rect 19444 18584 21180 18612
rect 21174 18572 21180 18584
rect 21232 18572 21238 18624
rect 21450 18572 21456 18624
rect 21508 18572 21514 18624
rect 21545 18615 21603 18621
rect 21545 18581 21557 18615
rect 21591 18612 21603 18615
rect 21634 18612 21640 18624
rect 21591 18584 21640 18612
rect 21591 18581 21603 18584
rect 21545 18575 21603 18581
rect 21634 18572 21640 18584
rect 21692 18612 21698 18624
rect 22370 18612 22376 18624
rect 21692 18584 22376 18612
rect 21692 18572 21698 18584
rect 22370 18572 22376 18584
rect 22428 18572 22434 18624
rect 22572 18612 22600 18643
rect 24118 18640 24124 18652
rect 24176 18680 24182 18692
rect 24762 18680 24768 18692
rect 24176 18652 24768 18680
rect 24176 18640 24182 18652
rect 24762 18640 24768 18652
rect 24820 18640 24826 18692
rect 25038 18640 25044 18692
rect 25096 18640 25102 18692
rect 25222 18640 25228 18692
rect 25280 18680 25286 18692
rect 26053 18683 26111 18689
rect 26053 18680 26065 18683
rect 25280 18652 26065 18680
rect 25280 18640 25286 18652
rect 26053 18649 26065 18652
rect 26099 18649 26111 18683
rect 27798 18680 27804 18692
rect 27278 18652 27804 18680
rect 26053 18643 26111 18649
rect 27798 18640 27804 18652
rect 27856 18640 27862 18692
rect 27908 18680 27936 18720
rect 28261 18717 28273 18751
rect 28307 18748 28319 18751
rect 28442 18748 28448 18760
rect 28307 18720 28448 18748
rect 28307 18717 28319 18720
rect 28261 18711 28319 18717
rect 28442 18708 28448 18720
rect 28500 18708 28506 18760
rect 29178 18708 29184 18760
rect 29236 18708 29242 18760
rect 29914 18708 29920 18760
rect 29972 18748 29978 18760
rect 30101 18751 30159 18757
rect 30101 18748 30113 18751
rect 29972 18720 30113 18748
rect 29972 18708 29978 18720
rect 30101 18717 30113 18720
rect 30147 18717 30159 18751
rect 30101 18711 30159 18717
rect 28994 18680 29000 18692
rect 27908 18652 29000 18680
rect 28994 18640 29000 18652
rect 29052 18640 29058 18692
rect 32140 18680 32168 18779
rect 34146 18776 34152 18788
rect 34204 18776 34210 18828
rect 34977 18819 35035 18825
rect 34977 18785 34989 18819
rect 35023 18816 35035 18819
rect 35986 18816 35992 18828
rect 35023 18788 35992 18816
rect 35023 18785 35035 18788
rect 34977 18779 35035 18785
rect 35986 18776 35992 18788
rect 36044 18776 36050 18828
rect 37476 18816 37504 18844
rect 37016 18788 37504 18816
rect 37016 18760 37044 18788
rect 37550 18776 37556 18828
rect 37608 18816 37614 18828
rect 37608 18788 38332 18816
rect 37608 18776 37614 18788
rect 32582 18708 32588 18760
rect 32640 18748 32646 18760
rect 35621 18751 35679 18757
rect 35621 18748 35633 18751
rect 32640 18720 35633 18748
rect 32640 18708 32646 18720
rect 35621 18717 35633 18720
rect 35667 18717 35679 18751
rect 35621 18711 35679 18717
rect 36998 18708 37004 18760
rect 37056 18708 37062 18760
rect 37200 18720 38148 18748
rect 35342 18680 35348 18692
rect 32140 18652 35348 18680
rect 35342 18640 35348 18652
rect 35400 18680 35406 18692
rect 35897 18683 35955 18689
rect 35897 18680 35909 18683
rect 35400 18652 35909 18680
rect 35400 18640 35406 18652
rect 35897 18649 35909 18652
rect 35943 18649 35955 18683
rect 35897 18643 35955 18649
rect 23934 18612 23940 18624
rect 22572 18584 23940 18612
rect 23934 18572 23940 18584
rect 23992 18572 23998 18624
rect 24394 18572 24400 18624
rect 24452 18612 24458 18624
rect 24949 18615 25007 18621
rect 24949 18612 24961 18615
rect 24452 18584 24961 18612
rect 24452 18572 24458 18584
rect 24949 18581 24961 18584
rect 24995 18581 25007 18615
rect 25056 18612 25084 18640
rect 27982 18612 27988 18624
rect 25056 18584 27988 18612
rect 24949 18575 25007 18581
rect 27982 18572 27988 18584
rect 28040 18572 28046 18624
rect 28445 18615 28503 18621
rect 28445 18581 28457 18615
rect 28491 18612 28503 18615
rect 28718 18612 28724 18624
rect 28491 18584 28724 18612
rect 28491 18581 28503 18584
rect 28445 18575 28503 18581
rect 28718 18572 28724 18584
rect 28776 18572 28782 18624
rect 29733 18615 29791 18621
rect 29733 18581 29745 18615
rect 29779 18612 29791 18615
rect 29914 18612 29920 18624
rect 29779 18584 29920 18612
rect 29779 18581 29791 18584
rect 29733 18575 29791 18581
rect 29914 18572 29920 18584
rect 29972 18572 29978 18624
rect 30466 18572 30472 18624
rect 30524 18612 30530 18624
rect 30745 18615 30803 18621
rect 30745 18612 30757 18615
rect 30524 18584 30757 18612
rect 30524 18572 30530 18584
rect 30745 18581 30757 18584
rect 30791 18612 30803 18615
rect 31662 18612 31668 18624
rect 30791 18584 31668 18612
rect 30791 18581 30803 18584
rect 30745 18575 30803 18581
rect 31662 18572 31668 18584
rect 31720 18572 31726 18624
rect 31846 18572 31852 18624
rect 31904 18572 31910 18624
rect 32030 18572 32036 18624
rect 32088 18612 32094 18624
rect 32950 18612 32956 18624
rect 32088 18584 32956 18612
rect 32088 18572 32094 18584
rect 32950 18572 32956 18584
rect 33008 18612 33014 18624
rect 33045 18615 33103 18621
rect 33045 18612 33057 18615
rect 33008 18584 33057 18612
rect 33008 18572 33014 18584
rect 33045 18581 33057 18584
rect 33091 18581 33103 18615
rect 33045 18575 33103 18581
rect 33134 18572 33140 18624
rect 33192 18612 33198 18624
rect 33686 18612 33692 18624
rect 33192 18584 33692 18612
rect 33192 18572 33198 18584
rect 33686 18572 33692 18584
rect 33744 18572 33750 18624
rect 33781 18615 33839 18621
rect 33781 18581 33793 18615
rect 33827 18612 33839 18615
rect 34146 18612 34152 18624
rect 33827 18584 34152 18612
rect 33827 18581 33839 18584
rect 33781 18575 33839 18581
rect 34146 18572 34152 18584
rect 34204 18572 34210 18624
rect 34238 18572 34244 18624
rect 34296 18572 34302 18624
rect 34698 18572 34704 18624
rect 34756 18612 34762 18624
rect 37200 18612 37228 18720
rect 34756 18584 37228 18612
rect 34756 18572 34762 18584
rect 38010 18572 38016 18624
rect 38068 18572 38074 18624
rect 38120 18612 38148 18720
rect 38304 18680 38332 18788
rect 38562 18776 38568 18828
rect 38620 18776 38626 18828
rect 38378 18708 38384 18760
rect 38436 18748 38442 18760
rect 40037 18751 40095 18757
rect 40037 18748 40049 18751
rect 38436 18720 40049 18748
rect 38436 18708 38442 18720
rect 40037 18717 40049 18720
rect 40083 18717 40095 18751
rect 40037 18711 40095 18717
rect 48593 18751 48651 18757
rect 48593 18717 48605 18751
rect 48639 18748 48651 18751
rect 48774 18748 48780 18760
rect 48639 18720 48780 18748
rect 48639 18717 48651 18720
rect 48593 18711 48651 18717
rect 48774 18708 48780 18720
rect 48832 18708 48838 18760
rect 49053 18751 49111 18757
rect 49053 18717 49065 18751
rect 49099 18748 49111 18751
rect 49142 18748 49148 18760
rect 49099 18720 49148 18748
rect 49099 18717 49111 18720
rect 49053 18711 49111 18717
rect 49142 18708 49148 18720
rect 49200 18708 49206 18760
rect 39758 18680 39764 18692
rect 38304 18652 39764 18680
rect 39758 18640 39764 18652
rect 39816 18680 39822 18692
rect 40313 18683 40371 18689
rect 40313 18680 40325 18683
rect 39816 18652 40325 18680
rect 39816 18640 39822 18652
rect 40313 18649 40325 18652
rect 40359 18649 40371 18683
rect 41598 18680 41604 18692
rect 41538 18652 41604 18680
rect 40313 18643 40371 18649
rect 41598 18640 41604 18652
rect 41656 18680 41662 18692
rect 42061 18683 42119 18689
rect 42061 18680 42073 18683
rect 41656 18652 42073 18680
rect 41656 18640 41662 18652
rect 42061 18649 42073 18652
rect 42107 18649 42119 18683
rect 42061 18643 42119 18649
rect 38381 18615 38439 18621
rect 38381 18612 38393 18615
rect 38120 18584 38393 18612
rect 38381 18581 38393 18584
rect 38427 18581 38439 18615
rect 38381 18575 38439 18581
rect 38473 18615 38531 18621
rect 38473 18581 38485 18615
rect 38519 18612 38531 18615
rect 40494 18612 40500 18624
rect 38519 18584 40500 18612
rect 38519 18581 38531 18584
rect 38473 18575 38531 18581
rect 40494 18572 40500 18584
rect 40552 18572 40558 18624
rect 40586 18572 40592 18624
rect 40644 18612 40650 18624
rect 41785 18615 41843 18621
rect 41785 18612 41797 18615
rect 40644 18584 41797 18612
rect 40644 18572 40650 18584
rect 41785 18581 41797 18584
rect 41831 18581 41843 18615
rect 41785 18575 41843 18581
rect 48406 18572 48412 18624
rect 48464 18572 48470 18624
rect 1104 18522 49864 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 27950 18522
rect 28002 18470 28014 18522
rect 28066 18470 28078 18522
rect 28130 18470 28142 18522
rect 28194 18470 28206 18522
rect 28258 18470 37950 18522
rect 38002 18470 38014 18522
rect 38066 18470 38078 18522
rect 38130 18470 38142 18522
rect 38194 18470 38206 18522
rect 38258 18470 47950 18522
rect 48002 18470 48014 18522
rect 48066 18470 48078 18522
rect 48130 18470 48142 18522
rect 48194 18470 48206 18522
rect 48258 18470 49864 18522
rect 1104 18448 49864 18470
rect 3421 18411 3479 18417
rect 3421 18377 3433 18411
rect 3467 18408 3479 18411
rect 5074 18408 5080 18420
rect 3467 18380 5080 18408
rect 3467 18377 3479 18380
rect 3421 18371 3479 18377
rect 5074 18368 5080 18380
rect 5132 18368 5138 18420
rect 5626 18368 5632 18420
rect 5684 18408 5690 18420
rect 7837 18411 7895 18417
rect 7837 18408 7849 18411
rect 5684 18380 7849 18408
rect 5684 18368 5690 18380
rect 7837 18377 7849 18380
rect 7883 18377 7895 18411
rect 7837 18371 7895 18377
rect 9674 18368 9680 18420
rect 9732 18408 9738 18420
rect 10781 18411 10839 18417
rect 10781 18408 10793 18411
rect 9732 18380 10793 18408
rect 9732 18368 9738 18380
rect 10781 18377 10793 18380
rect 10827 18377 10839 18411
rect 12710 18408 12716 18420
rect 10781 18371 10839 18377
rect 11716 18380 12716 18408
rect 4982 18340 4988 18352
rect 3620 18312 4988 18340
rect 3620 18281 3648 18312
rect 4982 18300 4988 18312
rect 5040 18300 5046 18352
rect 11606 18340 11612 18352
rect 9968 18312 11612 18340
rect 1765 18275 1823 18281
rect 1765 18241 1777 18275
rect 1811 18272 1823 18275
rect 3605 18275 3663 18281
rect 1811 18244 3556 18272
rect 1811 18241 1823 18244
rect 1765 18235 1823 18241
rect 2774 18164 2780 18216
rect 2832 18164 2838 18216
rect 3528 18136 3556 18244
rect 3605 18241 3617 18275
rect 3651 18241 3663 18275
rect 3605 18235 3663 18241
rect 3694 18232 3700 18284
rect 3752 18272 3758 18284
rect 9968 18281 9996 18312
rect 11606 18300 11612 18312
rect 11664 18300 11670 18352
rect 4433 18275 4491 18281
rect 4433 18272 4445 18275
rect 3752 18244 4445 18272
rect 3752 18232 3758 18244
rect 4433 18241 4445 18244
rect 4479 18241 4491 18275
rect 4433 18235 4491 18241
rect 7745 18275 7803 18281
rect 7745 18241 7757 18275
rect 7791 18241 7803 18275
rect 7745 18235 7803 18241
rect 9953 18275 10011 18281
rect 9953 18241 9965 18275
rect 9999 18241 10011 18275
rect 9953 18235 10011 18241
rect 10873 18275 10931 18281
rect 10873 18241 10885 18275
rect 10919 18272 10931 18275
rect 11422 18272 11428 18284
rect 10919 18244 11428 18272
rect 10919 18241 10931 18244
rect 10873 18235 10931 18241
rect 4154 18164 4160 18216
rect 4212 18164 4218 18216
rect 7760 18204 7788 18235
rect 11422 18232 11428 18244
rect 11480 18232 11486 18284
rect 10965 18207 11023 18213
rect 7760 18176 10548 18204
rect 9769 18139 9827 18145
rect 3528 18108 7972 18136
rect 7944 18068 7972 18108
rect 9769 18105 9781 18139
rect 9815 18136 9827 18139
rect 10226 18136 10232 18148
rect 9815 18108 10232 18136
rect 9815 18105 9827 18108
rect 9769 18099 9827 18105
rect 10226 18096 10232 18108
rect 10284 18096 10290 18148
rect 10410 18096 10416 18148
rect 10468 18096 10474 18148
rect 10318 18068 10324 18080
rect 7944 18040 10324 18068
rect 10318 18028 10324 18040
rect 10376 18028 10382 18080
rect 10520 18068 10548 18176
rect 10965 18173 10977 18207
rect 11011 18204 11023 18207
rect 11054 18204 11060 18216
rect 11011 18176 11060 18204
rect 11011 18173 11023 18176
rect 10965 18167 11023 18173
rect 11054 18164 11060 18176
rect 11112 18164 11118 18216
rect 11716 18213 11744 18380
rect 12710 18368 12716 18380
rect 12768 18408 12774 18420
rect 13538 18408 13544 18420
rect 12768 18380 13544 18408
rect 12768 18368 12774 18380
rect 13538 18368 13544 18380
rect 13596 18368 13602 18420
rect 13630 18368 13636 18420
rect 13688 18408 13694 18420
rect 14277 18411 14335 18417
rect 14277 18408 14289 18411
rect 13688 18380 14289 18408
rect 13688 18368 13694 18380
rect 14277 18377 14289 18380
rect 14323 18377 14335 18411
rect 14277 18371 14335 18377
rect 15010 18368 15016 18420
rect 15068 18368 15074 18420
rect 17957 18411 18015 18417
rect 17957 18408 17969 18411
rect 15212 18380 17969 18408
rect 11882 18300 11888 18352
rect 11940 18340 11946 18352
rect 11940 18312 12466 18340
rect 11940 18300 11946 18312
rect 13446 18300 13452 18352
rect 13504 18340 13510 18352
rect 15212 18340 15240 18380
rect 17957 18377 17969 18380
rect 18003 18377 18015 18411
rect 17957 18371 18015 18377
rect 18417 18411 18475 18417
rect 18417 18377 18429 18411
rect 18463 18408 18475 18411
rect 22097 18411 22155 18417
rect 22097 18408 22109 18411
rect 18463 18380 22109 18408
rect 18463 18377 18475 18380
rect 18417 18371 18475 18377
rect 22097 18377 22109 18380
rect 22143 18377 22155 18411
rect 22097 18371 22155 18377
rect 22465 18411 22523 18417
rect 22465 18377 22477 18411
rect 22511 18408 22523 18411
rect 25774 18408 25780 18420
rect 22511 18380 25780 18408
rect 22511 18377 22523 18380
rect 22465 18371 22523 18377
rect 25774 18368 25780 18380
rect 25832 18368 25838 18420
rect 26237 18411 26295 18417
rect 26237 18377 26249 18411
rect 26283 18408 26295 18411
rect 27246 18408 27252 18420
rect 26283 18380 27252 18408
rect 26283 18377 26295 18380
rect 26237 18371 26295 18377
rect 27246 18368 27252 18380
rect 27304 18368 27310 18420
rect 27525 18411 27583 18417
rect 27525 18377 27537 18411
rect 27571 18408 27583 18411
rect 28994 18408 29000 18420
rect 27571 18380 29000 18408
rect 27571 18377 27583 18380
rect 27525 18371 27583 18377
rect 28994 18368 29000 18380
rect 29052 18368 29058 18420
rect 29178 18368 29184 18420
rect 29236 18408 29242 18420
rect 35897 18411 35955 18417
rect 35897 18408 35909 18411
rect 29236 18380 35909 18408
rect 29236 18368 29242 18380
rect 35897 18377 35909 18380
rect 35943 18377 35955 18411
rect 35897 18371 35955 18377
rect 36170 18368 36176 18420
rect 36228 18408 36234 18420
rect 39206 18408 39212 18420
rect 36228 18380 39212 18408
rect 36228 18368 36234 18380
rect 39206 18368 39212 18380
rect 39264 18368 39270 18420
rect 39758 18368 39764 18420
rect 39816 18368 39822 18420
rect 40034 18368 40040 18420
rect 40092 18408 40098 18420
rect 40865 18411 40923 18417
rect 40865 18408 40877 18411
rect 40092 18380 40877 18408
rect 40092 18368 40098 18380
rect 40865 18377 40877 18380
rect 40911 18377 40923 18411
rect 40865 18371 40923 18377
rect 48774 18368 48780 18420
rect 48832 18368 48838 18420
rect 13504 18312 15240 18340
rect 15304 18312 16436 18340
rect 13504 18300 13510 18312
rect 14182 18232 14188 18284
rect 14240 18272 14246 18284
rect 15304 18272 15332 18312
rect 14240 18244 15332 18272
rect 16301 18275 16359 18281
rect 14240 18232 14246 18244
rect 16301 18241 16313 18275
rect 16347 18241 16359 18275
rect 16408 18272 16436 18312
rect 16666 18300 16672 18352
rect 16724 18300 16730 18352
rect 17313 18343 17371 18349
rect 17313 18309 17325 18343
rect 17359 18340 17371 18343
rect 19886 18340 19892 18352
rect 17359 18312 18276 18340
rect 17359 18309 17371 18312
rect 17313 18303 17371 18309
rect 17497 18275 17555 18281
rect 17497 18272 17509 18275
rect 16408 18244 17509 18272
rect 16301 18235 16359 18241
rect 17497 18241 17509 18244
rect 17543 18241 17555 18275
rect 17497 18235 17555 18241
rect 11701 18207 11759 18213
rect 11701 18173 11713 18207
rect 11747 18173 11759 18207
rect 11701 18167 11759 18173
rect 11977 18207 12035 18213
rect 11977 18173 11989 18207
rect 12023 18204 12035 18207
rect 13354 18204 13360 18216
rect 12023 18176 13360 18204
rect 12023 18173 12035 18176
rect 11977 18167 12035 18173
rect 10594 18096 10600 18148
rect 10652 18136 10658 18148
rect 11716 18136 11744 18167
rect 13354 18164 13360 18176
rect 13412 18164 13418 18216
rect 14369 18207 14427 18213
rect 14369 18173 14381 18207
rect 14415 18173 14427 18207
rect 14369 18167 14427 18173
rect 14553 18207 14611 18213
rect 14553 18173 14565 18207
rect 14599 18204 14611 18207
rect 15286 18204 15292 18216
rect 14599 18176 15292 18204
rect 14599 18173 14611 18176
rect 14553 18167 14611 18173
rect 10652 18108 11744 18136
rect 10652 18096 10658 18108
rect 13262 18096 13268 18148
rect 13320 18136 13326 18148
rect 13909 18139 13967 18145
rect 13909 18136 13921 18139
rect 13320 18108 13921 18136
rect 13320 18096 13326 18108
rect 13909 18105 13921 18108
rect 13955 18105 13967 18139
rect 14384 18136 14412 18167
rect 15286 18164 15292 18176
rect 15344 18164 15350 18216
rect 15473 18207 15531 18213
rect 15473 18173 15485 18207
rect 15519 18204 15531 18207
rect 16206 18204 16212 18216
rect 15519 18176 16212 18204
rect 15519 18173 15531 18176
rect 15473 18167 15531 18173
rect 16206 18164 16212 18176
rect 16264 18164 16270 18216
rect 16316 18204 16344 18235
rect 17770 18204 17776 18216
rect 16316 18176 17776 18204
rect 17770 18164 17776 18176
rect 17828 18164 17834 18216
rect 15197 18139 15255 18145
rect 14384 18108 15148 18136
rect 13909 18099 13967 18105
rect 12158 18068 12164 18080
rect 10520 18040 12164 18068
rect 12158 18028 12164 18040
rect 12216 18028 12222 18080
rect 12342 18028 12348 18080
rect 12400 18068 12406 18080
rect 13449 18071 13507 18077
rect 13449 18068 13461 18071
rect 12400 18040 13461 18068
rect 12400 18028 12406 18040
rect 13449 18037 13461 18040
rect 13495 18037 13507 18071
rect 15120 18068 15148 18108
rect 15197 18105 15209 18139
rect 15243 18136 15255 18139
rect 15378 18136 15384 18148
rect 15243 18108 15384 18136
rect 15243 18105 15255 18108
rect 15197 18099 15255 18105
rect 15378 18096 15384 18108
rect 15436 18096 15442 18148
rect 16114 18096 16120 18148
rect 16172 18096 16178 18148
rect 18248 18136 18276 18312
rect 19628 18312 19892 18340
rect 18325 18275 18383 18281
rect 18325 18241 18337 18275
rect 18371 18272 18383 18275
rect 19518 18272 19524 18284
rect 18371 18244 19524 18272
rect 18371 18241 18383 18244
rect 18325 18235 18383 18241
rect 19518 18232 19524 18244
rect 19576 18232 19582 18284
rect 19628 18281 19656 18312
rect 19886 18300 19892 18312
rect 19944 18300 19950 18352
rect 21542 18340 21548 18352
rect 21114 18312 21548 18340
rect 21542 18300 21548 18312
rect 21600 18300 21606 18352
rect 22830 18300 22836 18352
rect 22888 18340 22894 18352
rect 23293 18343 23351 18349
rect 23293 18340 23305 18343
rect 22888 18312 23305 18340
rect 22888 18300 22894 18312
rect 23293 18309 23305 18312
rect 23339 18309 23351 18343
rect 23293 18303 23351 18309
rect 19613 18275 19671 18281
rect 19613 18241 19625 18275
rect 19659 18241 19671 18275
rect 19613 18235 19671 18241
rect 22557 18275 22615 18281
rect 22557 18241 22569 18275
rect 22603 18272 22615 18275
rect 23308 18272 23336 18303
rect 23474 18300 23480 18352
rect 23532 18340 23538 18352
rect 24029 18343 24087 18349
rect 24029 18340 24041 18343
rect 23532 18312 24041 18340
rect 23532 18300 23538 18312
rect 24029 18309 24041 18312
rect 24075 18309 24087 18343
rect 27614 18340 27620 18352
rect 24029 18303 24087 18309
rect 24964 18312 27620 18340
rect 24670 18272 24676 18284
rect 22603 18244 23244 18272
rect 23308 18244 24676 18272
rect 22603 18241 22615 18244
rect 22557 18235 22615 18241
rect 18601 18207 18659 18213
rect 18601 18173 18613 18207
rect 18647 18204 18659 18207
rect 19889 18207 19947 18213
rect 19889 18204 19901 18207
rect 18647 18176 19901 18204
rect 18647 18173 18659 18176
rect 18601 18167 18659 18173
rect 19889 18173 19901 18176
rect 19935 18204 19947 18207
rect 20898 18204 20904 18216
rect 19935 18176 20904 18204
rect 19935 18173 19947 18176
rect 19889 18167 19947 18173
rect 20898 18164 20904 18176
rect 20956 18164 20962 18216
rect 22738 18164 22744 18216
rect 22796 18164 22802 18216
rect 23216 18204 23244 18244
rect 24670 18232 24676 18244
rect 24728 18232 24734 18284
rect 24964 18204 24992 18312
rect 27614 18300 27620 18312
rect 27672 18300 27678 18352
rect 28813 18343 28871 18349
rect 28813 18309 28825 18343
rect 28859 18340 28871 18343
rect 32122 18340 32128 18352
rect 28859 18312 32128 18340
rect 28859 18309 28871 18312
rect 28813 18303 28871 18309
rect 32122 18300 32128 18312
rect 32180 18300 32186 18352
rect 32582 18300 32588 18352
rect 32640 18340 32646 18352
rect 33134 18340 33140 18352
rect 32640 18312 33140 18340
rect 32640 18300 32646 18312
rect 33134 18300 33140 18312
rect 33192 18300 33198 18352
rect 34422 18300 34428 18352
rect 34480 18300 34486 18352
rect 35710 18300 35716 18352
rect 35768 18340 35774 18352
rect 38378 18340 38384 18352
rect 35768 18312 38384 18340
rect 35768 18300 35774 18312
rect 25038 18232 25044 18284
rect 25096 18232 25102 18284
rect 25130 18232 25136 18284
rect 25188 18232 25194 18284
rect 26329 18275 26387 18281
rect 26329 18241 26341 18275
rect 26375 18272 26387 18275
rect 27430 18272 27436 18284
rect 26375 18244 27436 18272
rect 26375 18241 26387 18244
rect 26329 18235 26387 18241
rect 27430 18232 27436 18244
rect 27488 18232 27494 18284
rect 28721 18275 28779 18281
rect 27724 18244 28396 18272
rect 23216 18176 24992 18204
rect 25314 18164 25320 18216
rect 25372 18164 25378 18216
rect 26234 18204 26240 18216
rect 25424 18176 26240 18204
rect 19610 18136 19616 18148
rect 18248 18108 19616 18136
rect 19610 18096 19616 18108
rect 19668 18096 19674 18148
rect 23750 18096 23756 18148
rect 23808 18136 23814 18148
rect 24673 18139 24731 18145
rect 24673 18136 24685 18139
rect 23808 18108 24685 18136
rect 23808 18096 23814 18108
rect 24673 18105 24685 18108
rect 24719 18105 24731 18139
rect 25424 18136 25452 18176
rect 26234 18164 26240 18176
rect 26292 18164 26298 18216
rect 26418 18164 26424 18216
rect 26476 18164 26482 18216
rect 27246 18164 27252 18216
rect 27304 18204 27310 18216
rect 27617 18207 27675 18213
rect 27617 18204 27629 18207
rect 27304 18176 27629 18204
rect 27304 18164 27310 18176
rect 27617 18173 27629 18176
rect 27663 18173 27675 18207
rect 27617 18167 27675 18173
rect 24673 18099 24731 18105
rect 24964 18108 25452 18136
rect 16574 18068 16580 18080
rect 15120 18040 16580 18068
rect 13449 18031 13507 18037
rect 16574 18028 16580 18040
rect 16632 18028 16638 18080
rect 18966 18028 18972 18080
rect 19024 18028 19030 18080
rect 21361 18071 21419 18077
rect 21361 18037 21373 18071
rect 21407 18068 21419 18071
rect 21910 18068 21916 18080
rect 21407 18040 21916 18068
rect 21407 18037 21419 18040
rect 21361 18031 21419 18037
rect 21910 18028 21916 18040
rect 21968 18028 21974 18080
rect 22278 18028 22284 18080
rect 22336 18068 22342 18080
rect 24964 18068 24992 18108
rect 25498 18096 25504 18148
rect 25556 18136 25562 18148
rect 27724 18136 27752 18244
rect 27801 18207 27859 18213
rect 27801 18173 27813 18207
rect 27847 18173 27859 18207
rect 27801 18167 27859 18173
rect 25556 18108 27752 18136
rect 25556 18096 25562 18108
rect 22336 18040 24992 18068
rect 22336 18028 22342 18040
rect 25038 18028 25044 18080
rect 25096 18068 25102 18080
rect 25869 18071 25927 18077
rect 25869 18068 25881 18071
rect 25096 18040 25881 18068
rect 25096 18028 25102 18040
rect 25869 18037 25881 18040
rect 25915 18037 25927 18071
rect 25869 18031 25927 18037
rect 27154 18028 27160 18080
rect 27212 18028 27218 18080
rect 27430 18028 27436 18080
rect 27488 18068 27494 18080
rect 27816 18068 27844 18167
rect 28368 18145 28396 18244
rect 28721 18241 28733 18275
rect 28767 18272 28779 18275
rect 29730 18272 29736 18284
rect 28767 18244 29736 18272
rect 28767 18241 28779 18244
rect 28721 18235 28779 18241
rect 29730 18232 29736 18244
rect 29788 18232 29794 18284
rect 30469 18275 30527 18281
rect 30469 18241 30481 18275
rect 30515 18272 30527 18275
rect 31297 18275 31355 18281
rect 31297 18272 31309 18275
rect 30515 18244 31309 18272
rect 30515 18241 30527 18244
rect 30469 18235 30527 18241
rect 31297 18241 31309 18244
rect 31343 18241 31355 18275
rect 31297 18235 31355 18241
rect 32674 18232 32680 18284
rect 32732 18272 32738 18284
rect 33042 18272 33048 18284
rect 32732 18244 33048 18272
rect 32732 18232 32738 18244
rect 33042 18232 33048 18244
rect 33100 18232 33106 18284
rect 35986 18232 35992 18284
rect 36044 18272 36050 18284
rect 36265 18275 36323 18281
rect 36265 18272 36277 18275
rect 36044 18244 36277 18272
rect 36044 18232 36050 18244
rect 36265 18241 36277 18244
rect 36311 18241 36323 18275
rect 36265 18235 36323 18241
rect 36357 18275 36415 18281
rect 36357 18241 36369 18275
rect 36403 18272 36415 18275
rect 37366 18272 37372 18284
rect 36403 18244 37372 18272
rect 36403 18241 36415 18244
rect 36357 18235 36415 18241
rect 37366 18232 37372 18244
rect 37424 18232 37430 18284
rect 37458 18232 37464 18284
rect 37516 18272 37522 18284
rect 38028 18281 38056 18312
rect 38378 18300 38384 18312
rect 38436 18300 38442 18352
rect 40129 18343 40187 18349
rect 40129 18340 40141 18343
rect 39514 18312 40141 18340
rect 40129 18309 40141 18312
rect 40175 18340 40187 18343
rect 40218 18340 40224 18352
rect 40175 18312 40224 18340
rect 40175 18309 40187 18312
rect 40129 18303 40187 18309
rect 40218 18300 40224 18312
rect 40276 18300 40282 18352
rect 37645 18275 37703 18281
rect 37645 18272 37657 18275
rect 37516 18244 37657 18272
rect 37516 18232 37522 18244
rect 37645 18241 37657 18244
rect 37691 18241 37703 18275
rect 37645 18235 37703 18241
rect 38013 18275 38071 18281
rect 38013 18241 38025 18275
rect 38059 18241 38071 18275
rect 38013 18235 38071 18241
rect 40773 18275 40831 18281
rect 40773 18241 40785 18275
rect 40819 18272 40831 18275
rect 48406 18272 48412 18284
rect 40819 18244 48412 18272
rect 40819 18241 40831 18244
rect 40773 18235 40831 18241
rect 48406 18232 48412 18244
rect 48464 18232 48470 18284
rect 48593 18275 48651 18281
rect 48593 18241 48605 18275
rect 48639 18272 48651 18275
rect 49050 18272 49056 18284
rect 48639 18244 49056 18272
rect 48639 18241 48651 18244
rect 48593 18235 48651 18241
rect 49050 18232 49056 18244
rect 49108 18232 49114 18284
rect 28810 18164 28816 18216
rect 28868 18204 28874 18216
rect 28905 18207 28963 18213
rect 28905 18204 28917 18207
rect 28868 18176 28917 18204
rect 28868 18164 28874 18176
rect 28905 18173 28917 18176
rect 28951 18173 28963 18207
rect 30561 18207 30619 18213
rect 30561 18204 30573 18207
rect 28905 18167 28963 18173
rect 29748 18176 30573 18204
rect 28353 18139 28411 18145
rect 28353 18105 28365 18139
rect 28399 18105 28411 18139
rect 28353 18099 28411 18105
rect 29362 18096 29368 18148
rect 29420 18136 29426 18148
rect 29748 18145 29776 18176
rect 30561 18173 30573 18176
rect 30607 18173 30619 18207
rect 30561 18167 30619 18173
rect 30745 18207 30803 18213
rect 30745 18173 30757 18207
rect 30791 18204 30803 18207
rect 31386 18204 31392 18216
rect 30791 18176 31392 18204
rect 30791 18173 30803 18176
rect 30745 18167 30803 18173
rect 31386 18164 31392 18176
rect 31444 18164 31450 18216
rect 32769 18207 32827 18213
rect 32769 18204 32781 18207
rect 31726 18176 32781 18204
rect 29733 18139 29791 18145
rect 29733 18136 29745 18139
rect 29420 18108 29745 18136
rect 29420 18096 29426 18108
rect 29733 18105 29745 18108
rect 29779 18105 29791 18139
rect 29733 18099 29791 18105
rect 30098 18096 30104 18148
rect 30156 18096 30162 18148
rect 27488 18040 27844 18068
rect 27488 18028 27494 18040
rect 28534 18028 28540 18080
rect 28592 18068 28598 18080
rect 31726 18068 31754 18176
rect 32769 18173 32781 18176
rect 32815 18173 32827 18207
rect 32769 18167 32827 18173
rect 32953 18207 33011 18213
rect 32953 18173 32965 18207
rect 32999 18204 33011 18207
rect 33410 18204 33416 18216
rect 32999 18176 33416 18204
rect 32999 18173 33011 18176
rect 32953 18167 33011 18173
rect 33410 18164 33416 18176
rect 33468 18164 33474 18216
rect 33597 18207 33655 18213
rect 33597 18173 33609 18207
rect 33643 18173 33655 18207
rect 33597 18167 33655 18173
rect 32490 18096 32496 18148
rect 32548 18136 32554 18148
rect 33612 18136 33640 18167
rect 33870 18164 33876 18216
rect 33928 18164 33934 18216
rect 34330 18164 34336 18216
rect 34388 18204 34394 18216
rect 34388 18176 34928 18204
rect 34388 18164 34394 18176
rect 32548 18108 33640 18136
rect 34900 18136 34928 18176
rect 35342 18164 35348 18216
rect 35400 18164 35406 18216
rect 36541 18207 36599 18213
rect 36541 18173 36553 18207
rect 36587 18204 36599 18207
rect 37826 18204 37832 18216
rect 36587 18176 37832 18204
rect 36587 18173 36599 18176
rect 36541 18167 36599 18173
rect 37826 18164 37832 18176
rect 37884 18164 37890 18216
rect 38286 18164 38292 18216
rect 38344 18204 38350 18216
rect 40957 18207 41015 18213
rect 40957 18204 40969 18207
rect 38344 18176 40969 18204
rect 38344 18164 38350 18176
rect 40957 18173 40969 18176
rect 41003 18173 41015 18207
rect 40957 18167 41015 18173
rect 34900 18108 36400 18136
rect 32548 18096 32554 18108
rect 28592 18040 31754 18068
rect 32309 18071 32367 18077
rect 28592 18028 28598 18040
rect 32309 18037 32321 18071
rect 32355 18068 32367 18071
rect 36262 18068 36268 18080
rect 32355 18040 36268 18068
rect 32355 18037 32367 18040
rect 32309 18031 32367 18037
rect 36262 18028 36268 18040
rect 36320 18028 36326 18080
rect 36372 18068 36400 18108
rect 36630 18096 36636 18148
rect 36688 18136 36694 18148
rect 40405 18139 40463 18145
rect 40405 18136 40417 18139
rect 36688 18108 38148 18136
rect 36688 18096 36694 18108
rect 37274 18068 37280 18080
rect 36372 18040 37280 18068
rect 37274 18028 37280 18040
rect 37332 18028 37338 18080
rect 38120 18068 38148 18108
rect 39316 18108 40417 18136
rect 39316 18068 39344 18108
rect 40405 18105 40417 18108
rect 40451 18105 40463 18139
rect 40405 18099 40463 18105
rect 38120 18040 39344 18068
rect 48314 18028 48320 18080
rect 48372 18068 48378 18080
rect 49237 18071 49295 18077
rect 49237 18068 49249 18071
rect 48372 18040 49249 18068
rect 48372 18028 48378 18040
rect 49237 18037 49249 18040
rect 49283 18037 49295 18071
rect 49237 18031 49295 18037
rect 1104 17978 49864 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 32950 17978
rect 33002 17926 33014 17978
rect 33066 17926 33078 17978
rect 33130 17926 33142 17978
rect 33194 17926 33206 17978
rect 33258 17926 42950 17978
rect 43002 17926 43014 17978
rect 43066 17926 43078 17978
rect 43130 17926 43142 17978
rect 43194 17926 43206 17978
rect 43258 17926 49864 17978
rect 1104 17904 49864 17926
rect 11054 17824 11060 17876
rect 11112 17864 11118 17876
rect 12250 17864 12256 17876
rect 11112 17836 12256 17864
rect 11112 17824 11118 17836
rect 12250 17824 12256 17836
rect 12308 17864 12314 17876
rect 12345 17867 12403 17873
rect 12345 17864 12357 17867
rect 12308 17836 12357 17864
rect 12308 17824 12314 17836
rect 12345 17833 12357 17836
rect 12391 17833 12403 17867
rect 12345 17827 12403 17833
rect 12526 17824 12532 17876
rect 12584 17864 12590 17876
rect 12897 17867 12955 17873
rect 12897 17864 12909 17867
rect 12584 17836 12909 17864
rect 12584 17824 12590 17836
rect 12897 17833 12909 17836
rect 12943 17833 12955 17867
rect 15010 17864 15016 17876
rect 12897 17827 12955 17833
rect 13004 17836 15016 17864
rect 11974 17756 11980 17808
rect 12032 17796 12038 17808
rect 12032 17768 12204 17796
rect 12032 17756 12038 17768
rect 1210 17688 1216 17740
rect 1268 17728 1274 17740
rect 2041 17731 2099 17737
rect 2041 17728 2053 17731
rect 1268 17700 2053 17728
rect 1268 17688 1274 17700
rect 2041 17697 2053 17700
rect 2087 17697 2099 17731
rect 2041 17691 2099 17697
rect 10594 17688 10600 17740
rect 10652 17688 10658 17740
rect 1765 17663 1823 17669
rect 1765 17629 1777 17663
rect 1811 17660 1823 17663
rect 8570 17660 8576 17672
rect 1811 17632 8576 17660
rect 1811 17629 1823 17632
rect 1765 17623 1823 17629
rect 8570 17620 8576 17632
rect 8628 17620 8634 17672
rect 12176 17660 12204 17768
rect 12406 17768 12940 17796
rect 12250 17688 12256 17740
rect 12308 17728 12314 17740
rect 12406 17728 12434 17768
rect 12912 17740 12940 17768
rect 12308 17700 12434 17728
rect 12308 17688 12314 17700
rect 12894 17688 12900 17740
rect 12952 17688 12958 17740
rect 13004 17660 13032 17836
rect 15010 17824 15016 17836
rect 15068 17824 15074 17876
rect 15286 17824 15292 17876
rect 15344 17864 15350 17876
rect 16025 17867 16083 17873
rect 16025 17864 16037 17867
rect 15344 17836 16037 17864
rect 15344 17824 15350 17836
rect 16025 17833 16037 17836
rect 16071 17833 16083 17867
rect 16025 17827 16083 17833
rect 16761 17867 16819 17873
rect 16761 17833 16773 17867
rect 16807 17864 16819 17867
rect 17218 17864 17224 17876
rect 16807 17836 17224 17864
rect 16807 17833 16819 17836
rect 16761 17827 16819 17833
rect 17218 17824 17224 17836
rect 17276 17824 17282 17876
rect 17310 17824 17316 17876
rect 17368 17864 17374 17876
rect 19429 17867 19487 17873
rect 19429 17864 19441 17867
rect 17368 17836 19441 17864
rect 17368 17824 17374 17836
rect 19429 17833 19441 17836
rect 19475 17833 19487 17867
rect 19429 17827 19487 17833
rect 19610 17824 19616 17876
rect 19668 17864 19674 17876
rect 19668 17836 21588 17864
rect 19668 17824 19674 17836
rect 16114 17756 16120 17808
rect 16172 17796 16178 17808
rect 16485 17799 16543 17805
rect 16485 17796 16497 17799
rect 16172 17768 16497 17796
rect 16172 17756 16178 17768
rect 16485 17765 16497 17768
rect 16531 17796 16543 17799
rect 21560 17796 21588 17836
rect 21726 17824 21732 17876
rect 21784 17864 21790 17876
rect 23293 17867 23351 17873
rect 23293 17864 23305 17867
rect 21784 17836 23305 17864
rect 21784 17824 21790 17836
rect 23293 17833 23305 17836
rect 23339 17833 23351 17867
rect 23293 17827 23351 17833
rect 24670 17824 24676 17876
rect 24728 17864 24734 17876
rect 28902 17864 28908 17876
rect 24728 17836 28908 17864
rect 24728 17824 24734 17836
rect 28902 17824 28908 17836
rect 28960 17864 28966 17876
rect 29273 17867 29331 17873
rect 29273 17864 29285 17867
rect 28960 17836 29285 17864
rect 28960 17824 28966 17836
rect 29273 17833 29285 17836
rect 29319 17833 29331 17867
rect 29273 17827 29331 17833
rect 29454 17824 29460 17876
rect 29512 17864 29518 17876
rect 32582 17864 32588 17876
rect 29512 17836 32588 17864
rect 29512 17824 29518 17836
rect 32582 17824 32588 17836
rect 32640 17824 32646 17876
rect 34146 17824 34152 17876
rect 34204 17864 34210 17876
rect 34333 17867 34391 17873
rect 34333 17864 34345 17867
rect 34204 17836 34345 17864
rect 34204 17824 34210 17836
rect 34333 17833 34345 17836
rect 34379 17864 34391 17867
rect 34882 17864 34888 17876
rect 34379 17836 34888 17864
rect 34379 17833 34391 17836
rect 34333 17827 34391 17833
rect 34882 17824 34888 17836
rect 34940 17824 34946 17876
rect 34974 17824 34980 17876
rect 35032 17864 35038 17876
rect 35158 17864 35164 17876
rect 35032 17836 35164 17864
rect 35032 17824 35038 17836
rect 35158 17824 35164 17836
rect 35216 17824 35222 17876
rect 48590 17864 48596 17876
rect 35268 17836 48596 17864
rect 24581 17799 24639 17805
rect 24581 17796 24593 17799
rect 16531 17768 20392 17796
rect 21560 17768 24593 17796
rect 16531 17765 16543 17768
rect 16485 17759 16543 17765
rect 13538 17688 13544 17740
rect 13596 17728 13602 17740
rect 14277 17731 14335 17737
rect 14277 17728 14289 17731
rect 13596 17700 14289 17728
rect 13596 17688 13602 17700
rect 14277 17697 14289 17700
rect 14323 17728 14335 17731
rect 15194 17728 15200 17740
rect 14323 17700 15200 17728
rect 14323 17697 14335 17700
rect 14277 17691 14335 17697
rect 15194 17688 15200 17700
rect 15252 17728 15258 17740
rect 16298 17728 16304 17740
rect 15252 17700 16304 17728
rect 15252 17688 15258 17700
rect 16298 17688 16304 17700
rect 16356 17688 16362 17740
rect 17405 17731 17463 17737
rect 17405 17697 17417 17731
rect 17451 17728 17463 17731
rect 17678 17728 17684 17740
rect 17451 17700 17684 17728
rect 17451 17697 17463 17700
rect 17405 17691 17463 17697
rect 17678 17688 17684 17700
rect 17736 17688 17742 17740
rect 18782 17688 18788 17740
rect 18840 17728 18846 17740
rect 19886 17728 19892 17740
rect 18840 17700 19892 17728
rect 18840 17688 18846 17700
rect 19886 17688 19892 17700
rect 19944 17688 19950 17740
rect 20254 17688 20260 17740
rect 20312 17688 20318 17740
rect 20364 17728 20392 17768
rect 24581 17765 24593 17768
rect 24627 17765 24639 17799
rect 24581 17759 24639 17765
rect 25590 17756 25596 17808
rect 25648 17796 25654 17808
rect 25777 17799 25835 17805
rect 25777 17796 25789 17799
rect 25648 17768 25789 17796
rect 25648 17756 25654 17768
rect 25777 17765 25789 17768
rect 25823 17765 25835 17799
rect 25777 17759 25835 17765
rect 26326 17756 26332 17808
rect 26384 17756 26390 17808
rect 28534 17756 28540 17808
rect 28592 17796 28598 17808
rect 29089 17799 29147 17805
rect 29089 17796 29101 17799
rect 28592 17768 29101 17796
rect 28592 17756 28598 17768
rect 29089 17765 29101 17768
rect 29135 17765 29147 17799
rect 29089 17759 29147 17765
rect 30374 17756 30380 17808
rect 30432 17796 30438 17808
rect 34517 17799 34575 17805
rect 34517 17796 34529 17799
rect 30432 17768 34529 17796
rect 30432 17756 30438 17768
rect 34517 17765 34529 17768
rect 34563 17796 34575 17799
rect 34606 17796 34612 17808
rect 34563 17768 34612 17796
rect 34563 17765 34575 17768
rect 34517 17759 34575 17765
rect 34606 17756 34612 17768
rect 34664 17756 34670 17808
rect 22005 17731 22063 17737
rect 20364 17700 21772 17728
rect 12176 17632 13032 17660
rect 13078 17620 13084 17672
rect 13136 17620 13142 17672
rect 13725 17663 13783 17669
rect 13725 17629 13737 17663
rect 13771 17629 13783 17663
rect 13725 17623 13783 17629
rect 10873 17595 10931 17601
rect 10873 17561 10885 17595
rect 10919 17561 10931 17595
rect 10873 17555 10931 17561
rect 10888 17524 10916 17555
rect 11514 17552 11520 17604
rect 11572 17552 11578 17604
rect 12250 17524 12256 17536
rect 10888 17496 12256 17524
rect 12250 17484 12256 17496
rect 12308 17484 12314 17536
rect 12894 17484 12900 17536
rect 12952 17524 12958 17536
rect 13541 17527 13599 17533
rect 13541 17524 13553 17527
rect 12952 17496 13553 17524
rect 12952 17484 12958 17496
rect 13541 17493 13553 17496
rect 13587 17524 13599 17527
rect 13630 17524 13636 17536
rect 13587 17496 13636 17524
rect 13587 17493 13599 17496
rect 13541 17487 13599 17493
rect 13630 17484 13636 17496
rect 13688 17484 13694 17536
rect 13740 17524 13768 17623
rect 16206 17620 16212 17672
rect 16264 17660 16270 17672
rect 17129 17663 17187 17669
rect 17129 17660 17141 17663
rect 16264 17632 17141 17660
rect 16264 17620 16270 17632
rect 17129 17629 17141 17632
rect 17175 17629 17187 17663
rect 17129 17623 17187 17629
rect 17957 17663 18015 17669
rect 17957 17629 17969 17663
rect 18003 17660 18015 17663
rect 18322 17660 18328 17672
rect 18003 17632 18328 17660
rect 18003 17629 18015 17632
rect 17957 17623 18015 17629
rect 18322 17620 18328 17632
rect 18380 17660 18386 17672
rect 18966 17660 18972 17672
rect 18380 17632 18972 17660
rect 18380 17620 18386 17632
rect 18966 17620 18972 17632
rect 19024 17620 19030 17672
rect 19613 17663 19671 17669
rect 19613 17629 19625 17663
rect 19659 17660 19671 17663
rect 20162 17660 20168 17672
rect 19659 17632 20168 17660
rect 19659 17629 19671 17632
rect 19613 17623 19671 17629
rect 20162 17620 20168 17632
rect 20220 17620 20226 17672
rect 21744 17660 21772 17700
rect 22005 17697 22017 17731
rect 22051 17728 22063 17731
rect 22186 17728 22192 17740
rect 22051 17700 22192 17728
rect 22051 17697 22063 17700
rect 22005 17691 22063 17697
rect 22186 17688 22192 17700
rect 22244 17688 22250 17740
rect 23750 17688 23756 17740
rect 23808 17688 23814 17740
rect 23845 17731 23903 17737
rect 23845 17697 23857 17731
rect 23891 17728 23903 17731
rect 24026 17728 24032 17740
rect 23891 17700 24032 17728
rect 23891 17697 23903 17700
rect 23845 17691 23903 17697
rect 24026 17688 24032 17700
rect 24084 17688 24090 17740
rect 25038 17688 25044 17740
rect 25096 17688 25102 17740
rect 25133 17731 25191 17737
rect 25133 17697 25145 17731
rect 25179 17697 25191 17731
rect 27065 17731 27123 17737
rect 27065 17728 27077 17731
rect 25133 17691 25191 17697
rect 25608 17700 27077 17728
rect 21744 17632 22508 17660
rect 14553 17595 14611 17601
rect 14553 17561 14565 17595
rect 14599 17592 14611 17595
rect 14642 17592 14648 17604
rect 14599 17564 14648 17592
rect 14599 17561 14611 17564
rect 14553 17555 14611 17561
rect 14642 17552 14648 17564
rect 14700 17552 14706 17604
rect 15102 17552 15108 17604
rect 15160 17552 15166 17604
rect 19702 17592 19708 17604
rect 15856 17564 19708 17592
rect 15856 17524 15884 17564
rect 19702 17552 19708 17564
rect 19760 17552 19766 17604
rect 19886 17552 19892 17604
rect 19944 17592 19950 17604
rect 19944 17564 20484 17592
rect 19944 17552 19950 17564
rect 13740 17496 15884 17524
rect 17221 17527 17279 17533
rect 17221 17493 17233 17527
rect 17267 17524 17279 17527
rect 17494 17524 17500 17536
rect 17267 17496 17500 17524
rect 17267 17493 17279 17496
rect 17221 17487 17279 17493
rect 17494 17484 17500 17496
rect 17552 17484 17558 17536
rect 18506 17484 18512 17536
rect 18564 17524 18570 17536
rect 20346 17524 20352 17536
rect 18564 17496 20352 17524
rect 18564 17484 18570 17496
rect 20346 17484 20352 17496
rect 20404 17484 20410 17536
rect 20456 17524 20484 17564
rect 20530 17552 20536 17604
rect 20588 17552 20594 17604
rect 21542 17552 21548 17604
rect 21600 17552 21606 17604
rect 20714 17524 20720 17536
rect 20456 17496 20720 17524
rect 20714 17484 20720 17496
rect 20772 17484 20778 17536
rect 21174 17484 21180 17536
rect 21232 17524 21238 17536
rect 21450 17524 21456 17536
rect 21232 17496 21456 17524
rect 21232 17484 21238 17496
rect 21450 17484 21456 17496
rect 21508 17524 21514 17536
rect 22281 17527 22339 17533
rect 22281 17524 22293 17527
rect 21508 17496 22293 17524
rect 21508 17484 21514 17496
rect 22281 17493 22293 17496
rect 22327 17493 22339 17527
rect 22480 17524 22508 17632
rect 23934 17620 23940 17672
rect 23992 17660 23998 17672
rect 25148 17660 25176 17691
rect 25608 17672 25636 17700
rect 27065 17697 27077 17700
rect 27111 17728 27123 17731
rect 28350 17728 28356 17740
rect 27111 17700 28356 17728
rect 27111 17697 27123 17700
rect 27065 17691 27123 17697
rect 28350 17688 28356 17700
rect 28408 17728 28414 17740
rect 28408 17700 30788 17728
rect 28408 17688 28414 17700
rect 23992 17632 25176 17660
rect 23992 17620 23998 17632
rect 25590 17620 25596 17672
rect 25648 17620 25654 17672
rect 25961 17663 26019 17669
rect 25961 17629 25973 17663
rect 26007 17629 26019 17663
rect 25961 17623 26019 17629
rect 22649 17595 22707 17601
rect 22649 17561 22661 17595
rect 22695 17592 22707 17595
rect 23661 17595 23719 17601
rect 23661 17592 23673 17595
rect 22695 17564 23673 17592
rect 22695 17561 22707 17564
rect 22649 17555 22707 17561
rect 23661 17561 23673 17564
rect 23707 17561 23719 17595
rect 23661 17555 23719 17561
rect 24394 17552 24400 17604
rect 24452 17592 24458 17604
rect 25976 17592 26004 17623
rect 28902 17620 28908 17672
rect 28960 17660 28966 17672
rect 29917 17663 29975 17669
rect 29917 17660 29929 17663
rect 28960 17632 29929 17660
rect 28960 17620 28966 17632
rect 29917 17629 29929 17632
rect 29963 17660 29975 17663
rect 30374 17660 30380 17672
rect 29963 17632 30380 17660
rect 29963 17629 29975 17632
rect 29917 17623 29975 17629
rect 30374 17620 30380 17632
rect 30432 17620 30438 17672
rect 24452 17564 25912 17592
rect 25976 17564 27292 17592
rect 24452 17552 24458 17564
rect 24762 17524 24768 17536
rect 22480 17496 24768 17524
rect 22281 17487 22339 17493
rect 24762 17484 24768 17496
rect 24820 17484 24826 17536
rect 24854 17484 24860 17536
rect 24912 17524 24918 17536
rect 24949 17527 25007 17533
rect 24949 17524 24961 17527
rect 24912 17496 24961 17524
rect 24912 17484 24918 17496
rect 24949 17493 24961 17496
rect 24995 17493 25007 17527
rect 25884 17524 25912 17564
rect 26421 17527 26479 17533
rect 26421 17524 26433 17527
rect 25884 17496 26433 17524
rect 24949 17487 25007 17493
rect 26421 17493 26433 17496
rect 26467 17524 26479 17527
rect 26602 17524 26608 17536
rect 26467 17496 26608 17524
rect 26467 17493 26479 17496
rect 26421 17487 26479 17493
rect 26602 17484 26608 17496
rect 26660 17484 26666 17536
rect 27264 17524 27292 17564
rect 27338 17552 27344 17604
rect 27396 17552 27402 17604
rect 27614 17552 27620 17604
rect 27672 17592 27678 17604
rect 30098 17592 30104 17604
rect 27672 17564 27830 17592
rect 28736 17564 30104 17592
rect 27672 17552 27678 17564
rect 28736 17524 28764 17564
rect 30098 17552 30104 17564
rect 30156 17552 30162 17604
rect 30760 17601 30788 17700
rect 30926 17688 30932 17740
rect 30984 17728 30990 17740
rect 30984 17700 31800 17728
rect 30984 17688 30990 17700
rect 30834 17620 30840 17672
rect 30892 17660 30898 17672
rect 31665 17663 31723 17669
rect 31665 17660 31677 17663
rect 30892 17632 31677 17660
rect 30892 17620 30898 17632
rect 31665 17629 31677 17632
rect 31711 17629 31723 17663
rect 31772 17660 31800 17700
rect 31938 17688 31944 17740
rect 31996 17688 32002 17740
rect 33226 17688 33232 17740
rect 33284 17688 33290 17740
rect 33413 17731 33471 17737
rect 33413 17697 33425 17731
rect 33459 17728 33471 17731
rect 35158 17728 35164 17740
rect 33459 17700 35164 17728
rect 33459 17697 33471 17700
rect 33413 17691 33471 17697
rect 35158 17688 35164 17700
rect 35216 17688 35222 17740
rect 35268 17660 35296 17836
rect 48590 17824 48596 17836
rect 48648 17824 48654 17876
rect 38013 17799 38071 17805
rect 38013 17765 38025 17799
rect 38059 17796 38071 17799
rect 39850 17796 39856 17808
rect 38059 17768 39856 17796
rect 38059 17765 38071 17768
rect 38013 17759 38071 17765
rect 39850 17756 39856 17768
rect 39908 17756 39914 17808
rect 40494 17756 40500 17808
rect 40552 17756 40558 17808
rect 35710 17688 35716 17740
rect 35768 17728 35774 17740
rect 35805 17731 35863 17737
rect 35805 17728 35817 17731
rect 35768 17700 35817 17728
rect 35768 17688 35774 17700
rect 35805 17697 35817 17700
rect 35851 17697 35863 17731
rect 35805 17691 35863 17697
rect 36081 17731 36139 17737
rect 36081 17697 36093 17731
rect 36127 17728 36139 17731
rect 36170 17728 36176 17740
rect 36127 17700 36176 17728
rect 36127 17697 36139 17700
rect 36081 17691 36139 17697
rect 36170 17688 36176 17700
rect 36228 17688 36234 17740
rect 36538 17688 36544 17740
rect 36596 17728 36602 17740
rect 37553 17731 37611 17737
rect 37553 17728 37565 17731
rect 36596 17700 37565 17728
rect 36596 17688 36602 17700
rect 37553 17697 37565 17700
rect 37599 17697 37611 17731
rect 37553 17691 37611 17697
rect 38470 17688 38476 17740
rect 38528 17688 38534 17740
rect 38565 17731 38623 17737
rect 38565 17697 38577 17731
rect 38611 17697 38623 17731
rect 38565 17691 38623 17697
rect 37458 17660 37464 17672
rect 31772 17632 35296 17660
rect 37214 17632 37464 17660
rect 31665 17623 31723 17629
rect 37458 17620 37464 17632
rect 37516 17620 37522 17672
rect 30745 17595 30803 17601
rect 30745 17561 30757 17595
rect 30791 17592 30803 17595
rect 32490 17592 32496 17604
rect 30791 17564 32496 17592
rect 30791 17561 30803 17564
rect 30745 17555 30803 17561
rect 32490 17552 32496 17564
rect 32548 17552 32554 17604
rect 38580 17592 38608 17691
rect 39942 17688 39948 17740
rect 40000 17728 40006 17740
rect 40957 17731 41015 17737
rect 40957 17728 40969 17731
rect 40000 17700 40969 17728
rect 40000 17688 40006 17700
rect 40957 17697 40969 17700
rect 41003 17697 41015 17731
rect 40957 17691 41015 17697
rect 41046 17688 41052 17740
rect 41104 17688 41110 17740
rect 48593 17663 48651 17669
rect 48593 17629 48605 17663
rect 48639 17660 48651 17663
rect 49050 17660 49056 17672
rect 48639 17632 49056 17660
rect 48639 17629 48651 17632
rect 48593 17623 48651 17629
rect 49050 17620 49056 17632
rect 49108 17620 49114 17672
rect 32784 17564 36032 17592
rect 27264 17496 28764 17524
rect 28810 17484 28816 17536
rect 28868 17484 28874 17536
rect 29638 17484 29644 17536
rect 29696 17484 29702 17536
rect 30374 17484 30380 17536
rect 30432 17524 30438 17536
rect 31202 17524 31208 17536
rect 30432 17496 31208 17524
rect 30432 17484 30438 17496
rect 31202 17484 31208 17496
rect 31260 17484 31266 17536
rect 31297 17527 31355 17533
rect 31297 17493 31309 17527
rect 31343 17524 31355 17527
rect 31386 17524 31392 17536
rect 31343 17496 31392 17524
rect 31343 17493 31355 17496
rect 31297 17487 31355 17493
rect 31386 17484 31392 17496
rect 31444 17484 31450 17536
rect 31478 17484 31484 17536
rect 31536 17524 31542 17536
rect 31757 17527 31815 17533
rect 31757 17524 31769 17527
rect 31536 17496 31769 17524
rect 31536 17484 31542 17496
rect 31757 17493 31769 17496
rect 31803 17493 31815 17527
rect 31757 17487 31815 17493
rect 32122 17484 32128 17536
rect 32180 17524 32186 17536
rect 32401 17527 32459 17533
rect 32401 17524 32413 17527
rect 32180 17496 32413 17524
rect 32180 17484 32186 17496
rect 32401 17493 32413 17496
rect 32447 17524 32459 17527
rect 32674 17524 32680 17536
rect 32447 17496 32680 17524
rect 32447 17493 32459 17496
rect 32401 17487 32459 17493
rect 32674 17484 32680 17496
rect 32732 17484 32738 17536
rect 32784 17533 32812 17564
rect 32769 17527 32827 17533
rect 32769 17493 32781 17527
rect 32815 17493 32827 17527
rect 32769 17487 32827 17493
rect 33137 17527 33195 17533
rect 33137 17493 33149 17527
rect 33183 17524 33195 17527
rect 33410 17524 33416 17536
rect 33183 17496 33416 17524
rect 33183 17493 33195 17496
rect 33137 17487 33195 17493
rect 33410 17484 33416 17496
rect 33468 17524 33474 17536
rect 33781 17527 33839 17533
rect 33781 17524 33793 17527
rect 33468 17496 33793 17524
rect 33468 17484 33474 17496
rect 33781 17493 33793 17496
rect 33827 17493 33839 17527
rect 33781 17487 33839 17493
rect 34882 17484 34888 17536
rect 34940 17484 34946 17536
rect 35250 17484 35256 17536
rect 35308 17524 35314 17536
rect 35434 17524 35440 17536
rect 35308 17496 35440 17524
rect 35308 17484 35314 17496
rect 35434 17484 35440 17496
rect 35492 17484 35498 17536
rect 35529 17527 35587 17533
rect 35529 17493 35541 17527
rect 35575 17524 35587 17527
rect 35894 17524 35900 17536
rect 35575 17496 35900 17524
rect 35575 17493 35587 17496
rect 35529 17487 35587 17493
rect 35894 17484 35900 17496
rect 35952 17484 35958 17536
rect 36004 17524 36032 17564
rect 37384 17564 38608 17592
rect 40865 17595 40923 17601
rect 36170 17524 36176 17536
rect 36004 17496 36176 17524
rect 36170 17484 36176 17496
rect 36228 17484 36234 17536
rect 36814 17484 36820 17536
rect 36872 17524 36878 17536
rect 37384 17524 37412 17564
rect 40865 17561 40877 17595
rect 40911 17592 40923 17595
rect 48406 17592 48412 17604
rect 40911 17564 48412 17592
rect 40911 17561 40923 17564
rect 40865 17555 40923 17561
rect 48406 17552 48412 17564
rect 48464 17552 48470 17604
rect 48498 17552 48504 17604
rect 48556 17592 48562 17604
rect 48556 17564 49280 17592
rect 48556 17552 48562 17564
rect 36872 17496 37412 17524
rect 36872 17484 36878 17496
rect 38378 17484 38384 17536
rect 38436 17484 38442 17536
rect 48777 17527 48835 17533
rect 48777 17493 48789 17527
rect 48823 17524 48835 17527
rect 49142 17524 49148 17536
rect 48823 17496 49148 17524
rect 48823 17493 48835 17496
rect 48777 17487 48835 17493
rect 49142 17484 49148 17496
rect 49200 17484 49206 17536
rect 49252 17533 49280 17564
rect 49237 17527 49295 17533
rect 49237 17493 49249 17527
rect 49283 17493 49295 17527
rect 49237 17487 49295 17493
rect 1104 17434 49864 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 27950 17434
rect 28002 17382 28014 17434
rect 28066 17382 28078 17434
rect 28130 17382 28142 17434
rect 28194 17382 28206 17434
rect 28258 17382 37950 17434
rect 38002 17382 38014 17434
rect 38066 17382 38078 17434
rect 38130 17382 38142 17434
rect 38194 17382 38206 17434
rect 38258 17382 47950 17434
rect 48002 17382 48014 17434
rect 48066 17382 48078 17434
rect 48130 17382 48142 17434
rect 48194 17382 48206 17434
rect 48258 17382 49864 17434
rect 1104 17360 49864 17382
rect 10413 17323 10471 17329
rect 10413 17289 10425 17323
rect 10459 17320 10471 17323
rect 13446 17320 13452 17332
rect 10459 17292 13452 17320
rect 10459 17289 10471 17292
rect 10413 17283 10471 17289
rect 13446 17280 13452 17292
rect 13504 17280 13510 17332
rect 13998 17280 14004 17332
rect 14056 17320 14062 17332
rect 14921 17323 14979 17329
rect 14921 17320 14933 17323
rect 14056 17292 14933 17320
rect 14056 17280 14062 17292
rect 14921 17289 14933 17292
rect 14967 17289 14979 17323
rect 14921 17283 14979 17289
rect 15562 17280 15568 17332
rect 15620 17280 15626 17332
rect 16025 17323 16083 17329
rect 16025 17289 16037 17323
rect 16071 17320 16083 17323
rect 16114 17320 16120 17332
rect 16071 17292 16120 17320
rect 16071 17289 16083 17292
rect 16025 17283 16083 17289
rect 16114 17280 16120 17292
rect 16172 17280 16178 17332
rect 16482 17280 16488 17332
rect 16540 17320 16546 17332
rect 18414 17320 18420 17332
rect 16540 17292 18420 17320
rect 16540 17280 16546 17292
rect 18414 17280 18420 17292
rect 18472 17280 18478 17332
rect 20254 17320 20260 17332
rect 19168 17292 20260 17320
rect 10137 17255 10195 17261
rect 10137 17221 10149 17255
rect 10183 17252 10195 17255
rect 11790 17252 11796 17264
rect 10183 17224 11796 17252
rect 10183 17221 10195 17224
rect 10137 17215 10195 17221
rect 11790 17212 11796 17224
rect 11848 17212 11854 17264
rect 12437 17255 12495 17261
rect 12437 17221 12449 17255
rect 12483 17252 12495 17255
rect 13081 17255 13139 17261
rect 13081 17252 13093 17255
rect 12483 17224 13093 17252
rect 12483 17221 12495 17224
rect 12437 17215 12495 17221
rect 13081 17221 13093 17224
rect 13127 17252 13139 17255
rect 13722 17252 13728 17264
rect 13127 17224 13728 17252
rect 13127 17221 13139 17224
rect 13081 17215 13139 17221
rect 13722 17212 13728 17224
rect 13780 17212 13786 17264
rect 14185 17255 14243 17261
rect 14185 17221 14197 17255
rect 14231 17252 14243 17255
rect 14274 17252 14280 17264
rect 14231 17224 14280 17252
rect 14231 17221 14243 17224
rect 14185 17215 14243 17221
rect 14274 17212 14280 17224
rect 14332 17212 14338 17264
rect 15010 17212 15016 17264
rect 15068 17252 15074 17264
rect 17773 17255 17831 17261
rect 15068 17224 17724 17252
rect 15068 17212 15074 17224
rect 1765 17187 1823 17193
rect 1765 17153 1777 17187
rect 1811 17184 1823 17187
rect 8294 17184 8300 17196
rect 1811 17156 8300 17184
rect 1811 17153 1823 17156
rect 1765 17147 1823 17153
rect 8294 17144 8300 17156
rect 8352 17144 8358 17196
rect 9950 17144 9956 17196
rect 10008 17184 10014 17196
rect 10781 17187 10839 17193
rect 10781 17184 10793 17187
rect 10008 17156 10793 17184
rect 10008 17144 10014 17156
rect 10781 17153 10793 17156
rect 10827 17153 10839 17187
rect 12912 17184 13032 17188
rect 14366 17184 14372 17196
rect 10781 17147 10839 17153
rect 11900 17160 14372 17184
rect 11900 17156 12940 17160
rect 13004 17156 14372 17160
rect 1302 17076 1308 17128
rect 1360 17116 1366 17128
rect 2041 17119 2099 17125
rect 2041 17116 2053 17119
rect 1360 17088 2053 17116
rect 1360 17076 1366 17088
rect 2041 17085 2053 17088
rect 2087 17085 2099 17119
rect 10686 17116 10692 17128
rect 2041 17079 2099 17085
rect 9876 17088 10692 17116
rect 9876 16992 9904 17088
rect 10686 17076 10692 17088
rect 10744 17116 10750 17128
rect 10873 17119 10931 17125
rect 10873 17116 10885 17119
rect 10744 17088 10885 17116
rect 10744 17076 10750 17088
rect 10873 17085 10885 17088
rect 10919 17085 10931 17119
rect 10873 17079 10931 17085
rect 10965 17119 11023 17125
rect 10965 17085 10977 17119
rect 11011 17116 11023 17119
rect 11900 17116 11928 17156
rect 11011 17088 11928 17116
rect 11011 17085 11023 17088
rect 10965 17079 11023 17085
rect 11974 17076 11980 17128
rect 12032 17116 12038 17128
rect 13280 17125 13308 17156
rect 14366 17144 14372 17156
rect 14424 17144 14430 17196
rect 15102 17144 15108 17196
rect 15160 17144 15166 17196
rect 15746 17144 15752 17196
rect 15804 17184 15810 17196
rect 15933 17187 15991 17193
rect 15933 17184 15945 17187
rect 15804 17156 15945 17184
rect 15804 17144 15810 17156
rect 15933 17153 15945 17156
rect 15979 17153 15991 17187
rect 15933 17147 15991 17153
rect 16945 17187 17003 17193
rect 16945 17153 16957 17187
rect 16991 17153 17003 17187
rect 17696 17184 17724 17224
rect 17773 17221 17785 17255
rect 17819 17252 17831 17255
rect 18322 17252 18328 17264
rect 17819 17224 18328 17252
rect 17819 17221 17831 17224
rect 17773 17215 17831 17221
rect 18322 17212 18328 17224
rect 18380 17212 18386 17264
rect 18506 17184 18512 17196
rect 17696 17156 18512 17184
rect 16945 17147 17003 17153
rect 13173 17119 13231 17125
rect 13173 17116 13185 17119
rect 12032 17088 13185 17116
rect 12032 17076 12038 17088
rect 13173 17085 13185 17088
rect 13219 17085 13231 17119
rect 13173 17079 13231 17085
rect 13265 17119 13323 17125
rect 13265 17085 13277 17119
rect 13311 17085 13323 17119
rect 13265 17079 13323 17085
rect 13817 17119 13875 17125
rect 13817 17085 13829 17119
rect 13863 17116 13875 17119
rect 15764 17116 15792 17144
rect 13863 17088 15792 17116
rect 13863 17085 13875 17088
rect 13817 17079 13875 17085
rect 16022 17076 16028 17128
rect 16080 17116 16086 17128
rect 16117 17119 16175 17125
rect 16117 17116 16129 17119
rect 16080 17088 16129 17116
rect 16080 17076 16086 17088
rect 16117 17085 16129 17088
rect 16163 17085 16175 17119
rect 16117 17079 16175 17085
rect 11054 17008 11060 17060
rect 11112 17048 11118 17060
rect 14369 17051 14427 17057
rect 14369 17048 14381 17051
rect 11112 17020 14381 17048
rect 11112 17008 11118 17020
rect 14369 17017 14381 17020
rect 14415 17017 14427 17051
rect 16960 17048 16988 17147
rect 18506 17144 18512 17156
rect 18564 17144 18570 17196
rect 19168 17193 19196 17292
rect 20254 17280 20260 17292
rect 20312 17280 20318 17332
rect 20346 17280 20352 17332
rect 20404 17320 20410 17332
rect 20404 17292 20760 17320
rect 20404 17280 20410 17292
rect 19153 17187 19211 17193
rect 19153 17153 19165 17187
rect 19199 17153 19211 17187
rect 19153 17147 19211 17153
rect 20530 17144 20536 17196
rect 20588 17144 20594 17196
rect 17034 17076 17040 17128
rect 17092 17116 17098 17128
rect 17129 17119 17187 17125
rect 17129 17116 17141 17119
rect 17092 17088 17141 17116
rect 17092 17076 17098 17088
rect 17129 17085 17141 17088
rect 17175 17085 17187 17119
rect 17129 17079 17187 17085
rect 18598 17076 18604 17128
rect 18656 17076 18662 17128
rect 19429 17119 19487 17125
rect 19429 17085 19441 17119
rect 19475 17116 19487 17119
rect 20070 17116 20076 17128
rect 19475 17088 20076 17116
rect 19475 17085 19487 17088
rect 19429 17079 19487 17085
rect 20070 17076 20076 17088
rect 20128 17116 20134 17128
rect 20732 17116 20760 17292
rect 20898 17280 20904 17332
rect 20956 17280 20962 17332
rect 20990 17280 20996 17332
rect 21048 17320 21054 17332
rect 22186 17320 22192 17332
rect 21048 17292 22192 17320
rect 21048 17280 21054 17292
rect 22186 17280 22192 17292
rect 22244 17280 22250 17332
rect 23934 17280 23940 17332
rect 23992 17320 23998 17332
rect 24397 17323 24455 17329
rect 24397 17320 24409 17323
rect 23992 17292 24409 17320
rect 23992 17280 23998 17292
rect 24397 17289 24409 17292
rect 24443 17289 24455 17323
rect 24397 17283 24455 17289
rect 24857 17323 24915 17329
rect 24857 17289 24869 17323
rect 24903 17320 24915 17323
rect 24946 17320 24952 17332
rect 24903 17292 24952 17320
rect 24903 17289 24915 17292
rect 24857 17283 24915 17289
rect 24946 17280 24952 17292
rect 25004 17280 25010 17332
rect 25317 17323 25375 17329
rect 25317 17289 25329 17323
rect 25363 17320 25375 17323
rect 27341 17323 27399 17329
rect 27341 17320 27353 17323
rect 25363 17292 27353 17320
rect 25363 17289 25375 17292
rect 25317 17283 25375 17289
rect 27341 17289 27353 17292
rect 27387 17289 27399 17323
rect 27341 17283 27399 17289
rect 27801 17323 27859 17329
rect 27801 17289 27813 17323
rect 27847 17320 27859 17323
rect 28534 17320 28540 17332
rect 27847 17292 28540 17320
rect 27847 17289 27859 17292
rect 27801 17283 27859 17289
rect 24762 17212 24768 17264
rect 24820 17252 24826 17264
rect 24820 17224 25360 17252
rect 24820 17212 24826 17224
rect 22646 17144 22652 17196
rect 22704 17144 22710 17196
rect 24026 17144 24032 17196
rect 24084 17144 24090 17196
rect 25222 17144 25228 17196
rect 25280 17144 25286 17196
rect 25332 17184 25360 17224
rect 25958 17212 25964 17264
rect 26016 17212 26022 17264
rect 27816 17252 27844 17283
rect 28534 17280 28540 17292
rect 28592 17280 28598 17332
rect 28629 17323 28687 17329
rect 28629 17289 28641 17323
rect 28675 17320 28687 17323
rect 32306 17320 32312 17332
rect 28675 17292 32312 17320
rect 28675 17289 28687 17292
rect 28629 17283 28687 17289
rect 32306 17280 32312 17292
rect 32364 17280 32370 17332
rect 32398 17280 32404 17332
rect 32456 17320 32462 17332
rect 33318 17320 33324 17332
rect 32456 17292 33324 17320
rect 32456 17280 32462 17292
rect 33318 17280 33324 17292
rect 33376 17320 33382 17332
rect 34057 17323 34115 17329
rect 34057 17320 34069 17323
rect 33376 17292 34069 17320
rect 33376 17280 33382 17292
rect 34057 17289 34069 17292
rect 34103 17289 34115 17323
rect 34057 17283 34115 17289
rect 34882 17280 34888 17332
rect 34940 17320 34946 17332
rect 37829 17323 37887 17329
rect 37829 17320 37841 17323
rect 34940 17292 37841 17320
rect 34940 17280 34946 17292
rect 37829 17289 37841 17292
rect 37875 17289 37887 17323
rect 40126 17320 40132 17332
rect 37829 17283 37887 17289
rect 39592 17292 40132 17320
rect 27080 17224 27844 17252
rect 27080 17184 27108 17224
rect 27890 17212 27896 17264
rect 27948 17252 27954 17264
rect 28997 17255 29055 17261
rect 28997 17252 29009 17255
rect 27948 17224 29009 17252
rect 27948 17212 27954 17224
rect 28997 17221 29009 17224
rect 29043 17221 29055 17255
rect 28997 17215 29055 17221
rect 29089 17255 29147 17261
rect 29089 17221 29101 17255
rect 29135 17252 29147 17255
rect 29270 17252 29276 17264
rect 29135 17224 29276 17252
rect 29135 17221 29147 17224
rect 29089 17215 29147 17221
rect 29270 17212 29276 17224
rect 29328 17212 29334 17264
rect 30193 17255 30251 17261
rect 30193 17221 30205 17255
rect 30239 17252 30251 17255
rect 32490 17252 32496 17264
rect 30239 17224 31754 17252
rect 30239 17221 30251 17224
rect 30193 17215 30251 17221
rect 25332 17156 27108 17184
rect 27338 17144 27344 17196
rect 27396 17184 27402 17196
rect 27522 17184 27528 17196
rect 27396 17156 27528 17184
rect 27396 17144 27402 17156
rect 27522 17144 27528 17156
rect 27580 17144 27586 17196
rect 27709 17187 27767 17193
rect 27709 17153 27721 17187
rect 27755 17153 27767 17187
rect 27709 17147 27767 17153
rect 22925 17119 22983 17125
rect 20128 17088 20668 17116
rect 20732 17088 22784 17116
rect 20128 17076 20134 17088
rect 20640 17048 20668 17088
rect 22646 17048 22652 17060
rect 16960 17020 19288 17048
rect 20640 17020 22652 17048
rect 14369 17011 14427 17017
rect 9858 16940 9864 16992
rect 9916 16940 9922 16992
rect 11698 16940 11704 16992
rect 11756 16980 11762 16992
rect 11885 16983 11943 16989
rect 11885 16980 11897 16983
rect 11756 16952 11897 16980
rect 11756 16940 11762 16952
rect 11885 16949 11897 16952
rect 11931 16949 11943 16983
rect 11885 16943 11943 16949
rect 12710 16940 12716 16992
rect 12768 16940 12774 16992
rect 13078 16940 13084 16992
rect 13136 16980 13142 16992
rect 17402 16980 17408 16992
rect 13136 16952 17408 16980
rect 13136 16940 13142 16952
rect 17402 16940 17408 16952
rect 17460 16940 17466 16992
rect 17494 16940 17500 16992
rect 17552 16940 17558 16992
rect 19260 16980 19288 17020
rect 22646 17008 22652 17020
rect 22704 17008 22710 17060
rect 19886 16980 19892 16992
rect 19260 16952 19892 16980
rect 19886 16940 19892 16952
rect 19944 16940 19950 16992
rect 21269 16983 21327 16989
rect 21269 16949 21281 16983
rect 21315 16980 21327 16983
rect 21542 16980 21548 16992
rect 21315 16952 21548 16980
rect 21315 16949 21327 16952
rect 21269 16943 21327 16949
rect 21542 16940 21548 16952
rect 21600 16980 21606 16992
rect 21637 16983 21695 16989
rect 21637 16980 21649 16983
rect 21600 16952 21649 16980
rect 21600 16940 21606 16952
rect 21637 16949 21649 16952
rect 21683 16980 21695 16983
rect 22189 16983 22247 16989
rect 22189 16980 22201 16983
rect 21683 16952 22201 16980
rect 21683 16949 21695 16952
rect 21637 16943 21695 16949
rect 22189 16949 22201 16952
rect 22235 16980 22247 16983
rect 22554 16980 22560 16992
rect 22235 16952 22560 16980
rect 22235 16949 22247 16952
rect 22189 16943 22247 16949
rect 22554 16940 22560 16952
rect 22612 16940 22618 16992
rect 22756 16980 22784 17088
rect 22925 17085 22937 17119
rect 22971 17116 22983 17119
rect 23658 17116 23664 17128
rect 22971 17088 23664 17116
rect 22971 17085 22983 17088
rect 22925 17079 22983 17085
rect 23658 17076 23664 17088
rect 23716 17076 23722 17128
rect 25130 17076 25136 17128
rect 25188 17116 25194 17128
rect 25409 17119 25467 17125
rect 25409 17116 25421 17119
rect 25188 17088 25421 17116
rect 25188 17076 25194 17088
rect 25409 17085 25421 17088
rect 25455 17085 25467 17119
rect 25409 17079 25467 17085
rect 27246 17076 27252 17128
rect 27304 17116 27310 17128
rect 27724 17116 27752 17147
rect 28074 17144 28080 17196
rect 28132 17184 28138 17196
rect 29454 17184 29460 17196
rect 28132 17156 29460 17184
rect 28132 17144 28138 17156
rect 29454 17144 29460 17156
rect 29512 17144 29518 17196
rect 29638 17144 29644 17196
rect 29696 17184 29702 17196
rect 30285 17187 30343 17193
rect 30285 17184 30297 17187
rect 29696 17156 30297 17184
rect 29696 17144 29702 17156
rect 30285 17153 30297 17156
rect 30331 17153 30343 17187
rect 30926 17184 30932 17196
rect 30285 17147 30343 17153
rect 30484 17156 30932 17184
rect 27304 17088 27752 17116
rect 27985 17119 28043 17125
rect 27304 17076 27310 17088
rect 27985 17085 27997 17119
rect 28031 17116 28043 17119
rect 28534 17116 28540 17128
rect 28031 17088 28540 17116
rect 28031 17085 28043 17088
rect 27985 17079 28043 17085
rect 28534 17076 28540 17088
rect 28592 17076 28598 17128
rect 29178 17076 29184 17128
rect 29236 17076 29242 17128
rect 29822 17076 29828 17128
rect 29880 17116 29886 17128
rect 30374 17116 30380 17128
rect 29880 17088 30380 17116
rect 29880 17076 29886 17088
rect 30374 17076 30380 17088
rect 30432 17076 30438 17128
rect 25866 17008 25872 17060
rect 25924 17048 25930 17060
rect 28810 17048 28816 17060
rect 25924 17020 28816 17048
rect 25924 17008 25930 17020
rect 28810 17008 28816 17020
rect 28868 17008 28874 17060
rect 30484 17048 30512 17156
rect 30926 17144 30932 17156
rect 30984 17144 30990 17196
rect 31202 17144 31208 17196
rect 31260 17184 31266 17196
rect 31389 17187 31447 17193
rect 31389 17184 31401 17187
rect 31260 17156 31401 17184
rect 31260 17144 31266 17156
rect 31389 17153 31401 17156
rect 31435 17153 31447 17187
rect 31726 17184 31754 17224
rect 32324 17224 32496 17252
rect 32122 17184 32128 17196
rect 31726 17156 32128 17184
rect 31389 17147 31447 17153
rect 32122 17144 32128 17156
rect 32180 17144 32186 17196
rect 32324 17193 32352 17224
rect 32490 17212 32496 17224
rect 32548 17212 32554 17264
rect 32582 17212 32588 17264
rect 32640 17212 32646 17264
rect 34146 17252 34152 17264
rect 33810 17224 34152 17252
rect 34146 17212 34152 17224
rect 34204 17212 34210 17264
rect 34606 17212 34612 17264
rect 34664 17212 34670 17264
rect 35342 17212 35348 17264
rect 35400 17252 35406 17264
rect 35618 17252 35624 17264
rect 35400 17224 35624 17252
rect 35400 17212 35406 17224
rect 35618 17212 35624 17224
rect 35676 17212 35682 17264
rect 36446 17212 36452 17264
rect 36504 17212 36510 17264
rect 37734 17212 37740 17264
rect 37792 17252 37798 17264
rect 39592 17252 39620 17292
rect 40126 17280 40132 17292
rect 40184 17280 40190 17332
rect 40218 17280 40224 17332
rect 40276 17320 40282 17332
rect 48314 17320 48320 17332
rect 40276 17292 48320 17320
rect 40276 17280 40282 17292
rect 48314 17280 48320 17292
rect 48372 17280 48378 17332
rect 48406 17280 48412 17332
rect 48464 17280 48470 17332
rect 48590 17280 48596 17332
rect 48648 17320 48654 17332
rect 49237 17323 49295 17329
rect 49237 17320 49249 17323
rect 48648 17292 49249 17320
rect 48648 17280 48654 17292
rect 49237 17289 49249 17292
rect 49283 17289 49295 17323
rect 49237 17283 49295 17289
rect 41049 17255 41107 17261
rect 41049 17252 41061 17255
rect 37792 17224 39620 17252
rect 40434 17224 41061 17252
rect 37792 17212 37798 17224
rect 41049 17221 41061 17224
rect 41095 17252 41107 17255
rect 41138 17252 41144 17264
rect 41095 17224 41144 17252
rect 41095 17221 41107 17224
rect 41049 17215 41107 17221
rect 41138 17212 41144 17224
rect 41196 17212 41202 17264
rect 32309 17187 32367 17193
rect 32309 17153 32321 17187
rect 32355 17153 32367 17187
rect 36078 17184 36084 17196
rect 32309 17147 32367 17153
rect 33888 17156 36084 17184
rect 33888 17128 33916 17156
rect 36078 17144 36084 17156
rect 36136 17184 36142 17196
rect 36136 17156 36216 17184
rect 36136 17144 36142 17156
rect 30558 17076 30564 17128
rect 30616 17116 30622 17128
rect 31481 17119 31539 17125
rect 31481 17116 31493 17119
rect 30616 17088 31493 17116
rect 30616 17076 30622 17088
rect 31481 17085 31493 17088
rect 31527 17085 31539 17119
rect 31481 17079 31539 17085
rect 31573 17119 31631 17125
rect 31573 17085 31585 17119
rect 31619 17085 31631 17119
rect 31573 17079 31631 17085
rect 29748 17020 30512 17048
rect 25958 16980 25964 16992
rect 22756 16952 25964 16980
rect 25958 16940 25964 16952
rect 26016 16940 26022 16992
rect 26326 16940 26332 16992
rect 26384 16980 26390 16992
rect 27798 16980 27804 16992
rect 26384 16952 27804 16980
rect 26384 16940 26390 16952
rect 27798 16940 27804 16952
rect 27856 16980 27862 16992
rect 29748 16980 29776 17020
rect 30742 17008 30748 17060
rect 30800 17048 30806 17060
rect 31588 17048 31616 17079
rect 31662 17076 31668 17128
rect 31720 17116 31726 17128
rect 33870 17116 33876 17128
rect 31720 17088 33876 17116
rect 31720 17076 31726 17088
rect 33870 17076 33876 17088
rect 33928 17076 33934 17128
rect 34882 17076 34888 17128
rect 34940 17116 34946 17128
rect 35345 17119 35403 17125
rect 35345 17116 35357 17119
rect 34940 17088 35357 17116
rect 34940 17076 34946 17088
rect 35345 17085 35357 17088
rect 35391 17085 35403 17119
rect 36188 17116 36216 17156
rect 36262 17144 36268 17196
rect 36320 17184 36326 17196
rect 36357 17187 36415 17193
rect 36357 17184 36369 17187
rect 36320 17156 36369 17184
rect 36320 17144 36326 17156
rect 36357 17153 36369 17156
rect 36403 17153 36415 17187
rect 36357 17147 36415 17153
rect 37921 17187 37979 17193
rect 37921 17153 37933 17187
rect 37967 17184 37979 17187
rect 48593 17187 48651 17193
rect 37967 17156 38516 17184
rect 37967 17153 37979 17156
rect 37921 17147 37979 17153
rect 38488 17128 38516 17156
rect 48593 17153 48605 17187
rect 48639 17184 48651 17187
rect 48774 17184 48780 17196
rect 48639 17156 48780 17184
rect 48639 17153 48651 17156
rect 48593 17147 48651 17153
rect 48774 17144 48780 17156
rect 48832 17144 48838 17196
rect 49145 17187 49203 17193
rect 49145 17153 49157 17187
rect 49191 17184 49203 17187
rect 49234 17184 49240 17196
rect 49191 17156 49240 17184
rect 49191 17153 49203 17156
rect 49145 17147 49203 17153
rect 49234 17144 49240 17156
rect 49292 17144 49298 17196
rect 36538 17116 36544 17128
rect 36188 17088 36544 17116
rect 35345 17079 35403 17085
rect 36538 17076 36544 17088
rect 36596 17076 36602 17128
rect 36630 17076 36636 17128
rect 36688 17076 36694 17128
rect 38105 17119 38163 17125
rect 38105 17085 38117 17119
rect 38151 17116 38163 17119
rect 38286 17116 38292 17128
rect 38151 17088 38292 17116
rect 38151 17085 38163 17088
rect 38105 17079 38163 17085
rect 38286 17076 38292 17088
rect 38344 17076 38350 17128
rect 38470 17076 38476 17128
rect 38528 17076 38534 17128
rect 38933 17119 38991 17125
rect 38933 17085 38945 17119
rect 38979 17085 38991 17119
rect 38933 17079 38991 17085
rect 39209 17119 39267 17125
rect 39209 17085 39221 17119
rect 39255 17116 39267 17119
rect 40586 17116 40592 17128
rect 39255 17088 40592 17116
rect 39255 17085 39267 17088
rect 39209 17079 39267 17085
rect 30800 17020 31616 17048
rect 35989 17051 36047 17057
rect 30800 17008 30806 17020
rect 35989 17017 36001 17051
rect 36035 17048 36047 17051
rect 36035 17020 37136 17048
rect 36035 17017 36047 17020
rect 35989 17011 36047 17017
rect 27856 16952 29776 16980
rect 29825 16983 29883 16989
rect 27856 16940 27862 16952
rect 29825 16949 29837 16983
rect 29871 16980 29883 16983
rect 30926 16980 30932 16992
rect 29871 16952 30932 16980
rect 29871 16949 29883 16952
rect 29825 16943 29883 16949
rect 30926 16940 30932 16952
rect 30984 16940 30990 16992
rect 31021 16983 31079 16989
rect 31021 16949 31033 16983
rect 31067 16980 31079 16983
rect 33962 16980 33968 16992
rect 31067 16952 33968 16980
rect 31067 16949 31079 16952
rect 31021 16943 31079 16949
rect 33962 16940 33968 16952
rect 34020 16940 34026 16992
rect 36538 16940 36544 16992
rect 36596 16980 36602 16992
rect 37001 16983 37059 16989
rect 37001 16980 37013 16983
rect 36596 16952 37013 16980
rect 36596 16940 36602 16952
rect 37001 16949 37013 16952
rect 37047 16949 37059 16983
rect 37108 16980 37136 17020
rect 37182 17008 37188 17060
rect 37240 17048 37246 17060
rect 37461 17051 37519 17057
rect 37461 17048 37473 17051
rect 37240 17020 37473 17048
rect 37240 17008 37246 17020
rect 37461 17017 37473 17020
rect 37507 17017 37519 17051
rect 37461 17011 37519 17017
rect 37734 17008 37740 17060
rect 37792 17048 37798 17060
rect 38948 17048 38976 17079
rect 40586 17076 40592 17088
rect 40644 17076 40650 17128
rect 37792 17020 38976 17048
rect 37792 17008 37798 17020
rect 40402 17008 40408 17060
rect 40460 17048 40466 17060
rect 41322 17048 41328 17060
rect 40460 17020 41328 17048
rect 40460 17008 40466 17020
rect 41322 17008 41328 17020
rect 41380 17008 41386 17060
rect 37642 16980 37648 16992
rect 37108 16952 37648 16980
rect 37001 16943 37059 16949
rect 37642 16940 37648 16952
rect 37700 16940 37706 16992
rect 38286 16940 38292 16992
rect 38344 16980 38350 16992
rect 40681 16983 40739 16989
rect 40681 16980 40693 16983
rect 38344 16952 40693 16980
rect 38344 16940 38350 16952
rect 40681 16949 40693 16952
rect 40727 16980 40739 16983
rect 41046 16980 41052 16992
rect 40727 16952 41052 16980
rect 40727 16949 40739 16952
rect 40681 16943 40739 16949
rect 41046 16940 41052 16952
rect 41104 16940 41110 16992
rect 1104 16890 49864 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 32950 16890
rect 33002 16838 33014 16890
rect 33066 16838 33078 16890
rect 33130 16838 33142 16890
rect 33194 16838 33206 16890
rect 33258 16838 42950 16890
rect 43002 16838 43014 16890
rect 43066 16838 43078 16890
rect 43130 16838 43142 16890
rect 43194 16838 43206 16890
rect 43258 16838 49864 16890
rect 1104 16816 49864 16838
rect 5350 16736 5356 16788
rect 5408 16776 5414 16788
rect 11974 16776 11980 16788
rect 5408 16748 11980 16776
rect 5408 16736 5414 16748
rect 11974 16736 11980 16748
rect 12032 16736 12038 16788
rect 14185 16779 14243 16785
rect 14185 16745 14197 16779
rect 14231 16776 14243 16779
rect 14274 16776 14280 16788
rect 14231 16748 14280 16776
rect 14231 16745 14243 16748
rect 14185 16739 14243 16745
rect 14274 16736 14280 16748
rect 14332 16736 14338 16788
rect 14734 16736 14740 16788
rect 14792 16776 14798 16788
rect 17218 16776 17224 16788
rect 14792 16748 17224 16776
rect 14792 16736 14798 16748
rect 17218 16736 17224 16748
rect 17276 16736 17282 16788
rect 17392 16779 17450 16785
rect 17392 16745 17404 16779
rect 17438 16776 17450 16779
rect 18782 16776 18788 16788
rect 17438 16748 18788 16776
rect 17438 16745 17450 16748
rect 17392 16739 17450 16745
rect 18782 16736 18788 16748
rect 18840 16776 18846 16788
rect 20990 16776 20996 16788
rect 18840 16748 20996 16776
rect 18840 16736 18846 16748
rect 20990 16736 20996 16748
rect 21048 16736 21054 16788
rect 23934 16776 23940 16788
rect 21100 16748 23940 16776
rect 15194 16708 15200 16720
rect 15028 16680 15200 16708
rect 4522 16600 4528 16652
rect 4580 16640 4586 16652
rect 5442 16640 5448 16652
rect 4580 16612 5448 16640
rect 4580 16600 4586 16612
rect 5442 16600 5448 16612
rect 5500 16640 5506 16652
rect 8205 16643 8263 16649
rect 8205 16640 8217 16643
rect 5500 16612 8217 16640
rect 5500 16600 5506 16612
rect 8205 16609 8217 16612
rect 8251 16609 8263 16643
rect 8205 16603 8263 16609
rect 8389 16643 8447 16649
rect 8389 16609 8401 16643
rect 8435 16640 8447 16643
rect 8478 16640 8484 16652
rect 8435 16612 8484 16640
rect 8435 16609 8447 16612
rect 8389 16603 8447 16609
rect 8478 16600 8484 16612
rect 8536 16600 8542 16652
rect 8570 16600 8576 16652
rect 8628 16640 8634 16652
rect 10597 16643 10655 16649
rect 10597 16640 10609 16643
rect 8628 16612 10609 16640
rect 8628 16600 8634 16612
rect 10597 16609 10609 16612
rect 10643 16609 10655 16643
rect 10597 16603 10655 16609
rect 10870 16600 10876 16652
rect 10928 16640 10934 16652
rect 11609 16643 11667 16649
rect 11609 16640 11621 16643
rect 10928 16612 11621 16640
rect 10928 16600 10934 16612
rect 11609 16609 11621 16612
rect 11655 16609 11667 16643
rect 11609 16603 11667 16609
rect 13633 16643 13691 16649
rect 13633 16609 13645 16643
rect 13679 16640 13691 16643
rect 13906 16640 13912 16652
rect 13679 16612 13912 16640
rect 13679 16609 13691 16612
rect 13633 16603 13691 16609
rect 13906 16600 13912 16612
rect 13964 16640 13970 16652
rect 15028 16649 15056 16680
rect 15194 16668 15200 16680
rect 15252 16668 15258 16720
rect 16942 16708 16948 16720
rect 16132 16680 16948 16708
rect 16132 16652 16160 16680
rect 16942 16668 16948 16680
rect 17000 16668 17006 16720
rect 18414 16668 18420 16720
rect 18472 16708 18478 16720
rect 21100 16708 21128 16748
rect 23934 16736 23940 16748
rect 23992 16736 23998 16788
rect 27338 16776 27344 16788
rect 24044 16748 27344 16776
rect 18472 16680 21128 16708
rect 18472 16668 18478 16680
rect 22738 16668 22744 16720
rect 22796 16668 22802 16720
rect 24044 16708 24072 16748
rect 27338 16736 27344 16748
rect 27396 16736 27402 16788
rect 28626 16736 28632 16788
rect 28684 16736 28690 16788
rect 34517 16779 34575 16785
rect 28736 16748 34468 16776
rect 25498 16708 25504 16720
rect 23952 16680 24072 16708
rect 24228 16680 25504 16708
rect 15013 16643 15071 16649
rect 13964 16612 14964 16640
rect 13964 16600 13970 16612
rect 1765 16575 1823 16581
rect 1765 16541 1777 16575
rect 1811 16572 1823 16575
rect 11054 16572 11060 16584
rect 1811 16544 11060 16572
rect 1811 16541 1823 16544
rect 1765 16535 1823 16541
rect 11054 16532 11060 16544
rect 11112 16532 11118 16584
rect 11514 16532 11520 16584
rect 11572 16572 11578 16584
rect 11698 16572 11704 16584
rect 11572 16544 11704 16572
rect 11572 16532 11578 16544
rect 11698 16532 11704 16544
rect 11756 16532 11762 16584
rect 12529 16575 12587 16581
rect 12529 16541 12541 16575
rect 12575 16572 12587 16575
rect 13354 16572 13360 16584
rect 12575 16544 13360 16572
rect 12575 16541 12587 16544
rect 12529 16535 12587 16541
rect 13354 16532 13360 16544
rect 13412 16532 13418 16584
rect 14182 16532 14188 16584
rect 14240 16572 14246 16584
rect 14829 16575 14887 16581
rect 14829 16572 14841 16575
rect 14240 16544 14841 16572
rect 14240 16532 14246 16544
rect 14829 16541 14841 16544
rect 14875 16541 14887 16575
rect 14829 16535 14887 16541
rect 14936 16572 14964 16612
rect 15013 16609 15025 16643
rect 15059 16609 15071 16643
rect 15013 16603 15071 16609
rect 15120 16612 16068 16640
rect 15120 16572 15148 16612
rect 14936 16544 15148 16572
rect 16040 16572 16068 16612
rect 16114 16600 16120 16652
rect 16172 16600 16178 16652
rect 16209 16643 16267 16649
rect 16209 16609 16221 16643
rect 16255 16609 16267 16643
rect 16209 16603 16267 16609
rect 16224 16572 16252 16603
rect 16298 16600 16304 16652
rect 16356 16640 16362 16652
rect 17129 16643 17187 16649
rect 17129 16640 17141 16643
rect 16356 16612 17141 16640
rect 16356 16600 16362 16612
rect 17129 16609 17141 16612
rect 17175 16640 17187 16643
rect 18598 16640 18604 16652
rect 17175 16612 18604 16640
rect 17175 16609 17187 16612
rect 17129 16603 17187 16609
rect 18598 16600 18604 16612
rect 18656 16600 18662 16652
rect 20346 16600 20352 16652
rect 20404 16640 20410 16652
rect 20404 16612 20944 16640
rect 20404 16600 20410 16612
rect 16040 16544 16252 16572
rect 1302 16464 1308 16516
rect 1360 16504 1366 16516
rect 2501 16507 2559 16513
rect 2501 16504 2513 16507
rect 1360 16476 2513 16504
rect 1360 16464 1366 16476
rect 2501 16473 2513 16476
rect 2547 16473 2559 16507
rect 9582 16504 9588 16516
rect 2501 16467 2559 16473
rect 7760 16476 9588 16504
rect 7760 16445 7788 16476
rect 9582 16464 9588 16476
rect 9640 16464 9646 16516
rect 10045 16507 10103 16513
rect 10045 16473 10057 16507
rect 10091 16504 10103 16507
rect 10413 16507 10471 16513
rect 10413 16504 10425 16507
rect 10091 16476 10425 16504
rect 10091 16473 10103 16476
rect 10045 16467 10103 16473
rect 10413 16473 10425 16476
rect 10459 16504 10471 16507
rect 10502 16504 10508 16516
rect 10459 16476 10508 16504
rect 10459 16473 10471 16476
rect 10413 16467 10471 16473
rect 10502 16464 10508 16476
rect 10560 16464 10566 16516
rect 11425 16507 11483 16513
rect 11425 16473 11437 16507
rect 11471 16504 11483 16507
rect 12618 16504 12624 16516
rect 11471 16476 12624 16504
rect 11471 16473 11483 16476
rect 11425 16467 11483 16473
rect 12618 16464 12624 16476
rect 12676 16464 12682 16516
rect 14200 16504 14228 16532
rect 14936 16504 14964 16544
rect 16482 16532 16488 16584
rect 16540 16572 16546 16584
rect 16669 16575 16727 16581
rect 16669 16572 16681 16575
rect 16540 16544 16681 16572
rect 16540 16532 16546 16544
rect 16669 16541 16681 16544
rect 16715 16541 16727 16575
rect 20257 16575 20315 16581
rect 18538 16544 20208 16572
rect 16669 16535 16727 16541
rect 15010 16504 15016 16516
rect 13372 16476 14228 16504
rect 14292 16476 14872 16504
rect 14936 16476 15016 16504
rect 7745 16439 7803 16445
rect 7745 16405 7757 16439
rect 7791 16405 7803 16439
rect 7745 16399 7803 16405
rect 7834 16396 7840 16448
rect 7892 16436 7898 16448
rect 8113 16439 8171 16445
rect 8113 16436 8125 16439
rect 7892 16408 8125 16436
rect 7892 16396 7898 16408
rect 8113 16405 8125 16408
rect 8159 16405 8171 16439
rect 8113 16399 8171 16405
rect 11057 16439 11115 16445
rect 11057 16405 11069 16439
rect 11103 16436 11115 16439
rect 11330 16436 11336 16448
rect 11103 16408 11336 16436
rect 11103 16405 11115 16408
rect 11057 16399 11115 16405
rect 11330 16396 11336 16408
rect 11388 16396 11394 16448
rect 11514 16396 11520 16448
rect 11572 16396 11578 16448
rect 12345 16439 12403 16445
rect 12345 16405 12357 16439
rect 12391 16436 12403 16439
rect 12526 16436 12532 16448
rect 12391 16408 12532 16436
rect 12391 16405 12403 16408
rect 12345 16399 12403 16405
rect 12526 16396 12532 16408
rect 12584 16396 12590 16448
rect 12986 16396 12992 16448
rect 13044 16396 13050 16448
rect 13372 16445 13400 16476
rect 13357 16439 13415 16445
rect 13357 16405 13369 16439
rect 13403 16405 13415 16439
rect 13357 16399 13415 16405
rect 13449 16439 13507 16445
rect 13449 16405 13461 16439
rect 13495 16436 13507 16439
rect 13630 16436 13636 16448
rect 13495 16408 13636 16436
rect 13495 16405 13507 16408
rect 13449 16399 13507 16405
rect 13630 16396 13636 16408
rect 13688 16436 13694 16448
rect 14292 16436 14320 16476
rect 14844 16448 14872 16476
rect 15010 16464 15016 16476
rect 15068 16464 15074 16516
rect 15470 16464 15476 16516
rect 15528 16504 15534 16516
rect 16025 16507 16083 16513
rect 16025 16504 16037 16507
rect 15528 16476 16037 16504
rect 15528 16464 15534 16476
rect 16025 16473 16037 16476
rect 16071 16504 16083 16507
rect 16500 16504 16528 16532
rect 16071 16476 16528 16504
rect 18708 16476 20116 16504
rect 16071 16473 16083 16476
rect 16025 16467 16083 16473
rect 13688 16408 14320 16436
rect 14461 16439 14519 16445
rect 13688 16396 13694 16408
rect 14461 16405 14473 16439
rect 14507 16436 14519 16439
rect 14734 16436 14740 16448
rect 14507 16408 14740 16436
rect 14507 16405 14519 16408
rect 14461 16399 14519 16405
rect 14734 16396 14740 16408
rect 14792 16396 14798 16448
rect 14826 16396 14832 16448
rect 14884 16436 14890 16448
rect 14921 16439 14979 16445
rect 14921 16436 14933 16439
rect 14884 16408 14933 16436
rect 14884 16396 14890 16408
rect 14921 16405 14933 16408
rect 14967 16405 14979 16439
rect 14921 16399 14979 16405
rect 15654 16396 15660 16448
rect 15712 16396 15718 16448
rect 17218 16396 17224 16448
rect 17276 16436 17282 16448
rect 18708 16436 18736 16476
rect 17276 16408 18736 16436
rect 17276 16396 17282 16408
rect 18874 16396 18880 16448
rect 18932 16396 18938 16448
rect 18966 16396 18972 16448
rect 19024 16436 19030 16448
rect 20088 16445 20116 16476
rect 19429 16439 19487 16445
rect 19429 16436 19441 16439
rect 19024 16408 19441 16436
rect 19024 16396 19030 16408
rect 19429 16405 19441 16408
rect 19475 16405 19487 16439
rect 19429 16399 19487 16405
rect 20073 16439 20131 16445
rect 20073 16405 20085 16439
rect 20119 16405 20131 16439
rect 20180 16436 20208 16544
rect 20257 16541 20269 16575
rect 20303 16541 20315 16575
rect 20916 16572 20944 16612
rect 21266 16600 21272 16652
rect 21324 16600 21330 16652
rect 23952 16649 23980 16680
rect 23753 16643 23811 16649
rect 23753 16609 23765 16643
rect 23799 16640 23811 16643
rect 23937 16643 23995 16649
rect 23799 16612 23888 16640
rect 23799 16609 23811 16612
rect 23753 16603 23811 16609
rect 20993 16575 21051 16581
rect 20993 16572 21005 16575
rect 20916 16544 21005 16572
rect 20257 16535 20315 16541
rect 20993 16541 21005 16544
rect 21039 16541 21051 16575
rect 23860 16572 23888 16612
rect 23937 16609 23949 16643
rect 23983 16609 23995 16643
rect 24228 16640 24256 16680
rect 25498 16668 25504 16680
rect 25556 16668 25562 16720
rect 27614 16668 27620 16720
rect 27672 16708 27678 16720
rect 28169 16711 28227 16717
rect 28169 16708 28181 16711
rect 27672 16680 28181 16708
rect 27672 16668 27678 16680
rect 28169 16677 28181 16680
rect 28215 16677 28227 16711
rect 28169 16671 28227 16677
rect 23937 16603 23995 16609
rect 24044 16612 24256 16640
rect 24044 16572 24072 16612
rect 24578 16600 24584 16652
rect 24636 16640 24642 16652
rect 25590 16640 25596 16652
rect 24636 16612 25596 16640
rect 24636 16600 24642 16612
rect 25590 16600 25596 16612
rect 25648 16600 25654 16652
rect 25866 16600 25872 16652
rect 25924 16600 25930 16652
rect 26602 16600 26608 16652
rect 26660 16640 26666 16652
rect 27985 16643 28043 16649
rect 27985 16640 27997 16643
rect 26660 16612 27997 16640
rect 26660 16600 26666 16612
rect 27985 16609 27997 16612
rect 28031 16609 28043 16643
rect 27985 16603 28043 16609
rect 23860 16544 24072 16572
rect 20993 16535 21051 16541
rect 20272 16504 20300 16535
rect 26970 16532 26976 16584
rect 27028 16572 27034 16584
rect 27522 16572 27528 16584
rect 27028 16544 27528 16572
rect 27028 16532 27034 16544
rect 27522 16532 27528 16544
rect 27580 16572 27586 16584
rect 27617 16575 27675 16581
rect 27617 16572 27629 16575
rect 27580 16544 27629 16572
rect 27580 16532 27586 16544
rect 27617 16541 27629 16544
rect 27663 16541 27675 16575
rect 28000 16572 28028 16603
rect 28736 16572 28764 16748
rect 34146 16708 34152 16720
rect 29288 16680 31432 16708
rect 29288 16652 29316 16680
rect 29270 16600 29276 16652
rect 29328 16600 29334 16652
rect 29454 16600 29460 16652
rect 29512 16640 29518 16652
rect 31404 16649 31432 16680
rect 33612 16680 34152 16708
rect 30285 16643 30343 16649
rect 30285 16640 30297 16643
rect 29512 16612 30297 16640
rect 29512 16600 29518 16612
rect 30285 16609 30297 16612
rect 30331 16609 30343 16643
rect 30285 16603 30343 16609
rect 31389 16643 31447 16649
rect 31389 16609 31401 16643
rect 31435 16609 31447 16643
rect 31389 16603 31447 16609
rect 31573 16643 31631 16649
rect 31573 16609 31585 16643
rect 31619 16640 31631 16643
rect 31662 16640 31668 16652
rect 31619 16612 31668 16640
rect 31619 16609 31631 16612
rect 31573 16603 31631 16609
rect 31662 16600 31668 16612
rect 31720 16600 31726 16652
rect 32217 16643 32275 16649
rect 32217 16609 32229 16643
rect 32263 16640 32275 16643
rect 32490 16640 32496 16652
rect 32263 16612 32496 16640
rect 32263 16609 32275 16612
rect 32217 16603 32275 16609
rect 32490 16600 32496 16612
rect 32548 16600 32554 16652
rect 28000 16544 28764 16572
rect 27617 16535 27675 16541
rect 28810 16532 28816 16584
rect 28868 16572 28874 16584
rect 28868 16544 32076 16572
rect 33612 16558 33640 16680
rect 34146 16668 34152 16680
rect 34204 16708 34210 16720
rect 34241 16711 34299 16717
rect 34241 16708 34253 16711
rect 34204 16680 34253 16708
rect 34204 16668 34210 16680
rect 34241 16677 34253 16680
rect 34287 16677 34299 16711
rect 34440 16708 34468 16748
rect 34517 16745 34529 16779
rect 34563 16776 34575 16779
rect 34606 16776 34612 16788
rect 34563 16748 34612 16776
rect 34563 16745 34575 16748
rect 34517 16739 34575 16745
rect 34606 16736 34612 16748
rect 34664 16736 34670 16788
rect 48498 16776 48504 16788
rect 34716 16748 48504 16776
rect 34716 16708 34744 16748
rect 48498 16736 48504 16748
rect 48556 16736 48562 16788
rect 48774 16736 48780 16788
rect 48832 16736 48838 16788
rect 34440 16680 34744 16708
rect 34808 16680 35848 16708
rect 34241 16671 34299 16677
rect 34422 16600 34428 16652
rect 34480 16640 34486 16652
rect 34808 16640 34836 16680
rect 34480 16612 34836 16640
rect 34480 16600 34486 16612
rect 35710 16600 35716 16652
rect 35768 16600 35774 16652
rect 35820 16640 35848 16680
rect 36262 16668 36268 16720
rect 36320 16668 36326 16720
rect 36372 16680 36952 16708
rect 36372 16640 36400 16680
rect 35820 16612 36400 16640
rect 36722 16600 36728 16652
rect 36780 16600 36786 16652
rect 36817 16643 36875 16649
rect 36817 16609 36829 16643
rect 36863 16609 36875 16643
rect 36924 16640 36952 16680
rect 36998 16668 37004 16720
rect 37056 16708 37062 16720
rect 37369 16711 37427 16717
rect 37369 16708 37381 16711
rect 37056 16680 37381 16708
rect 37056 16668 37062 16680
rect 37369 16677 37381 16680
rect 37415 16708 37427 16711
rect 37458 16708 37464 16720
rect 37415 16680 37464 16708
rect 37415 16677 37427 16680
rect 37369 16671 37427 16677
rect 37458 16668 37464 16680
rect 37516 16668 37522 16720
rect 41230 16708 41236 16720
rect 40420 16680 41236 16708
rect 40218 16640 40224 16652
rect 36924 16612 40224 16640
rect 36817 16603 36875 16609
rect 34514 16572 34520 16584
rect 28868 16532 28874 16544
rect 22554 16504 22560 16516
rect 20272 16476 21220 16504
rect 22494 16476 22560 16504
rect 20530 16436 20536 16448
rect 20180 16408 20536 16436
rect 20073 16399 20131 16405
rect 20530 16396 20536 16408
rect 20588 16436 20594 16448
rect 20625 16439 20683 16445
rect 20625 16436 20637 16439
rect 20588 16408 20637 16436
rect 20588 16396 20594 16408
rect 20625 16405 20637 16408
rect 20671 16436 20683 16439
rect 20806 16436 20812 16448
rect 20671 16408 20812 16436
rect 20671 16405 20683 16408
rect 20625 16399 20683 16405
rect 20806 16396 20812 16408
rect 20864 16396 20870 16448
rect 21192 16436 21220 16476
rect 22554 16464 22560 16476
rect 22612 16504 22618 16516
rect 22830 16504 22836 16516
rect 22612 16476 22836 16504
rect 22612 16464 22618 16476
rect 22830 16464 22836 16476
rect 22888 16464 22894 16516
rect 24670 16464 24676 16516
rect 24728 16464 24734 16516
rect 25958 16504 25964 16516
rect 24780 16476 25964 16504
rect 22646 16436 22652 16448
rect 21192 16408 22652 16436
rect 22646 16396 22652 16408
rect 22704 16396 22710 16448
rect 23290 16396 23296 16448
rect 23348 16396 23354 16448
rect 23382 16396 23388 16448
rect 23440 16436 23446 16448
rect 23661 16439 23719 16445
rect 23661 16436 23673 16439
rect 23440 16408 23673 16436
rect 23440 16396 23446 16408
rect 23661 16405 23673 16408
rect 23707 16405 23719 16439
rect 23661 16399 23719 16405
rect 24026 16396 24032 16448
rect 24084 16436 24090 16448
rect 24581 16439 24639 16445
rect 24581 16436 24593 16439
rect 24084 16408 24593 16436
rect 24084 16396 24090 16408
rect 24581 16405 24593 16408
rect 24627 16436 24639 16439
rect 24780 16436 24808 16476
rect 25958 16464 25964 16476
rect 26016 16464 26022 16516
rect 27246 16464 27252 16516
rect 27304 16504 27310 16516
rect 28258 16504 28264 16516
rect 27304 16476 28264 16504
rect 27304 16464 27310 16476
rect 28258 16464 28264 16476
rect 28316 16504 28322 16516
rect 28353 16507 28411 16513
rect 28353 16504 28365 16507
rect 28316 16476 28365 16504
rect 28316 16464 28322 16476
rect 28353 16473 28365 16476
rect 28399 16473 28411 16507
rect 28353 16467 28411 16473
rect 28994 16464 29000 16516
rect 29052 16504 29058 16516
rect 30101 16507 30159 16513
rect 30101 16504 30113 16507
rect 29052 16476 30113 16504
rect 29052 16464 29058 16476
rect 30101 16473 30113 16476
rect 30147 16473 30159 16507
rect 30101 16467 30159 16473
rect 30190 16464 30196 16516
rect 30248 16464 30254 16516
rect 31846 16504 31852 16516
rect 30944 16476 31852 16504
rect 24627 16408 24808 16436
rect 24627 16405 24639 16408
rect 24581 16399 24639 16405
rect 25038 16396 25044 16448
rect 25096 16436 25102 16448
rect 28074 16436 28080 16448
rect 25096 16408 28080 16436
rect 25096 16396 25102 16408
rect 28074 16396 28080 16408
rect 28132 16396 28138 16448
rect 29733 16439 29791 16445
rect 29733 16405 29745 16439
rect 29779 16436 29791 16439
rect 30834 16436 30840 16448
rect 29779 16408 30840 16436
rect 29779 16405 29791 16408
rect 29733 16399 29791 16405
rect 30834 16396 30840 16408
rect 30892 16396 30898 16448
rect 30944 16445 30972 16476
rect 31846 16464 31852 16476
rect 31904 16464 31910 16516
rect 30929 16439 30987 16445
rect 30929 16405 30941 16439
rect 30975 16405 30987 16439
rect 30929 16399 30987 16405
rect 31294 16396 31300 16448
rect 31352 16396 31358 16448
rect 32048 16436 32076 16544
rect 33888 16544 34520 16572
rect 32122 16464 32128 16516
rect 32180 16504 32186 16516
rect 32398 16504 32404 16516
rect 32180 16476 32404 16504
rect 32180 16464 32186 16476
rect 32398 16464 32404 16476
rect 32456 16504 32462 16516
rect 32493 16507 32551 16513
rect 32493 16504 32505 16507
rect 32456 16476 32505 16504
rect 32456 16464 32462 16476
rect 32493 16473 32505 16476
rect 32539 16473 32551 16507
rect 32493 16467 32551 16473
rect 33888 16436 33916 16544
rect 34514 16532 34520 16544
rect 34572 16532 34578 16584
rect 34606 16532 34612 16584
rect 34664 16572 34670 16584
rect 34885 16575 34943 16581
rect 34885 16572 34897 16575
rect 34664 16544 34897 16572
rect 34664 16532 34670 16544
rect 34885 16541 34897 16544
rect 34931 16541 34943 16575
rect 34885 16535 34943 16541
rect 35894 16532 35900 16584
rect 35952 16572 35958 16584
rect 36832 16572 36860 16603
rect 40218 16600 40224 16612
rect 40276 16600 40282 16652
rect 36906 16572 36912 16584
rect 35952 16544 36492 16572
rect 36832 16544 36912 16572
rect 35952 16532 35958 16544
rect 36464 16516 36492 16544
rect 36906 16532 36912 16544
rect 36964 16532 36970 16584
rect 37458 16532 37464 16584
rect 37516 16572 37522 16584
rect 37734 16572 37740 16584
rect 37516 16544 37740 16572
rect 37516 16532 37522 16544
rect 37734 16532 37740 16544
rect 37792 16532 37798 16584
rect 40420 16581 40448 16680
rect 41230 16668 41236 16680
rect 41288 16668 41294 16720
rect 41322 16668 41328 16720
rect 41380 16708 41386 16720
rect 41509 16711 41567 16717
rect 41509 16708 41521 16711
rect 41380 16680 41521 16708
rect 41380 16668 41386 16680
rect 41509 16677 41521 16680
rect 41555 16708 41567 16711
rect 46106 16708 46112 16720
rect 41555 16680 46112 16708
rect 41555 16677 41567 16680
rect 41509 16671 41567 16677
rect 46106 16668 46112 16680
rect 46164 16668 46170 16720
rect 40494 16600 40500 16652
rect 40552 16600 40558 16652
rect 40586 16600 40592 16652
rect 40644 16600 40650 16652
rect 41049 16643 41107 16649
rect 41049 16609 41061 16643
rect 41095 16640 41107 16643
rect 41138 16640 41144 16652
rect 41095 16612 41144 16640
rect 41095 16609 41107 16612
rect 41049 16603 41107 16609
rect 41138 16600 41144 16612
rect 41196 16640 41202 16652
rect 41196 16612 41414 16640
rect 41196 16600 41202 16612
rect 40405 16575 40463 16581
rect 40405 16541 40417 16575
rect 40451 16541 40463 16575
rect 40405 16535 40463 16541
rect 41386 16572 41414 16612
rect 41598 16572 41604 16584
rect 41386 16544 41604 16572
rect 34054 16504 34060 16516
rect 33980 16476 34060 16504
rect 33980 16445 34008 16476
rect 34054 16464 34060 16476
rect 34112 16504 34118 16516
rect 36354 16504 36360 16516
rect 34112 16476 36360 16504
rect 34112 16464 34118 16476
rect 36354 16464 36360 16476
rect 36412 16464 36418 16516
rect 36446 16464 36452 16516
rect 36504 16504 36510 16516
rect 36998 16504 37004 16516
rect 36504 16476 37004 16504
rect 36504 16464 36510 16476
rect 36998 16464 37004 16476
rect 37056 16464 37062 16516
rect 38013 16507 38071 16513
rect 38013 16473 38025 16507
rect 38059 16504 38071 16507
rect 38286 16504 38292 16516
rect 38059 16476 38292 16504
rect 38059 16473 38071 16476
rect 38013 16467 38071 16473
rect 38286 16464 38292 16476
rect 38344 16464 38350 16516
rect 39758 16504 39764 16516
rect 39238 16476 39764 16504
rect 39758 16464 39764 16476
rect 39816 16464 39822 16516
rect 41386 16448 41414 16544
rect 41598 16532 41604 16544
rect 41656 16532 41662 16584
rect 48593 16575 48651 16581
rect 48593 16541 48605 16575
rect 48639 16572 48651 16575
rect 49053 16575 49111 16581
rect 49053 16572 49065 16575
rect 48639 16544 49065 16572
rect 48639 16541 48651 16544
rect 48593 16535 48651 16541
rect 49053 16541 49065 16544
rect 49099 16572 49111 16575
rect 49142 16572 49148 16584
rect 49099 16544 49148 16572
rect 49099 16541 49111 16544
rect 49053 16535 49111 16541
rect 49142 16532 49148 16544
rect 49200 16532 49206 16584
rect 32048 16408 33916 16436
rect 33965 16439 34023 16445
rect 33965 16405 33977 16439
rect 34011 16405 34023 16439
rect 33965 16399 34023 16405
rect 34514 16396 34520 16448
rect 34572 16436 34578 16448
rect 34974 16436 34980 16448
rect 34572 16408 34980 16436
rect 34572 16396 34578 16408
rect 34974 16396 34980 16408
rect 35032 16396 35038 16448
rect 36538 16396 36544 16448
rect 36596 16436 36602 16448
rect 36633 16439 36691 16445
rect 36633 16436 36645 16439
rect 36596 16408 36645 16436
rect 36596 16396 36602 16408
rect 36633 16405 36645 16408
rect 36679 16405 36691 16439
rect 36633 16399 36691 16405
rect 36722 16396 36728 16448
rect 36780 16436 36786 16448
rect 38378 16436 38384 16448
rect 36780 16408 38384 16436
rect 36780 16396 36786 16408
rect 38378 16396 38384 16408
rect 38436 16396 38442 16448
rect 38654 16396 38660 16448
rect 38712 16436 38718 16448
rect 39485 16439 39543 16445
rect 39485 16436 39497 16439
rect 38712 16408 39497 16436
rect 38712 16396 38718 16408
rect 39485 16405 39497 16408
rect 39531 16405 39543 16439
rect 39485 16399 39543 16405
rect 40034 16396 40040 16448
rect 40092 16396 40098 16448
rect 41322 16396 41328 16448
rect 41380 16408 41414 16448
rect 41380 16396 41386 16408
rect 48774 16396 48780 16448
rect 48832 16436 48838 16448
rect 49237 16439 49295 16445
rect 49237 16436 49249 16439
rect 48832 16408 49249 16436
rect 48832 16396 48838 16408
rect 49237 16405 49249 16408
rect 49283 16405 49295 16439
rect 49237 16399 49295 16405
rect 1104 16346 49864 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 27950 16346
rect 28002 16294 28014 16346
rect 28066 16294 28078 16346
rect 28130 16294 28142 16346
rect 28194 16294 28206 16346
rect 28258 16294 37950 16346
rect 38002 16294 38014 16346
rect 38066 16294 38078 16346
rect 38130 16294 38142 16346
rect 38194 16294 38206 16346
rect 38258 16294 47950 16346
rect 48002 16294 48014 16346
rect 48066 16294 48078 16346
rect 48130 16294 48142 16346
rect 48194 16294 48206 16346
rect 48258 16294 49864 16346
rect 1104 16272 49864 16294
rect 8297 16235 8355 16241
rect 8297 16201 8309 16235
rect 8343 16232 8355 16235
rect 8386 16232 8392 16244
rect 8343 16204 8392 16232
rect 8343 16201 8355 16204
rect 8297 16195 8355 16201
rect 8386 16192 8392 16204
rect 8444 16192 8450 16244
rect 9306 16192 9312 16244
rect 9364 16192 9370 16244
rect 10318 16192 10324 16244
rect 10376 16232 10382 16244
rect 11057 16235 11115 16241
rect 11057 16232 11069 16235
rect 10376 16204 11069 16232
rect 10376 16192 10382 16204
rect 11057 16201 11069 16204
rect 11103 16201 11115 16235
rect 11057 16195 11115 16201
rect 11514 16192 11520 16244
rect 11572 16232 11578 16244
rect 11977 16235 12035 16241
rect 11977 16232 11989 16235
rect 11572 16204 11989 16232
rect 11572 16192 11578 16204
rect 11977 16201 11989 16204
rect 12023 16201 12035 16235
rect 11977 16195 12035 16201
rect 12437 16235 12495 16241
rect 12437 16201 12449 16235
rect 12483 16232 12495 16235
rect 13173 16235 13231 16241
rect 13173 16232 13185 16235
rect 12483 16204 13185 16232
rect 12483 16201 12495 16204
rect 12437 16195 12495 16201
rect 13173 16201 13185 16204
rect 13219 16201 13231 16235
rect 13173 16195 13231 16201
rect 13541 16235 13599 16241
rect 13541 16201 13553 16235
rect 13587 16232 13599 16235
rect 14369 16235 14427 16241
rect 14369 16232 14381 16235
rect 13587 16204 14381 16232
rect 13587 16201 13599 16204
rect 13541 16195 13599 16201
rect 14369 16201 14381 16204
rect 14415 16201 14427 16235
rect 14369 16195 14427 16201
rect 14550 16192 14556 16244
rect 14608 16232 14614 16244
rect 14737 16235 14795 16241
rect 14737 16232 14749 16235
rect 14608 16204 14749 16232
rect 14608 16192 14614 16204
rect 14737 16201 14749 16204
rect 14783 16201 14795 16235
rect 14737 16195 14795 16201
rect 11146 16164 11152 16176
rect 1780 16136 11152 16164
rect 1780 16105 1808 16136
rect 11146 16124 11152 16136
rect 11204 16124 11210 16176
rect 11238 16124 11244 16176
rect 11296 16164 11302 16176
rect 11296 16136 12572 16164
rect 11296 16124 11302 16136
rect 1765 16099 1823 16105
rect 1765 16065 1777 16099
rect 1811 16065 1823 16099
rect 1765 16059 1823 16065
rect 9217 16099 9275 16105
rect 9217 16065 9229 16099
rect 9263 16096 9275 16099
rect 10778 16096 10784 16108
rect 9263 16068 10784 16096
rect 9263 16065 9275 16068
rect 9217 16059 9275 16065
rect 10778 16056 10784 16068
rect 10836 16056 10842 16108
rect 10870 16056 10876 16108
rect 10928 16096 10934 16108
rect 10965 16099 11023 16105
rect 10965 16096 10977 16099
rect 10928 16068 10977 16096
rect 10928 16056 10934 16068
rect 10965 16065 10977 16068
rect 11011 16065 11023 16099
rect 10965 16059 11023 16065
rect 12345 16099 12403 16105
rect 12345 16065 12357 16099
rect 12391 16096 12403 16099
rect 12434 16096 12440 16108
rect 12391 16068 12440 16096
rect 12391 16065 12403 16068
rect 12345 16059 12403 16065
rect 12434 16056 12440 16068
rect 12492 16056 12498 16108
rect 1302 15988 1308 16040
rect 1360 16028 1366 16040
rect 2041 16031 2099 16037
rect 2041 16028 2053 16031
rect 1360 16000 2053 16028
rect 1360 15988 1366 16000
rect 2041 15997 2053 16000
rect 2087 15997 2099 16031
rect 2041 15991 2099 15997
rect 4154 15988 4160 16040
rect 4212 16028 4218 16040
rect 8389 16031 8447 16037
rect 8389 16028 8401 16031
rect 4212 16000 8401 16028
rect 4212 15988 4218 16000
rect 8389 15997 8401 16000
rect 8435 15997 8447 16031
rect 8389 15991 8447 15997
rect 8478 15988 8484 16040
rect 8536 15988 8542 16040
rect 10413 16031 10471 16037
rect 10413 15997 10425 16031
rect 10459 16028 10471 16031
rect 10888 16028 10916 16056
rect 12544 16040 12572 16136
rect 12986 16124 12992 16176
rect 13044 16164 13050 16176
rect 13633 16167 13691 16173
rect 13633 16164 13645 16167
rect 13044 16136 13645 16164
rect 13044 16124 13050 16136
rect 13633 16133 13645 16136
rect 13679 16133 13691 16167
rect 13633 16127 13691 16133
rect 14752 16096 14780 16195
rect 14918 16192 14924 16244
rect 14976 16232 14982 16244
rect 17405 16235 17463 16241
rect 17405 16232 17417 16235
rect 14976 16204 17417 16232
rect 14976 16192 14982 16204
rect 17405 16201 17417 16204
rect 17451 16201 17463 16235
rect 17405 16195 17463 16201
rect 18322 16192 18328 16244
rect 18380 16232 18386 16244
rect 18785 16235 18843 16241
rect 18785 16232 18797 16235
rect 18380 16204 18797 16232
rect 18380 16192 18386 16204
rect 18785 16201 18797 16204
rect 18831 16201 18843 16235
rect 18785 16195 18843 16201
rect 19058 16192 19064 16244
rect 19116 16232 19122 16244
rect 22002 16232 22008 16244
rect 19116 16204 22008 16232
rect 19116 16192 19122 16204
rect 22002 16192 22008 16204
rect 22060 16192 22066 16244
rect 23109 16235 23167 16241
rect 23109 16201 23121 16235
rect 23155 16232 23167 16235
rect 24854 16232 24860 16244
rect 23155 16204 24860 16232
rect 23155 16201 23167 16204
rect 23109 16195 23167 16201
rect 24854 16192 24860 16204
rect 24912 16192 24918 16244
rect 26329 16235 26387 16241
rect 26329 16232 26341 16235
rect 24964 16204 26341 16232
rect 15930 16124 15936 16176
rect 15988 16124 15994 16176
rect 18874 16164 18880 16176
rect 18524 16136 18880 16164
rect 17034 16096 17040 16108
rect 14752 16068 17040 16096
rect 15948 16040 15976 16068
rect 17034 16056 17040 16068
rect 17092 16056 17098 16108
rect 17773 16099 17831 16105
rect 17773 16065 17785 16099
rect 17819 16096 17831 16099
rect 18414 16096 18420 16108
rect 17819 16068 18420 16096
rect 17819 16065 17831 16068
rect 17773 16059 17831 16065
rect 18414 16056 18420 16068
rect 18472 16056 18478 16108
rect 10459 16000 10916 16028
rect 10459 15997 10471 16000
rect 10413 15991 10471 15997
rect 11054 15988 11060 16040
rect 11112 16028 11118 16040
rect 11112 16000 12480 16028
rect 11112 15988 11118 16000
rect 8496 15960 8524 15988
rect 11974 15960 11980 15972
rect 8496 15932 11980 15960
rect 11974 15920 11980 15932
rect 12032 15920 12038 15972
rect 12452 15960 12480 16000
rect 12526 15988 12532 16040
rect 12584 15988 12590 16040
rect 12894 15988 12900 16040
rect 12952 16028 12958 16040
rect 13725 16031 13783 16037
rect 13725 16028 13737 16031
rect 12952 16000 13737 16028
rect 12952 15988 12958 16000
rect 13725 15997 13737 16000
rect 13771 16028 13783 16031
rect 14550 16028 14556 16040
rect 13771 16000 14556 16028
rect 13771 15997 13783 16000
rect 13725 15991 13783 15997
rect 14550 15988 14556 16000
rect 14608 15988 14614 16040
rect 14826 15988 14832 16040
rect 14884 15988 14890 16040
rect 15010 15988 15016 16040
rect 15068 15988 15074 16040
rect 15194 15988 15200 16040
rect 15252 16028 15258 16040
rect 15749 16031 15807 16037
rect 15749 16028 15761 16031
rect 15252 16000 15761 16028
rect 15252 15988 15258 16000
rect 15749 15997 15761 16000
rect 15795 15997 15807 16031
rect 15749 15991 15807 15997
rect 13630 15960 13636 15972
rect 12452 15932 13636 15960
rect 13630 15920 13636 15932
rect 13688 15920 13694 15972
rect 15764 15960 15792 15991
rect 15838 15988 15844 16040
rect 15896 15988 15902 16040
rect 15930 15988 15936 16040
rect 15988 15988 15994 16040
rect 17865 16031 17923 16037
rect 17865 15997 17877 16031
rect 17911 15997 17923 16031
rect 17865 15991 17923 15997
rect 18049 16031 18107 16037
rect 18049 15997 18061 16031
rect 18095 16028 18107 16031
rect 18524 16028 18552 16136
rect 18874 16124 18880 16136
rect 18932 16164 18938 16176
rect 19429 16167 19487 16173
rect 19429 16164 19441 16167
rect 18932 16136 19441 16164
rect 18932 16124 18938 16136
rect 19429 16133 19441 16136
rect 19475 16133 19487 16167
rect 20806 16164 20812 16176
rect 20654 16136 20812 16164
rect 19429 16127 19487 16133
rect 20806 16124 20812 16136
rect 20864 16164 20870 16176
rect 21361 16167 21419 16173
rect 21361 16164 21373 16167
rect 20864 16136 21373 16164
rect 20864 16124 20870 16136
rect 21361 16133 21373 16136
rect 21407 16164 21419 16167
rect 21542 16164 21548 16176
rect 21407 16136 21548 16164
rect 21407 16133 21419 16136
rect 21361 16127 21419 16133
rect 21542 16124 21548 16136
rect 21600 16124 21606 16176
rect 23477 16167 23535 16173
rect 23477 16133 23489 16167
rect 23523 16164 23535 16167
rect 23566 16164 23572 16176
rect 23523 16136 23572 16164
rect 23523 16133 23535 16136
rect 23477 16127 23535 16133
rect 23566 16124 23572 16136
rect 23624 16124 23630 16176
rect 23658 16124 23664 16176
rect 23716 16164 23722 16176
rect 24964 16164 24992 16204
rect 26329 16201 26341 16204
rect 26375 16232 26387 16235
rect 26418 16232 26424 16244
rect 26375 16204 26424 16232
rect 26375 16201 26387 16204
rect 26329 16195 26387 16201
rect 26418 16192 26424 16204
rect 26476 16192 26482 16244
rect 26878 16192 26884 16244
rect 26936 16232 26942 16244
rect 30101 16235 30159 16241
rect 26936 16204 29960 16232
rect 26936 16192 26942 16204
rect 23716 16136 24992 16164
rect 23716 16124 23722 16136
rect 18598 16056 18604 16108
rect 18656 16096 18662 16108
rect 19153 16099 19211 16105
rect 19153 16096 19165 16099
rect 18656 16068 19165 16096
rect 18656 16056 18662 16068
rect 19153 16065 19165 16068
rect 19199 16065 19211 16099
rect 19153 16059 19211 16065
rect 18095 16000 18552 16028
rect 18095 15997 18107 16000
rect 18049 15991 18107 15997
rect 16482 15960 16488 15972
rect 15764 15932 16488 15960
rect 16482 15920 16488 15932
rect 16540 15920 16546 15972
rect 16761 15963 16819 15969
rect 16761 15929 16773 15963
rect 16807 15960 16819 15963
rect 16942 15960 16948 15972
rect 16807 15932 16948 15960
rect 16807 15929 16819 15932
rect 16761 15923 16819 15929
rect 16942 15920 16948 15932
rect 17000 15920 17006 15972
rect 17880 15960 17908 15991
rect 22738 15988 22744 16040
rect 22796 16028 22802 16040
rect 23768 16037 23796 16136
rect 26786 16124 26792 16176
rect 26844 16164 26850 16176
rect 27614 16164 27620 16176
rect 26844 16136 27620 16164
rect 26844 16124 26850 16136
rect 27614 16124 27620 16136
rect 27672 16124 27678 16176
rect 29932 16164 29960 16204
rect 30101 16201 30113 16235
rect 30147 16232 30159 16235
rect 30742 16232 30748 16244
rect 30147 16204 30748 16232
rect 30147 16201 30159 16204
rect 30101 16195 30159 16201
rect 30742 16192 30748 16204
rect 30800 16192 30806 16244
rect 30926 16192 30932 16244
rect 30984 16192 30990 16244
rect 31018 16192 31024 16244
rect 31076 16192 31082 16244
rect 33962 16192 33968 16244
rect 34020 16192 34026 16244
rect 34514 16192 34520 16244
rect 34572 16232 34578 16244
rect 34572 16204 34836 16232
rect 34572 16192 34578 16204
rect 32769 16167 32827 16173
rect 32769 16164 32781 16167
rect 29932 16136 32781 16164
rect 32769 16133 32781 16136
rect 32815 16133 32827 16167
rect 33410 16164 33416 16176
rect 32769 16127 32827 16133
rect 33244 16136 33416 16164
rect 24578 16056 24584 16108
rect 24636 16056 24642 16108
rect 25958 16056 25964 16108
rect 26016 16056 26022 16108
rect 26602 16056 26608 16108
rect 26660 16096 26666 16108
rect 27525 16099 27583 16105
rect 27525 16096 27537 16099
rect 26660 16068 27537 16096
rect 26660 16056 26666 16068
rect 27525 16065 27537 16068
rect 27571 16065 27583 16099
rect 27525 16059 27583 16065
rect 28350 16056 28356 16108
rect 28408 16056 28414 16108
rect 31478 16096 31484 16108
rect 29762 16082 31484 16096
rect 29748 16068 31484 16082
rect 23569 16031 23627 16037
rect 23569 16028 23581 16031
rect 22796 16000 23581 16028
rect 22796 15988 22802 16000
rect 23569 15997 23581 16000
rect 23615 15997 23627 16031
rect 23569 15991 23627 15997
rect 23753 16031 23811 16037
rect 23753 15997 23765 16031
rect 23799 15997 23811 16031
rect 23753 15991 23811 15997
rect 24118 15988 24124 16040
rect 24176 16028 24182 16040
rect 24857 16031 24915 16037
rect 24857 16028 24869 16031
rect 24176 16000 24869 16028
rect 24176 15988 24182 16000
rect 24857 15997 24869 16000
rect 24903 16028 24915 16031
rect 26050 16028 26056 16040
rect 24903 16000 26056 16028
rect 24903 15997 24915 16000
rect 24857 15991 24915 15997
rect 26050 15988 26056 16000
rect 26108 15988 26114 16040
rect 26234 15988 26240 16040
rect 26292 16028 26298 16040
rect 27430 16028 27436 16040
rect 26292 16000 27436 16028
rect 26292 15988 26298 16000
rect 27430 15988 27436 16000
rect 27488 15988 27494 16040
rect 27709 16031 27767 16037
rect 27709 15997 27721 16031
rect 27755 15997 27767 16031
rect 27709 15991 27767 15997
rect 19058 15960 19064 15972
rect 17880 15932 19064 15960
rect 19058 15920 19064 15932
rect 19116 15920 19122 15972
rect 20901 15963 20959 15969
rect 20901 15929 20913 15963
rect 20947 15960 20959 15963
rect 20947 15932 21680 15960
rect 20947 15929 20959 15932
rect 20901 15923 20959 15929
rect 7929 15895 7987 15901
rect 7929 15861 7941 15895
rect 7975 15892 7987 15895
rect 9214 15892 9220 15904
rect 7975 15864 9220 15892
rect 7975 15861 7987 15864
rect 7929 15855 7987 15861
rect 9214 15852 9220 15864
rect 9272 15852 9278 15904
rect 10226 15852 10232 15904
rect 10284 15892 10290 15904
rect 10597 15895 10655 15901
rect 10597 15892 10609 15895
rect 10284 15864 10609 15892
rect 10284 15852 10290 15864
rect 10597 15861 10609 15864
rect 10643 15892 10655 15895
rect 11054 15892 11060 15904
rect 10643 15864 11060 15892
rect 10643 15861 10655 15864
rect 10597 15855 10655 15861
rect 11054 15852 11060 15864
rect 11112 15852 11118 15904
rect 11701 15895 11759 15901
rect 11701 15861 11713 15895
rect 11747 15892 11759 15895
rect 11882 15892 11888 15904
rect 11747 15864 11888 15892
rect 11747 15861 11759 15864
rect 11701 15855 11759 15861
rect 11882 15852 11888 15864
rect 11940 15852 11946 15904
rect 15381 15895 15439 15901
rect 15381 15861 15393 15895
rect 15427 15892 15439 15895
rect 15838 15892 15844 15904
rect 15427 15864 15844 15892
rect 15427 15861 15439 15864
rect 15381 15855 15439 15861
rect 15838 15852 15844 15864
rect 15896 15852 15902 15904
rect 16301 15895 16359 15901
rect 16301 15861 16313 15895
rect 16347 15892 16359 15895
rect 16666 15892 16672 15904
rect 16347 15864 16672 15892
rect 16347 15861 16359 15864
rect 16301 15855 16359 15861
rect 16666 15852 16672 15864
rect 16724 15852 16730 15904
rect 16850 15852 16856 15904
rect 16908 15852 16914 15904
rect 17126 15852 17132 15904
rect 17184 15892 17190 15904
rect 20530 15892 20536 15904
rect 17184 15864 20536 15892
rect 17184 15852 17190 15864
rect 20530 15852 20536 15864
rect 20588 15852 20594 15904
rect 21652 15892 21680 15932
rect 22830 15920 22836 15972
rect 22888 15960 22894 15972
rect 24026 15960 24032 15972
rect 22888 15932 24032 15960
rect 22888 15920 22894 15932
rect 24026 15920 24032 15932
rect 24084 15920 24090 15972
rect 26418 15920 26424 15972
rect 26476 15960 26482 15972
rect 27724 15960 27752 15991
rect 28626 15988 28632 16040
rect 28684 16028 28690 16040
rect 29086 16028 29092 16040
rect 28684 16000 29092 16028
rect 28684 15988 28690 16000
rect 29086 15988 29092 16000
rect 29144 15988 29150 16040
rect 29270 15988 29276 16040
rect 29328 16028 29334 16040
rect 29748 16028 29776 16068
rect 31478 16056 31484 16068
rect 31536 16056 31542 16108
rect 32677 16099 32735 16105
rect 32677 16065 32689 16099
rect 32723 16096 32735 16099
rect 33244 16096 33272 16136
rect 33410 16124 33416 16136
rect 33468 16164 33474 16176
rect 34808 16173 34836 16204
rect 35158 16192 35164 16244
rect 35216 16232 35222 16244
rect 36817 16235 36875 16241
rect 36817 16232 36829 16235
rect 35216 16204 36829 16232
rect 35216 16192 35222 16204
rect 36817 16201 36829 16204
rect 36863 16232 36875 16235
rect 36906 16232 36912 16244
rect 36863 16204 36912 16232
rect 36863 16201 36875 16204
rect 36817 16195 36875 16201
rect 36906 16192 36912 16204
rect 36964 16192 36970 16244
rect 40034 16192 40040 16244
rect 40092 16232 40098 16244
rect 40957 16235 41015 16241
rect 40957 16232 40969 16235
rect 40092 16204 40969 16232
rect 40092 16192 40098 16204
rect 40957 16201 40969 16204
rect 41003 16201 41015 16235
rect 40957 16195 41015 16201
rect 34793 16167 34851 16173
rect 33468 16136 34652 16164
rect 33468 16124 33474 16136
rect 32723 16068 33272 16096
rect 32723 16065 32735 16068
rect 32677 16059 32735 16065
rect 33318 16056 33324 16108
rect 33376 16096 33382 16108
rect 33873 16099 33931 16105
rect 33873 16096 33885 16099
rect 33376 16068 33885 16096
rect 33376 16056 33382 16068
rect 33873 16065 33885 16068
rect 33919 16065 33931 16099
rect 33873 16059 33931 16065
rect 31113 16031 31171 16037
rect 31113 16028 31125 16031
rect 29328 16000 29776 16028
rect 30484 16000 31125 16028
rect 29328 15988 29334 16000
rect 26476 15932 27752 15960
rect 26476 15920 26482 15932
rect 22278 15892 22284 15904
rect 21652 15864 22284 15892
rect 22278 15852 22284 15864
rect 22336 15892 22342 15904
rect 25314 15892 25320 15904
rect 22336 15864 25320 15892
rect 22336 15852 22342 15864
rect 25314 15852 25320 15864
rect 25372 15852 25378 15904
rect 25958 15852 25964 15904
rect 26016 15892 26022 15904
rect 26602 15892 26608 15904
rect 26016 15864 26608 15892
rect 26016 15852 26022 15864
rect 26602 15852 26608 15864
rect 26660 15852 26666 15904
rect 26694 15852 26700 15904
rect 26752 15892 26758 15904
rect 27157 15895 27215 15901
rect 27157 15892 27169 15895
rect 26752 15864 27169 15892
rect 26752 15852 26758 15864
rect 27157 15861 27169 15864
rect 27203 15861 27215 15895
rect 27157 15855 27215 15861
rect 29730 15852 29736 15904
rect 29788 15892 29794 15904
rect 30484 15892 30512 16000
rect 31113 15997 31125 16000
rect 31159 15997 31171 16031
rect 31113 15991 31171 15997
rect 31846 15988 31852 16040
rect 31904 16028 31910 16040
rect 32766 16028 32772 16040
rect 31904 16000 32772 16028
rect 31904 15988 31910 16000
rect 32766 15988 32772 16000
rect 32824 16028 32830 16040
rect 34624 16037 34652 16136
rect 34793 16133 34805 16167
rect 34839 16164 34851 16167
rect 35434 16164 35440 16176
rect 34839 16136 35440 16164
rect 34839 16133 34851 16136
rect 34793 16127 34851 16133
rect 35434 16124 35440 16136
rect 35492 16124 35498 16176
rect 37458 16124 37464 16176
rect 37516 16164 37522 16176
rect 38473 16167 38531 16173
rect 37516 16136 38240 16164
rect 37516 16124 37522 16136
rect 36446 16056 36452 16108
rect 36504 16056 36510 16108
rect 38212 16105 38240 16136
rect 38473 16133 38485 16167
rect 38519 16164 38531 16167
rect 38562 16164 38568 16176
rect 38519 16136 38568 16164
rect 38519 16133 38531 16136
rect 38473 16127 38531 16133
rect 38562 16124 38568 16136
rect 38620 16124 38626 16176
rect 39758 16164 39764 16176
rect 39698 16136 39764 16164
rect 39758 16124 39764 16136
rect 39816 16164 39822 16176
rect 41322 16164 41328 16176
rect 39816 16136 41328 16164
rect 39816 16124 39822 16136
rect 41322 16124 41328 16136
rect 41380 16124 41386 16176
rect 38197 16099 38255 16105
rect 38197 16065 38209 16099
rect 38243 16065 38255 16099
rect 38197 16059 38255 16065
rect 40865 16099 40923 16105
rect 40865 16065 40877 16099
rect 40911 16096 40923 16099
rect 48682 16096 48688 16108
rect 40911 16068 48688 16096
rect 40911 16065 40923 16068
rect 40865 16059 40923 16065
rect 48682 16056 48688 16068
rect 48740 16056 48746 16108
rect 48777 16099 48835 16105
rect 48777 16065 48789 16099
rect 48823 16096 48835 16099
rect 49050 16096 49056 16108
rect 48823 16068 49056 16096
rect 48823 16065 48835 16068
rect 48777 16059 48835 16065
rect 49050 16056 49056 16068
rect 49108 16056 49114 16108
rect 32861 16031 32919 16037
rect 32861 16028 32873 16031
rect 32824 16000 32873 16028
rect 32824 15988 32830 16000
rect 32861 15997 32873 16000
rect 32907 15997 32919 16031
rect 32861 15991 32919 15997
rect 34057 16031 34115 16037
rect 34057 15997 34069 16031
rect 34103 15997 34115 16031
rect 34057 15991 34115 15997
rect 34609 16031 34667 16037
rect 34609 15997 34621 16031
rect 34655 16028 34667 16031
rect 34790 16028 34796 16040
rect 34655 16000 34796 16028
rect 34655 15997 34667 16000
rect 34609 15991 34667 15997
rect 30834 15920 30840 15972
rect 30892 15960 30898 15972
rect 32398 15960 32404 15972
rect 30892 15932 32404 15960
rect 30892 15920 30898 15932
rect 32398 15920 32404 15932
rect 32456 15920 32462 15972
rect 32582 15920 32588 15972
rect 32640 15960 32646 15972
rect 34072 15960 34100 15991
rect 34790 15988 34796 16000
rect 34848 15988 34854 16040
rect 34882 15988 34888 16040
rect 34940 16028 34946 16040
rect 35069 16031 35127 16037
rect 35069 16028 35081 16031
rect 34940 16000 35081 16028
rect 34940 15988 34946 16000
rect 35069 15997 35081 16000
rect 35115 15997 35127 16031
rect 35069 15991 35127 15997
rect 35345 16031 35403 16037
rect 35345 15997 35357 16031
rect 35391 16028 35403 16031
rect 36814 16028 36820 16040
rect 35391 16000 36820 16028
rect 35391 15997 35403 16000
rect 35345 15991 35403 15997
rect 36814 15988 36820 16000
rect 36872 15988 36878 16040
rect 37274 15988 37280 16040
rect 37332 16028 37338 16040
rect 37461 16031 37519 16037
rect 37461 16028 37473 16031
rect 37332 16000 37473 16028
rect 37332 15988 37338 16000
rect 37461 15997 37473 16000
rect 37507 15997 37519 16031
rect 37461 15991 37519 15997
rect 39945 16031 40003 16037
rect 39945 15997 39957 16031
rect 39991 16028 40003 16031
rect 40310 16028 40316 16040
rect 39991 16000 40316 16028
rect 39991 15997 40003 16000
rect 39945 15991 40003 15997
rect 40310 15988 40316 16000
rect 40368 16028 40374 16040
rect 40586 16028 40592 16040
rect 40368 16000 40592 16028
rect 40368 15988 40374 16000
rect 40586 15988 40592 16000
rect 40644 15988 40650 16040
rect 41046 15988 41052 16040
rect 41104 15988 41110 16040
rect 37734 15960 37740 15972
rect 32640 15932 34100 15960
rect 34440 15932 35204 15960
rect 32640 15920 32646 15932
rect 29788 15864 30512 15892
rect 29788 15852 29794 15864
rect 30558 15852 30564 15904
rect 30616 15852 30622 15904
rect 31478 15852 31484 15904
rect 31536 15892 31542 15904
rect 31573 15895 31631 15901
rect 31573 15892 31585 15895
rect 31536 15864 31585 15892
rect 31536 15852 31542 15864
rect 31573 15861 31585 15864
rect 31619 15861 31631 15895
rect 31573 15855 31631 15861
rect 31662 15852 31668 15904
rect 31720 15892 31726 15904
rect 31757 15895 31815 15901
rect 31757 15892 31769 15895
rect 31720 15864 31769 15892
rect 31720 15852 31726 15864
rect 31757 15861 31769 15864
rect 31803 15861 31815 15895
rect 31757 15855 31815 15861
rect 32309 15895 32367 15901
rect 32309 15861 32321 15895
rect 32355 15892 32367 15895
rect 33410 15892 33416 15904
rect 32355 15864 33416 15892
rect 32355 15861 32367 15864
rect 32309 15855 32367 15861
rect 33410 15852 33416 15864
rect 33468 15852 33474 15904
rect 33505 15895 33563 15901
rect 33505 15861 33517 15895
rect 33551 15892 33563 15895
rect 34440 15892 34468 15932
rect 33551 15864 34468 15892
rect 35176 15892 35204 15932
rect 36740 15932 37740 15960
rect 36740 15892 36768 15932
rect 37734 15920 37740 15932
rect 37792 15920 37798 15972
rect 49234 15920 49240 15972
rect 49292 15920 49298 15972
rect 35176 15864 36768 15892
rect 33551 15861 33563 15864
rect 33505 15855 33563 15861
rect 37366 15852 37372 15904
rect 37424 15892 37430 15904
rect 40497 15895 40555 15901
rect 40497 15892 40509 15895
rect 37424 15864 40509 15892
rect 37424 15852 37430 15864
rect 40497 15861 40509 15864
rect 40543 15861 40555 15895
rect 40497 15855 40555 15861
rect 41598 15852 41604 15904
rect 41656 15852 41662 15904
rect 1104 15802 49864 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 32950 15802
rect 33002 15750 33014 15802
rect 33066 15750 33078 15802
rect 33130 15750 33142 15802
rect 33194 15750 33206 15802
rect 33258 15750 42950 15802
rect 43002 15750 43014 15802
rect 43066 15750 43078 15802
rect 43130 15750 43142 15802
rect 43194 15750 43206 15802
rect 43258 15750 49864 15802
rect 1104 15728 49864 15750
rect 10778 15648 10784 15700
rect 10836 15688 10842 15700
rect 10836 15660 14780 15688
rect 10836 15648 10842 15660
rect 12066 15580 12072 15632
rect 12124 15620 12130 15632
rect 14277 15623 14335 15629
rect 14277 15620 14289 15623
rect 12124 15592 14289 15620
rect 12124 15580 12130 15592
rect 14277 15589 14289 15592
rect 14323 15589 14335 15623
rect 14752 15620 14780 15660
rect 14826 15648 14832 15700
rect 14884 15688 14890 15700
rect 14884 15660 16068 15688
rect 14884 15648 14890 15660
rect 15470 15620 15476 15632
rect 14752 15592 15476 15620
rect 14277 15583 14335 15589
rect 15470 15580 15476 15592
rect 15528 15580 15534 15632
rect 15565 15623 15623 15629
rect 15565 15589 15577 15623
rect 15611 15589 15623 15623
rect 15565 15583 15623 15589
rect 1302 15512 1308 15564
rect 1360 15552 1366 15564
rect 2041 15555 2099 15561
rect 2041 15552 2053 15555
rect 1360 15524 2053 15552
rect 1360 15512 1366 15524
rect 2041 15521 2053 15524
rect 2087 15521 2099 15555
rect 2041 15515 2099 15521
rect 10594 15512 10600 15564
rect 10652 15552 10658 15564
rect 10781 15555 10839 15561
rect 10781 15552 10793 15555
rect 10652 15524 10793 15552
rect 10652 15512 10658 15524
rect 10781 15521 10793 15524
rect 10827 15521 10839 15555
rect 10781 15515 10839 15521
rect 11057 15555 11115 15561
rect 11057 15521 11069 15555
rect 11103 15552 11115 15555
rect 12802 15552 12808 15564
rect 11103 15524 12808 15552
rect 11103 15521 11115 15524
rect 11057 15515 11115 15521
rect 12802 15512 12808 15524
rect 12860 15512 12866 15564
rect 13446 15512 13452 15564
rect 13504 15512 13510 15564
rect 13633 15555 13691 15561
rect 13633 15521 13645 15555
rect 13679 15521 13691 15555
rect 13633 15515 13691 15521
rect 1765 15487 1823 15493
rect 1765 15453 1777 15487
rect 1811 15484 1823 15487
rect 10410 15484 10416 15496
rect 1811 15456 10416 15484
rect 1811 15453 1823 15456
rect 1765 15447 1823 15453
rect 10410 15444 10416 15456
rect 10468 15444 10474 15496
rect 12710 15444 12716 15496
rect 12768 15484 12774 15496
rect 13357 15487 13415 15493
rect 13357 15484 13369 15487
rect 12768 15456 13369 15484
rect 12768 15444 12774 15456
rect 13357 15453 13369 15456
rect 13403 15453 13415 15487
rect 13648 15484 13676 15515
rect 14826 15512 14832 15564
rect 14884 15512 14890 15564
rect 15378 15512 15384 15564
rect 15436 15552 15442 15564
rect 15580 15552 15608 15583
rect 15930 15580 15936 15632
rect 15988 15580 15994 15632
rect 16040 15620 16068 15660
rect 16574 15648 16580 15700
rect 16632 15688 16638 15700
rect 16761 15691 16819 15697
rect 16761 15688 16773 15691
rect 16632 15660 16773 15688
rect 16632 15648 16638 15660
rect 16761 15657 16773 15660
rect 16807 15657 16819 15691
rect 17126 15688 17132 15700
rect 16761 15651 16819 15657
rect 16868 15660 17132 15688
rect 16868 15620 16896 15660
rect 17126 15648 17132 15660
rect 17184 15648 17190 15700
rect 18506 15648 18512 15700
rect 18564 15688 18570 15700
rect 18969 15691 19027 15697
rect 18969 15688 18981 15691
rect 18564 15660 18981 15688
rect 18564 15648 18570 15660
rect 18969 15657 18981 15660
rect 19015 15657 19027 15691
rect 18969 15651 19027 15657
rect 19337 15691 19395 15697
rect 19337 15657 19349 15691
rect 19383 15688 19395 15691
rect 19426 15688 19432 15700
rect 19383 15660 19432 15688
rect 19383 15657 19395 15660
rect 19337 15651 19395 15657
rect 19426 15648 19432 15660
rect 19484 15648 19490 15700
rect 19886 15648 19892 15700
rect 19944 15648 19950 15700
rect 21177 15691 21235 15697
rect 21177 15688 21189 15691
rect 19996 15660 21189 15688
rect 16040 15592 16896 15620
rect 15436 15524 15608 15552
rect 15436 15512 15442 15524
rect 15838 15484 15844 15496
rect 13648 15456 15844 15484
rect 13357 15447 13415 15453
rect 15838 15444 15844 15456
rect 15896 15444 15902 15496
rect 15948 15493 15976 15580
rect 16040 15561 16068 15592
rect 16942 15580 16948 15632
rect 17000 15620 17006 15632
rect 17000 15592 17172 15620
rect 17000 15580 17006 15592
rect 16025 15555 16083 15561
rect 16025 15521 16037 15555
rect 16071 15521 16083 15555
rect 16025 15515 16083 15521
rect 16209 15555 16267 15561
rect 16209 15521 16221 15555
rect 16255 15552 16267 15555
rect 16482 15552 16488 15564
rect 16255 15524 16488 15552
rect 16255 15521 16267 15524
rect 16209 15515 16267 15521
rect 16482 15512 16488 15524
rect 16540 15512 16546 15564
rect 17144 15493 17172 15592
rect 19150 15580 19156 15632
rect 19208 15620 19214 15632
rect 19996 15620 20024 15660
rect 21177 15657 21189 15660
rect 21223 15657 21235 15691
rect 21177 15651 21235 15657
rect 21726 15648 21732 15700
rect 21784 15688 21790 15700
rect 22462 15688 22468 15700
rect 21784 15660 22468 15688
rect 21784 15648 21790 15660
rect 22462 15648 22468 15660
rect 22520 15648 22526 15700
rect 23474 15648 23480 15700
rect 23532 15688 23538 15700
rect 25869 15691 25927 15697
rect 25869 15688 25881 15691
rect 23532 15660 25881 15688
rect 23532 15648 23538 15660
rect 25869 15657 25881 15660
rect 25915 15657 25927 15691
rect 25869 15651 25927 15657
rect 26602 15648 26608 15700
rect 26660 15688 26666 15700
rect 26878 15688 26884 15700
rect 26660 15660 26884 15688
rect 26660 15648 26666 15660
rect 26878 15648 26884 15660
rect 26936 15648 26942 15700
rect 27157 15691 27215 15697
rect 27157 15657 27169 15691
rect 27203 15688 27215 15691
rect 27338 15688 27344 15700
rect 27203 15660 27344 15688
rect 27203 15657 27215 15660
rect 27157 15651 27215 15657
rect 27338 15648 27344 15660
rect 27396 15648 27402 15700
rect 32217 15691 32275 15697
rect 32217 15657 32229 15691
rect 32263 15688 32275 15691
rect 32582 15688 32588 15700
rect 32263 15660 32588 15688
rect 32263 15657 32275 15660
rect 32217 15651 32275 15657
rect 32582 15648 32588 15660
rect 32640 15648 32646 15700
rect 34146 15648 34152 15700
rect 34204 15688 34210 15700
rect 34333 15691 34391 15697
rect 34333 15688 34345 15691
rect 34204 15660 34345 15688
rect 34204 15648 34210 15660
rect 34333 15657 34345 15660
rect 34379 15657 34391 15691
rect 34333 15651 34391 15657
rect 36633 15691 36691 15697
rect 36633 15657 36645 15691
rect 36679 15688 36691 15691
rect 36814 15688 36820 15700
rect 36679 15660 36820 15688
rect 36679 15657 36691 15660
rect 36633 15651 36691 15657
rect 36814 15648 36820 15660
rect 36872 15648 36878 15700
rect 36998 15648 37004 15700
rect 37056 15688 37062 15700
rect 37826 15688 37832 15700
rect 37056 15660 37832 15688
rect 37056 15648 37062 15660
rect 37826 15648 37832 15660
rect 37884 15688 37890 15700
rect 39485 15691 39543 15697
rect 39485 15688 39497 15691
rect 37884 15660 39497 15688
rect 37884 15648 37890 15660
rect 39485 15657 39497 15660
rect 39531 15657 39543 15691
rect 39485 15651 39543 15657
rect 41598 15648 41604 15700
rect 41656 15688 41662 15700
rect 42061 15691 42119 15697
rect 42061 15688 42073 15691
rect 41656 15660 42073 15688
rect 41656 15648 41662 15660
rect 42061 15657 42073 15660
rect 42107 15657 42119 15691
rect 42061 15651 42119 15657
rect 48682 15648 48688 15700
rect 48740 15688 48746 15700
rect 49145 15691 49203 15697
rect 49145 15688 49157 15691
rect 48740 15660 49157 15688
rect 48740 15648 48746 15660
rect 49145 15657 49157 15660
rect 49191 15657 49203 15691
rect 49145 15651 49203 15657
rect 28810 15620 28816 15632
rect 19208 15592 20024 15620
rect 20272 15592 28816 15620
rect 19208 15580 19214 15592
rect 17221 15555 17279 15561
rect 17221 15521 17233 15555
rect 17267 15521 17279 15555
rect 17221 15515 17279 15521
rect 15933 15487 15991 15493
rect 15933 15453 15945 15487
rect 15979 15453 15991 15487
rect 15933 15447 15991 15453
rect 17129 15487 17187 15493
rect 17129 15453 17141 15487
rect 17175 15453 17187 15487
rect 17236 15484 17264 15515
rect 17310 15512 17316 15564
rect 17368 15512 17374 15564
rect 17773 15487 17831 15493
rect 17773 15484 17785 15487
rect 17236 15456 17785 15484
rect 17129 15447 17187 15453
rect 17773 15453 17785 15456
rect 17819 15484 17831 15487
rect 18601 15487 18659 15493
rect 17819 15456 18552 15484
rect 17819 15453 17831 15456
rect 17773 15447 17831 15453
rect 6457 15419 6515 15425
rect 6457 15385 6469 15419
rect 6503 15416 6515 15419
rect 6503 15388 10364 15416
rect 6503 15385 6515 15388
rect 6457 15379 6515 15385
rect 6546 15308 6552 15360
rect 6604 15308 6610 15360
rect 10336 15348 10364 15388
rect 11698 15376 11704 15428
rect 11756 15376 11762 15428
rect 13630 15416 13636 15428
rect 13004 15388 13636 15416
rect 11790 15348 11796 15360
rect 10336 15320 11796 15348
rect 11790 15308 11796 15320
rect 11848 15308 11854 15360
rect 12526 15308 12532 15360
rect 12584 15308 12590 15360
rect 13004 15357 13032 15388
rect 13630 15376 13636 15388
rect 13688 15376 13694 15428
rect 14737 15419 14795 15425
rect 14737 15385 14749 15419
rect 14783 15416 14795 15419
rect 17862 15416 17868 15428
rect 14783 15388 17868 15416
rect 14783 15385 14795 15388
rect 14737 15379 14795 15385
rect 17862 15376 17868 15388
rect 17920 15376 17926 15428
rect 18524 15416 18552 15456
rect 18601 15453 18613 15487
rect 18647 15484 18659 15487
rect 19794 15484 19800 15496
rect 18647 15456 19800 15484
rect 18647 15453 18659 15456
rect 18601 15447 18659 15453
rect 19794 15444 19800 15456
rect 19852 15444 19858 15496
rect 20272 15416 20300 15592
rect 28810 15580 28816 15592
rect 28868 15580 28874 15632
rect 34164 15620 34192 15648
rect 31864 15592 34192 15620
rect 20533 15555 20591 15561
rect 20533 15521 20545 15555
rect 20579 15552 20591 15555
rect 21358 15552 21364 15564
rect 20579 15524 21364 15552
rect 20579 15521 20591 15524
rect 20533 15515 20591 15521
rect 21358 15512 21364 15524
rect 21416 15512 21422 15564
rect 21637 15555 21695 15561
rect 21637 15552 21649 15555
rect 21468 15524 21649 15552
rect 21082 15444 21088 15496
rect 21140 15484 21146 15496
rect 21468 15484 21496 15524
rect 21637 15521 21649 15524
rect 21683 15552 21695 15555
rect 21726 15552 21732 15564
rect 21683 15524 21732 15552
rect 21683 15521 21695 15524
rect 21637 15515 21695 15521
rect 21726 15512 21732 15524
rect 21784 15512 21790 15564
rect 21821 15555 21879 15561
rect 21821 15521 21833 15555
rect 21867 15552 21879 15555
rect 21910 15552 21916 15564
rect 21867 15524 21916 15552
rect 21867 15521 21879 15524
rect 21821 15515 21879 15521
rect 21910 15512 21916 15524
rect 21968 15512 21974 15564
rect 23753 15555 23811 15561
rect 23753 15521 23765 15555
rect 23799 15552 23811 15555
rect 23842 15552 23848 15564
rect 23799 15524 23848 15552
rect 23799 15521 23811 15524
rect 23753 15515 23811 15521
rect 23842 15512 23848 15524
rect 23900 15512 23906 15564
rect 23934 15512 23940 15564
rect 23992 15552 23998 15564
rect 25038 15552 25044 15564
rect 23992 15524 25044 15552
rect 23992 15512 23998 15524
rect 25038 15512 25044 15524
rect 25096 15552 25102 15564
rect 25133 15555 25191 15561
rect 25133 15552 25145 15555
rect 25096 15524 25145 15552
rect 25096 15512 25102 15524
rect 25133 15521 25145 15524
rect 25179 15521 25191 15555
rect 25133 15515 25191 15521
rect 25314 15512 25320 15564
rect 25372 15552 25378 15564
rect 26234 15552 26240 15564
rect 25372 15524 26240 15552
rect 25372 15512 25378 15524
rect 26234 15512 26240 15524
rect 26292 15512 26298 15564
rect 26510 15512 26516 15564
rect 26568 15512 26574 15564
rect 26602 15512 26608 15564
rect 26660 15552 26666 15564
rect 27985 15555 28043 15561
rect 27985 15552 27997 15555
rect 26660 15524 27997 15552
rect 26660 15512 26666 15524
rect 27985 15521 27997 15524
rect 28031 15521 28043 15555
rect 27985 15515 28043 15521
rect 30742 15512 30748 15564
rect 30800 15512 30806 15564
rect 31478 15512 31484 15564
rect 31536 15552 31542 15564
rect 31864 15552 31892 15592
rect 31536 15524 31892 15552
rect 31536 15512 31542 15524
rect 21140 15456 21496 15484
rect 21140 15444 21146 15456
rect 21542 15444 21548 15496
rect 21600 15484 21606 15496
rect 22189 15487 22247 15493
rect 22189 15484 22201 15487
rect 21600 15456 22201 15484
rect 21600 15444 21606 15456
rect 22189 15453 22201 15456
rect 22235 15453 22247 15487
rect 22189 15447 22247 15453
rect 23569 15487 23627 15493
rect 23569 15453 23581 15487
rect 23615 15484 23627 15487
rect 27154 15484 27160 15496
rect 23615 15456 27160 15484
rect 23615 15453 23627 15456
rect 23569 15447 23627 15453
rect 27154 15444 27160 15456
rect 27212 15444 27218 15496
rect 27798 15444 27804 15496
rect 27856 15484 27862 15496
rect 28445 15487 28503 15493
rect 28445 15484 28457 15487
rect 27856 15456 28457 15484
rect 27856 15444 27862 15456
rect 28445 15453 28457 15456
rect 28491 15453 28503 15487
rect 28445 15447 28503 15453
rect 30466 15444 30472 15496
rect 30524 15444 30530 15496
rect 31864 15470 31892 15524
rect 32214 15512 32220 15564
rect 32272 15552 32278 15564
rect 33137 15555 33195 15561
rect 33137 15552 33149 15555
rect 32272 15524 33149 15552
rect 32272 15512 32278 15524
rect 33137 15521 33149 15524
rect 33183 15521 33195 15555
rect 33137 15515 33195 15521
rect 33321 15555 33379 15561
rect 33321 15521 33333 15555
rect 33367 15552 33379 15555
rect 33502 15552 33508 15564
rect 33367 15524 33508 15552
rect 33367 15521 33379 15524
rect 33321 15515 33379 15521
rect 33502 15512 33508 15524
rect 33560 15552 33566 15564
rect 34146 15552 34152 15564
rect 33560 15524 34152 15552
rect 33560 15512 33566 15524
rect 34146 15512 34152 15524
rect 34204 15512 34210 15564
rect 35161 15555 35219 15561
rect 35161 15521 35173 15555
rect 35207 15552 35219 15555
rect 36354 15552 36360 15564
rect 35207 15524 36360 15552
rect 35207 15521 35219 15524
rect 35161 15515 35219 15521
rect 36354 15512 36360 15524
rect 36412 15512 36418 15564
rect 40037 15555 40095 15561
rect 40037 15552 40049 15555
rect 37752 15524 40049 15552
rect 32674 15444 32680 15496
rect 32732 15484 32738 15496
rect 33045 15487 33103 15493
rect 33045 15484 33057 15487
rect 32732 15456 33057 15484
rect 32732 15444 32738 15456
rect 33045 15453 33057 15456
rect 33091 15484 33103 15487
rect 34514 15484 34520 15496
rect 33091 15456 34520 15484
rect 33091 15453 33103 15456
rect 33045 15447 33103 15453
rect 34514 15444 34520 15456
rect 34572 15444 34578 15496
rect 34882 15444 34888 15496
rect 34940 15444 34946 15496
rect 37458 15444 37464 15496
rect 37516 15484 37522 15496
rect 37752 15493 37780 15524
rect 40037 15521 40049 15524
rect 40083 15521 40095 15555
rect 40037 15515 40095 15521
rect 40310 15512 40316 15564
rect 40368 15512 40374 15564
rect 37737 15487 37795 15493
rect 37737 15484 37749 15487
rect 37516 15456 37749 15484
rect 37516 15444 37522 15456
rect 37737 15453 37749 15456
rect 37783 15453 37795 15487
rect 37737 15447 37795 15453
rect 48869 15487 48927 15493
rect 48869 15453 48881 15487
rect 48915 15484 48927 15487
rect 49326 15484 49332 15496
rect 48915 15456 49332 15484
rect 48915 15453 48927 15456
rect 48869 15447 48927 15453
rect 49326 15444 49332 15456
rect 49384 15444 49390 15496
rect 18524 15388 20300 15416
rect 20349 15419 20407 15425
rect 20349 15385 20361 15419
rect 20395 15416 20407 15419
rect 23477 15419 23535 15425
rect 20395 15388 23152 15416
rect 20395 15385 20407 15388
rect 20349 15379 20407 15385
rect 12989 15351 13047 15357
rect 12989 15317 13001 15351
rect 13035 15317 13047 15351
rect 12989 15311 13047 15317
rect 14458 15308 14464 15360
rect 14516 15348 14522 15360
rect 14645 15351 14703 15357
rect 14645 15348 14657 15351
rect 14516 15320 14657 15348
rect 14516 15308 14522 15320
rect 14645 15317 14657 15320
rect 14691 15317 14703 15351
rect 14645 15311 14703 15317
rect 15470 15308 15476 15360
rect 15528 15348 15534 15360
rect 16022 15348 16028 15360
rect 15528 15320 16028 15348
rect 15528 15308 15534 15320
rect 16022 15308 16028 15320
rect 16080 15348 16086 15360
rect 18417 15351 18475 15357
rect 18417 15348 18429 15351
rect 16080 15320 18429 15348
rect 16080 15308 16086 15320
rect 18417 15317 18429 15320
rect 18463 15317 18475 15351
rect 18417 15311 18475 15317
rect 20254 15308 20260 15360
rect 20312 15308 20318 15360
rect 23124 15357 23152 15388
rect 23477 15385 23489 15419
rect 23523 15416 23535 15419
rect 25041 15419 25099 15425
rect 23523 15388 24716 15416
rect 23523 15385 23535 15388
rect 23477 15379 23535 15385
rect 24688 15357 24716 15388
rect 25041 15385 25053 15419
rect 25087 15416 25099 15419
rect 25590 15416 25596 15428
rect 25087 15388 25596 15416
rect 25087 15385 25099 15388
rect 25041 15379 25099 15385
rect 25590 15376 25596 15388
rect 25648 15376 25654 15428
rect 26326 15376 26332 15428
rect 26384 15416 26390 15428
rect 27338 15416 27344 15428
rect 26384 15388 27344 15416
rect 26384 15376 26390 15388
rect 27338 15376 27344 15388
rect 27396 15376 27402 15428
rect 27706 15376 27712 15428
rect 27764 15416 27770 15428
rect 27893 15419 27951 15425
rect 27893 15416 27905 15419
rect 27764 15388 27905 15416
rect 27764 15376 27770 15388
rect 27893 15385 27905 15388
rect 27939 15416 27951 15419
rect 28629 15419 28687 15425
rect 28629 15416 28641 15419
rect 27939 15388 28641 15416
rect 27939 15385 27951 15388
rect 27893 15379 27951 15385
rect 28629 15385 28641 15388
rect 28675 15385 28687 15419
rect 28629 15379 28687 15385
rect 29181 15419 29239 15425
rect 29181 15385 29193 15419
rect 29227 15416 29239 15419
rect 30374 15416 30380 15428
rect 29227 15388 30380 15416
rect 29227 15385 29239 15388
rect 29181 15379 29239 15385
rect 30374 15376 30380 15388
rect 30432 15376 30438 15428
rect 36446 15416 36452 15428
rect 32600 15388 35572 15416
rect 36386 15388 36452 15416
rect 23109 15351 23167 15357
rect 23109 15317 23121 15351
rect 23155 15317 23167 15351
rect 23109 15311 23167 15317
rect 24673 15351 24731 15357
rect 24673 15317 24685 15351
rect 24719 15317 24731 15351
rect 24673 15311 24731 15317
rect 26237 15351 26295 15357
rect 26237 15317 26249 15351
rect 26283 15348 26295 15351
rect 26970 15348 26976 15360
rect 26283 15320 26976 15348
rect 26283 15317 26295 15320
rect 26237 15311 26295 15317
rect 26970 15308 26976 15320
rect 27028 15308 27034 15360
rect 27430 15308 27436 15360
rect 27488 15308 27494 15360
rect 29270 15308 29276 15360
rect 29328 15308 29334 15360
rect 29825 15351 29883 15357
rect 29825 15317 29837 15351
rect 29871 15348 29883 15351
rect 31110 15348 31116 15360
rect 29871 15320 31116 15348
rect 29871 15317 29883 15320
rect 29825 15311 29883 15317
rect 31110 15308 31116 15320
rect 31168 15308 31174 15360
rect 31478 15308 31484 15360
rect 31536 15348 31542 15360
rect 31662 15348 31668 15360
rect 31536 15320 31668 15348
rect 31536 15308 31542 15320
rect 31662 15308 31668 15320
rect 31720 15348 31726 15360
rect 32600 15348 32628 15388
rect 31720 15320 32628 15348
rect 31720 15308 31726 15320
rect 32674 15308 32680 15360
rect 32732 15308 32738 15360
rect 33870 15308 33876 15360
rect 33928 15308 33934 15360
rect 35544 15348 35572 15388
rect 36446 15376 36452 15388
rect 36504 15376 36510 15428
rect 37366 15376 37372 15428
rect 37424 15416 37430 15428
rect 38013 15419 38071 15425
rect 38013 15416 38025 15419
rect 37424 15388 38025 15416
rect 37424 15376 37430 15388
rect 38013 15385 38025 15388
rect 38059 15385 38071 15419
rect 39758 15416 39764 15428
rect 39238 15388 39764 15416
rect 38013 15379 38071 15385
rect 36078 15348 36084 15360
rect 35544 15320 36084 15348
rect 36078 15308 36084 15320
rect 36136 15348 36142 15360
rect 36538 15348 36544 15360
rect 36136 15320 36544 15348
rect 36136 15308 36142 15320
rect 36538 15308 36544 15320
rect 36596 15308 36602 15360
rect 37090 15308 37096 15360
rect 37148 15308 37154 15360
rect 38028 15348 38056 15379
rect 39758 15376 39764 15388
rect 39816 15376 39822 15428
rect 41322 15376 41328 15428
rect 41380 15376 41386 15428
rect 41046 15348 41052 15360
rect 38028 15320 41052 15348
rect 41046 15308 41052 15320
rect 41104 15348 41110 15360
rect 41785 15351 41843 15357
rect 41785 15348 41797 15351
rect 41104 15320 41797 15348
rect 41104 15308 41110 15320
rect 41785 15317 41797 15320
rect 41831 15317 41843 15351
rect 41785 15311 41843 15317
rect 1104 15258 49864 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 27950 15258
rect 28002 15206 28014 15258
rect 28066 15206 28078 15258
rect 28130 15206 28142 15258
rect 28194 15206 28206 15258
rect 28258 15206 37950 15258
rect 38002 15206 38014 15258
rect 38066 15206 38078 15258
rect 38130 15206 38142 15258
rect 38194 15206 38206 15258
rect 38258 15206 47950 15258
rect 48002 15206 48014 15258
rect 48066 15206 48078 15258
rect 48130 15206 48142 15258
rect 48194 15206 48206 15258
rect 48258 15206 49864 15258
rect 1104 15184 49864 15206
rect 9214 15104 9220 15156
rect 9272 15144 9278 15156
rect 9769 15147 9827 15153
rect 9769 15144 9781 15147
rect 9272 15116 9781 15144
rect 9272 15104 9278 15116
rect 9769 15113 9781 15116
rect 9815 15113 9827 15147
rect 9769 15107 9827 15113
rect 10980 15116 12940 15144
rect 9582 15036 9588 15088
rect 9640 15076 9646 15088
rect 10980 15085 11008 15116
rect 9861 15079 9919 15085
rect 9861 15076 9873 15079
rect 9640 15048 9873 15076
rect 9640 15036 9646 15048
rect 9861 15045 9873 15048
rect 9907 15045 9919 15079
rect 9861 15039 9919 15045
rect 10597 15079 10655 15085
rect 10597 15045 10609 15079
rect 10643 15076 10655 15079
rect 10965 15079 11023 15085
rect 10965 15076 10977 15079
rect 10643 15048 10977 15076
rect 10643 15045 10655 15048
rect 10597 15039 10655 15045
rect 10965 15045 10977 15048
rect 11011 15045 11023 15079
rect 10965 15039 11023 15045
rect 11146 15036 11152 15088
rect 11204 15036 11210 15088
rect 12342 15036 12348 15088
rect 12400 15076 12406 15088
rect 12912 15076 12940 15116
rect 12986 15104 12992 15156
rect 13044 15144 13050 15156
rect 13044 15116 13676 15144
rect 13044 15104 13050 15116
rect 13538 15076 13544 15088
rect 12400 15036 12434 15076
rect 12912 15048 13124 15076
rect 1765 15011 1823 15017
rect 1765 14977 1777 15011
rect 1811 15008 1823 15011
rect 6546 15008 6552 15020
rect 1811 14980 6552 15008
rect 1811 14977 1823 14980
rect 1765 14971 1823 14977
rect 6546 14968 6552 14980
rect 6604 14968 6610 15020
rect 12253 15011 12311 15017
rect 12253 15008 12265 15011
rect 11164 14980 12265 15008
rect 11164 14952 11192 14980
rect 12253 14977 12265 14980
rect 12299 14977 12311 15011
rect 12406 15008 12434 15036
rect 12406 14980 12480 15008
rect 12253 14971 12311 14977
rect 1302 14900 1308 14952
rect 1360 14940 1366 14952
rect 2041 14943 2099 14949
rect 2041 14940 2053 14943
rect 1360 14912 2053 14940
rect 1360 14900 1366 14912
rect 2041 14909 2053 14912
rect 2087 14909 2099 14943
rect 2041 14903 2099 14909
rect 10042 14900 10048 14952
rect 10100 14900 10106 14952
rect 11146 14900 11152 14952
rect 11204 14900 11210 14952
rect 11609 14943 11667 14949
rect 11609 14909 11621 14943
rect 11655 14940 11667 14943
rect 12342 14940 12348 14952
rect 11655 14912 12348 14940
rect 11655 14909 11667 14912
rect 11609 14903 11667 14909
rect 12342 14900 12348 14912
rect 12400 14900 12406 14952
rect 12452 14949 12480 14980
rect 12437 14943 12495 14949
rect 12437 14909 12449 14943
rect 12483 14909 12495 14943
rect 12437 14903 12495 14909
rect 11422 14832 11428 14884
rect 11480 14872 11486 14884
rect 11885 14875 11943 14881
rect 11885 14872 11897 14875
rect 11480 14844 11897 14872
rect 11480 14832 11486 14844
rect 11885 14841 11897 14844
rect 11931 14841 11943 14875
rect 11885 14835 11943 14841
rect 11974 14832 11980 14884
rect 12032 14872 12038 14884
rect 12802 14872 12808 14884
rect 12032 14844 12808 14872
rect 12032 14832 12038 14844
rect 12802 14832 12808 14844
rect 12860 14832 12866 14884
rect 9401 14807 9459 14813
rect 9401 14773 9413 14807
rect 9447 14804 9459 14807
rect 10962 14804 10968 14816
rect 9447 14776 10968 14804
rect 9447 14773 9459 14776
rect 9401 14767 9459 14773
rect 10962 14764 10968 14776
rect 11020 14764 11026 14816
rect 11698 14764 11704 14816
rect 11756 14804 11762 14816
rect 12897 14807 12955 14813
rect 12897 14804 12909 14807
rect 11756 14776 12909 14804
rect 11756 14764 11762 14776
rect 12897 14773 12909 14776
rect 12943 14804 12955 14807
rect 12986 14804 12992 14816
rect 12943 14776 12992 14804
rect 12943 14773 12955 14776
rect 12897 14767 12955 14773
rect 12986 14764 12992 14776
rect 13044 14764 13050 14816
rect 13096 14804 13124 15048
rect 13280 15048 13544 15076
rect 13280 15017 13308 15048
rect 13538 15036 13544 15048
rect 13596 15036 13602 15088
rect 13648 15076 13676 15116
rect 14550 15104 14556 15156
rect 14608 15144 14614 15156
rect 15013 15147 15071 15153
rect 15013 15144 15025 15147
rect 14608 15116 15025 15144
rect 14608 15104 14614 15116
rect 15013 15113 15025 15116
rect 15059 15113 15071 15147
rect 15013 15107 15071 15113
rect 13998 15076 14004 15088
rect 13648 15048 14004 15076
rect 13998 15036 14004 15048
rect 14056 15036 14062 15088
rect 13265 15011 13323 15017
rect 13265 14977 13277 15011
rect 13311 14977 13323 15011
rect 13265 14971 13323 14977
rect 13541 14943 13599 14949
rect 13541 14909 13553 14943
rect 13587 14940 13599 14943
rect 13906 14940 13912 14952
rect 13587 14912 13912 14940
rect 13587 14909 13599 14912
rect 13541 14903 13599 14909
rect 13906 14900 13912 14912
rect 13964 14900 13970 14952
rect 15028 14940 15056 15107
rect 15562 15104 15568 15156
rect 15620 15104 15626 15156
rect 15933 15147 15991 15153
rect 15933 15113 15945 15147
rect 15979 15144 15991 15147
rect 18325 15147 18383 15153
rect 18325 15144 18337 15147
rect 15979 15116 18337 15144
rect 15979 15113 15991 15116
rect 15933 15107 15991 15113
rect 18325 15113 18337 15116
rect 18371 15113 18383 15147
rect 18325 15107 18383 15113
rect 18693 15147 18751 15153
rect 18693 15113 18705 15147
rect 18739 15144 18751 15147
rect 19426 15144 19432 15156
rect 18739 15116 19432 15144
rect 18739 15113 18751 15116
rect 18693 15107 18751 15113
rect 19426 15104 19432 15116
rect 19484 15104 19490 15156
rect 19518 15104 19524 15156
rect 19576 15104 19582 15156
rect 19978 15144 19984 15156
rect 19628 15116 19984 15144
rect 15654 15036 15660 15088
rect 15712 15076 15718 15088
rect 16025 15079 16083 15085
rect 16025 15076 16037 15079
rect 15712 15048 16037 15076
rect 15712 15036 15718 15048
rect 16025 15045 16037 15048
rect 16071 15045 16083 15079
rect 16025 15039 16083 15045
rect 16482 15036 16488 15088
rect 16540 15076 16546 15088
rect 19628 15076 19656 15116
rect 19978 15104 19984 15116
rect 20036 15144 20042 15156
rect 21818 15144 21824 15156
rect 20036 15116 21036 15144
rect 20036 15104 20042 15116
rect 16540 15048 19656 15076
rect 19889 15079 19947 15085
rect 16540 15036 16546 15048
rect 19889 15045 19901 15079
rect 19935 15076 19947 15079
rect 20806 15076 20812 15088
rect 19935 15048 20812 15076
rect 19935 15045 19947 15048
rect 19889 15039 19947 15045
rect 20806 15036 20812 15048
rect 20864 15036 20870 15088
rect 17218 14968 17224 15020
rect 17276 14968 17282 15020
rect 18598 15008 18604 15020
rect 17420 14980 18604 15008
rect 16114 14940 16120 14952
rect 15028 14912 16120 14940
rect 16114 14900 16120 14912
rect 16172 14900 16178 14952
rect 16758 14900 16764 14952
rect 16816 14940 16822 14952
rect 17420 14949 17448 14980
rect 18598 14968 18604 14980
rect 18656 14968 18662 15020
rect 18785 15011 18843 15017
rect 18785 14977 18797 15011
rect 18831 15008 18843 15011
rect 19242 15008 19248 15020
rect 18831 14980 19248 15008
rect 18831 14977 18843 14980
rect 18785 14971 18843 14977
rect 17313 14943 17371 14949
rect 17313 14940 17325 14943
rect 16816 14912 17325 14940
rect 16816 14900 16822 14912
rect 17313 14909 17325 14912
rect 17359 14909 17371 14943
rect 17313 14903 17371 14909
rect 17405 14943 17463 14949
rect 17405 14909 17417 14943
rect 17451 14909 17463 14943
rect 17405 14903 17463 14909
rect 18049 14943 18107 14949
rect 18049 14909 18061 14943
rect 18095 14940 18107 14943
rect 18800 14940 18828 14971
rect 19242 14968 19248 14980
rect 19300 14968 19306 15020
rect 19981 15011 20039 15017
rect 19981 14977 19993 15011
rect 20027 15008 20039 15011
rect 20898 15008 20904 15020
rect 20027 14980 20904 15008
rect 20027 14977 20039 14980
rect 19981 14971 20039 14977
rect 20898 14968 20904 14980
rect 20956 14968 20962 15020
rect 21008 15008 21036 15116
rect 21100 15116 21824 15144
rect 21100 15085 21128 15116
rect 21818 15104 21824 15116
rect 21876 15104 21882 15156
rect 22646 15104 22652 15156
rect 22704 15144 22710 15156
rect 22925 15147 22983 15153
rect 22925 15144 22937 15147
rect 22704 15116 22937 15144
rect 22704 15104 22710 15116
rect 22925 15113 22937 15116
rect 22971 15113 22983 15147
rect 22925 15107 22983 15113
rect 23385 15147 23443 15153
rect 23385 15113 23397 15147
rect 23431 15144 23443 15147
rect 23474 15144 23480 15156
rect 23431 15116 23480 15144
rect 23431 15113 23443 15116
rect 23385 15107 23443 15113
rect 23474 15104 23480 15116
rect 23532 15104 23538 15156
rect 23750 15104 23756 15156
rect 23808 15144 23814 15156
rect 24121 15147 24179 15153
rect 24121 15144 24133 15147
rect 23808 15116 24133 15144
rect 23808 15104 23814 15116
rect 24121 15113 24133 15116
rect 24167 15113 24179 15147
rect 24121 15107 24179 15113
rect 24228 15116 29592 15144
rect 21085 15079 21143 15085
rect 21085 15045 21097 15079
rect 21131 15045 21143 15079
rect 21085 15039 21143 15045
rect 21266 15036 21272 15088
rect 21324 15076 21330 15088
rect 24228 15076 24256 15116
rect 21324 15048 24256 15076
rect 21324 15036 21330 15048
rect 25038 15036 25044 15088
rect 25096 15076 25102 15088
rect 25317 15079 25375 15085
rect 25317 15076 25329 15079
rect 25096 15048 25329 15076
rect 25096 15036 25102 15048
rect 25317 15045 25329 15048
rect 25363 15045 25375 15079
rect 25317 15039 25375 15045
rect 26329 15079 26387 15085
rect 26329 15045 26341 15079
rect 26375 15076 26387 15079
rect 26375 15048 27292 15076
rect 26375 15045 26387 15048
rect 26329 15039 26387 15045
rect 21008 14980 21312 15008
rect 18095 14912 18828 14940
rect 18095 14909 18107 14912
rect 18049 14903 18107 14909
rect 15930 14872 15936 14884
rect 14568 14844 15936 14872
rect 14568 14804 14596 14844
rect 15930 14832 15936 14844
rect 15988 14832 15994 14884
rect 16574 14832 16580 14884
rect 16632 14872 16638 14884
rect 17420 14872 17448 14903
rect 18874 14900 18880 14952
rect 18932 14900 18938 14952
rect 20070 14900 20076 14952
rect 20128 14900 20134 14952
rect 20530 14900 20536 14952
rect 20588 14940 20594 14952
rect 21284 14949 21312 14980
rect 23290 14968 23296 15020
rect 23348 14968 23354 15020
rect 24489 15011 24547 15017
rect 24489 14977 24501 15011
rect 24535 15008 24547 15011
rect 25225 15011 25283 15017
rect 25225 15008 25237 15011
rect 24535 14980 25237 15008
rect 24535 14977 24547 14980
rect 24489 14971 24547 14977
rect 25225 14977 25237 14980
rect 25271 15008 25283 15011
rect 25406 15008 25412 15020
rect 25271 14980 25412 15008
rect 25271 14977 25283 14980
rect 25225 14971 25283 14977
rect 25406 14968 25412 14980
rect 25464 14968 25470 15020
rect 25498 14968 25504 15020
rect 25556 15008 25562 15020
rect 26237 15011 26295 15017
rect 26237 15008 26249 15011
rect 25556 14980 26249 15008
rect 25556 14968 25562 14980
rect 26237 14977 26249 14980
rect 26283 15008 26295 15011
rect 26973 15011 27031 15017
rect 26973 15008 26985 15011
rect 26283 14980 26985 15008
rect 26283 14977 26295 14980
rect 26237 14971 26295 14977
rect 26973 14977 26985 14980
rect 27019 15008 27031 15011
rect 27062 15008 27068 15020
rect 27019 14980 27068 15008
rect 27019 14977 27031 14980
rect 26973 14971 27031 14977
rect 27062 14968 27068 14980
rect 27120 14968 27126 15020
rect 21177 14943 21235 14949
rect 21177 14940 21189 14943
rect 20588 14912 21189 14940
rect 20588 14900 20594 14912
rect 21177 14909 21189 14912
rect 21223 14909 21235 14943
rect 21177 14903 21235 14909
rect 21269 14943 21327 14949
rect 21269 14909 21281 14943
rect 21315 14909 21327 14943
rect 21269 14903 21327 14909
rect 23569 14943 23627 14949
rect 23569 14909 23581 14943
rect 23615 14909 23627 14943
rect 23569 14903 23627 14909
rect 16632 14844 17448 14872
rect 16632 14832 16638 14844
rect 17494 14832 17500 14884
rect 17552 14872 17558 14884
rect 20717 14875 20775 14881
rect 20717 14872 20729 14875
rect 17552 14844 20729 14872
rect 17552 14832 17558 14844
rect 20717 14841 20729 14844
rect 20763 14841 20775 14875
rect 21192 14872 21220 14903
rect 21726 14872 21732 14884
rect 21192 14844 21732 14872
rect 20717 14835 20775 14841
rect 21726 14832 21732 14844
rect 21784 14832 21790 14884
rect 13096 14776 14596 14804
rect 15838 14764 15844 14816
rect 15896 14804 15902 14816
rect 16853 14807 16911 14813
rect 16853 14804 16865 14807
rect 15896 14776 16865 14804
rect 15896 14764 15902 14776
rect 16853 14773 16865 14776
rect 16899 14773 16911 14807
rect 16853 14767 16911 14773
rect 17402 14764 17408 14816
rect 17460 14804 17466 14816
rect 19334 14804 19340 14816
rect 17460 14776 19340 14804
rect 17460 14764 17466 14776
rect 19334 14764 19340 14776
rect 19392 14764 19398 14816
rect 19610 14764 19616 14816
rect 19668 14804 19674 14816
rect 19886 14804 19892 14816
rect 19668 14776 19892 14804
rect 19668 14764 19674 14776
rect 19886 14764 19892 14776
rect 19944 14804 19950 14816
rect 22005 14807 22063 14813
rect 22005 14804 22017 14807
rect 19944 14776 22017 14804
rect 19944 14764 19950 14776
rect 22005 14773 22017 14776
rect 22051 14773 22063 14807
rect 23584 14804 23612 14903
rect 24578 14900 24584 14952
rect 24636 14900 24642 14952
rect 24670 14900 24676 14952
rect 24728 14900 24734 14952
rect 24762 14900 24768 14952
rect 24820 14940 24826 14952
rect 26421 14943 26479 14949
rect 24820 14912 25912 14940
rect 24820 14900 24826 14912
rect 24302 14832 24308 14884
rect 24360 14872 24366 14884
rect 25884 14881 25912 14912
rect 26421 14909 26433 14943
rect 26467 14909 26479 14943
rect 26421 14903 26479 14909
rect 25869 14875 25927 14881
rect 24360 14844 25728 14872
rect 24360 14832 24366 14844
rect 25038 14804 25044 14816
rect 23584 14776 25044 14804
rect 22005 14767 22063 14773
rect 25038 14764 25044 14776
rect 25096 14764 25102 14816
rect 25590 14764 25596 14816
rect 25648 14764 25654 14816
rect 25700 14804 25728 14844
rect 25869 14841 25881 14875
rect 25915 14841 25927 14875
rect 25869 14835 25927 14841
rect 26436 14804 26464 14903
rect 27264 14881 27292 15048
rect 27522 15036 27528 15088
rect 27580 15076 27586 15088
rect 27617 15079 27675 15085
rect 27617 15076 27629 15079
rect 27580 15048 27629 15076
rect 27580 15036 27586 15048
rect 27617 15045 27629 15048
rect 27663 15045 27675 15079
rect 28350 15076 28356 15088
rect 27617 15039 27675 15045
rect 28000 15048 28356 15076
rect 28000 15017 28028 15048
rect 28350 15036 28356 15048
rect 28408 15036 28414 15088
rect 29270 15036 29276 15088
rect 29328 15036 29334 15088
rect 29564 15076 29592 15116
rect 29730 15104 29736 15156
rect 29788 15104 29794 15156
rect 30282 15104 30288 15156
rect 30340 15144 30346 15156
rect 30340 15116 30512 15144
rect 30340 15104 30346 15116
rect 30006 15076 30012 15088
rect 29564 15048 30012 15076
rect 30006 15036 30012 15048
rect 30064 15036 30070 15088
rect 30190 15036 30196 15088
rect 30248 15076 30254 15088
rect 30248 15048 30420 15076
rect 30248 15036 30254 15048
rect 27985 15011 28043 15017
rect 27985 14977 27997 15011
rect 28031 14977 28043 15011
rect 27985 14971 28043 14977
rect 27338 14900 27344 14952
rect 27396 14940 27402 14952
rect 28261 14943 28319 14949
rect 28261 14940 28273 14943
rect 27396 14912 28273 14940
rect 27396 14900 27402 14912
rect 28261 14909 28273 14912
rect 28307 14940 28319 14943
rect 29822 14940 29828 14952
rect 28307 14912 29828 14940
rect 28307 14909 28319 14912
rect 28261 14903 28319 14909
rect 29822 14900 29828 14912
rect 29880 14940 29886 14952
rect 29880 14912 30328 14940
rect 29880 14900 29886 14912
rect 27249 14875 27307 14881
rect 27249 14841 27261 14875
rect 27295 14872 27307 14875
rect 27295 14844 28120 14872
rect 27295 14841 27307 14844
rect 27249 14835 27307 14841
rect 25700 14776 26464 14804
rect 26878 14764 26884 14816
rect 26936 14804 26942 14816
rect 27433 14807 27491 14813
rect 27433 14804 27445 14807
rect 26936 14776 27445 14804
rect 26936 14764 26942 14776
rect 27433 14773 27445 14776
rect 27479 14773 27491 14807
rect 28092 14804 28120 14844
rect 28442 14804 28448 14816
rect 28092 14776 28448 14804
rect 27433 14767 27491 14773
rect 28442 14764 28448 14776
rect 28500 14764 28506 14816
rect 29822 14764 29828 14816
rect 29880 14804 29886 14816
rect 30193 14807 30251 14813
rect 30193 14804 30205 14807
rect 29880 14776 30205 14804
rect 29880 14764 29886 14776
rect 30193 14773 30205 14776
rect 30239 14773 30251 14807
rect 30300 14804 30328 14912
rect 30392 14872 30420 15048
rect 30484 14940 30512 15116
rect 30650 15104 30656 15156
rect 30708 15144 30714 15156
rect 30926 15144 30932 15156
rect 30708 15116 30932 15144
rect 30708 15104 30714 15116
rect 30926 15104 30932 15116
rect 30984 15104 30990 15156
rect 31294 15104 31300 15156
rect 31352 15144 31358 15156
rect 31389 15147 31447 15153
rect 31389 15144 31401 15147
rect 31352 15116 31401 15144
rect 31352 15104 31358 15116
rect 31389 15113 31401 15116
rect 31435 15113 31447 15147
rect 31389 15107 31447 15113
rect 31570 15104 31576 15156
rect 31628 15144 31634 15156
rect 32677 15147 32735 15153
rect 32677 15144 32689 15147
rect 31628 15116 32689 15144
rect 31628 15104 31634 15116
rect 32677 15113 32689 15116
rect 32723 15113 32735 15147
rect 32677 15107 32735 15113
rect 33870 15104 33876 15156
rect 33928 15104 33934 15156
rect 34698 15104 34704 15156
rect 34756 15104 34762 15156
rect 35069 15147 35127 15153
rect 35069 15113 35081 15147
rect 35115 15144 35127 15147
rect 37274 15144 37280 15156
rect 35115 15116 37280 15144
rect 35115 15113 35127 15116
rect 35069 15107 35127 15113
rect 37274 15104 37280 15116
rect 37332 15104 37338 15156
rect 37660 15116 37872 15144
rect 30561 15079 30619 15085
rect 30561 15045 30573 15079
rect 30607 15076 30619 15079
rect 31478 15076 31484 15088
rect 30607 15048 31484 15076
rect 30607 15045 30619 15048
rect 30561 15039 30619 15045
rect 31478 15036 31484 15048
rect 31536 15036 31542 15088
rect 31849 15079 31907 15085
rect 31849 15076 31861 15079
rect 31726 15048 31861 15076
rect 30926 14968 30932 15020
rect 30984 15008 30990 15020
rect 31726 15008 31754 15048
rect 31849 15045 31861 15048
rect 31895 15045 31907 15079
rect 31849 15039 31907 15045
rect 32769 15079 32827 15085
rect 32769 15045 32781 15079
rect 32815 15076 32827 15079
rect 37182 15076 37188 15088
rect 32815 15048 37188 15076
rect 32815 15045 32827 15048
rect 32769 15039 32827 15045
rect 37182 15036 37188 15048
rect 37240 15036 37246 15088
rect 37660 15076 37688 15116
rect 37844 15088 37872 15116
rect 38562 15104 38568 15156
rect 38620 15144 38626 15156
rect 39669 15147 39727 15153
rect 39669 15144 39681 15147
rect 38620 15116 39681 15144
rect 38620 15104 38626 15116
rect 39669 15113 39681 15116
rect 39715 15113 39727 15147
rect 39669 15107 39727 15113
rect 40126 15104 40132 15156
rect 40184 15104 40190 15156
rect 40310 15104 40316 15156
rect 40368 15144 40374 15156
rect 49237 15147 49295 15153
rect 49237 15144 49249 15147
rect 40368 15116 49249 15144
rect 40368 15104 40374 15116
rect 49237 15113 49249 15116
rect 49283 15113 49295 15147
rect 49237 15107 49295 15113
rect 37292 15048 37688 15076
rect 30984 14980 31754 15008
rect 30984 14968 30990 14980
rect 35894 14968 35900 15020
rect 35952 14968 35958 15020
rect 36170 14968 36176 15020
rect 36228 15008 36234 15020
rect 36265 15011 36323 15017
rect 36265 15008 36277 15011
rect 36228 14980 36277 15008
rect 36228 14968 36234 14980
rect 36265 14977 36277 14980
rect 36311 14977 36323 15011
rect 36265 14971 36323 14977
rect 36446 14968 36452 15020
rect 36504 15008 36510 15020
rect 36909 15011 36967 15017
rect 36909 15008 36921 15011
rect 36504 14980 36921 15008
rect 36504 14968 36510 14980
rect 36909 14977 36921 14980
rect 36955 15008 36967 15011
rect 37292 15008 37320 15048
rect 37826 15036 37832 15088
rect 37884 15076 37890 15088
rect 40037 15079 40095 15085
rect 37884 15048 38226 15076
rect 37884 15036 37890 15048
rect 40037 15045 40049 15079
rect 40083 15076 40095 15079
rect 48406 15076 48412 15088
rect 40083 15048 48412 15076
rect 40083 15045 40095 15048
rect 40037 15039 40095 15045
rect 48406 15036 48412 15048
rect 48464 15036 48470 15088
rect 36955 14980 37320 15008
rect 36955 14977 36967 14980
rect 36909 14971 36967 14977
rect 37458 14968 37464 15020
rect 37516 14968 37522 15020
rect 39850 14968 39856 15020
rect 39908 15008 39914 15020
rect 41049 15011 41107 15017
rect 41049 15008 41061 15011
rect 39908 14980 41061 15008
rect 39908 14968 39914 14980
rect 41049 14977 41061 14980
rect 41095 14977 41107 15011
rect 41049 14971 41107 14977
rect 48777 15011 48835 15017
rect 48777 14977 48789 15011
rect 48823 15008 48835 15011
rect 49050 15008 49056 15020
rect 48823 14980 49056 15008
rect 48823 14977 48835 14980
rect 48777 14971 48835 14977
rect 49050 14968 49056 14980
rect 49108 14968 49114 15020
rect 30745 14943 30803 14949
rect 30745 14940 30757 14943
rect 30484 14912 30757 14940
rect 30745 14909 30757 14912
rect 30791 14909 30803 14943
rect 30745 14903 30803 14909
rect 30834 14900 30840 14952
rect 30892 14940 30898 14952
rect 32953 14943 33011 14949
rect 32953 14940 32965 14943
rect 30892 14912 32965 14940
rect 30892 14900 30898 14912
rect 32953 14909 32965 14912
rect 32999 14940 33011 14943
rect 33870 14940 33876 14952
rect 32999 14912 33876 14940
rect 32999 14909 33011 14912
rect 32953 14903 33011 14909
rect 33870 14900 33876 14912
rect 33928 14900 33934 14952
rect 33962 14900 33968 14952
rect 34020 14900 34026 14952
rect 34054 14900 34060 14952
rect 34112 14900 34118 14952
rect 34606 14900 34612 14952
rect 34664 14940 34670 14952
rect 35161 14943 35219 14949
rect 35161 14940 35173 14943
rect 34664 14912 35173 14940
rect 34664 14900 34670 14912
rect 35161 14909 35173 14912
rect 35207 14909 35219 14943
rect 35161 14903 35219 14909
rect 35342 14900 35348 14952
rect 35400 14900 35406 14952
rect 35912 14940 35940 14968
rect 36357 14943 36415 14949
rect 36357 14940 36369 14943
rect 35912 14912 36369 14940
rect 36357 14909 36369 14912
rect 36403 14909 36415 14943
rect 36357 14903 36415 14909
rect 36538 14900 36544 14952
rect 36596 14900 36602 14952
rect 36998 14900 37004 14952
rect 37056 14940 37062 14952
rect 37737 14943 37795 14949
rect 37737 14940 37749 14943
rect 37056 14912 37749 14940
rect 37056 14900 37062 14912
rect 37737 14909 37749 14912
rect 37783 14909 37795 14943
rect 37737 14903 37795 14909
rect 38470 14900 38476 14952
rect 38528 14940 38534 14952
rect 38528 14912 38792 14940
rect 38528 14900 38534 14912
rect 32309 14875 32367 14881
rect 32309 14872 32321 14875
rect 30392 14844 32321 14872
rect 32309 14841 32321 14844
rect 32355 14841 32367 14875
rect 32309 14835 32367 14841
rect 35897 14875 35955 14881
rect 35897 14841 35909 14875
rect 35943 14872 35955 14875
rect 37274 14872 37280 14884
rect 35943 14844 37280 14872
rect 35943 14841 35955 14844
rect 35897 14835 35955 14841
rect 37274 14832 37280 14844
rect 37332 14832 37338 14884
rect 38764 14872 38792 14912
rect 38930 14900 38936 14952
rect 38988 14940 38994 14952
rect 40221 14943 40279 14949
rect 40221 14940 40233 14943
rect 38988 14912 40233 14940
rect 38988 14900 38994 14912
rect 40221 14909 40233 14912
rect 40267 14909 40279 14943
rect 40221 14903 40279 14909
rect 40310 14872 40316 14884
rect 38764 14844 40316 14872
rect 40310 14832 40316 14844
rect 40368 14832 40374 14884
rect 32766 14804 32772 14816
rect 30300 14776 32772 14804
rect 30193 14767 30251 14773
rect 32766 14764 32772 14776
rect 32824 14764 32830 14816
rect 33505 14807 33563 14813
rect 33505 14773 33517 14807
rect 33551 14804 33563 14807
rect 36722 14804 36728 14816
rect 33551 14776 36728 14804
rect 33551 14773 33563 14776
rect 33505 14767 33563 14773
rect 36722 14764 36728 14776
rect 36780 14764 36786 14816
rect 37550 14764 37556 14816
rect 37608 14804 37614 14816
rect 39209 14807 39267 14813
rect 39209 14804 39221 14807
rect 37608 14776 39221 14804
rect 37608 14764 37614 14776
rect 39209 14773 39221 14776
rect 39255 14773 39267 14807
rect 39209 14767 39267 14773
rect 40865 14807 40923 14813
rect 40865 14773 40877 14807
rect 40911 14804 40923 14807
rect 45830 14804 45836 14816
rect 40911 14776 45836 14804
rect 40911 14773 40923 14776
rect 40865 14767 40923 14773
rect 45830 14764 45836 14776
rect 45888 14764 45894 14816
rect 1104 14714 49864 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 32950 14714
rect 33002 14662 33014 14714
rect 33066 14662 33078 14714
rect 33130 14662 33142 14714
rect 33194 14662 33206 14714
rect 33258 14662 42950 14714
rect 43002 14662 43014 14714
rect 43066 14662 43078 14714
rect 43130 14662 43142 14714
rect 43194 14662 43206 14714
rect 43258 14662 49864 14714
rect 1104 14640 49864 14662
rect 10410 14560 10416 14612
rect 10468 14560 10474 14612
rect 11606 14560 11612 14612
rect 11664 14600 11670 14612
rect 11793 14603 11851 14609
rect 11793 14600 11805 14603
rect 11664 14572 11805 14600
rect 11664 14560 11670 14572
rect 11793 14569 11805 14572
rect 11839 14569 11851 14603
rect 11793 14563 11851 14569
rect 12618 14560 12624 14612
rect 12676 14600 12682 14612
rect 12989 14603 13047 14609
rect 12989 14600 13001 14603
rect 12676 14572 13001 14600
rect 12676 14560 12682 14572
rect 12989 14569 13001 14572
rect 13035 14569 13047 14603
rect 12989 14563 13047 14569
rect 13170 14560 13176 14612
rect 13228 14600 13234 14612
rect 17126 14600 17132 14612
rect 13228 14572 17132 14600
rect 13228 14560 13234 14572
rect 17126 14560 17132 14572
rect 17184 14560 17190 14612
rect 17218 14560 17224 14612
rect 17276 14600 17282 14612
rect 17681 14603 17739 14609
rect 17681 14600 17693 14603
rect 17276 14572 17693 14600
rect 17276 14560 17282 14572
rect 17681 14569 17693 14572
rect 17727 14569 17739 14603
rect 17681 14563 17739 14569
rect 17862 14560 17868 14612
rect 17920 14600 17926 14612
rect 18141 14603 18199 14609
rect 18141 14600 18153 14603
rect 17920 14572 18153 14600
rect 17920 14560 17926 14572
rect 18141 14569 18153 14572
rect 18187 14569 18199 14603
rect 18141 14563 18199 14569
rect 18598 14560 18604 14612
rect 18656 14600 18662 14612
rect 18656 14572 19012 14600
rect 18656 14560 18662 14572
rect 13262 14532 13268 14544
rect 12360 14504 13268 14532
rect 1302 14424 1308 14476
rect 1360 14464 1366 14476
rect 12360 14473 12388 14504
rect 13262 14492 13268 14504
rect 13320 14492 13326 14544
rect 14458 14492 14464 14544
rect 14516 14492 14522 14544
rect 14918 14492 14924 14544
rect 14976 14532 14982 14544
rect 18874 14532 18880 14544
rect 14976 14504 18880 14532
rect 14976 14492 14982 14504
rect 18874 14492 18880 14504
rect 18932 14492 18938 14544
rect 2041 14467 2099 14473
rect 2041 14464 2053 14467
rect 1360 14436 2053 14464
rect 1360 14424 1366 14436
rect 2041 14433 2053 14436
rect 2087 14433 2099 14467
rect 2041 14427 2099 14433
rect 12345 14467 12403 14473
rect 12345 14433 12357 14467
rect 12391 14433 12403 14467
rect 12345 14427 12403 14433
rect 12526 14424 12532 14476
rect 12584 14464 12590 14476
rect 13541 14467 13599 14473
rect 13541 14464 13553 14467
rect 12584 14436 13553 14464
rect 12584 14424 12590 14436
rect 13541 14433 13553 14436
rect 13587 14433 13599 14467
rect 15013 14467 15071 14473
rect 15013 14464 15025 14467
rect 13541 14427 13599 14433
rect 14108 14436 15025 14464
rect 1765 14399 1823 14405
rect 1765 14365 1777 14399
rect 1811 14396 1823 14399
rect 9769 14399 9827 14405
rect 9769 14396 9781 14399
rect 1811 14368 9781 14396
rect 1811 14365 1823 14368
rect 1765 14359 1823 14365
rect 9769 14365 9781 14368
rect 9815 14365 9827 14399
rect 9769 14359 9827 14365
rect 10318 14356 10324 14408
rect 10376 14356 10382 14408
rect 10686 14356 10692 14408
rect 10744 14396 10750 14408
rect 11149 14399 11207 14405
rect 11149 14396 11161 14399
rect 10744 14368 11161 14396
rect 10744 14356 10750 14368
rect 11149 14365 11161 14368
rect 11195 14396 11207 14399
rect 11195 14368 12756 14396
rect 11195 14365 11207 14368
rect 11149 14359 11207 14365
rect 9582 14288 9588 14340
rect 9640 14288 9646 14340
rect 12161 14331 12219 14337
rect 12161 14297 12173 14331
rect 12207 14328 12219 14331
rect 12526 14328 12532 14340
rect 12207 14300 12532 14328
rect 12207 14297 12219 14300
rect 12161 14291 12219 14297
rect 12526 14288 12532 14300
rect 12584 14288 12590 14340
rect 12728 14328 12756 14368
rect 12802 14356 12808 14408
rect 12860 14396 12866 14408
rect 14108 14396 14136 14436
rect 15013 14433 15025 14436
rect 15059 14433 15071 14467
rect 15013 14427 15071 14433
rect 12860 14368 14136 14396
rect 12860 14356 12866 14368
rect 14182 14356 14188 14408
rect 14240 14396 14246 14408
rect 14921 14399 14979 14405
rect 14921 14396 14933 14399
rect 14240 14368 14933 14396
rect 14240 14356 14246 14368
rect 14921 14365 14933 14368
rect 14967 14365 14979 14399
rect 15028 14396 15056 14427
rect 16114 14424 16120 14476
rect 16172 14464 16178 14476
rect 16945 14467 17003 14473
rect 16945 14464 16957 14467
rect 16172 14436 16957 14464
rect 16172 14424 16178 14436
rect 16945 14433 16957 14436
rect 16991 14433 17003 14467
rect 16945 14427 17003 14433
rect 17126 14424 17132 14476
rect 17184 14464 17190 14476
rect 17586 14464 17592 14476
rect 17184 14436 17592 14464
rect 17184 14424 17190 14436
rect 17586 14424 17592 14436
rect 17644 14424 17650 14476
rect 18693 14467 18751 14473
rect 18693 14433 18705 14467
rect 18739 14433 18751 14467
rect 18984 14464 19012 14572
rect 19058 14560 19064 14612
rect 19116 14600 19122 14612
rect 21082 14600 21088 14612
rect 19116 14572 21088 14600
rect 19116 14560 19122 14572
rect 21082 14560 21088 14572
rect 21140 14560 21146 14612
rect 21450 14560 21456 14612
rect 21508 14600 21514 14612
rect 22833 14603 22891 14609
rect 22833 14600 22845 14603
rect 21508 14572 22845 14600
rect 21508 14560 21514 14572
rect 22833 14569 22845 14572
rect 22879 14569 22891 14603
rect 22833 14563 22891 14569
rect 23198 14560 23204 14612
rect 23256 14600 23262 14612
rect 23293 14603 23351 14609
rect 23293 14600 23305 14603
rect 23256 14572 23305 14600
rect 23256 14560 23262 14572
rect 23293 14569 23305 14572
rect 23339 14600 23351 14603
rect 23569 14603 23627 14609
rect 23569 14600 23581 14603
rect 23339 14572 23581 14600
rect 23339 14569 23351 14572
rect 23293 14563 23351 14569
rect 23569 14569 23581 14572
rect 23615 14600 23627 14603
rect 24026 14600 24032 14612
rect 23615 14572 24032 14600
rect 23615 14569 23627 14572
rect 23569 14563 23627 14569
rect 24026 14560 24032 14572
rect 24084 14560 24090 14612
rect 25130 14560 25136 14612
rect 25188 14600 25194 14612
rect 27341 14603 27399 14609
rect 27341 14600 27353 14603
rect 25188 14572 27353 14600
rect 25188 14560 25194 14572
rect 27341 14569 27353 14572
rect 27387 14569 27399 14603
rect 27341 14563 27399 14569
rect 29733 14603 29791 14609
rect 29733 14569 29745 14603
rect 29779 14600 29791 14603
rect 33962 14600 33968 14612
rect 29779 14572 33968 14600
rect 29779 14569 29791 14572
rect 29733 14563 29791 14569
rect 33962 14560 33968 14572
rect 34020 14560 34026 14612
rect 35342 14560 35348 14612
rect 35400 14600 35406 14612
rect 35400 14572 36584 14600
rect 35400 14560 35406 14572
rect 24578 14492 24584 14544
rect 24636 14532 24642 14544
rect 25498 14532 25504 14544
rect 24636 14504 25504 14532
rect 24636 14492 24642 14504
rect 25498 14492 25504 14504
rect 25556 14492 25562 14544
rect 27801 14535 27859 14541
rect 27801 14501 27813 14535
rect 27847 14532 27859 14535
rect 27847 14504 30328 14532
rect 27847 14501 27859 14504
rect 27801 14495 27859 14501
rect 20073 14467 20131 14473
rect 20073 14464 20085 14467
rect 18984 14436 20085 14464
rect 18693 14427 18751 14433
rect 20073 14433 20085 14436
rect 20119 14433 20131 14467
rect 20073 14427 20131 14433
rect 17310 14396 17316 14408
rect 15028 14368 17316 14396
rect 14921 14359 14979 14365
rect 17310 14356 17316 14368
rect 17368 14396 17374 14408
rect 18708 14396 18736 14427
rect 20714 14424 20720 14476
rect 20772 14464 20778 14476
rect 21085 14467 21143 14473
rect 21085 14464 21097 14467
rect 20772 14436 21097 14464
rect 20772 14424 20778 14436
rect 21085 14433 21097 14436
rect 21131 14433 21143 14467
rect 21085 14427 21143 14433
rect 21358 14424 21364 14476
rect 21416 14424 21422 14476
rect 21726 14424 21732 14476
rect 21784 14464 21790 14476
rect 21784 14436 23704 14464
rect 21784 14424 21790 14436
rect 23676 14396 23704 14436
rect 24854 14424 24860 14476
rect 24912 14464 24918 14476
rect 25593 14467 25651 14473
rect 25593 14464 25605 14467
rect 24912 14436 25605 14464
rect 24912 14424 24918 14436
rect 25593 14433 25605 14436
rect 25639 14464 25651 14467
rect 27154 14464 27160 14476
rect 25639 14436 27160 14464
rect 25639 14433 25651 14436
rect 25593 14427 25651 14433
rect 27154 14424 27160 14436
rect 27212 14424 27218 14476
rect 27522 14424 27528 14476
rect 27580 14464 27586 14476
rect 28258 14464 28264 14476
rect 27580 14436 28264 14464
rect 27580 14424 27586 14436
rect 28258 14424 28264 14436
rect 28316 14424 28322 14476
rect 28445 14467 28503 14473
rect 28445 14433 28457 14467
rect 28491 14464 28503 14467
rect 28626 14464 28632 14476
rect 28491 14436 28632 14464
rect 28491 14433 28503 14436
rect 28445 14427 28503 14433
rect 28626 14424 28632 14436
rect 28684 14424 28690 14476
rect 25314 14396 25320 14408
rect 17368 14368 18736 14396
rect 19306 14368 21128 14396
rect 23676 14368 25320 14396
rect 17368 14356 17374 14368
rect 13170 14328 13176 14340
rect 12728 14300 13176 14328
rect 13170 14288 13176 14300
rect 13228 14288 13234 14340
rect 13357 14331 13415 14337
rect 13357 14297 13369 14331
rect 13403 14328 13415 14331
rect 15749 14331 15807 14337
rect 13403 14300 15056 14328
rect 13403 14297 13415 14300
rect 13357 14291 13415 14297
rect 11238 14220 11244 14272
rect 11296 14220 11302 14272
rect 12253 14263 12311 14269
rect 12253 14229 12265 14263
rect 12299 14260 12311 14263
rect 12618 14260 12624 14272
rect 12299 14232 12624 14260
rect 12299 14229 12311 14232
rect 12253 14223 12311 14229
rect 12618 14220 12624 14232
rect 12676 14220 12682 14272
rect 13446 14220 13452 14272
rect 13504 14220 13510 14272
rect 13722 14220 13728 14272
rect 13780 14260 13786 14272
rect 14829 14263 14887 14269
rect 14829 14260 14841 14263
rect 13780 14232 14841 14260
rect 13780 14220 13786 14232
rect 14829 14229 14841 14232
rect 14875 14229 14887 14263
rect 15028 14260 15056 14300
rect 15749 14297 15761 14331
rect 15795 14328 15807 14331
rect 16761 14331 16819 14337
rect 16761 14328 16773 14331
rect 15795 14300 16773 14328
rect 15795 14297 15807 14300
rect 15749 14291 15807 14297
rect 16761 14297 16773 14300
rect 16807 14297 16819 14331
rect 18601 14331 18659 14337
rect 18601 14328 18613 14331
rect 16761 14291 16819 14297
rect 17512 14300 18613 14328
rect 16393 14263 16451 14269
rect 16393 14260 16405 14263
rect 15028 14232 16405 14260
rect 14829 14223 14887 14229
rect 16393 14229 16405 14232
rect 16439 14229 16451 14263
rect 16393 14223 16451 14229
rect 16482 14220 16488 14272
rect 16540 14260 16546 14272
rect 16853 14263 16911 14269
rect 16853 14260 16865 14263
rect 16540 14232 16865 14260
rect 16540 14220 16546 14232
rect 16853 14229 16865 14232
rect 16899 14229 16911 14263
rect 16853 14223 16911 14229
rect 16942 14220 16948 14272
rect 17000 14260 17006 14272
rect 17512 14269 17540 14300
rect 18601 14297 18613 14300
rect 18647 14328 18659 14331
rect 19306 14328 19334 14368
rect 18647 14300 19334 14328
rect 18647 14297 18659 14300
rect 18601 14291 18659 14297
rect 19886 14288 19892 14340
rect 19944 14288 19950 14340
rect 21100 14328 21128 14368
rect 25314 14356 25320 14368
rect 25372 14356 25378 14408
rect 30101 14399 30159 14405
rect 30101 14365 30113 14399
rect 30147 14396 30159 14399
rect 30300 14396 30328 14504
rect 30392 14504 31892 14532
rect 30392 14473 30420 14504
rect 30377 14467 30435 14473
rect 30377 14433 30389 14467
rect 30423 14433 30435 14467
rect 30377 14427 30435 14433
rect 30742 14424 30748 14476
rect 30800 14464 30806 14476
rect 31481 14467 31539 14473
rect 31481 14464 31493 14467
rect 30800 14436 31493 14464
rect 30800 14424 30806 14436
rect 31481 14433 31493 14436
rect 31527 14433 31539 14467
rect 31864 14464 31892 14504
rect 31938 14492 31944 14544
rect 31996 14532 32002 14544
rect 31996 14504 32720 14532
rect 31996 14492 32002 14504
rect 32122 14464 32128 14476
rect 31864 14436 32128 14464
rect 31481 14427 31539 14433
rect 32122 14424 32128 14436
rect 32180 14424 32186 14476
rect 32490 14424 32496 14476
rect 32548 14464 32554 14476
rect 32692 14473 32720 14504
rect 32858 14492 32864 14544
rect 32916 14532 32922 14544
rect 36556 14532 36584 14572
rect 36630 14560 36636 14612
rect 36688 14560 36694 14612
rect 38102 14600 38108 14612
rect 37200 14572 38108 14600
rect 37200 14532 37228 14572
rect 38102 14560 38108 14572
rect 38160 14560 38166 14612
rect 38378 14560 38384 14612
rect 38436 14600 38442 14612
rect 38841 14603 38899 14609
rect 38841 14600 38853 14603
rect 38436 14572 38853 14600
rect 38436 14560 38442 14572
rect 38841 14569 38853 14572
rect 38887 14600 38899 14603
rect 38930 14600 38936 14612
rect 38887 14572 38936 14600
rect 38887 14569 38899 14572
rect 38841 14563 38899 14569
rect 38930 14560 38936 14572
rect 38988 14560 38994 14612
rect 39758 14560 39764 14612
rect 39816 14600 39822 14612
rect 39853 14603 39911 14609
rect 39853 14600 39865 14603
rect 39816 14572 39865 14600
rect 39816 14560 39822 14572
rect 39853 14569 39865 14572
rect 39899 14600 39911 14603
rect 40037 14603 40095 14609
rect 40037 14600 40049 14603
rect 39899 14572 40049 14600
rect 39899 14569 39911 14572
rect 39853 14563 39911 14569
rect 40037 14569 40049 14572
rect 40083 14569 40095 14603
rect 40037 14563 40095 14569
rect 32916 14504 34008 14532
rect 36556 14504 37228 14532
rect 32916 14492 32922 14504
rect 32585 14467 32643 14473
rect 32585 14464 32597 14467
rect 32548 14436 32597 14464
rect 32548 14424 32554 14436
rect 32585 14433 32597 14436
rect 32631 14433 32643 14467
rect 32585 14427 32643 14433
rect 32677 14467 32735 14473
rect 32677 14433 32689 14467
rect 32723 14433 32735 14467
rect 33873 14467 33931 14473
rect 33873 14464 33885 14467
rect 32677 14427 32735 14433
rect 32784 14436 33885 14464
rect 31389 14399 31447 14405
rect 31389 14396 31401 14399
rect 30147 14368 30236 14396
rect 30300 14368 31401 14396
rect 30147 14365 30159 14368
rect 30101 14359 30159 14365
rect 21266 14328 21272 14340
rect 21100 14300 21272 14328
rect 21266 14288 21272 14300
rect 21324 14288 21330 14340
rect 22646 14328 22652 14340
rect 22586 14300 22652 14328
rect 22646 14288 22652 14300
rect 22704 14328 22710 14340
rect 23198 14328 23204 14340
rect 22704 14300 23204 14328
rect 22704 14288 22710 14300
rect 23198 14288 23204 14300
rect 23256 14288 23262 14340
rect 25498 14328 25504 14340
rect 23584 14300 25504 14328
rect 17497 14263 17555 14269
rect 17497 14260 17509 14263
rect 17000 14232 17509 14260
rect 17000 14220 17006 14232
rect 17497 14229 17509 14232
rect 17543 14229 17555 14263
rect 17497 14223 17555 14229
rect 18506 14220 18512 14272
rect 18564 14220 18570 14272
rect 19518 14220 19524 14272
rect 19576 14220 19582 14272
rect 19794 14220 19800 14272
rect 19852 14260 19858 14272
rect 19981 14263 20039 14269
rect 19981 14260 19993 14263
rect 19852 14232 19993 14260
rect 19852 14220 19858 14232
rect 19981 14229 19993 14232
rect 20027 14229 20039 14263
rect 19981 14223 20039 14229
rect 20530 14220 20536 14272
rect 20588 14220 20594 14272
rect 20714 14220 20720 14272
rect 20772 14220 20778 14272
rect 22370 14220 22376 14272
rect 22428 14260 22434 14272
rect 23584 14260 23612 14300
rect 25498 14288 25504 14300
rect 25556 14288 25562 14340
rect 25876 14331 25934 14337
rect 25876 14297 25888 14331
rect 25922 14297 25934 14331
rect 25876 14291 25934 14297
rect 22428 14232 23612 14260
rect 22428 14220 22434 14232
rect 23658 14220 23664 14272
rect 23716 14260 23722 14272
rect 23845 14263 23903 14269
rect 23845 14260 23857 14263
rect 23716 14232 23857 14260
rect 23716 14220 23722 14232
rect 23845 14229 23857 14232
rect 23891 14229 23903 14263
rect 23845 14223 23903 14229
rect 24394 14220 24400 14272
rect 24452 14220 24458 14272
rect 24578 14220 24584 14272
rect 24636 14220 24642 14272
rect 24946 14220 24952 14272
rect 25004 14220 25010 14272
rect 25884 14260 25912 14291
rect 26878 14288 26884 14340
rect 26936 14288 26942 14340
rect 28169 14331 28227 14337
rect 28169 14297 28181 14331
rect 28215 14328 28227 14331
rect 28442 14328 28448 14340
rect 28215 14300 28448 14328
rect 28215 14297 28227 14300
rect 28169 14291 28227 14297
rect 28442 14288 28448 14300
rect 28500 14288 28506 14340
rect 28534 14288 28540 14340
rect 28592 14328 28598 14340
rect 29730 14328 29736 14340
rect 28592 14300 29736 14328
rect 28592 14288 28598 14300
rect 29730 14288 29736 14300
rect 29788 14288 29794 14340
rect 30208 14328 30236 14368
rect 31389 14365 31401 14368
rect 31435 14365 31447 14399
rect 31389 14359 31447 14365
rect 31754 14356 31760 14408
rect 31812 14396 31818 14408
rect 32784 14396 32812 14436
rect 33873 14433 33885 14436
rect 33919 14433 33931 14467
rect 33873 14427 33931 14433
rect 31812 14368 32812 14396
rect 31812 14356 31818 14368
rect 33410 14356 33416 14408
rect 33468 14396 33474 14408
rect 33689 14399 33747 14405
rect 33689 14396 33701 14399
rect 33468 14368 33701 14396
rect 33468 14356 33474 14368
rect 33689 14365 33701 14368
rect 33735 14365 33747 14399
rect 33689 14359 33747 14365
rect 33781 14399 33839 14405
rect 33781 14365 33793 14399
rect 33827 14396 33839 14399
rect 33980 14396 34008 14504
rect 34882 14424 34888 14476
rect 34940 14464 34946 14476
rect 37093 14467 37151 14473
rect 37093 14464 37105 14467
rect 34940 14436 37105 14464
rect 34940 14424 34946 14436
rect 37093 14433 37105 14436
rect 37139 14464 37151 14467
rect 37458 14464 37464 14476
rect 37139 14436 37464 14464
rect 37139 14433 37151 14436
rect 37093 14427 37151 14433
rect 37458 14424 37464 14436
rect 37516 14424 37522 14476
rect 37734 14424 37740 14476
rect 37792 14464 37798 14476
rect 49329 14467 49387 14473
rect 49329 14464 49341 14467
rect 37792 14436 39528 14464
rect 37792 14424 37798 14436
rect 39500 14405 39528 14436
rect 41386 14436 49341 14464
rect 33827 14368 34008 14396
rect 39485 14399 39543 14405
rect 33827 14365 33839 14368
rect 33781 14359 33839 14365
rect 39485 14365 39497 14399
rect 39531 14365 39543 14399
rect 39485 14359 39543 14365
rect 39574 14356 39580 14408
rect 39632 14396 39638 14408
rect 41386 14396 41414 14436
rect 49329 14433 49341 14436
rect 49375 14433 49387 14467
rect 49329 14427 49387 14433
rect 39632 14368 41414 14396
rect 48593 14399 48651 14405
rect 39632 14356 39638 14368
rect 48593 14365 48605 14399
rect 48639 14396 48651 14399
rect 49142 14396 49148 14408
rect 48639 14368 49148 14396
rect 48639 14365 48651 14368
rect 48593 14359 48651 14365
rect 49142 14356 49148 14368
rect 49200 14356 49206 14408
rect 30374 14328 30380 14340
rect 30208 14300 30380 14328
rect 30374 14288 30380 14300
rect 30432 14288 30438 14340
rect 32493 14331 32551 14337
rect 30944 14300 32260 14328
rect 25958 14260 25964 14272
rect 25884 14232 25964 14260
rect 25958 14220 25964 14232
rect 26016 14260 26022 14272
rect 28552 14260 28580 14288
rect 26016 14232 28580 14260
rect 26016 14220 26022 14232
rect 28994 14220 29000 14272
rect 29052 14220 29058 14272
rect 29546 14220 29552 14272
rect 29604 14260 29610 14272
rect 30944 14269 30972 14300
rect 30193 14263 30251 14269
rect 30193 14260 30205 14263
rect 29604 14232 30205 14260
rect 29604 14220 29610 14232
rect 30193 14229 30205 14232
rect 30239 14229 30251 14263
rect 30193 14223 30251 14229
rect 30929 14263 30987 14269
rect 30929 14229 30941 14263
rect 30975 14229 30987 14263
rect 30929 14223 30987 14229
rect 31110 14220 31116 14272
rect 31168 14260 31174 14272
rect 31297 14263 31355 14269
rect 31297 14260 31309 14263
rect 31168 14232 31309 14260
rect 31168 14220 31174 14232
rect 31297 14229 31309 14232
rect 31343 14229 31355 14263
rect 31297 14223 31355 14229
rect 32122 14220 32128 14272
rect 32180 14220 32186 14272
rect 32232 14260 32260 14300
rect 32493 14297 32505 14331
rect 32539 14328 32551 14331
rect 33594 14328 33600 14340
rect 32539 14300 33600 14328
rect 32539 14297 32551 14300
rect 32493 14291 32551 14297
rect 33594 14288 33600 14300
rect 33652 14288 33658 14340
rect 34440 14300 35112 14328
rect 33226 14260 33232 14272
rect 32232 14232 33232 14260
rect 33226 14220 33232 14232
rect 33284 14220 33290 14272
rect 33321 14263 33379 14269
rect 33321 14229 33333 14263
rect 33367 14260 33379 14263
rect 34440 14260 34468 14300
rect 33367 14232 34468 14260
rect 34517 14263 34575 14269
rect 33367 14229 33379 14232
rect 33321 14223 33379 14229
rect 34517 14229 34529 14263
rect 34563 14260 34575 14263
rect 34606 14260 34612 14272
rect 34563 14232 34612 14260
rect 34563 14229 34575 14232
rect 34517 14223 34575 14229
rect 34606 14220 34612 14232
rect 34664 14220 34670 14272
rect 35084 14260 35112 14300
rect 35158 14288 35164 14340
rect 35216 14288 35222 14340
rect 36446 14328 36452 14340
rect 36386 14300 36452 14328
rect 36446 14288 36452 14300
rect 36504 14288 36510 14340
rect 37369 14331 37427 14337
rect 37369 14297 37381 14331
rect 37415 14328 37427 14331
rect 37458 14328 37464 14340
rect 37415 14300 37464 14328
rect 37415 14297 37427 14300
rect 37369 14291 37427 14297
rect 37458 14288 37464 14300
rect 37516 14288 37522 14340
rect 37826 14288 37832 14340
rect 37884 14288 37890 14340
rect 37550 14260 37556 14272
rect 35084 14232 37556 14260
rect 37550 14220 37556 14232
rect 37608 14220 37614 14272
rect 39298 14220 39304 14272
rect 39356 14220 39362 14272
rect 48314 14220 48320 14272
rect 48372 14260 48378 14272
rect 48685 14263 48743 14269
rect 48685 14260 48697 14263
rect 48372 14232 48697 14260
rect 48372 14220 48378 14232
rect 48685 14229 48697 14232
rect 48731 14229 48743 14263
rect 48685 14223 48743 14229
rect 1104 14170 49864 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 27950 14170
rect 28002 14118 28014 14170
rect 28066 14118 28078 14170
rect 28130 14118 28142 14170
rect 28194 14118 28206 14170
rect 28258 14118 37950 14170
rect 38002 14118 38014 14170
rect 38066 14118 38078 14170
rect 38130 14118 38142 14170
rect 38194 14118 38206 14170
rect 38258 14118 47950 14170
rect 48002 14118 48014 14170
rect 48066 14118 48078 14170
rect 48130 14118 48142 14170
rect 48194 14118 48206 14170
rect 48258 14118 49864 14170
rect 1104 14096 49864 14118
rect 3605 14059 3663 14065
rect 3605 14025 3617 14059
rect 3651 14056 3663 14059
rect 10226 14056 10232 14068
rect 3651 14028 10232 14056
rect 3651 14025 3663 14028
rect 3605 14019 3663 14025
rect 10226 14016 10232 14028
rect 10284 14016 10290 14068
rect 10318 14016 10324 14068
rect 10376 14056 10382 14068
rect 10413 14059 10471 14065
rect 10413 14056 10425 14059
rect 10376 14028 10425 14056
rect 10376 14016 10382 14028
rect 10413 14025 10425 14028
rect 10459 14025 10471 14059
rect 10413 14019 10471 14025
rect 10686 14016 10692 14068
rect 10744 14016 10750 14068
rect 11701 14059 11759 14065
rect 11701 14025 11713 14059
rect 11747 14056 11759 14059
rect 12158 14056 12164 14068
rect 11747 14028 12164 14056
rect 11747 14025 11759 14028
rect 11701 14019 11759 14025
rect 12158 14016 12164 14028
rect 12216 14016 12222 14068
rect 14642 14016 14648 14068
rect 14700 14056 14706 14068
rect 14737 14059 14795 14065
rect 14737 14056 14749 14059
rect 14700 14028 14749 14056
rect 14700 14016 14706 14028
rect 14737 14025 14749 14028
rect 14783 14025 14795 14059
rect 14737 14019 14795 14025
rect 15194 14016 15200 14068
rect 15252 14056 15258 14068
rect 15565 14059 15623 14065
rect 15565 14056 15577 14059
rect 15252 14028 15577 14056
rect 15252 14016 15258 14028
rect 15565 14025 15577 14028
rect 15611 14025 15623 14059
rect 15565 14019 15623 14025
rect 16574 14016 16580 14068
rect 16632 14056 16638 14068
rect 17129 14059 17187 14065
rect 17129 14056 17141 14059
rect 16632 14028 17141 14056
rect 16632 14016 16638 14028
rect 17129 14025 17141 14028
rect 17175 14025 17187 14059
rect 17129 14019 17187 14025
rect 17494 14016 17500 14068
rect 17552 14016 17558 14068
rect 18325 14059 18383 14065
rect 18325 14025 18337 14059
rect 18371 14056 18383 14059
rect 18414 14056 18420 14068
rect 18371 14028 18420 14056
rect 18371 14025 18383 14028
rect 18325 14019 18383 14025
rect 18414 14016 18420 14028
rect 18472 14016 18478 14068
rect 18693 14059 18751 14065
rect 18693 14025 18705 14059
rect 18739 14056 18751 14059
rect 18966 14056 18972 14068
rect 18739 14028 18972 14056
rect 18739 14025 18751 14028
rect 18693 14019 18751 14025
rect 18966 14016 18972 14028
rect 19024 14016 19030 14068
rect 19794 14016 19800 14068
rect 19852 14056 19858 14068
rect 22370 14056 22376 14068
rect 19852 14028 22376 14056
rect 19852 14016 19858 14028
rect 22370 14016 22376 14028
rect 22428 14016 22434 14068
rect 22646 14016 22652 14068
rect 22704 14016 22710 14068
rect 23753 14059 23811 14065
rect 23753 14025 23765 14059
rect 23799 14056 23811 14059
rect 23842 14056 23848 14068
rect 23799 14028 23848 14056
rect 23799 14025 23811 14028
rect 23753 14019 23811 14025
rect 23842 14016 23848 14028
rect 23900 14016 23906 14068
rect 25498 14016 25504 14068
rect 25556 14056 25562 14068
rect 25556 14028 26464 14056
rect 25556 14016 25562 14028
rect 11238 13988 11244 14000
rect 1780 13960 11244 13988
rect 1780 13929 1808 13960
rect 11238 13948 11244 13960
rect 11296 13948 11302 14000
rect 13998 13948 14004 14000
rect 14056 13948 14062 14000
rect 19518 13988 19524 14000
rect 16132 13960 19524 13988
rect 1765 13923 1823 13929
rect 1765 13889 1777 13923
rect 1811 13889 1823 13923
rect 1765 13883 1823 13889
rect 3510 13880 3516 13932
rect 3568 13920 3574 13932
rect 3973 13923 4031 13929
rect 3973 13920 3985 13923
rect 3568 13892 3985 13920
rect 3568 13880 3574 13892
rect 3973 13889 3985 13892
rect 4019 13889 4031 13923
rect 3973 13883 4031 13889
rect 10965 13923 11023 13929
rect 10965 13889 10977 13923
rect 11011 13920 11023 13923
rect 12069 13923 12127 13929
rect 11011 13892 11652 13920
rect 11011 13889 11023 13892
rect 10965 13883 11023 13889
rect 1302 13812 1308 13864
rect 1360 13852 1366 13864
rect 2041 13855 2099 13861
rect 2041 13852 2053 13855
rect 1360 13824 2053 13852
rect 1360 13812 1366 13824
rect 2041 13821 2053 13824
rect 2087 13821 2099 13855
rect 2041 13815 2099 13821
rect 9582 13812 9588 13864
rect 9640 13852 9646 13864
rect 9861 13855 9919 13861
rect 9861 13852 9873 13855
rect 9640 13824 9873 13852
rect 9640 13812 9646 13824
rect 9861 13821 9873 13824
rect 9907 13852 9919 13855
rect 11514 13852 11520 13864
rect 9907 13824 11520 13852
rect 9907 13821 9919 13824
rect 9861 13815 9919 13821
rect 11514 13812 11520 13824
rect 11572 13812 11578 13864
rect 11624 13852 11652 13892
rect 12069 13889 12081 13923
rect 12115 13889 12127 13923
rect 12069 13883 12127 13889
rect 12161 13923 12219 13929
rect 12161 13889 12173 13923
rect 12207 13920 12219 13923
rect 12342 13920 12348 13932
rect 12207 13892 12348 13920
rect 12207 13889 12219 13892
rect 12161 13883 12219 13889
rect 12084 13852 12112 13883
rect 12342 13880 12348 13892
rect 12400 13880 12406 13932
rect 15838 13880 15844 13932
rect 15896 13920 15902 13932
rect 15933 13923 15991 13929
rect 15933 13920 15945 13923
rect 15896 13892 15945 13920
rect 15896 13880 15902 13892
rect 15933 13889 15945 13892
rect 15979 13889 15991 13923
rect 16132 13920 16160 13960
rect 19518 13948 19524 13960
rect 19576 13948 19582 14000
rect 22664 13988 22692 14016
rect 24026 13988 24032 14000
rect 21206 13974 22692 13988
rect 21192 13960 22692 13974
rect 23506 13960 24032 13988
rect 15933 13883 15991 13889
rect 16040 13892 16160 13920
rect 11624 13824 12112 13852
rect 12253 13855 12311 13861
rect 12253 13821 12265 13855
rect 12299 13852 12311 13855
rect 12299 13824 12333 13852
rect 12299 13821 12311 13824
rect 12253 13815 12311 13821
rect 10042 13744 10048 13796
rect 10100 13784 10106 13796
rect 12268 13784 12296 13815
rect 12802 13812 12808 13864
rect 12860 13852 12866 13864
rect 12989 13855 13047 13861
rect 12989 13852 13001 13855
rect 12860 13824 13001 13852
rect 12860 13812 12866 13824
rect 12989 13821 13001 13824
rect 13035 13821 13047 13855
rect 12989 13815 13047 13821
rect 13265 13855 13323 13861
rect 13265 13821 13277 13855
rect 13311 13852 13323 13855
rect 13354 13852 13360 13864
rect 13311 13824 13360 13852
rect 13311 13821 13323 13824
rect 13265 13815 13323 13821
rect 13354 13812 13360 13824
rect 13412 13812 13418 13864
rect 13998 13812 14004 13864
rect 14056 13852 14062 13864
rect 14918 13852 14924 13864
rect 14056 13824 14924 13852
rect 14056 13812 14062 13824
rect 14918 13812 14924 13824
rect 14976 13852 14982 13864
rect 16040 13861 16068 13892
rect 16666 13880 16672 13932
rect 16724 13920 16730 13932
rect 17589 13923 17647 13929
rect 17589 13920 17601 13923
rect 16724 13892 17601 13920
rect 16724 13880 16730 13892
rect 17589 13889 17601 13892
rect 17635 13889 17647 13923
rect 17589 13883 17647 13889
rect 18785 13923 18843 13929
rect 18785 13889 18797 13923
rect 18831 13920 18843 13923
rect 19426 13920 19432 13932
rect 18831 13892 19432 13920
rect 18831 13889 18843 13892
rect 18785 13883 18843 13889
rect 19426 13880 19432 13892
rect 19484 13880 19490 13932
rect 15013 13855 15071 13861
rect 15013 13852 15025 13855
rect 14976 13824 15025 13852
rect 14976 13812 14982 13824
rect 15013 13821 15025 13824
rect 15059 13852 15071 13855
rect 15197 13855 15255 13861
rect 15197 13852 15209 13855
rect 15059 13824 15209 13852
rect 15059 13821 15071 13824
rect 15013 13815 15071 13821
rect 15197 13821 15209 13824
rect 15243 13821 15255 13855
rect 15197 13815 15255 13821
rect 16025 13855 16083 13861
rect 16025 13821 16037 13855
rect 16071 13821 16083 13855
rect 16025 13815 16083 13821
rect 16206 13812 16212 13864
rect 16264 13812 16270 13864
rect 16482 13812 16488 13864
rect 16540 13852 16546 13864
rect 16761 13855 16819 13861
rect 16761 13852 16773 13855
rect 16540 13824 16773 13852
rect 16540 13812 16546 13824
rect 16761 13821 16773 13824
rect 16807 13821 16819 13855
rect 16761 13815 16819 13821
rect 17678 13812 17684 13864
rect 17736 13812 17742 13864
rect 18877 13855 18935 13861
rect 18877 13821 18889 13855
rect 18923 13821 18935 13855
rect 18877 13815 18935 13821
rect 12526 13784 12532 13796
rect 10100 13756 12532 13784
rect 10100 13744 10106 13756
rect 12526 13744 12532 13756
rect 12584 13744 12590 13796
rect 15746 13784 15752 13796
rect 14292 13756 15752 13784
rect 10870 13676 10876 13728
rect 10928 13716 10934 13728
rect 14292 13716 14320 13756
rect 15746 13744 15752 13756
rect 15804 13744 15810 13796
rect 16776 13756 17448 13784
rect 10928 13688 14320 13716
rect 10928 13676 10934 13688
rect 15378 13676 15384 13728
rect 15436 13716 15442 13728
rect 16776 13716 16804 13756
rect 15436 13688 16804 13716
rect 17420 13716 17448 13756
rect 18782 13744 18788 13796
rect 18840 13784 18846 13796
rect 18892 13784 18920 13815
rect 18966 13812 18972 13864
rect 19024 13852 19030 13864
rect 19705 13855 19763 13861
rect 19705 13852 19717 13855
rect 19024 13824 19717 13852
rect 19024 13812 19030 13824
rect 19705 13821 19717 13824
rect 19751 13821 19763 13855
rect 19705 13815 19763 13821
rect 20714 13812 20720 13864
rect 20772 13852 20778 13864
rect 21192 13852 21220 13960
rect 24026 13948 24032 13960
rect 24084 13948 24090 14000
rect 25130 13948 25136 14000
rect 25188 13948 25194 14000
rect 26436 13988 26464 14028
rect 26510 14016 26516 14068
rect 26568 14056 26574 14068
rect 26605 14059 26663 14065
rect 26605 14056 26617 14059
rect 26568 14028 26617 14056
rect 26568 14016 26574 14028
rect 26605 14025 26617 14028
rect 26651 14025 26663 14059
rect 30006 14056 30012 14068
rect 26605 14019 26663 14025
rect 29380 14028 30012 14056
rect 26436 13960 28856 13988
rect 24854 13880 24860 13932
rect 24912 13880 24918 13932
rect 26786 13920 26792 13932
rect 26266 13892 26792 13920
rect 26786 13880 26792 13892
rect 26844 13880 26850 13932
rect 27157 13923 27215 13929
rect 27157 13889 27169 13923
rect 27203 13920 27215 13923
rect 28074 13920 28080 13932
rect 27203 13892 28080 13920
rect 27203 13889 27215 13892
rect 27157 13883 27215 13889
rect 28074 13880 28080 13892
rect 28132 13880 28138 13932
rect 28828 13920 28856 13960
rect 28902 13948 28908 14000
rect 28960 13948 28966 14000
rect 29270 13920 29276 13932
rect 28828 13892 29276 13920
rect 29270 13880 29276 13892
rect 29328 13880 29334 13932
rect 29380 13929 29408 14028
rect 30006 14016 30012 14028
rect 30064 14056 30070 14068
rect 30466 14056 30472 14068
rect 30064 14028 30472 14056
rect 30064 14016 30070 14028
rect 30466 14016 30472 14028
rect 30524 14016 30530 14068
rect 31110 14016 31116 14068
rect 31168 14016 31174 14068
rect 31573 14059 31631 14065
rect 31573 14025 31585 14059
rect 31619 14056 31631 14059
rect 36081 14059 36139 14065
rect 36081 14056 36093 14059
rect 31619 14028 36093 14056
rect 31619 14025 31631 14028
rect 31573 14019 31631 14025
rect 36081 14025 36093 14028
rect 36127 14025 36139 14059
rect 36081 14019 36139 14025
rect 36446 14016 36452 14068
rect 36504 14056 36510 14068
rect 36725 14059 36783 14065
rect 36725 14056 36737 14059
rect 36504 14028 36737 14056
rect 36504 14016 36510 14028
rect 36725 14025 36737 14028
rect 36771 14025 36783 14059
rect 36725 14019 36783 14025
rect 37461 14059 37519 14065
rect 37461 14025 37473 14059
rect 37507 14056 37519 14059
rect 41506 14056 41512 14068
rect 37507 14028 41512 14056
rect 37507 14025 37519 14028
rect 37461 14019 37519 14025
rect 41506 14016 41512 14028
rect 41564 14016 41570 14068
rect 45649 14059 45707 14065
rect 45649 14025 45661 14059
rect 45695 14056 45707 14059
rect 47026 14056 47032 14068
rect 45695 14028 47032 14056
rect 45695 14025 45707 14028
rect 45649 14019 45707 14025
rect 47026 14016 47032 14028
rect 47084 14016 47090 14068
rect 48406 14016 48412 14068
rect 48464 14016 48470 14068
rect 49234 14016 49240 14068
rect 49292 14016 49298 14068
rect 31386 13988 31392 14000
rect 30866 13960 31392 13988
rect 31386 13948 31392 13960
rect 31444 13948 31450 14000
rect 32858 13988 32864 14000
rect 31726 13960 32864 13988
rect 29365 13923 29423 13929
rect 29365 13889 29377 13923
rect 29411 13889 29423 13923
rect 29365 13883 29423 13889
rect 20772 13824 21220 13852
rect 20772 13812 20778 13824
rect 21358 13812 21364 13864
rect 21416 13852 21422 13864
rect 21453 13855 21511 13861
rect 21453 13852 21465 13855
rect 21416 13824 21465 13852
rect 21416 13812 21422 13824
rect 21453 13821 21465 13824
rect 21499 13821 21511 13855
rect 21453 13815 21511 13821
rect 22002 13812 22008 13864
rect 22060 13812 22066 13864
rect 22278 13812 22284 13864
rect 22336 13812 22342 13864
rect 24210 13812 24216 13864
rect 24268 13812 24274 13864
rect 28626 13812 28632 13864
rect 28684 13852 28690 13864
rect 31726 13852 31754 13960
rect 32858 13948 32864 13960
rect 32916 13948 32922 14000
rect 34330 13988 34336 14000
rect 33810 13960 34336 13988
rect 34330 13948 34336 13960
rect 34388 13948 34394 14000
rect 37550 13988 37556 14000
rect 35084 13960 37556 13988
rect 34885 13923 34943 13929
rect 34885 13920 34897 13923
rect 34440 13892 34897 13920
rect 28684 13824 31754 13852
rect 28684 13812 28690 13824
rect 32306 13812 32312 13864
rect 32364 13812 32370 13864
rect 32585 13855 32643 13861
rect 32585 13852 32597 13855
rect 32416 13824 32597 13852
rect 18840 13756 18920 13784
rect 18840 13744 18846 13756
rect 31294 13744 31300 13796
rect 31352 13784 31358 13796
rect 32214 13784 32220 13796
rect 31352 13756 32220 13784
rect 31352 13744 31358 13756
rect 32214 13744 32220 13756
rect 32272 13784 32278 13796
rect 32416 13784 32444 13824
rect 32585 13821 32597 13824
rect 32631 13821 32643 13855
rect 32585 13815 32643 13821
rect 32674 13812 32680 13864
rect 32732 13852 32738 13864
rect 34440 13852 34468 13892
rect 34885 13889 34897 13892
rect 34931 13889 34943 13923
rect 34885 13883 34943 13889
rect 34974 13880 34980 13932
rect 35032 13880 35038 13932
rect 35084 13852 35112 13960
rect 37550 13948 37556 13960
rect 37608 13948 37614 14000
rect 37642 13948 37648 14000
rect 37700 13988 37706 14000
rect 37921 13991 37979 13997
rect 37921 13988 37933 13991
rect 37700 13960 37933 13988
rect 37700 13948 37706 13960
rect 37921 13957 37933 13960
rect 37967 13957 37979 13991
rect 37921 13951 37979 13957
rect 39298 13948 39304 14000
rect 39356 13988 39362 14000
rect 45005 13991 45063 13997
rect 45005 13988 45017 13991
rect 39356 13960 45017 13988
rect 39356 13948 39362 13960
rect 45005 13957 45017 13960
rect 45051 13957 45063 13991
rect 45005 13951 45063 13957
rect 48133 13991 48191 13997
rect 48133 13957 48145 13991
rect 48179 13988 48191 13991
rect 49142 13988 49148 14000
rect 48179 13960 49148 13988
rect 48179 13957 48191 13960
rect 48133 13951 48191 13957
rect 49142 13948 49148 13960
rect 49200 13948 49206 14000
rect 37829 13923 37887 13929
rect 37829 13920 37841 13923
rect 35728 13892 37841 13920
rect 32732 13824 34468 13852
rect 34624 13824 35112 13852
rect 35161 13855 35219 13861
rect 32732 13812 32738 13824
rect 32272 13756 32444 13784
rect 32272 13744 32278 13756
rect 33870 13744 33876 13796
rect 33928 13784 33934 13796
rect 34057 13787 34115 13793
rect 34057 13784 34069 13787
rect 33928 13756 34069 13784
rect 33928 13744 33934 13756
rect 34057 13753 34069 13756
rect 34103 13753 34115 13787
rect 34057 13747 34115 13753
rect 34517 13787 34575 13793
rect 34517 13753 34529 13787
rect 34563 13784 34575 13787
rect 34624 13784 34652 13824
rect 35161 13821 35173 13855
rect 35207 13821 35219 13855
rect 35161 13815 35219 13821
rect 34563 13756 34652 13784
rect 35176 13784 35204 13815
rect 35342 13784 35348 13796
rect 35176 13756 35348 13784
rect 34563 13753 34575 13756
rect 34517 13747 34575 13753
rect 35342 13744 35348 13756
rect 35400 13744 35406 13796
rect 35728 13793 35756 13892
rect 37829 13889 37841 13892
rect 37875 13889 37887 13923
rect 37829 13883 37887 13889
rect 39025 13923 39083 13929
rect 39025 13889 39037 13923
rect 39071 13920 39083 13923
rect 39390 13920 39396 13932
rect 39071 13892 39396 13920
rect 39071 13889 39083 13892
rect 39025 13883 39083 13889
rect 39390 13880 39396 13892
rect 39448 13920 39454 13932
rect 39758 13920 39764 13932
rect 39448 13892 39764 13920
rect 39448 13880 39454 13892
rect 39758 13880 39764 13892
rect 39816 13880 39822 13932
rect 45830 13880 45836 13932
rect 45888 13880 45894 13932
rect 48222 13880 48228 13932
rect 48280 13920 48286 13932
rect 48593 13923 48651 13929
rect 48593 13920 48605 13923
rect 48280 13892 48605 13920
rect 48280 13880 48286 13892
rect 48593 13889 48605 13892
rect 48639 13889 48651 13923
rect 48593 13883 48651 13889
rect 36170 13812 36176 13864
rect 36228 13812 36234 13864
rect 36357 13855 36415 13861
rect 36357 13821 36369 13855
rect 36403 13852 36415 13855
rect 36630 13852 36636 13864
rect 36403 13824 36636 13852
rect 36403 13821 36415 13824
rect 36357 13815 36415 13821
rect 36630 13812 36636 13824
rect 36688 13812 36694 13864
rect 38013 13855 38071 13861
rect 38013 13821 38025 13855
rect 38059 13821 38071 13855
rect 38013 13815 38071 13821
rect 45189 13855 45247 13861
rect 45189 13821 45201 13855
rect 45235 13852 45247 13855
rect 46474 13852 46480 13864
rect 45235 13824 46480 13852
rect 45235 13821 45247 13824
rect 45189 13815 45247 13821
rect 35713 13787 35771 13793
rect 35713 13753 35725 13787
rect 35759 13753 35771 13787
rect 35713 13747 35771 13753
rect 37734 13744 37740 13796
rect 37792 13784 37798 13796
rect 38028 13784 38056 13815
rect 46474 13812 46480 13824
rect 46532 13812 46538 13864
rect 37792 13756 38056 13784
rect 37792 13744 37798 13756
rect 19337 13719 19395 13725
rect 19337 13716 19349 13719
rect 17420 13688 19349 13716
rect 15436 13676 15442 13688
rect 19337 13685 19349 13688
rect 19383 13716 19395 13719
rect 19794 13716 19800 13728
rect 19383 13688 19800 13716
rect 19383 13685 19395 13688
rect 19337 13679 19395 13685
rect 19794 13676 19800 13688
rect 19852 13676 19858 13728
rect 19968 13719 20026 13725
rect 19968 13685 19980 13719
rect 20014 13716 20026 13719
rect 20438 13716 20444 13728
rect 20014 13688 20444 13716
rect 20014 13685 20026 13688
rect 19968 13679 20026 13685
rect 20438 13676 20444 13688
rect 20496 13716 20502 13728
rect 23842 13716 23848 13728
rect 20496 13688 23848 13716
rect 20496 13676 20502 13688
rect 23842 13676 23848 13688
rect 23900 13676 23906 13728
rect 29628 13719 29686 13725
rect 29628 13685 29640 13719
rect 29674 13716 29686 13719
rect 30834 13716 30840 13728
rect 29674 13688 30840 13716
rect 29674 13685 29686 13688
rect 29628 13679 29686 13685
rect 30834 13676 30840 13688
rect 30892 13676 30898 13728
rect 31202 13676 31208 13728
rect 31260 13716 31266 13728
rect 33318 13716 33324 13728
rect 31260 13688 33324 13716
rect 31260 13676 31266 13688
rect 33318 13676 33324 13688
rect 33376 13676 33382 13728
rect 33686 13676 33692 13728
rect 33744 13716 33750 13728
rect 38378 13716 38384 13728
rect 33744 13688 38384 13716
rect 33744 13676 33750 13688
rect 38378 13676 38384 13688
rect 38436 13676 38442 13728
rect 1104 13626 49864 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 32950 13626
rect 33002 13574 33014 13626
rect 33066 13574 33078 13626
rect 33130 13574 33142 13626
rect 33194 13574 33206 13626
rect 33258 13574 42950 13626
rect 43002 13574 43014 13626
rect 43066 13574 43078 13626
rect 43130 13574 43142 13626
rect 43194 13574 43206 13626
rect 43258 13574 49864 13626
rect 1104 13552 49864 13574
rect 14461 13515 14519 13521
rect 14461 13512 14473 13515
rect 2746 13484 14473 13512
rect 2746 13376 2774 13484
rect 14461 13481 14473 13484
rect 14507 13481 14519 13515
rect 14461 13475 14519 13481
rect 14918 13472 14924 13524
rect 14976 13512 14982 13524
rect 15102 13512 15108 13524
rect 14976 13484 15108 13512
rect 14976 13472 14982 13484
rect 15102 13472 15108 13484
rect 15160 13472 15166 13524
rect 17402 13512 17408 13524
rect 16500 13484 17408 13512
rect 12526 13404 12532 13456
rect 12584 13444 12590 13456
rect 14826 13444 14832 13456
rect 12584 13416 14832 13444
rect 12584 13404 12590 13416
rect 14826 13404 14832 13416
rect 14884 13404 14890 13456
rect 15197 13447 15255 13453
rect 15197 13413 15209 13447
rect 15243 13444 15255 13447
rect 15470 13444 15476 13456
rect 15243 13416 15476 13444
rect 15243 13413 15255 13416
rect 15197 13407 15255 13413
rect 15470 13404 15476 13416
rect 15528 13404 15534 13456
rect 16500 13444 16528 13484
rect 17402 13472 17408 13484
rect 17460 13512 17466 13524
rect 17678 13512 17684 13524
rect 17460 13484 17684 13512
rect 17460 13472 17466 13484
rect 17678 13472 17684 13484
rect 17736 13512 17742 13524
rect 18141 13515 18199 13521
rect 18141 13512 18153 13515
rect 17736 13484 18153 13512
rect 17736 13472 17742 13484
rect 18141 13481 18153 13484
rect 18187 13481 18199 13515
rect 18141 13475 18199 13481
rect 19705 13515 19763 13521
rect 19705 13481 19717 13515
rect 19751 13512 19763 13515
rect 20254 13512 20260 13524
rect 19751 13484 20260 13512
rect 19751 13481 19763 13484
rect 19705 13475 19763 13481
rect 20254 13472 20260 13484
rect 20312 13472 20318 13524
rect 20346 13472 20352 13524
rect 20404 13512 20410 13524
rect 22097 13515 22155 13521
rect 22097 13512 22109 13515
rect 20404 13484 22109 13512
rect 20404 13472 20410 13484
rect 22097 13481 22109 13484
rect 22143 13481 22155 13515
rect 22097 13475 22155 13481
rect 23293 13515 23351 13521
rect 23293 13481 23305 13515
rect 23339 13512 23351 13515
rect 23382 13512 23388 13524
rect 23339 13484 23388 13512
rect 23339 13481 23351 13484
rect 23293 13475 23351 13481
rect 23382 13472 23388 13484
rect 23440 13472 23446 13524
rect 23474 13472 23480 13524
rect 23532 13512 23538 13524
rect 24118 13512 24124 13524
rect 23532 13484 24124 13512
rect 23532 13472 23538 13484
rect 24118 13472 24124 13484
rect 24176 13472 24182 13524
rect 24857 13515 24915 13521
rect 24857 13481 24869 13515
rect 24903 13512 24915 13515
rect 25222 13512 25228 13524
rect 24903 13484 25228 13512
rect 24903 13481 24915 13484
rect 24857 13475 24915 13481
rect 25222 13472 25228 13484
rect 25280 13472 25286 13524
rect 28074 13472 28080 13524
rect 28132 13512 28138 13524
rect 28350 13512 28356 13524
rect 28132 13484 28356 13512
rect 28132 13472 28138 13484
rect 28350 13472 28356 13484
rect 28408 13472 28414 13524
rect 28445 13515 28503 13521
rect 28445 13481 28457 13515
rect 28491 13512 28503 13515
rect 28491 13484 32444 13512
rect 28491 13481 28503 13484
rect 28445 13475 28503 13481
rect 16316 13416 16528 13444
rect 1780 13348 2774 13376
rect 10781 13379 10839 13385
rect 1780 13317 1808 13348
rect 10781 13345 10793 13379
rect 10827 13376 10839 13379
rect 11054 13376 11060 13388
rect 10827 13348 11060 13376
rect 10827 13345 10839 13348
rect 10781 13339 10839 13345
rect 11054 13336 11060 13348
rect 11112 13336 11118 13388
rect 14734 13336 14740 13388
rect 14792 13376 14798 13388
rect 15657 13379 15715 13385
rect 15657 13376 15669 13379
rect 14792 13348 15669 13376
rect 14792 13336 14798 13348
rect 15657 13345 15669 13348
rect 15703 13345 15715 13379
rect 15657 13339 15715 13345
rect 15841 13379 15899 13385
rect 15841 13345 15853 13379
rect 15887 13376 15899 13379
rect 16316 13376 16344 13416
rect 17770 13404 17776 13456
rect 17828 13444 17834 13456
rect 17828 13416 19380 13444
rect 17828 13404 17834 13416
rect 15887 13348 16344 13376
rect 16393 13379 16451 13385
rect 15887 13345 15899 13348
rect 15841 13339 15899 13345
rect 16393 13345 16405 13379
rect 16439 13376 16451 13379
rect 18966 13376 18972 13388
rect 16439 13348 18972 13376
rect 16439 13345 16451 13348
rect 16393 13339 16451 13345
rect 1765 13311 1823 13317
rect 1765 13277 1777 13311
rect 1811 13277 1823 13311
rect 1765 13271 1823 13277
rect 2774 13268 2780 13320
rect 2832 13268 2838 13320
rect 12802 13268 12808 13320
rect 12860 13308 12866 13320
rect 13078 13308 13084 13320
rect 12860 13280 13084 13308
rect 12860 13268 12866 13280
rect 13078 13268 13084 13280
rect 13136 13308 13142 13320
rect 16408 13308 16436 13339
rect 18966 13336 18972 13348
rect 19024 13336 19030 13388
rect 19352 13376 19380 13416
rect 19426 13404 19432 13456
rect 19484 13444 19490 13456
rect 19886 13444 19892 13456
rect 19484 13416 19892 13444
rect 19484 13404 19490 13416
rect 19886 13404 19892 13416
rect 19944 13404 19950 13456
rect 27430 13444 27436 13456
rect 20088 13416 21956 13444
rect 20088 13376 20116 13416
rect 19352 13348 20116 13376
rect 20162 13336 20168 13388
rect 20220 13336 20226 13388
rect 20257 13379 20315 13385
rect 20257 13345 20269 13379
rect 20303 13345 20315 13379
rect 20257 13339 20315 13345
rect 19978 13308 19984 13320
rect 13136 13280 16436 13308
rect 17972 13280 19984 13308
rect 13136 13268 13142 13280
rect 11057 13243 11115 13249
rect 11057 13209 11069 13243
rect 11103 13209 11115 13243
rect 11057 13203 11115 13209
rect 11072 13172 11100 13203
rect 11698 13200 11704 13252
rect 11756 13200 11762 13252
rect 13725 13243 13783 13249
rect 13725 13209 13737 13243
rect 13771 13240 13783 13243
rect 14369 13243 14427 13249
rect 14369 13240 14381 13243
rect 13771 13212 14381 13240
rect 13771 13209 13783 13212
rect 13725 13203 13783 13209
rect 14369 13209 14381 13212
rect 14415 13240 14427 13243
rect 14415 13212 15516 13240
rect 14415 13209 14427 13212
rect 14369 13203 14427 13209
rect 11974 13172 11980 13184
rect 11072 13144 11980 13172
rect 11974 13132 11980 13144
rect 12032 13132 12038 13184
rect 12710 13132 12716 13184
rect 12768 13172 12774 13184
rect 13081 13175 13139 13181
rect 13081 13172 13093 13175
rect 12768 13144 13093 13172
rect 12768 13132 12774 13144
rect 13081 13141 13093 13144
rect 13127 13141 13139 13175
rect 13081 13135 13139 13141
rect 13909 13175 13967 13181
rect 13909 13141 13921 13175
rect 13955 13172 13967 13175
rect 14090 13172 14096 13184
rect 13955 13144 14096 13172
rect 13955 13141 13967 13144
rect 13909 13135 13967 13141
rect 14090 13132 14096 13144
rect 14148 13132 14154 13184
rect 14182 13132 14188 13184
rect 14240 13172 14246 13184
rect 15378 13172 15384 13184
rect 14240 13144 15384 13172
rect 14240 13132 14246 13144
rect 15378 13132 15384 13144
rect 15436 13132 15442 13184
rect 15488 13172 15516 13212
rect 15562 13200 15568 13252
rect 15620 13200 15626 13252
rect 16390 13200 16396 13252
rect 16448 13240 16454 13252
rect 16669 13243 16727 13249
rect 16669 13240 16681 13243
rect 16448 13212 16681 13240
rect 16448 13200 16454 13212
rect 16669 13209 16681 13212
rect 16715 13209 16727 13243
rect 16669 13203 16727 13209
rect 17126 13200 17132 13252
rect 17184 13200 17190 13252
rect 17972 13172 18000 13280
rect 19978 13268 19984 13280
rect 20036 13268 20042 13320
rect 18693 13243 18751 13249
rect 18693 13209 18705 13243
rect 18739 13240 18751 13243
rect 20073 13243 20131 13249
rect 20073 13240 20085 13243
rect 18739 13212 20085 13240
rect 18739 13209 18751 13212
rect 18693 13203 18751 13209
rect 20073 13209 20085 13212
rect 20119 13209 20131 13243
rect 20073 13203 20131 13209
rect 15488 13144 18000 13172
rect 19058 13132 19064 13184
rect 19116 13172 19122 13184
rect 19702 13172 19708 13184
rect 19116 13144 19708 13172
rect 19116 13132 19122 13144
rect 19702 13132 19708 13144
rect 19760 13132 19766 13184
rect 20272 13172 20300 13339
rect 21450 13336 21456 13388
rect 21508 13336 21514 13388
rect 21928 13376 21956 13416
rect 22572 13416 27436 13444
rect 22572 13385 22600 13416
rect 27430 13404 27436 13416
rect 27488 13404 27494 13456
rect 29733 13447 29791 13453
rect 29733 13413 29745 13447
rect 29779 13444 29791 13447
rect 30834 13444 30840 13456
rect 29779 13416 30840 13444
rect 29779 13413 29791 13416
rect 29733 13407 29791 13413
rect 30834 13404 30840 13416
rect 30892 13404 30898 13456
rect 32416 13444 32444 13484
rect 32766 13472 32772 13524
rect 32824 13472 32830 13524
rect 33318 13472 33324 13524
rect 33376 13472 33382 13524
rect 34885 13515 34943 13521
rect 34885 13481 34897 13515
rect 34931 13512 34943 13515
rect 35986 13512 35992 13524
rect 34931 13484 35992 13512
rect 34931 13481 34943 13484
rect 34885 13475 34943 13481
rect 35986 13472 35992 13484
rect 36044 13472 36050 13524
rect 37366 13512 37372 13524
rect 36556 13484 37372 13512
rect 33686 13444 33692 13456
rect 32416 13416 33692 13444
rect 33686 13404 33692 13416
rect 33744 13404 33750 13456
rect 36556 13444 36584 13484
rect 37366 13472 37372 13484
rect 37424 13472 37430 13524
rect 37826 13472 37832 13524
rect 37884 13512 37890 13524
rect 38473 13515 38531 13521
rect 38473 13512 38485 13515
rect 37884 13484 38485 13512
rect 37884 13472 37890 13484
rect 38473 13481 38485 13484
rect 38519 13512 38531 13515
rect 38746 13512 38752 13524
rect 38519 13484 38752 13512
rect 38519 13481 38531 13484
rect 38473 13475 38531 13481
rect 38746 13472 38752 13484
rect 38804 13472 38810 13524
rect 35544 13416 36584 13444
rect 22557 13379 22615 13385
rect 21928 13348 22094 13376
rect 22066 13308 22094 13348
rect 22557 13345 22569 13379
rect 22603 13345 22615 13379
rect 22557 13339 22615 13345
rect 22741 13379 22799 13385
rect 22741 13345 22753 13379
rect 22787 13376 22799 13379
rect 23750 13376 23756 13388
rect 22787 13348 23756 13376
rect 22787 13345 22799 13348
rect 22741 13339 22799 13345
rect 23750 13336 23756 13348
rect 23808 13336 23814 13388
rect 23937 13379 23995 13385
rect 23937 13345 23949 13379
rect 23983 13376 23995 13379
rect 25501 13379 25559 13385
rect 23983 13348 25452 13376
rect 23983 13345 23995 13348
rect 23937 13339 23995 13345
rect 22830 13308 22836 13320
rect 22066 13280 22836 13308
rect 22830 13268 22836 13280
rect 22888 13268 22894 13320
rect 23658 13268 23664 13320
rect 23716 13268 23722 13320
rect 24946 13268 24952 13320
rect 25004 13308 25010 13320
rect 25225 13311 25283 13317
rect 25225 13308 25237 13311
rect 25004 13280 25237 13308
rect 25004 13268 25010 13280
rect 25225 13277 25237 13280
rect 25271 13277 25283 13311
rect 25424 13308 25452 13348
rect 25501 13345 25513 13379
rect 25547 13376 25559 13379
rect 25958 13376 25964 13388
rect 25547 13348 25964 13376
rect 25547 13345 25559 13348
rect 25501 13339 25559 13345
rect 25958 13336 25964 13348
rect 26016 13336 26022 13388
rect 29089 13379 29147 13385
rect 29089 13345 29101 13379
rect 29135 13376 29147 13379
rect 29638 13376 29644 13388
rect 29135 13348 29644 13376
rect 29135 13345 29147 13348
rect 29089 13339 29147 13345
rect 29638 13336 29644 13348
rect 29696 13336 29702 13388
rect 30282 13336 30288 13388
rect 30340 13336 30346 13388
rect 31021 13379 31079 13385
rect 31021 13345 31033 13379
rect 31067 13376 31079 13379
rect 32306 13376 32312 13388
rect 31067 13348 32312 13376
rect 31067 13345 31079 13348
rect 31021 13339 31079 13345
rect 32306 13336 32312 13348
rect 32364 13336 32370 13388
rect 32490 13336 32496 13388
rect 32548 13376 32554 13388
rect 32766 13376 32772 13388
rect 32548 13348 32772 13376
rect 32548 13336 32554 13348
rect 32766 13336 32772 13348
rect 32824 13336 32830 13388
rect 32858 13336 32864 13388
rect 32916 13376 32922 13388
rect 33873 13379 33931 13385
rect 33873 13376 33885 13379
rect 32916 13348 33885 13376
rect 32916 13336 32922 13348
rect 33873 13345 33885 13348
rect 33919 13345 33931 13379
rect 33873 13339 33931 13345
rect 35066 13336 35072 13388
rect 35124 13376 35130 13388
rect 35342 13376 35348 13388
rect 35124 13348 35348 13376
rect 35124 13336 35130 13348
rect 35342 13336 35348 13348
rect 35400 13336 35406 13388
rect 35544 13385 35572 13416
rect 35529 13379 35587 13385
rect 35529 13345 35541 13379
rect 35575 13345 35587 13379
rect 37090 13376 37096 13388
rect 35529 13339 35587 13345
rect 36188 13348 37096 13376
rect 25774 13308 25780 13320
rect 25424 13280 25780 13308
rect 25225 13271 25283 13277
rect 25774 13268 25780 13280
rect 25832 13268 25838 13320
rect 28810 13268 28816 13320
rect 28868 13308 28874 13320
rect 28905 13311 28963 13317
rect 28905 13308 28917 13311
rect 28868 13280 28917 13308
rect 28868 13268 28874 13280
rect 28905 13277 28917 13280
rect 28951 13277 28963 13311
rect 28905 13271 28963 13277
rect 29822 13268 29828 13320
rect 29880 13308 29886 13320
rect 30101 13311 30159 13317
rect 30101 13308 30113 13311
rect 29880 13280 30113 13308
rect 29880 13268 29886 13280
rect 30101 13277 30113 13280
rect 30147 13277 30159 13311
rect 33318 13308 33324 13320
rect 32430 13280 33324 13308
rect 30101 13271 30159 13277
rect 33318 13268 33324 13280
rect 33376 13268 33382 13320
rect 33594 13268 33600 13320
rect 33652 13308 33658 13320
rect 33689 13311 33747 13317
rect 33689 13308 33701 13311
rect 33652 13280 33701 13308
rect 33652 13268 33658 13280
rect 33689 13277 33701 13280
rect 33735 13277 33747 13311
rect 33689 13271 33747 13277
rect 35253 13311 35311 13317
rect 35253 13277 35265 13311
rect 35299 13308 35311 13311
rect 36188 13308 36216 13348
rect 37090 13336 37096 13348
rect 37148 13336 37154 13388
rect 35299 13280 36216 13308
rect 36449 13311 36507 13317
rect 35299 13277 35311 13280
rect 35253 13271 35311 13277
rect 36449 13277 36461 13311
rect 36495 13277 36507 13311
rect 36449 13271 36507 13277
rect 22465 13243 22523 13249
rect 22465 13209 22477 13243
rect 22511 13240 22523 13243
rect 23753 13243 23811 13249
rect 22511 13212 23704 13240
rect 22511 13209 22523 13212
rect 22465 13203 22523 13209
rect 23676 13184 23704 13212
rect 23753 13209 23765 13243
rect 23799 13240 23811 13243
rect 24026 13240 24032 13252
rect 23799 13212 24032 13240
rect 23799 13209 23811 13212
rect 23753 13203 23811 13209
rect 24026 13200 24032 13212
rect 24084 13240 24090 13252
rect 24394 13240 24400 13252
rect 24084 13212 24400 13240
rect 24084 13200 24090 13212
rect 24394 13200 24400 13212
rect 24452 13200 24458 13252
rect 26326 13240 26332 13252
rect 25332 13212 26332 13240
rect 20438 13172 20444 13184
rect 20272 13144 20444 13172
rect 20438 13132 20444 13144
rect 20496 13132 20502 13184
rect 20898 13132 20904 13184
rect 20956 13132 20962 13184
rect 21082 13132 21088 13184
rect 21140 13172 21146 13184
rect 21269 13175 21327 13181
rect 21269 13172 21281 13175
rect 21140 13144 21281 13172
rect 21140 13132 21146 13144
rect 21269 13141 21281 13144
rect 21315 13141 21327 13175
rect 21269 13135 21327 13141
rect 21358 13132 21364 13184
rect 21416 13172 21422 13184
rect 21818 13172 21824 13184
rect 21416 13144 21824 13172
rect 21416 13132 21422 13144
rect 21818 13132 21824 13144
rect 21876 13132 21882 13184
rect 23658 13132 23664 13184
rect 23716 13132 23722 13184
rect 24486 13132 24492 13184
rect 24544 13172 24550 13184
rect 25332 13181 25360 13212
rect 26326 13200 26332 13212
rect 26384 13200 26390 13252
rect 31297 13243 31355 13249
rect 31297 13209 31309 13243
rect 31343 13209 31355 13243
rect 33870 13240 33876 13252
rect 31297 13203 31355 13209
rect 32784 13212 33876 13240
rect 25317 13175 25375 13181
rect 25317 13172 25329 13175
rect 24544 13144 25329 13172
rect 24544 13132 24550 13144
rect 25317 13141 25329 13144
rect 25363 13141 25375 13175
rect 25317 13135 25375 13141
rect 26050 13132 26056 13184
rect 26108 13132 26114 13184
rect 26786 13132 26792 13184
rect 26844 13132 26850 13184
rect 27709 13175 27767 13181
rect 27709 13141 27721 13175
rect 27755 13172 27767 13175
rect 28534 13172 28540 13184
rect 27755 13144 28540 13172
rect 27755 13141 27767 13144
rect 27709 13135 27767 13141
rect 28534 13132 28540 13144
rect 28592 13132 28598 13184
rect 28813 13175 28871 13181
rect 28813 13141 28825 13175
rect 28859 13172 28871 13175
rect 28994 13172 29000 13184
rect 28859 13144 29000 13172
rect 28859 13141 28871 13144
rect 28813 13135 28871 13141
rect 28994 13132 29000 13144
rect 29052 13132 29058 13184
rect 29914 13132 29920 13184
rect 29972 13172 29978 13184
rect 30193 13175 30251 13181
rect 30193 13172 30205 13175
rect 29972 13144 30205 13172
rect 29972 13132 29978 13144
rect 30193 13141 30205 13144
rect 30239 13141 30251 13175
rect 31312 13172 31340 13203
rect 32784 13172 32812 13212
rect 33870 13200 33876 13212
rect 33928 13200 33934 13252
rect 34330 13200 34336 13252
rect 34388 13200 34394 13252
rect 35342 13200 35348 13252
rect 35400 13240 35406 13252
rect 36081 13243 36139 13249
rect 36081 13240 36093 13243
rect 35400 13212 36093 13240
rect 35400 13200 35406 13212
rect 36081 13209 36093 13212
rect 36127 13240 36139 13243
rect 36354 13240 36360 13252
rect 36127 13212 36360 13240
rect 36127 13209 36139 13212
rect 36081 13203 36139 13209
rect 36354 13200 36360 13212
rect 36412 13200 36418 13252
rect 36464 13184 36492 13271
rect 37826 13268 37832 13320
rect 37884 13268 37890 13320
rect 41506 13268 41512 13320
rect 41564 13268 41570 13320
rect 46474 13268 46480 13320
rect 46532 13308 46538 13320
rect 47949 13311 48007 13317
rect 47949 13308 47961 13311
rect 46532 13280 47961 13308
rect 46532 13268 46538 13280
rect 47949 13277 47961 13280
rect 47995 13277 48007 13311
rect 47949 13271 48007 13277
rect 36630 13200 36636 13252
rect 36688 13240 36694 13252
rect 36725 13243 36783 13249
rect 36725 13240 36737 13243
rect 36688 13212 36737 13240
rect 36688 13200 36694 13212
rect 36725 13209 36737 13212
rect 36771 13209 36783 13243
rect 36725 13203 36783 13209
rect 49142 13200 49148 13252
rect 49200 13200 49206 13252
rect 31312 13144 32812 13172
rect 33781 13175 33839 13181
rect 30193 13135 30251 13141
rect 33781 13141 33793 13175
rect 33827 13172 33839 13175
rect 34790 13172 34796 13184
rect 33827 13144 34796 13172
rect 33827 13141 33839 13144
rect 33781 13135 33839 13141
rect 34790 13132 34796 13144
rect 34848 13172 34854 13184
rect 35986 13172 35992 13184
rect 34848 13144 35992 13172
rect 34848 13132 34854 13144
rect 35986 13132 35992 13144
rect 36044 13132 36050 13184
rect 36446 13132 36452 13184
rect 36504 13172 36510 13184
rect 37366 13172 37372 13184
rect 36504 13144 37372 13172
rect 36504 13132 36510 13144
rect 37366 13132 37372 13144
rect 37424 13132 37430 13184
rect 37734 13132 37740 13184
rect 37792 13172 37798 13184
rect 38197 13175 38255 13181
rect 38197 13172 38209 13175
rect 37792 13144 38209 13172
rect 37792 13132 37798 13144
rect 38197 13141 38209 13144
rect 38243 13141 38255 13175
rect 38197 13135 38255 13141
rect 41325 13175 41383 13181
rect 41325 13141 41337 13175
rect 41371 13172 41383 13175
rect 46106 13172 46112 13184
rect 41371 13144 46112 13172
rect 41371 13141 41383 13144
rect 41325 13135 41383 13141
rect 46106 13132 46112 13144
rect 46164 13132 46170 13184
rect 1104 13082 49864 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 27950 13082
rect 28002 13030 28014 13082
rect 28066 13030 28078 13082
rect 28130 13030 28142 13082
rect 28194 13030 28206 13082
rect 28258 13030 37950 13082
rect 38002 13030 38014 13082
rect 38066 13030 38078 13082
rect 38130 13030 38142 13082
rect 38194 13030 38206 13082
rect 38258 13030 47950 13082
rect 48002 13030 48014 13082
rect 48066 13030 48078 13082
rect 48130 13030 48142 13082
rect 48194 13030 48206 13082
rect 48258 13030 49864 13082
rect 1104 13008 49864 13030
rect 2869 12971 2927 12977
rect 2869 12937 2881 12971
rect 2915 12968 2927 12971
rect 5442 12968 5448 12980
rect 2915 12940 5448 12968
rect 2915 12937 2927 12940
rect 2869 12931 2927 12937
rect 5442 12928 5448 12940
rect 5500 12928 5506 12980
rect 10962 12928 10968 12980
rect 11020 12968 11026 12980
rect 12161 12971 12219 12977
rect 12161 12968 12173 12971
rect 11020 12940 12173 12968
rect 11020 12928 11026 12940
rect 12161 12937 12173 12940
rect 12207 12937 12219 12971
rect 12161 12931 12219 12937
rect 13354 12928 13360 12980
rect 13412 12968 13418 12980
rect 14829 12971 14887 12977
rect 14829 12968 14841 12971
rect 13412 12940 14841 12968
rect 13412 12928 13418 12940
rect 14829 12937 14841 12940
rect 14875 12937 14887 12971
rect 14829 12931 14887 12937
rect 15933 12971 15991 12977
rect 15933 12937 15945 12971
rect 15979 12968 15991 12971
rect 16022 12968 16028 12980
rect 15979 12940 16028 12968
rect 15979 12937 15991 12940
rect 15933 12931 15991 12937
rect 16022 12928 16028 12940
rect 16080 12928 16086 12980
rect 16390 12928 16396 12980
rect 16448 12968 16454 12980
rect 16853 12971 16911 12977
rect 16853 12968 16865 12971
rect 16448 12940 16865 12968
rect 16448 12928 16454 12940
rect 16853 12937 16865 12940
rect 16899 12968 16911 12971
rect 17126 12968 17132 12980
rect 16899 12940 17132 12968
rect 16899 12937 16911 12940
rect 16853 12931 16911 12937
rect 17126 12928 17132 12940
rect 17184 12928 17190 12980
rect 20530 12968 20536 12980
rect 17788 12940 20536 12968
rect 1302 12860 1308 12912
rect 1360 12900 1366 12912
rect 1673 12903 1731 12909
rect 1673 12900 1685 12903
rect 1360 12872 1685 12900
rect 1360 12860 1366 12872
rect 1673 12869 1685 12872
rect 1719 12900 1731 12903
rect 2133 12903 2191 12909
rect 2133 12900 2145 12903
rect 1719 12872 2145 12900
rect 1719 12869 1731 12872
rect 1673 12863 1731 12869
rect 2133 12869 2145 12872
rect 2179 12869 2191 12903
rect 2133 12863 2191 12869
rect 11333 12903 11391 12909
rect 11333 12869 11345 12903
rect 11379 12900 11391 12903
rect 11698 12900 11704 12912
rect 11379 12872 11704 12900
rect 11379 12869 11391 12872
rect 11333 12863 11391 12869
rect 11698 12860 11704 12872
rect 11756 12860 11762 12912
rect 12066 12860 12072 12912
rect 12124 12860 12130 12912
rect 12805 12903 12863 12909
rect 12805 12900 12817 12903
rect 12636 12872 12817 12900
rect 1210 12792 1216 12844
rect 1268 12832 1274 12844
rect 3053 12835 3111 12841
rect 3053 12832 3065 12835
rect 1268 12804 3065 12832
rect 1268 12792 1274 12804
rect 3053 12801 3065 12804
rect 3099 12832 3111 12835
rect 3329 12835 3387 12841
rect 3329 12832 3341 12835
rect 3099 12804 3341 12832
rect 3099 12801 3111 12804
rect 3053 12795 3111 12801
rect 3329 12801 3341 12804
rect 3375 12801 3387 12835
rect 11716 12832 11744 12860
rect 12526 12832 12532 12844
rect 11716 12804 12532 12832
rect 3329 12795 3387 12801
rect 12526 12792 12532 12804
rect 12584 12832 12590 12844
rect 12636 12832 12664 12872
rect 12805 12869 12817 12872
rect 12851 12900 12863 12903
rect 12851 12872 13846 12900
rect 12851 12869 12863 12872
rect 12805 12863 12863 12869
rect 15102 12860 15108 12912
rect 15160 12900 15166 12912
rect 17788 12900 17816 12940
rect 20530 12928 20536 12940
rect 20588 12928 20594 12980
rect 20717 12971 20775 12977
rect 20717 12937 20729 12971
rect 20763 12937 20775 12971
rect 20717 12931 20775 12937
rect 15160 12872 17816 12900
rect 17865 12903 17923 12909
rect 15160 12860 15166 12872
rect 17865 12869 17877 12903
rect 17911 12900 17923 12903
rect 17954 12900 17960 12912
rect 17911 12872 17960 12900
rect 17911 12869 17923 12872
rect 17865 12863 17923 12869
rect 17954 12860 17960 12872
rect 18012 12900 18018 12912
rect 18322 12900 18328 12912
rect 18012 12872 18328 12900
rect 18012 12860 18018 12872
rect 18322 12860 18328 12872
rect 18380 12900 18386 12912
rect 18782 12900 18788 12912
rect 18380 12872 18788 12900
rect 18380 12860 18386 12872
rect 18782 12860 18788 12872
rect 18840 12860 18846 12912
rect 20732 12900 20760 12931
rect 20898 12928 20904 12980
rect 20956 12968 20962 12980
rect 21818 12968 21824 12980
rect 20956 12940 21824 12968
rect 20956 12928 20962 12940
rect 21818 12928 21824 12940
rect 21876 12928 21882 12980
rect 22649 12971 22707 12977
rect 22649 12937 22661 12971
rect 22695 12968 22707 12971
rect 22738 12968 22744 12980
rect 22695 12940 22744 12968
rect 22695 12937 22707 12940
rect 22649 12931 22707 12937
rect 22738 12928 22744 12940
rect 22796 12928 22802 12980
rect 23106 12928 23112 12980
rect 23164 12928 23170 12980
rect 23474 12928 23480 12980
rect 23532 12968 23538 12980
rect 23842 12968 23848 12980
rect 23532 12940 23848 12968
rect 23532 12928 23538 12940
rect 23842 12928 23848 12940
rect 23900 12928 23906 12980
rect 24762 12968 24768 12980
rect 23952 12940 24768 12968
rect 20990 12900 20996 12912
rect 20732 12872 20996 12900
rect 20990 12860 20996 12872
rect 21048 12860 21054 12912
rect 21177 12903 21235 12909
rect 21177 12869 21189 12903
rect 21223 12900 21235 12903
rect 23952 12900 23980 12940
rect 24762 12928 24768 12940
rect 24820 12928 24826 12980
rect 25038 12928 25044 12980
rect 25096 12968 25102 12980
rect 25593 12971 25651 12977
rect 25593 12968 25605 12971
rect 25096 12940 25605 12968
rect 25096 12928 25102 12940
rect 25593 12937 25605 12940
rect 25639 12937 25651 12971
rect 25593 12931 25651 12937
rect 26326 12928 26332 12980
rect 26384 12968 26390 12980
rect 26697 12971 26755 12977
rect 26697 12968 26709 12971
rect 26384 12940 26709 12968
rect 26384 12928 26390 12940
rect 26697 12937 26709 12940
rect 26743 12968 26755 12971
rect 27338 12968 27344 12980
rect 26743 12940 27344 12968
rect 26743 12937 26755 12940
rect 26697 12931 26755 12937
rect 27338 12928 27344 12940
rect 27396 12928 27402 12980
rect 28442 12968 28448 12980
rect 27448 12940 28448 12968
rect 26145 12903 26203 12909
rect 26145 12900 26157 12903
rect 21223 12872 23980 12900
rect 25346 12872 26157 12900
rect 21223 12869 21235 12872
rect 21177 12863 21235 12869
rect 26145 12869 26157 12872
rect 26191 12900 26203 12903
rect 26786 12900 26792 12912
rect 26191 12872 26792 12900
rect 26191 12869 26203 12872
rect 26145 12863 26203 12869
rect 26786 12860 26792 12872
rect 26844 12860 26850 12912
rect 27448 12909 27476 12940
rect 28442 12928 28448 12940
rect 28500 12968 28506 12980
rect 28500 12940 31616 12968
rect 28500 12928 28506 12940
rect 27433 12903 27491 12909
rect 27433 12869 27445 12903
rect 27479 12869 27491 12903
rect 28718 12900 28724 12912
rect 28658 12872 28724 12900
rect 27433 12863 27491 12869
rect 28718 12860 28724 12872
rect 28776 12860 28782 12912
rect 29546 12860 29552 12912
rect 29604 12860 29610 12912
rect 12584 12804 12664 12832
rect 12584 12792 12590 12804
rect 12710 12792 12716 12844
rect 12768 12832 12774 12844
rect 13078 12832 13084 12844
rect 12768 12804 13084 12832
rect 12768 12792 12774 12804
rect 13078 12792 13084 12804
rect 13136 12792 13142 12844
rect 16025 12835 16083 12841
rect 16025 12801 16037 12835
rect 16071 12832 16083 12835
rect 16206 12832 16212 12844
rect 16071 12804 16212 12832
rect 16071 12801 16083 12804
rect 16025 12795 16083 12801
rect 1857 12767 1915 12773
rect 1857 12733 1869 12767
rect 1903 12764 1915 12767
rect 9858 12764 9864 12776
rect 1903 12736 9864 12764
rect 1903 12733 1915 12736
rect 1857 12727 1915 12733
rect 9858 12724 9864 12736
rect 9916 12724 9922 12776
rect 12250 12724 12256 12776
rect 12308 12724 12314 12776
rect 13354 12724 13360 12776
rect 13412 12724 13418 12776
rect 14090 12724 14096 12776
rect 14148 12764 14154 12776
rect 16040 12764 16068 12795
rect 16206 12792 16212 12804
rect 16264 12792 16270 12844
rect 16482 12792 16488 12844
rect 16540 12792 16546 12844
rect 18693 12835 18751 12841
rect 18693 12801 18705 12835
rect 18739 12832 18751 12835
rect 18966 12832 18972 12844
rect 18739 12804 18972 12832
rect 18739 12801 18751 12804
rect 18693 12795 18751 12801
rect 18966 12792 18972 12804
rect 19024 12792 19030 12844
rect 19610 12792 19616 12844
rect 19668 12792 19674 12844
rect 21085 12835 21143 12841
rect 21085 12801 21097 12835
rect 21131 12832 21143 12835
rect 21910 12832 21916 12844
rect 21131 12804 21916 12832
rect 21131 12801 21143 12804
rect 21085 12795 21143 12801
rect 21910 12792 21916 12804
rect 21968 12792 21974 12844
rect 23014 12792 23020 12844
rect 23072 12792 23078 12844
rect 26234 12792 26240 12844
rect 26292 12832 26298 12844
rect 26329 12835 26387 12841
rect 26329 12832 26341 12835
rect 26292 12804 26341 12832
rect 26292 12792 26298 12804
rect 26329 12801 26341 12804
rect 26375 12832 26387 12835
rect 26970 12832 26976 12844
rect 26375 12804 26976 12832
rect 26375 12801 26387 12804
rect 26329 12795 26387 12801
rect 26970 12792 26976 12804
rect 27028 12792 27034 12844
rect 27154 12792 27160 12844
rect 27212 12792 27218 12844
rect 29362 12792 29368 12844
rect 29420 12832 29426 12844
rect 30006 12832 30012 12844
rect 29420 12804 30012 12832
rect 29420 12792 29426 12804
rect 30006 12792 30012 12804
rect 30064 12792 30070 12844
rect 31386 12792 31392 12844
rect 31444 12792 31450 12844
rect 14148 12736 16068 12764
rect 16117 12767 16175 12773
rect 14148 12724 14154 12736
rect 16117 12733 16129 12767
rect 16163 12764 16175 12767
rect 16500 12764 16528 12792
rect 16163 12736 16528 12764
rect 17221 12767 17279 12773
rect 16163 12733 16175 12736
rect 16117 12727 16175 12733
rect 17221 12733 17233 12767
rect 17267 12764 17279 12767
rect 19518 12764 19524 12776
rect 17267 12736 19524 12764
rect 17267 12733 17279 12736
rect 17221 12727 17279 12733
rect 19518 12724 19524 12736
rect 19576 12724 19582 12776
rect 19702 12724 19708 12776
rect 19760 12724 19766 12776
rect 19889 12767 19947 12773
rect 19889 12733 19901 12767
rect 19935 12764 19947 12767
rect 20898 12764 20904 12776
rect 19935 12736 20904 12764
rect 19935 12733 19947 12736
rect 19889 12727 19947 12733
rect 20898 12724 20904 12736
rect 20956 12724 20962 12776
rect 21174 12724 21180 12776
rect 21232 12764 21238 12776
rect 21269 12767 21327 12773
rect 21269 12764 21281 12767
rect 21232 12736 21281 12764
rect 21232 12724 21238 12736
rect 21269 12733 21281 12736
rect 21315 12733 21327 12767
rect 21269 12727 21327 12733
rect 21358 12724 21364 12776
rect 21416 12764 21422 12776
rect 22005 12767 22063 12773
rect 22005 12764 22017 12767
rect 21416 12736 22017 12764
rect 21416 12724 21422 12736
rect 22005 12733 22017 12736
rect 22051 12733 22063 12767
rect 22005 12727 22063 12733
rect 22094 12724 22100 12776
rect 22152 12764 22158 12776
rect 23201 12767 23259 12773
rect 23201 12764 23213 12767
rect 22152 12736 23213 12764
rect 22152 12724 22158 12736
rect 23201 12733 23213 12736
rect 23247 12764 23259 12767
rect 23382 12764 23388 12776
rect 23247 12736 23388 12764
rect 23247 12733 23259 12736
rect 23201 12727 23259 12733
rect 23382 12724 23388 12736
rect 23440 12724 23446 12776
rect 23842 12724 23848 12776
rect 23900 12724 23906 12776
rect 24118 12724 24124 12776
rect 24176 12764 24182 12776
rect 26510 12764 26516 12776
rect 24176 12736 26516 12764
rect 24176 12724 24182 12736
rect 26510 12724 26516 12736
rect 26568 12724 26574 12776
rect 29181 12767 29239 12773
rect 29181 12764 29193 12767
rect 26620 12736 29193 12764
rect 15289 12699 15347 12705
rect 15289 12665 15301 12699
rect 15335 12696 15347 12699
rect 15654 12696 15660 12708
rect 15335 12668 15660 12696
rect 15335 12665 15347 12668
rect 15289 12659 15347 12665
rect 15654 12656 15660 12668
rect 15712 12696 15718 12708
rect 16482 12696 16488 12708
rect 15712 12668 16488 12696
rect 15712 12656 15718 12668
rect 16482 12656 16488 12668
rect 16540 12656 16546 12708
rect 16761 12699 16819 12705
rect 16761 12665 16773 12699
rect 16807 12696 16819 12699
rect 17678 12696 17684 12708
rect 16807 12668 17684 12696
rect 16807 12665 16819 12668
rect 16761 12659 16819 12665
rect 17678 12656 17684 12668
rect 17736 12656 17742 12708
rect 20441 12699 20499 12705
rect 20441 12665 20453 12699
rect 20487 12696 20499 12699
rect 23400 12696 23428 12724
rect 20487 12668 20944 12696
rect 23400 12668 23980 12696
rect 20487 12665 20499 12668
rect 20441 12659 20499 12665
rect 11701 12631 11759 12637
rect 11701 12597 11713 12631
rect 11747 12628 11759 12631
rect 12618 12628 12624 12640
rect 11747 12600 12624 12628
rect 11747 12597 11759 12600
rect 11701 12591 11759 12597
rect 12618 12588 12624 12600
rect 12676 12588 12682 12640
rect 15565 12631 15623 12637
rect 15565 12597 15577 12631
rect 15611 12628 15623 12631
rect 17402 12628 17408 12640
rect 15611 12600 17408 12628
rect 15611 12597 15623 12600
rect 15565 12591 15623 12597
rect 17402 12588 17408 12600
rect 17460 12588 17466 12640
rect 18690 12588 18696 12640
rect 18748 12628 18754 12640
rect 19245 12631 19303 12637
rect 19245 12628 19257 12631
rect 18748 12600 19257 12628
rect 18748 12588 18754 12600
rect 19245 12597 19257 12600
rect 19291 12597 19303 12631
rect 20916 12628 20944 12668
rect 21450 12628 21456 12640
rect 20916 12600 21456 12628
rect 19245 12591 19303 12597
rect 21450 12588 21456 12600
rect 21508 12628 21514 12640
rect 23474 12628 23480 12640
rect 21508 12600 23480 12628
rect 21508 12588 21514 12600
rect 23474 12588 23480 12600
rect 23532 12588 23538 12640
rect 23952 12628 23980 12668
rect 25866 12656 25872 12708
rect 25924 12656 25930 12708
rect 26620 12628 26648 12736
rect 29181 12733 29193 12736
rect 29227 12733 29239 12767
rect 29181 12727 29239 12733
rect 29546 12724 29552 12776
rect 29604 12764 29610 12776
rect 30285 12767 30343 12773
rect 30285 12764 30297 12767
rect 29604 12736 30297 12764
rect 29604 12724 29610 12736
rect 30285 12733 30297 12736
rect 30331 12733 30343 12767
rect 31588 12764 31616 12940
rect 31754 12928 31760 12980
rect 31812 12968 31818 12980
rect 32398 12968 32404 12980
rect 31812 12940 32404 12968
rect 31812 12928 31818 12940
rect 32398 12928 32404 12940
rect 32456 12928 32462 12980
rect 32677 12971 32735 12977
rect 32677 12968 32689 12971
rect 32508 12940 32689 12968
rect 31754 12792 31760 12844
rect 31812 12832 31818 12844
rect 32508 12832 32536 12940
rect 32677 12937 32689 12940
rect 32723 12937 32735 12971
rect 32677 12931 32735 12937
rect 32766 12928 32772 12980
rect 32824 12928 32830 12980
rect 33778 12928 33784 12980
rect 33836 12968 33842 12980
rect 34054 12968 34060 12980
rect 33836 12940 34060 12968
rect 33836 12928 33842 12940
rect 34054 12928 34060 12940
rect 34112 12968 34118 12980
rect 34422 12968 34428 12980
rect 34112 12940 34428 12968
rect 34112 12928 34118 12940
rect 34422 12928 34428 12940
rect 34480 12928 34486 12980
rect 35526 12928 35532 12980
rect 35584 12968 35590 12980
rect 35802 12968 35808 12980
rect 35584 12940 35808 12968
rect 35584 12928 35590 12940
rect 35802 12928 35808 12940
rect 35860 12928 35866 12980
rect 35897 12971 35955 12977
rect 35897 12937 35909 12971
rect 35943 12968 35955 12971
rect 36078 12968 36084 12980
rect 35943 12940 36084 12968
rect 35943 12937 35955 12940
rect 35897 12931 35955 12937
rect 36078 12928 36084 12940
rect 36136 12968 36142 12980
rect 36633 12971 36691 12977
rect 36633 12968 36645 12971
rect 36136 12940 36645 12968
rect 36136 12928 36142 12940
rect 36633 12937 36645 12940
rect 36679 12968 36691 12971
rect 36814 12968 36820 12980
rect 36679 12940 36820 12968
rect 36679 12937 36691 12940
rect 36633 12931 36691 12937
rect 36814 12928 36820 12940
rect 36872 12928 36878 12980
rect 36909 12971 36967 12977
rect 36909 12937 36921 12971
rect 36955 12968 36967 12971
rect 37001 12971 37059 12977
rect 37001 12968 37013 12971
rect 36955 12940 37013 12968
rect 36955 12937 36967 12940
rect 36909 12931 36967 12937
rect 37001 12937 37013 12940
rect 37047 12968 37059 12971
rect 37826 12968 37832 12980
rect 37047 12940 37832 12968
rect 37047 12937 37059 12940
rect 37001 12931 37059 12937
rect 34882 12900 34888 12912
rect 31812 12804 32536 12832
rect 32600 12872 34888 12900
rect 31812 12792 31818 12804
rect 31588 12736 31754 12764
rect 30285 12727 30343 12733
rect 31726 12696 31754 12736
rect 32306 12724 32312 12776
rect 32364 12764 32370 12776
rect 32600 12764 32628 12872
rect 34882 12860 34888 12872
rect 34940 12900 34946 12912
rect 36446 12900 36452 12912
rect 34940 12872 36452 12900
rect 34940 12860 34946 12872
rect 36446 12860 36452 12872
rect 36504 12860 36510 12912
rect 36722 12860 36728 12912
rect 36780 12900 36786 12912
rect 36924 12900 36952 12931
rect 37826 12928 37832 12940
rect 37884 12928 37890 12980
rect 36780 12872 36952 12900
rect 36780 12860 36786 12872
rect 37734 12860 37740 12912
rect 37792 12860 37798 12912
rect 38746 12860 38752 12912
rect 38804 12860 38810 12912
rect 39942 12860 39948 12912
rect 40000 12900 40006 12912
rect 40037 12903 40095 12909
rect 40037 12900 40049 12903
rect 40000 12872 40049 12900
rect 40000 12860 40006 12872
rect 40037 12869 40049 12872
rect 40083 12900 40095 12903
rect 40497 12903 40555 12909
rect 40497 12900 40509 12903
rect 40083 12872 40509 12900
rect 40083 12869 40095 12872
rect 40037 12863 40095 12869
rect 40497 12869 40509 12872
rect 40543 12869 40555 12903
rect 40497 12863 40555 12869
rect 34054 12792 34060 12844
rect 34112 12792 34118 12844
rect 35158 12792 35164 12844
rect 35216 12832 35222 12844
rect 35216 12804 37136 12832
rect 35216 12792 35222 12804
rect 32364 12736 32628 12764
rect 32861 12767 32919 12773
rect 32364 12724 32370 12736
rect 32861 12733 32873 12767
rect 32907 12733 32919 12767
rect 32861 12727 32919 12733
rect 32876 12696 32904 12727
rect 33502 12724 33508 12776
rect 33560 12764 33566 12776
rect 35618 12764 35624 12776
rect 33560 12736 35624 12764
rect 33560 12724 33566 12736
rect 35618 12724 35624 12736
rect 35676 12724 35682 12776
rect 36081 12767 36139 12773
rect 36081 12733 36093 12767
rect 36127 12764 36139 12767
rect 36188 12764 36216 12804
rect 36127 12736 36216 12764
rect 37108 12764 37136 12804
rect 37366 12792 37372 12844
rect 37424 12832 37430 12844
rect 37461 12835 37519 12841
rect 37461 12832 37473 12835
rect 37424 12804 37473 12832
rect 37424 12792 37430 12804
rect 37461 12801 37473 12804
rect 37507 12801 37519 12835
rect 37461 12795 37519 12801
rect 46106 12792 46112 12844
rect 46164 12792 46170 12844
rect 47026 12792 47032 12844
rect 47084 12832 47090 12844
rect 47949 12835 48007 12841
rect 47949 12832 47961 12835
rect 47084 12804 47961 12832
rect 47084 12792 47090 12804
rect 47949 12801 47961 12804
rect 47995 12801 48007 12835
rect 47949 12795 48007 12801
rect 49142 12792 49148 12844
rect 49200 12792 49206 12844
rect 39485 12767 39543 12773
rect 39485 12764 39497 12767
rect 37108 12736 39497 12764
rect 36127 12733 36139 12736
rect 36081 12727 36139 12733
rect 39485 12733 39497 12736
rect 39531 12733 39543 12767
rect 39485 12727 39543 12733
rect 34514 12696 34520 12708
rect 31726 12668 32904 12696
rect 33244 12668 34520 12696
rect 23952 12600 26648 12628
rect 27154 12588 27160 12640
rect 27212 12628 27218 12640
rect 29362 12628 29368 12640
rect 27212 12600 29368 12628
rect 27212 12588 27218 12600
rect 29362 12588 29368 12600
rect 29420 12588 29426 12640
rect 32309 12631 32367 12637
rect 32309 12597 32321 12631
rect 32355 12628 32367 12631
rect 33244 12628 33272 12668
rect 34514 12656 34520 12668
rect 34572 12656 34578 12708
rect 35437 12699 35495 12705
rect 35437 12665 35449 12699
rect 35483 12696 35495 12699
rect 37366 12696 37372 12708
rect 35483 12668 37372 12696
rect 35483 12665 35495 12668
rect 35437 12659 35495 12665
rect 37366 12656 37372 12668
rect 37424 12656 37430 12708
rect 40221 12699 40279 12705
rect 40221 12665 40233 12699
rect 40267 12696 40279 12699
rect 47026 12696 47032 12708
rect 40267 12668 47032 12696
rect 40267 12665 40279 12668
rect 40221 12659 40279 12665
rect 47026 12656 47032 12668
rect 47084 12656 47090 12708
rect 32355 12600 33272 12628
rect 32355 12597 32367 12600
rect 32309 12591 32367 12597
rect 33318 12588 33324 12640
rect 33376 12628 33382 12640
rect 33413 12631 33471 12637
rect 33413 12628 33425 12631
rect 33376 12600 33425 12628
rect 33376 12588 33382 12600
rect 33413 12597 33425 12600
rect 33459 12628 33471 12631
rect 33597 12631 33655 12637
rect 33597 12628 33609 12631
rect 33459 12600 33609 12628
rect 33459 12597 33471 12600
rect 33413 12591 33471 12597
rect 33597 12597 33609 12600
rect 33643 12628 33655 12631
rect 34330 12628 34336 12640
rect 33643 12600 34336 12628
rect 33643 12597 33655 12600
rect 33597 12591 33655 12597
rect 34330 12588 34336 12600
rect 34388 12588 34394 12640
rect 36078 12588 36084 12640
rect 36136 12628 36142 12640
rect 36541 12631 36599 12637
rect 36541 12628 36553 12631
rect 36136 12600 36553 12628
rect 36136 12588 36142 12600
rect 36541 12597 36553 12600
rect 36587 12628 36599 12631
rect 39482 12628 39488 12640
rect 36587 12600 39488 12628
rect 36587 12597 36599 12600
rect 36541 12591 36599 12597
rect 39482 12588 39488 12600
rect 39540 12588 39546 12640
rect 45925 12631 45983 12637
rect 45925 12597 45937 12631
rect 45971 12628 45983 12631
rect 47946 12628 47952 12640
rect 45971 12600 47952 12628
rect 45971 12597 45983 12600
rect 45925 12591 45983 12597
rect 47946 12588 47952 12600
rect 48004 12588 48010 12640
rect 1104 12538 49864 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 32950 12538
rect 33002 12486 33014 12538
rect 33066 12486 33078 12538
rect 33130 12486 33142 12538
rect 33194 12486 33206 12538
rect 33258 12486 42950 12538
rect 43002 12486 43014 12538
rect 43066 12486 43078 12538
rect 43130 12486 43142 12538
rect 43194 12486 43206 12538
rect 43258 12486 49864 12538
rect 1104 12464 49864 12486
rect 12434 12384 12440 12436
rect 12492 12424 12498 12436
rect 13262 12424 13268 12436
rect 12492 12396 13268 12424
rect 12492 12384 12498 12396
rect 13262 12384 13268 12396
rect 13320 12424 13326 12436
rect 16025 12427 16083 12433
rect 13320 12396 15976 12424
rect 13320 12384 13326 12396
rect 15948 12368 15976 12396
rect 16025 12393 16037 12427
rect 16071 12424 16083 12427
rect 16114 12424 16120 12436
rect 16071 12396 16120 12424
rect 16071 12393 16083 12396
rect 16025 12387 16083 12393
rect 16114 12384 16120 12396
rect 16172 12384 16178 12436
rect 19334 12384 19340 12436
rect 19392 12424 19398 12436
rect 19429 12427 19487 12433
rect 19429 12424 19441 12427
rect 19392 12396 19441 12424
rect 19392 12384 19398 12396
rect 19429 12393 19441 12396
rect 19475 12393 19487 12427
rect 19429 12387 19487 12393
rect 20901 12427 20959 12433
rect 20901 12393 20913 12427
rect 20947 12424 20959 12427
rect 20947 12396 22876 12424
rect 20947 12393 20959 12396
rect 20901 12387 20959 12393
rect 15930 12316 15936 12368
rect 15988 12356 15994 12368
rect 22848 12356 22876 12396
rect 22922 12384 22928 12436
rect 22980 12424 22986 12436
rect 23293 12427 23351 12433
rect 23293 12424 23305 12427
rect 22980 12396 23305 12424
rect 22980 12384 22986 12396
rect 23293 12393 23305 12396
rect 23339 12393 23351 12427
rect 26050 12424 26056 12436
rect 23293 12387 23351 12393
rect 23676 12396 26056 12424
rect 23566 12356 23572 12368
rect 15988 12328 18828 12356
rect 15988 12316 15994 12328
rect 1857 12291 1915 12297
rect 1857 12257 1869 12291
rect 1903 12288 1915 12291
rect 5442 12288 5448 12300
rect 1903 12260 5448 12288
rect 1903 12257 1915 12260
rect 1857 12251 1915 12257
rect 5442 12248 5448 12260
rect 5500 12248 5506 12300
rect 9493 12291 9551 12297
rect 9493 12257 9505 12291
rect 9539 12288 9551 12291
rect 11054 12288 11060 12300
rect 9539 12260 11060 12288
rect 9539 12257 9551 12260
rect 9493 12251 9551 12257
rect 11054 12248 11060 12260
rect 11112 12288 11118 12300
rect 11701 12291 11759 12297
rect 11701 12288 11713 12291
rect 11112 12260 11713 12288
rect 11112 12248 11118 12260
rect 11701 12257 11713 12260
rect 11747 12288 11759 12291
rect 12710 12288 12716 12300
rect 11747 12260 12716 12288
rect 11747 12257 11759 12260
rect 11701 12251 11759 12257
rect 12710 12248 12716 12260
rect 12768 12288 12774 12300
rect 14277 12291 14335 12297
rect 14277 12288 14289 12291
rect 12768 12260 14289 12288
rect 12768 12248 12774 12260
rect 14277 12257 14289 12260
rect 14323 12257 14335 12291
rect 14277 12251 14335 12257
rect 14553 12291 14611 12297
rect 14553 12257 14565 12291
rect 14599 12288 14611 12291
rect 14918 12288 14924 12300
rect 14599 12260 14924 12288
rect 14599 12257 14611 12260
rect 14553 12251 14611 12257
rect 14918 12248 14924 12260
rect 14976 12248 14982 12300
rect 17218 12248 17224 12300
rect 17276 12288 17282 12300
rect 17313 12291 17371 12297
rect 17313 12288 17325 12291
rect 17276 12260 17325 12288
rect 17276 12248 17282 12260
rect 17313 12257 17325 12260
rect 17359 12257 17371 12291
rect 17313 12251 17371 12257
rect 1302 12180 1308 12232
rect 1360 12220 1366 12232
rect 1581 12223 1639 12229
rect 1581 12220 1593 12223
rect 1360 12192 1593 12220
rect 1360 12180 1366 12192
rect 1581 12189 1593 12192
rect 1627 12189 1639 12223
rect 1581 12183 1639 12189
rect 1596 12152 1624 12183
rect 15838 12180 15844 12232
rect 15896 12220 15902 12232
rect 16485 12223 16543 12229
rect 16485 12220 16497 12223
rect 15896 12192 16497 12220
rect 15896 12180 15902 12192
rect 16485 12189 16497 12192
rect 16531 12220 16543 12223
rect 17126 12220 17132 12232
rect 16531 12192 17132 12220
rect 16531 12189 16543 12192
rect 16485 12183 16543 12189
rect 17126 12180 17132 12192
rect 17184 12180 17190 12232
rect 17954 12180 17960 12232
rect 18012 12180 18018 12232
rect 2685 12155 2743 12161
rect 2685 12152 2697 12155
rect 1596 12124 2697 12152
rect 2685 12121 2697 12124
rect 2731 12121 2743 12155
rect 2685 12115 2743 12121
rect 9769 12155 9827 12161
rect 9769 12121 9781 12155
rect 9815 12152 9827 12155
rect 10042 12152 10048 12164
rect 9815 12124 10048 12152
rect 9815 12121 9827 12124
rect 9769 12115 9827 12121
rect 10042 12112 10048 12124
rect 10100 12112 10106 12164
rect 11698 12152 11704 12164
rect 10994 12124 11704 12152
rect 11698 12112 11704 12124
rect 11756 12112 11762 12164
rect 11977 12155 12035 12161
rect 11977 12121 11989 12155
rect 12023 12121 12035 12155
rect 11977 12115 12035 12121
rect 11238 12044 11244 12096
rect 11296 12044 11302 12096
rect 11992 12084 12020 12115
rect 12526 12112 12532 12164
rect 12584 12112 12590 12164
rect 13722 12112 13728 12164
rect 13780 12112 13786 12164
rect 15010 12152 15016 12164
rect 14936 12124 15016 12152
rect 12710 12084 12716 12096
rect 11992 12056 12716 12084
rect 12710 12044 12716 12056
rect 12768 12044 12774 12096
rect 13740 12084 13768 12112
rect 14734 12084 14740 12096
rect 13740 12056 14740 12084
rect 14734 12044 14740 12056
rect 14792 12044 14798 12096
rect 14936 12084 14964 12124
rect 15010 12112 15016 12124
rect 15068 12112 15074 12164
rect 16850 12112 16856 12164
rect 16908 12152 16914 12164
rect 18693 12155 18751 12161
rect 18693 12152 18705 12155
rect 16908 12124 18705 12152
rect 16908 12112 16914 12124
rect 18693 12121 18705 12124
rect 18739 12121 18751 12155
rect 18800 12152 18828 12328
rect 22572 12328 22784 12356
rect 22848 12328 23572 12356
rect 19334 12248 19340 12300
rect 19392 12288 19398 12300
rect 19392 12260 19932 12288
rect 19392 12248 19398 12260
rect 19518 12180 19524 12232
rect 19576 12220 19582 12232
rect 19797 12223 19855 12229
rect 19797 12220 19809 12223
rect 19576 12192 19809 12220
rect 19576 12180 19582 12192
rect 19797 12189 19809 12192
rect 19843 12189 19855 12223
rect 19904 12220 19932 12260
rect 19978 12248 19984 12300
rect 20036 12248 20042 12300
rect 20622 12248 20628 12300
rect 20680 12288 20686 12300
rect 21361 12291 21419 12297
rect 21361 12288 21373 12291
rect 20680 12260 21373 12288
rect 20680 12248 20686 12260
rect 21361 12257 21373 12260
rect 21407 12288 21419 12291
rect 21450 12288 21456 12300
rect 21407 12260 21456 12288
rect 21407 12257 21419 12260
rect 21361 12251 21419 12257
rect 21450 12248 21456 12260
rect 21508 12248 21514 12300
rect 21545 12291 21603 12297
rect 21545 12257 21557 12291
rect 21591 12288 21603 12291
rect 22094 12288 22100 12300
rect 21591 12260 22100 12288
rect 21591 12257 21603 12260
rect 21545 12251 21603 12257
rect 22094 12248 22100 12260
rect 22152 12248 22158 12300
rect 22572 12288 22600 12328
rect 22388 12260 22600 12288
rect 20990 12220 20996 12232
rect 19904 12192 20996 12220
rect 19797 12183 19855 12189
rect 20990 12180 20996 12192
rect 21048 12180 21054 12232
rect 21269 12223 21327 12229
rect 21269 12189 21281 12223
rect 21315 12220 21327 12223
rect 22388 12220 22416 12260
rect 22646 12248 22652 12300
rect 22704 12248 22710 12300
rect 22756 12288 22784 12328
rect 23566 12316 23572 12328
rect 23624 12316 23630 12368
rect 23676 12288 23704 12396
rect 26050 12384 26056 12396
rect 26108 12384 26114 12436
rect 26973 12427 27031 12433
rect 26973 12393 26985 12427
rect 27019 12424 27031 12427
rect 31754 12424 31760 12436
rect 27019 12396 31760 12424
rect 27019 12393 27031 12396
rect 26973 12387 27031 12393
rect 31754 12384 31760 12396
rect 31812 12384 31818 12436
rect 34698 12424 34704 12436
rect 32232 12396 34704 12424
rect 29178 12356 29184 12368
rect 27540 12328 29184 12356
rect 22756 12260 23704 12288
rect 23937 12291 23995 12297
rect 23937 12257 23949 12291
rect 23983 12288 23995 12291
rect 24486 12288 24492 12300
rect 23983 12260 24492 12288
rect 23983 12257 23995 12260
rect 23937 12251 23995 12257
rect 24486 12248 24492 12260
rect 24544 12248 24550 12300
rect 24857 12291 24915 12297
rect 24857 12257 24869 12291
rect 24903 12288 24915 12291
rect 24946 12288 24952 12300
rect 24903 12260 24952 12288
rect 24903 12257 24915 12260
rect 24857 12251 24915 12257
rect 24946 12248 24952 12260
rect 25004 12248 25010 12300
rect 25314 12248 25320 12300
rect 25372 12288 25378 12300
rect 27430 12288 27436 12300
rect 25372 12260 27436 12288
rect 25372 12248 25378 12260
rect 27430 12248 27436 12260
rect 27488 12248 27494 12300
rect 27540 12297 27568 12328
rect 29178 12316 29184 12328
rect 29236 12316 29242 12368
rect 31018 12316 31024 12368
rect 31076 12356 31082 12368
rect 32232 12356 32260 12396
rect 34698 12384 34704 12396
rect 34756 12384 34762 12436
rect 37642 12424 37648 12436
rect 34992 12396 37648 12424
rect 31076 12328 32260 12356
rect 31076 12316 31082 12328
rect 33870 12316 33876 12368
rect 33928 12356 33934 12368
rect 34992 12356 35020 12396
rect 37642 12384 37648 12396
rect 37700 12384 37706 12436
rect 38289 12427 38347 12433
rect 38289 12393 38301 12427
rect 38335 12424 38347 12427
rect 38335 12396 41414 12424
rect 38335 12393 38347 12396
rect 38289 12387 38347 12393
rect 33928 12328 35020 12356
rect 37093 12359 37151 12365
rect 33928 12316 33934 12328
rect 37093 12325 37105 12359
rect 37139 12356 37151 12359
rect 41386 12356 41414 12396
rect 37139 12328 41000 12356
rect 41386 12328 41644 12356
rect 37139 12325 37151 12328
rect 37093 12319 37151 12325
rect 27525 12291 27583 12297
rect 27525 12257 27537 12291
rect 27571 12257 27583 12291
rect 27525 12251 27583 12257
rect 29089 12291 29147 12297
rect 29089 12257 29101 12291
rect 29135 12288 29147 12291
rect 29362 12288 29368 12300
rect 29135 12260 29368 12288
rect 29135 12257 29147 12260
rect 29089 12251 29147 12257
rect 29362 12248 29368 12260
rect 29420 12288 29426 12300
rect 29733 12291 29791 12297
rect 29733 12288 29745 12291
rect 29420 12260 29745 12288
rect 29420 12248 29426 12260
rect 29733 12257 29745 12260
rect 29779 12257 29791 12291
rect 29733 12251 29791 12257
rect 32125 12291 32183 12297
rect 32125 12257 32137 12291
rect 32171 12288 32183 12291
rect 34054 12288 34060 12300
rect 32171 12260 34060 12288
rect 32171 12257 32183 12260
rect 32125 12251 32183 12257
rect 34054 12248 34060 12260
rect 34112 12248 34118 12300
rect 34790 12248 34796 12300
rect 34848 12288 34854 12300
rect 35161 12291 35219 12297
rect 35161 12288 35173 12291
rect 34848 12260 35173 12288
rect 34848 12248 34854 12260
rect 35161 12257 35173 12260
rect 35207 12257 35219 12291
rect 35161 12251 35219 12257
rect 35802 12248 35808 12300
rect 35860 12288 35866 12300
rect 35860 12260 37228 12288
rect 35860 12248 35866 12260
rect 21315 12192 22416 12220
rect 21315 12189 21327 12192
rect 21269 12183 21327 12189
rect 23566 12180 23572 12232
rect 23624 12220 23630 12232
rect 24302 12220 24308 12232
rect 23624 12192 24308 12220
rect 23624 12180 23630 12192
rect 24302 12180 24308 12192
rect 24360 12180 24366 12232
rect 24578 12180 24584 12232
rect 24636 12180 24642 12232
rect 26605 12223 26663 12229
rect 26605 12220 26617 12223
rect 25990 12192 26617 12220
rect 26605 12189 26617 12192
rect 26651 12220 26663 12223
rect 26786 12220 26792 12232
rect 26651 12192 26792 12220
rect 26651 12189 26663 12192
rect 26605 12183 26663 12189
rect 26786 12180 26792 12192
rect 26844 12220 26850 12232
rect 28261 12223 28319 12229
rect 26844 12192 27660 12220
rect 26844 12180 26850 12192
rect 21726 12152 21732 12164
rect 18800 12124 21732 12152
rect 18693 12115 18751 12121
rect 21726 12112 21732 12124
rect 21784 12112 21790 12164
rect 23661 12155 23719 12161
rect 23661 12152 23673 12155
rect 22112 12124 23673 12152
rect 15286 12084 15292 12096
rect 14936 12056 15292 12084
rect 15286 12044 15292 12056
rect 15344 12084 15350 12096
rect 16390 12084 16396 12096
rect 15344 12056 16396 12084
rect 15344 12044 15350 12056
rect 16390 12044 16396 12056
rect 16448 12044 16454 12096
rect 16482 12044 16488 12096
rect 16540 12084 16546 12096
rect 16761 12087 16819 12093
rect 16761 12084 16773 12087
rect 16540 12056 16773 12084
rect 16540 12044 16546 12056
rect 16761 12053 16773 12056
rect 16807 12053 16819 12087
rect 16761 12047 16819 12053
rect 17221 12087 17279 12093
rect 17221 12053 17233 12087
rect 17267 12084 17279 12087
rect 17310 12084 17316 12096
rect 17267 12056 17316 12084
rect 17267 12053 17279 12056
rect 17221 12047 17279 12053
rect 17310 12044 17316 12056
rect 17368 12044 17374 12096
rect 19889 12087 19947 12093
rect 19889 12053 19901 12087
rect 19935 12084 19947 12087
rect 20530 12084 20536 12096
rect 19935 12056 20536 12084
rect 19935 12053 19947 12056
rect 19889 12047 19947 12053
rect 20530 12044 20536 12056
rect 20588 12044 20594 12096
rect 21266 12044 21272 12096
rect 21324 12084 21330 12096
rect 21634 12084 21640 12096
rect 21324 12056 21640 12084
rect 21324 12044 21330 12056
rect 21634 12044 21640 12056
rect 21692 12044 21698 12096
rect 22112 12093 22140 12124
rect 23661 12121 23673 12124
rect 23707 12121 23719 12155
rect 26694 12152 26700 12164
rect 23661 12115 23719 12121
rect 26160 12124 26700 12152
rect 22097 12087 22155 12093
rect 22097 12053 22109 12087
rect 22143 12053 22155 12087
rect 22097 12047 22155 12053
rect 22462 12044 22468 12096
rect 22520 12044 22526 12096
rect 22554 12044 22560 12096
rect 22612 12044 22618 12096
rect 23753 12087 23811 12093
rect 23753 12053 23765 12087
rect 23799 12084 23811 12087
rect 26160 12084 26188 12124
rect 26694 12112 26700 12124
rect 26752 12112 26758 12164
rect 27154 12112 27160 12164
rect 27212 12152 27218 12164
rect 27433 12155 27491 12161
rect 27433 12152 27445 12155
rect 27212 12124 27445 12152
rect 27212 12112 27218 12124
rect 27433 12121 27445 12124
rect 27479 12152 27491 12155
rect 27522 12152 27528 12164
rect 27479 12124 27528 12152
rect 27479 12121 27491 12124
rect 27433 12115 27491 12121
rect 27522 12112 27528 12124
rect 27580 12112 27586 12164
rect 27632 12152 27660 12192
rect 28261 12189 28273 12223
rect 28307 12220 28319 12223
rect 28902 12220 28908 12232
rect 28307 12192 28908 12220
rect 28307 12189 28319 12192
rect 28261 12183 28319 12189
rect 28902 12180 28908 12192
rect 28960 12180 28966 12232
rect 31386 12180 31392 12232
rect 31444 12180 31450 12232
rect 34882 12180 34888 12232
rect 34940 12180 34946 12232
rect 28718 12152 28724 12164
rect 27632 12124 28724 12152
rect 28718 12112 28724 12124
rect 28776 12112 28782 12164
rect 29638 12112 29644 12164
rect 29696 12152 29702 12164
rect 30009 12155 30067 12161
rect 30009 12152 30021 12155
rect 29696 12124 30021 12152
rect 29696 12112 29702 12124
rect 30009 12121 30021 12124
rect 30055 12121 30067 12155
rect 31404 12152 31432 12180
rect 31234 12124 31800 12152
rect 30009 12115 30067 12121
rect 23799 12056 26188 12084
rect 23799 12053 23811 12056
rect 23753 12047 23811 12053
rect 26326 12044 26332 12096
rect 26384 12044 26390 12096
rect 27338 12044 27344 12096
rect 27396 12044 27402 12096
rect 30926 12044 30932 12096
rect 30984 12084 30990 12096
rect 31312 12084 31340 12124
rect 31772 12096 31800 12124
rect 32398 12112 32404 12164
rect 32456 12112 32462 12164
rect 34900 12152 34928 12180
rect 35066 12152 35072 12164
rect 33626 12124 34284 12152
rect 34900 12124 35072 12152
rect 30984 12056 31340 12084
rect 30984 12044 30990 12056
rect 31386 12044 31392 12096
rect 31444 12084 31450 12096
rect 31481 12087 31539 12093
rect 31481 12084 31493 12087
rect 31444 12056 31493 12084
rect 31444 12044 31450 12056
rect 31481 12053 31493 12056
rect 31527 12053 31539 12087
rect 31481 12047 31539 12053
rect 31754 12044 31760 12096
rect 31812 12084 31818 12096
rect 31849 12087 31907 12093
rect 31849 12084 31861 12087
rect 31812 12056 31861 12084
rect 31812 12044 31818 12056
rect 31849 12053 31861 12056
rect 31895 12084 31907 12087
rect 33318 12084 33324 12096
rect 31895 12056 33324 12084
rect 31895 12053 31907 12056
rect 31849 12047 31907 12053
rect 33318 12044 33324 12056
rect 33376 12084 33382 12096
rect 33704 12084 33732 12124
rect 34256 12093 34284 12124
rect 35066 12112 35072 12124
rect 35124 12112 35130 12164
rect 36722 12152 36728 12164
rect 36386 12124 36728 12152
rect 33376 12056 33732 12084
rect 34241 12087 34299 12093
rect 33376 12044 33382 12056
rect 34241 12053 34253 12087
rect 34287 12084 34299 12087
rect 34330 12084 34336 12096
rect 34287 12056 34336 12084
rect 34287 12053 34299 12056
rect 34241 12047 34299 12053
rect 34330 12044 34336 12056
rect 34388 12084 34394 12096
rect 34425 12087 34483 12093
rect 34425 12084 34437 12087
rect 34388 12056 34437 12084
rect 34388 12044 34394 12056
rect 34425 12053 34437 12056
rect 34471 12084 34483 12087
rect 36464 12084 36492 12124
rect 36722 12112 36728 12124
rect 36780 12112 36786 12164
rect 37200 12152 37228 12260
rect 37458 12248 37464 12300
rect 37516 12288 37522 12300
rect 37553 12291 37611 12297
rect 37553 12288 37565 12291
rect 37516 12260 37565 12288
rect 37516 12248 37522 12260
rect 37553 12257 37565 12260
rect 37599 12257 37611 12291
rect 37553 12251 37611 12257
rect 37642 12248 37648 12300
rect 37700 12248 37706 12300
rect 37734 12248 37740 12300
rect 37792 12288 37798 12300
rect 38841 12291 38899 12297
rect 38841 12288 38853 12291
rect 37792 12260 38853 12288
rect 37792 12248 37798 12260
rect 38841 12257 38853 12260
rect 38887 12257 38899 12291
rect 38841 12251 38899 12257
rect 37274 12180 37280 12232
rect 37332 12220 37338 12232
rect 40972 12229 41000 12328
rect 41616 12229 41644 12328
rect 49142 12248 49148 12300
rect 49200 12248 49206 12300
rect 38749 12223 38807 12229
rect 38749 12220 38761 12223
rect 37332 12192 38761 12220
rect 37332 12180 37338 12192
rect 38749 12189 38761 12192
rect 38795 12189 38807 12223
rect 39393 12223 39451 12229
rect 39393 12220 39405 12223
rect 38749 12183 38807 12189
rect 38856 12192 39405 12220
rect 38856 12152 38884 12192
rect 39393 12189 39405 12192
rect 39439 12220 39451 12223
rect 40129 12223 40187 12229
rect 40129 12220 40141 12223
rect 39439 12192 40141 12220
rect 39439 12189 39451 12192
rect 39393 12183 39451 12189
rect 40129 12189 40141 12192
rect 40175 12189 40187 12223
rect 40129 12183 40187 12189
rect 40957 12223 41015 12229
rect 40957 12189 40969 12223
rect 41003 12189 41015 12223
rect 40957 12183 41015 12189
rect 41601 12223 41659 12229
rect 41601 12189 41613 12223
rect 41647 12189 41659 12223
rect 46109 12223 46167 12229
rect 46109 12220 46121 12223
rect 41601 12183 41659 12189
rect 45526 12192 46121 12220
rect 37200 12124 38884 12152
rect 39298 12112 39304 12164
rect 39356 12152 39362 12164
rect 39577 12155 39635 12161
rect 39577 12152 39589 12155
rect 39356 12124 39589 12152
rect 39356 12112 39362 12124
rect 39577 12121 39589 12124
rect 39623 12121 39635 12155
rect 39577 12115 39635 12121
rect 40313 12155 40371 12161
rect 40313 12121 40325 12155
rect 40359 12152 40371 12155
rect 43346 12152 43352 12164
rect 40359 12124 43352 12152
rect 40359 12121 40371 12124
rect 40313 12115 40371 12121
rect 43346 12112 43352 12124
rect 43404 12112 43410 12164
rect 34471 12056 36492 12084
rect 34471 12053 34483 12056
rect 34425 12047 34483 12053
rect 36538 12044 36544 12096
rect 36596 12084 36602 12096
rect 36633 12087 36691 12093
rect 36633 12084 36645 12087
rect 36596 12056 36645 12084
rect 36596 12044 36602 12056
rect 36633 12053 36645 12056
rect 36679 12084 36691 12087
rect 36814 12084 36820 12096
rect 36679 12056 36820 12084
rect 36679 12053 36691 12056
rect 36633 12047 36691 12053
rect 36814 12044 36820 12056
rect 36872 12044 36878 12096
rect 37458 12044 37464 12096
rect 37516 12044 37522 12096
rect 38654 12044 38660 12096
rect 38712 12044 38718 12096
rect 40770 12044 40776 12096
rect 40828 12044 40834 12096
rect 41417 12087 41475 12093
rect 41417 12053 41429 12087
rect 41463 12084 41475 12087
rect 45526 12084 45554 12192
rect 46109 12189 46121 12192
rect 46155 12189 46167 12223
rect 46109 12183 46167 12189
rect 47946 12180 47952 12232
rect 48004 12180 48010 12232
rect 41463 12056 45554 12084
rect 41463 12053 41475 12056
rect 41417 12047 41475 12053
rect 45922 12044 45928 12096
rect 45980 12044 45986 12096
rect 1104 11994 49864 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 27950 11994
rect 28002 11942 28014 11994
rect 28066 11942 28078 11994
rect 28130 11942 28142 11994
rect 28194 11942 28206 11994
rect 28258 11942 37950 11994
rect 38002 11942 38014 11994
rect 38066 11942 38078 11994
rect 38130 11942 38142 11994
rect 38194 11942 38206 11994
rect 38258 11942 47950 11994
rect 48002 11942 48014 11994
rect 48066 11942 48078 11994
rect 48130 11942 48142 11994
rect 48194 11942 48206 11994
rect 48258 11942 49864 11994
rect 1104 11920 49864 11942
rect 2317 11883 2375 11889
rect 2317 11849 2329 11883
rect 2363 11880 2375 11883
rect 4154 11880 4160 11892
rect 2363 11852 4160 11880
rect 2363 11849 2375 11852
rect 2317 11843 2375 11849
rect 4154 11840 4160 11852
rect 4212 11840 4218 11892
rect 11609 11883 11667 11889
rect 11609 11849 11621 11883
rect 11655 11880 11667 11883
rect 11698 11880 11704 11892
rect 11655 11852 11704 11880
rect 11655 11849 11667 11852
rect 11609 11843 11667 11849
rect 11698 11840 11704 11852
rect 11756 11840 11762 11892
rect 12158 11840 12164 11892
rect 12216 11880 12222 11892
rect 12713 11883 12771 11889
rect 12713 11880 12725 11883
rect 12216 11852 12725 11880
rect 12216 11840 12222 11852
rect 12713 11849 12725 11852
rect 12759 11849 12771 11883
rect 12713 11843 12771 11849
rect 13262 11840 13268 11892
rect 13320 11880 13326 11892
rect 13541 11883 13599 11889
rect 13541 11880 13553 11883
rect 13320 11852 13553 11880
rect 13320 11840 13326 11852
rect 13541 11849 13553 11852
rect 13587 11849 13599 11883
rect 13541 11843 13599 11849
rect 13630 11840 13636 11892
rect 13688 11880 13694 11892
rect 14369 11883 14427 11889
rect 14369 11880 14381 11883
rect 13688 11852 14381 11880
rect 13688 11840 13694 11852
rect 14369 11849 14381 11852
rect 14415 11849 14427 11883
rect 15562 11880 15568 11892
rect 14369 11843 14427 11849
rect 15304 11852 15568 11880
rect 12805 11815 12863 11821
rect 12805 11781 12817 11815
rect 12851 11812 12863 11815
rect 14182 11812 14188 11824
rect 12851 11784 14188 11812
rect 12851 11781 12863 11784
rect 12805 11775 12863 11781
rect 14182 11772 14188 11784
rect 14240 11772 14246 11824
rect 14277 11815 14335 11821
rect 14277 11781 14289 11815
rect 14323 11812 14335 11815
rect 15194 11812 15200 11824
rect 14323 11784 15200 11812
rect 14323 11781 14335 11784
rect 14277 11775 14335 11781
rect 15194 11772 15200 11784
rect 15252 11772 15258 11824
rect 1210 11704 1216 11756
rect 1268 11744 1274 11756
rect 1581 11747 1639 11753
rect 1581 11744 1593 11747
rect 1268 11716 1593 11744
rect 1268 11704 1274 11716
rect 1581 11713 1593 11716
rect 1627 11713 1639 11747
rect 1581 11707 1639 11713
rect 2501 11747 2559 11753
rect 2501 11713 2513 11747
rect 2547 11713 2559 11747
rect 11882 11744 11888 11756
rect 2501 11707 2559 11713
rect 6886 11716 11888 11744
rect 1302 11636 1308 11688
rect 1360 11676 1366 11688
rect 2516 11676 2544 11707
rect 2777 11679 2835 11685
rect 2777 11676 2789 11679
rect 1360 11648 2789 11676
rect 1360 11636 1366 11648
rect 2777 11645 2789 11648
rect 2823 11645 2835 11679
rect 2777 11639 2835 11645
rect 1765 11611 1823 11617
rect 1765 11577 1777 11611
rect 1811 11608 1823 11611
rect 6886 11608 6914 11716
rect 11882 11704 11888 11716
rect 11940 11704 11946 11756
rect 15304 11744 15332 11852
rect 15562 11840 15568 11852
rect 15620 11840 15626 11892
rect 16390 11840 16396 11892
rect 16448 11840 16454 11892
rect 18782 11840 18788 11892
rect 18840 11880 18846 11892
rect 19242 11880 19248 11892
rect 18840 11852 19248 11880
rect 18840 11840 18846 11852
rect 19242 11840 19248 11852
rect 19300 11880 19306 11892
rect 19300 11852 22324 11880
rect 19300 11840 19306 11852
rect 16408 11812 16436 11840
rect 19153 11815 19211 11821
rect 16408 11784 17618 11812
rect 19153 11781 19165 11815
rect 19199 11812 19211 11815
rect 19334 11812 19340 11824
rect 19199 11784 19340 11812
rect 19199 11781 19211 11784
rect 19153 11775 19211 11781
rect 19334 11772 19340 11784
rect 19392 11772 19398 11824
rect 19886 11772 19892 11824
rect 19944 11772 19950 11824
rect 19981 11815 20039 11821
rect 19981 11781 19993 11815
rect 20027 11812 20039 11815
rect 20070 11812 20076 11824
rect 20027 11784 20076 11812
rect 20027 11781 20039 11784
rect 19981 11775 20039 11781
rect 12406 11716 12940 11744
rect 11238 11636 11244 11688
rect 11296 11676 11302 11688
rect 12250 11676 12256 11688
rect 11296 11648 12256 11676
rect 11296 11636 11302 11648
rect 12250 11636 12256 11648
rect 12308 11676 12314 11688
rect 12406 11676 12434 11716
rect 12912 11685 12940 11716
rect 14476 11716 15332 11744
rect 15473 11747 15531 11753
rect 12308 11648 12434 11676
rect 12897 11679 12955 11685
rect 12308 11636 12314 11648
rect 12897 11645 12909 11679
rect 12943 11645 12955 11679
rect 12897 11639 12955 11645
rect 13449 11679 13507 11685
rect 13449 11645 13461 11679
rect 13495 11676 13507 11679
rect 14476 11676 14504 11716
rect 15473 11713 15485 11747
rect 15519 11744 15531 11747
rect 15930 11744 15936 11756
rect 15519 11716 15936 11744
rect 15519 11713 15531 11716
rect 15473 11707 15531 11713
rect 15930 11704 15936 11716
rect 15988 11704 15994 11756
rect 19061 11747 19119 11753
rect 19061 11713 19073 11747
rect 19107 11744 19119 11747
rect 19996 11744 20024 11775
rect 20070 11772 20076 11784
rect 20128 11772 20134 11824
rect 22186 11812 22192 11824
rect 20548 11784 22192 11812
rect 19107 11716 20024 11744
rect 19107 11713 19119 11716
rect 19061 11707 19119 11713
rect 13495 11648 14504 11676
rect 14553 11679 14611 11685
rect 13495 11645 13507 11648
rect 13449 11639 13507 11645
rect 14553 11645 14565 11679
rect 14599 11645 14611 11679
rect 14553 11639 14611 11645
rect 1811 11580 6914 11608
rect 1811 11577 1823 11580
rect 1765 11571 1823 11577
rect 11790 11568 11796 11620
rect 11848 11608 11854 11620
rect 13464 11608 13492 11639
rect 11848 11580 13492 11608
rect 11848 11568 11854 11580
rect 14458 11568 14464 11620
rect 14516 11608 14522 11620
rect 14568 11608 14596 11639
rect 14734 11636 14740 11688
rect 14792 11676 14798 11688
rect 15657 11679 15715 11685
rect 15657 11676 15669 11679
rect 14792 11648 15669 11676
rect 14792 11636 14798 11648
rect 15657 11645 15669 11648
rect 15703 11645 15715 11679
rect 15657 11639 15715 11645
rect 16758 11636 16764 11688
rect 16816 11676 16822 11688
rect 16853 11679 16911 11685
rect 16853 11676 16865 11679
rect 16816 11648 16865 11676
rect 16816 11636 16822 11648
rect 16853 11645 16865 11648
rect 16899 11645 16911 11679
rect 16853 11639 16911 11645
rect 17129 11679 17187 11685
rect 17129 11645 17141 11679
rect 17175 11676 17187 11679
rect 20165 11679 20223 11685
rect 17175 11648 19472 11676
rect 17175 11645 17187 11648
rect 17129 11639 17187 11645
rect 14516 11580 14596 11608
rect 14752 11580 15608 11608
rect 14516 11568 14522 11580
rect 12345 11543 12403 11549
rect 12345 11509 12357 11543
rect 12391 11540 12403 11543
rect 12526 11540 12532 11552
rect 12391 11512 12532 11540
rect 12391 11509 12403 11512
rect 12345 11503 12403 11509
rect 12526 11500 12532 11512
rect 12584 11500 12590 11552
rect 13909 11543 13967 11549
rect 13909 11509 13921 11543
rect 13955 11540 13967 11543
rect 14752 11540 14780 11580
rect 13955 11512 14780 11540
rect 13955 11509 13967 11512
rect 13909 11503 13967 11509
rect 14826 11500 14832 11552
rect 14884 11540 14890 11552
rect 15105 11543 15163 11549
rect 15105 11540 15117 11543
rect 14884 11512 15117 11540
rect 14884 11500 14890 11512
rect 15105 11509 15117 11512
rect 15151 11509 15163 11543
rect 15580 11540 15608 11580
rect 16206 11568 16212 11620
rect 16264 11608 16270 11620
rect 16301 11611 16359 11617
rect 16301 11608 16313 11611
rect 16264 11580 16313 11608
rect 16264 11568 16270 11580
rect 16301 11577 16313 11580
rect 16347 11608 16359 11611
rect 16347 11580 16988 11608
rect 16347 11577 16359 11580
rect 16301 11571 16359 11577
rect 15654 11540 15660 11552
rect 15580 11512 15660 11540
rect 15105 11503 15163 11509
rect 15654 11500 15660 11512
rect 15712 11500 15718 11552
rect 16960 11540 16988 11580
rect 18138 11540 18144 11552
rect 16960 11512 18144 11540
rect 18138 11500 18144 11512
rect 18196 11500 18202 11552
rect 18230 11500 18236 11552
rect 18288 11540 18294 11552
rect 18601 11543 18659 11549
rect 18601 11540 18613 11543
rect 18288 11512 18613 11540
rect 18288 11500 18294 11512
rect 18601 11509 18613 11512
rect 18647 11509 18659 11543
rect 19444 11540 19472 11648
rect 20165 11645 20177 11679
rect 20211 11676 20223 11679
rect 20548 11676 20576 11784
rect 22186 11772 22192 11784
rect 22244 11772 22250 11824
rect 21085 11747 21143 11753
rect 21085 11713 21097 11747
rect 21131 11744 21143 11747
rect 21358 11744 21364 11756
rect 21131 11716 21364 11744
rect 21131 11713 21143 11716
rect 21085 11707 21143 11713
rect 21358 11704 21364 11716
rect 21416 11704 21422 11756
rect 21634 11704 21640 11756
rect 21692 11744 21698 11756
rect 21821 11747 21879 11753
rect 21821 11744 21833 11747
rect 21692 11716 21833 11744
rect 21692 11704 21698 11716
rect 21821 11713 21833 11716
rect 21867 11713 21879 11747
rect 21821 11707 21879 11713
rect 22094 11704 22100 11756
rect 22152 11704 22158 11756
rect 22296 11753 22324 11852
rect 24486 11840 24492 11892
rect 24544 11880 24550 11892
rect 25685 11883 25743 11889
rect 25685 11880 25697 11883
rect 24544 11852 25697 11880
rect 24544 11840 24550 11852
rect 25685 11849 25697 11852
rect 25731 11849 25743 11883
rect 25685 11843 25743 11849
rect 26421 11883 26479 11889
rect 26421 11849 26433 11883
rect 26467 11880 26479 11883
rect 27338 11880 27344 11892
rect 26467 11852 27344 11880
rect 26467 11849 26479 11852
rect 26421 11843 26479 11849
rect 27338 11840 27344 11852
rect 27396 11840 27402 11892
rect 27522 11840 27528 11892
rect 27580 11880 27586 11892
rect 27617 11883 27675 11889
rect 27617 11880 27629 11883
rect 27580 11852 27629 11880
rect 27580 11840 27586 11852
rect 27617 11849 27629 11852
rect 27663 11849 27675 11883
rect 27617 11843 27675 11849
rect 30745 11883 30803 11889
rect 30745 11849 30757 11883
rect 30791 11880 30803 11883
rect 31570 11880 31576 11892
rect 30791 11852 31576 11880
rect 30791 11849 30803 11852
rect 30745 11843 30803 11849
rect 31570 11840 31576 11852
rect 31628 11840 31634 11892
rect 31754 11840 31760 11892
rect 31812 11840 31818 11892
rect 32122 11840 32128 11892
rect 32180 11880 32186 11892
rect 32677 11883 32735 11889
rect 32677 11880 32689 11883
rect 32180 11852 32689 11880
rect 32180 11840 32186 11852
rect 32677 11849 32689 11852
rect 32723 11849 32735 11883
rect 32677 11843 32735 11849
rect 33686 11840 33692 11892
rect 33744 11880 33750 11892
rect 33873 11883 33931 11889
rect 33873 11880 33885 11883
rect 33744 11852 33885 11880
rect 33744 11840 33750 11852
rect 33873 11849 33885 11852
rect 33919 11849 33931 11883
rect 33873 11843 33931 11849
rect 34790 11840 34796 11892
rect 34848 11880 34854 11892
rect 35342 11880 35348 11892
rect 34848 11852 35348 11880
rect 34848 11840 34854 11852
rect 35342 11840 35348 11852
rect 35400 11840 35406 11892
rect 36078 11840 36084 11892
rect 36136 11880 36142 11892
rect 36909 11883 36967 11889
rect 36909 11880 36921 11883
rect 36136 11852 36921 11880
rect 36136 11840 36142 11852
rect 36909 11849 36921 11852
rect 36955 11880 36967 11883
rect 37734 11880 37740 11892
rect 36955 11852 37740 11880
rect 36955 11849 36967 11852
rect 36909 11843 36967 11849
rect 37734 11840 37740 11852
rect 37792 11840 37798 11892
rect 37826 11840 37832 11892
rect 37884 11880 37890 11892
rect 37921 11883 37979 11889
rect 37921 11880 37933 11883
rect 37884 11852 37933 11880
rect 37884 11840 37890 11852
rect 37921 11849 37933 11852
rect 37967 11849 37979 11883
rect 37921 11843 37979 11849
rect 38654 11840 38660 11892
rect 38712 11840 38718 11892
rect 22646 11772 22652 11824
rect 22704 11812 22710 11824
rect 24213 11815 24271 11821
rect 24213 11812 24225 11815
rect 22704 11784 24225 11812
rect 22704 11772 22710 11784
rect 24213 11781 24225 11784
rect 24259 11812 24271 11815
rect 24302 11812 24308 11824
rect 24259 11784 24308 11812
rect 24259 11781 24271 11784
rect 24213 11775 24271 11781
rect 24302 11772 24308 11784
rect 24360 11772 24366 11824
rect 25958 11812 25964 11824
rect 25438 11784 25964 11812
rect 25958 11772 25964 11784
rect 26016 11772 26022 11824
rect 28810 11812 28816 11824
rect 27632 11784 28816 11812
rect 22281 11747 22339 11753
rect 22281 11713 22293 11747
rect 22327 11744 22339 11747
rect 22554 11744 22560 11756
rect 22327 11716 22560 11744
rect 22327 11713 22339 11716
rect 22281 11707 22339 11713
rect 22554 11704 22560 11716
rect 22612 11704 22618 11756
rect 26142 11704 26148 11756
rect 26200 11744 26206 11756
rect 27338 11744 27344 11756
rect 26200 11716 27344 11744
rect 26200 11704 26206 11716
rect 27338 11704 27344 11716
rect 27396 11744 27402 11756
rect 27525 11747 27583 11753
rect 27525 11744 27537 11747
rect 27396 11716 27537 11744
rect 27396 11704 27402 11716
rect 27525 11713 27537 11716
rect 27571 11713 27583 11747
rect 27525 11707 27583 11713
rect 20211 11648 20576 11676
rect 20211 11645 20223 11648
rect 20165 11639 20223 11645
rect 20622 11636 20628 11688
rect 20680 11676 20686 11688
rect 21177 11679 21235 11685
rect 21177 11676 21189 11679
rect 20680 11648 21189 11676
rect 20680 11636 20686 11648
rect 21177 11645 21189 11648
rect 21223 11645 21235 11679
rect 21177 11639 21235 11645
rect 21269 11679 21327 11685
rect 21269 11645 21281 11679
rect 21315 11645 21327 11679
rect 21269 11639 21327 11645
rect 19521 11611 19579 11617
rect 19521 11577 19533 11611
rect 19567 11608 19579 11611
rect 20070 11608 20076 11620
rect 19567 11580 20076 11608
rect 19567 11577 19579 11580
rect 19521 11571 19579 11577
rect 20070 11568 20076 11580
rect 20128 11568 20134 11620
rect 20717 11611 20775 11617
rect 20717 11577 20729 11611
rect 20763 11608 20775 11611
rect 20806 11608 20812 11620
rect 20763 11580 20812 11608
rect 20763 11577 20775 11580
rect 20717 11571 20775 11577
rect 20806 11568 20812 11580
rect 20864 11568 20870 11620
rect 21284 11608 21312 11639
rect 21450 11636 21456 11688
rect 21508 11676 21514 11688
rect 22002 11676 22008 11688
rect 21508 11648 22008 11676
rect 21508 11636 21514 11648
rect 22002 11636 22008 11648
rect 22060 11676 22066 11688
rect 23385 11679 23443 11685
rect 23385 11676 23397 11679
rect 22060 11648 23397 11676
rect 22060 11636 22066 11648
rect 23385 11645 23397 11648
rect 23431 11676 23443 11679
rect 23474 11676 23480 11688
rect 23431 11648 23480 11676
rect 23431 11645 23443 11648
rect 23385 11639 23443 11645
rect 23474 11636 23480 11648
rect 23532 11676 23538 11688
rect 23842 11676 23848 11688
rect 23532 11648 23848 11676
rect 23532 11636 23538 11648
rect 23842 11636 23848 11648
rect 23900 11676 23906 11688
rect 23937 11679 23995 11685
rect 23937 11676 23949 11679
rect 23900 11648 23949 11676
rect 23900 11636 23906 11648
rect 23937 11645 23949 11648
rect 23983 11645 23995 11679
rect 23937 11639 23995 11645
rect 24302 11636 24308 11688
rect 24360 11676 24366 11688
rect 26326 11676 26332 11688
rect 24360 11648 26332 11676
rect 24360 11636 24366 11648
rect 26326 11636 26332 11648
rect 26384 11636 26390 11688
rect 27632 11676 27660 11784
rect 28810 11772 28816 11784
rect 28868 11772 28874 11824
rect 30006 11812 30012 11824
rect 29946 11784 30012 11812
rect 30006 11772 30012 11784
rect 30064 11812 30070 11824
rect 30926 11812 30932 11824
rect 30064 11784 30932 11812
rect 30064 11772 30070 11784
rect 30926 11772 30932 11784
rect 30984 11772 30990 11824
rect 31386 11812 31392 11824
rect 31036 11784 31392 11812
rect 27172 11648 27660 11676
rect 27709 11679 27767 11685
rect 21542 11608 21548 11620
rect 21284 11580 21548 11608
rect 21542 11568 21548 11580
rect 21600 11568 21606 11620
rect 21726 11568 21732 11620
rect 21784 11608 21790 11620
rect 23566 11608 23572 11620
rect 21784 11580 21956 11608
rect 21784 11568 21790 11580
rect 21174 11540 21180 11552
rect 19444 11512 21180 11540
rect 18601 11503 18659 11509
rect 21174 11500 21180 11512
rect 21232 11540 21238 11552
rect 21634 11540 21640 11552
rect 21232 11512 21640 11540
rect 21232 11500 21238 11512
rect 21634 11500 21640 11512
rect 21692 11500 21698 11552
rect 21928 11540 21956 11580
rect 22066 11580 23572 11608
rect 22066 11540 22094 11580
rect 23566 11568 23572 11580
rect 23624 11568 23630 11620
rect 27172 11617 27200 11648
rect 27709 11645 27721 11679
rect 27755 11645 27767 11679
rect 27709 11639 27767 11645
rect 28445 11679 28503 11685
rect 28445 11645 28457 11679
rect 28491 11645 28503 11679
rect 28445 11639 28503 11645
rect 28721 11679 28779 11685
rect 28721 11645 28733 11679
rect 28767 11676 28779 11679
rect 31036 11676 31064 11784
rect 31386 11772 31392 11784
rect 31444 11812 31450 11824
rect 36722 11812 36728 11824
rect 31444 11784 34100 11812
rect 36662 11784 36728 11812
rect 31444 11772 31450 11784
rect 31110 11704 31116 11756
rect 31168 11704 31174 11756
rect 28767 11648 31064 11676
rect 28767 11645 28779 11648
rect 28721 11639 28779 11645
rect 27157 11611 27215 11617
rect 27157 11577 27169 11611
rect 27203 11577 27215 11611
rect 27157 11571 27215 11577
rect 27246 11568 27252 11620
rect 27304 11608 27310 11620
rect 27724 11608 27752 11639
rect 27304 11580 27752 11608
rect 27304 11568 27310 11580
rect 21928 11512 22094 11540
rect 28460 11540 28488 11639
rect 31202 11636 31208 11688
rect 31260 11636 31266 11688
rect 31294 11636 31300 11688
rect 31352 11636 31358 11688
rect 31478 11636 31484 11688
rect 31536 11676 31542 11688
rect 32769 11679 32827 11685
rect 32769 11676 32781 11679
rect 31536 11648 32781 11676
rect 31536 11636 31542 11648
rect 32769 11645 32781 11648
rect 32815 11645 32827 11679
rect 32769 11639 32827 11645
rect 32858 11636 32864 11688
rect 32916 11636 32922 11688
rect 34072 11685 34100 11784
rect 36722 11772 36728 11784
rect 36780 11772 36786 11824
rect 37366 11772 37372 11824
rect 37424 11812 37430 11824
rect 39117 11815 39175 11821
rect 39117 11812 39129 11815
rect 37424 11784 39129 11812
rect 37424 11772 37430 11784
rect 39117 11781 39129 11784
rect 39163 11781 39175 11815
rect 39117 11775 39175 11781
rect 40770 11772 40776 11824
rect 40828 11812 40834 11824
rect 45097 11815 45155 11821
rect 45097 11812 45109 11815
rect 40828 11784 45109 11812
rect 40828 11772 40834 11784
rect 45097 11781 45109 11784
rect 45143 11781 45155 11815
rect 45097 11775 45155 11781
rect 49142 11772 49148 11824
rect 49200 11772 49206 11824
rect 36906 11704 36912 11756
rect 36964 11744 36970 11756
rect 37829 11747 37887 11753
rect 37829 11744 37841 11747
rect 36964 11716 37841 11744
rect 36964 11704 36970 11716
rect 37829 11713 37841 11716
rect 37875 11713 37887 11747
rect 37829 11707 37887 11713
rect 39022 11704 39028 11756
rect 39080 11704 39086 11756
rect 39942 11704 39948 11756
rect 40000 11744 40006 11756
rect 40405 11747 40463 11753
rect 40405 11744 40417 11747
rect 40000 11716 40417 11744
rect 40000 11704 40006 11716
rect 40405 11713 40417 11716
rect 40451 11713 40463 11747
rect 40405 11707 40463 11713
rect 45922 11704 45928 11756
rect 45980 11744 45986 11756
rect 47949 11747 48007 11753
rect 47949 11744 47961 11747
rect 45980 11716 47961 11744
rect 45980 11704 45986 11716
rect 47949 11713 47961 11716
rect 47995 11713 48007 11747
rect 47949 11707 48007 11713
rect 33965 11679 34023 11685
rect 33965 11645 33977 11679
rect 34011 11645 34023 11679
rect 33965 11639 34023 11645
rect 34057 11679 34115 11685
rect 34057 11645 34069 11679
rect 34103 11645 34115 11679
rect 34057 11639 34115 11645
rect 30558 11568 30564 11620
rect 30616 11608 30622 11620
rect 33980 11608 34008 11639
rect 35066 11636 35072 11688
rect 35124 11676 35130 11688
rect 35161 11679 35219 11685
rect 35161 11676 35173 11679
rect 35124 11648 35173 11676
rect 35124 11636 35130 11648
rect 35161 11645 35173 11648
rect 35207 11645 35219 11679
rect 35161 11639 35219 11645
rect 35437 11679 35495 11685
rect 35437 11645 35449 11679
rect 35483 11676 35495 11679
rect 35483 11648 36584 11676
rect 35483 11645 35495 11648
rect 35437 11639 35495 11645
rect 30616 11580 34008 11608
rect 36556 11608 36584 11648
rect 36630 11636 36636 11688
rect 36688 11676 36694 11688
rect 38013 11679 38071 11685
rect 38013 11676 38025 11679
rect 36688 11648 38025 11676
rect 36688 11636 36694 11648
rect 38013 11645 38025 11648
rect 38059 11645 38071 11679
rect 38013 11639 38071 11645
rect 39209 11679 39267 11685
rect 39209 11645 39221 11679
rect 39255 11645 39267 11679
rect 39209 11639 39267 11645
rect 36814 11608 36820 11620
rect 36556 11580 36820 11608
rect 30616 11568 30622 11580
rect 36814 11568 36820 11580
rect 36872 11608 36878 11620
rect 39224 11608 39252 11639
rect 36872 11580 39252 11608
rect 40129 11611 40187 11617
rect 36872 11568 36878 11580
rect 40129 11577 40141 11611
rect 40175 11608 40187 11611
rect 43714 11608 43720 11620
rect 40175 11580 43720 11608
rect 40175 11577 40187 11580
rect 40129 11571 40187 11577
rect 43714 11568 43720 11580
rect 43772 11568 43778 11620
rect 45281 11611 45339 11617
rect 45281 11577 45293 11611
rect 45327 11608 45339 11611
rect 46290 11608 46296 11620
rect 45327 11580 46296 11608
rect 45327 11577 45339 11580
rect 45281 11571 45339 11577
rect 46290 11568 46296 11580
rect 46348 11568 46354 11620
rect 29454 11540 29460 11552
rect 28460 11512 29460 11540
rect 29454 11500 29460 11512
rect 29512 11500 29518 11552
rect 30098 11500 30104 11552
rect 30156 11540 30162 11552
rect 30193 11543 30251 11549
rect 30193 11540 30205 11543
rect 30156 11512 30205 11540
rect 30156 11500 30162 11512
rect 30193 11509 30205 11512
rect 30239 11509 30251 11543
rect 30193 11503 30251 11509
rect 32309 11543 32367 11549
rect 32309 11509 32321 11543
rect 32355 11540 32367 11543
rect 33410 11540 33416 11552
rect 32355 11512 33416 11540
rect 32355 11509 32367 11512
rect 32309 11503 32367 11509
rect 33410 11500 33416 11512
rect 33468 11500 33474 11552
rect 33505 11543 33563 11549
rect 33505 11509 33517 11543
rect 33551 11540 33563 11543
rect 37366 11540 37372 11552
rect 33551 11512 37372 11540
rect 33551 11509 33563 11512
rect 33505 11503 33563 11509
rect 37366 11500 37372 11512
rect 37424 11500 37430 11552
rect 37461 11543 37519 11549
rect 37461 11509 37473 11543
rect 37507 11540 37519 11543
rect 40218 11540 40224 11552
rect 37507 11512 40224 11540
rect 37507 11509 37519 11512
rect 37461 11503 37519 11509
rect 40218 11500 40224 11512
rect 40276 11500 40282 11552
rect 1104 11450 49864 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 32950 11450
rect 33002 11398 33014 11450
rect 33066 11398 33078 11450
rect 33130 11398 33142 11450
rect 33194 11398 33206 11450
rect 33258 11398 42950 11450
rect 43002 11398 43014 11450
rect 43066 11398 43078 11450
rect 43130 11398 43142 11450
rect 43194 11398 43206 11450
rect 43258 11398 49864 11450
rect 1104 11376 49864 11398
rect 1210 11296 1216 11348
rect 1268 11336 1274 11348
rect 2133 11339 2191 11345
rect 2133 11336 2145 11339
rect 1268 11308 2145 11336
rect 1268 11296 1274 11308
rect 2133 11305 2145 11308
rect 2179 11305 2191 11339
rect 2133 11299 2191 11305
rect 12434 11296 12440 11348
rect 12492 11336 12498 11348
rect 13173 11339 13231 11345
rect 13173 11336 13185 11339
rect 12492 11308 13185 11336
rect 12492 11296 12498 11308
rect 13173 11305 13185 11308
rect 13219 11305 13231 11339
rect 13173 11299 13231 11305
rect 13446 11296 13452 11348
rect 13504 11336 13510 11348
rect 14369 11339 14427 11345
rect 14369 11336 14381 11339
rect 13504 11308 14381 11336
rect 13504 11296 13510 11308
rect 14369 11305 14381 11308
rect 14415 11305 14427 11339
rect 14369 11299 14427 11305
rect 16666 11296 16672 11348
rect 16724 11336 16730 11348
rect 16761 11339 16819 11345
rect 16761 11336 16773 11339
rect 16724 11308 16773 11336
rect 16724 11296 16730 11308
rect 16761 11305 16773 11308
rect 16807 11305 16819 11339
rect 16761 11299 16819 11305
rect 19061 11339 19119 11345
rect 19061 11305 19073 11339
rect 19107 11336 19119 11339
rect 19242 11336 19248 11348
rect 19107 11308 19248 11336
rect 19107 11305 19119 11308
rect 19061 11299 19119 11305
rect 19242 11296 19248 11308
rect 19300 11296 19306 11348
rect 19521 11339 19579 11345
rect 19521 11305 19533 11339
rect 19567 11336 19579 11339
rect 19886 11336 19892 11348
rect 19567 11308 19892 11336
rect 19567 11305 19579 11308
rect 19521 11299 19579 11305
rect 19886 11296 19892 11308
rect 19944 11296 19950 11348
rect 20704 11339 20762 11345
rect 20704 11305 20716 11339
rect 20750 11336 20762 11339
rect 21726 11336 21732 11348
rect 20750 11308 21732 11336
rect 20750 11305 20762 11308
rect 20704 11299 20762 11305
rect 21726 11296 21732 11308
rect 21784 11296 21790 11348
rect 22002 11296 22008 11348
rect 22060 11336 22066 11348
rect 22462 11336 22468 11348
rect 22060 11308 22468 11336
rect 22060 11296 22066 11308
rect 22462 11296 22468 11308
rect 22520 11296 22526 11348
rect 22554 11296 22560 11348
rect 22612 11336 22618 11348
rect 24394 11336 24400 11348
rect 22612 11308 24400 11336
rect 22612 11296 22618 11308
rect 24394 11296 24400 11308
rect 24452 11336 24458 11348
rect 28902 11336 28908 11348
rect 24452 11308 28908 11336
rect 24452 11296 24458 11308
rect 28902 11296 28908 11308
rect 28960 11296 28966 11348
rect 29733 11339 29791 11345
rect 29733 11305 29745 11339
rect 29779 11336 29791 11339
rect 29779 11308 33364 11336
rect 29779 11305 29791 11308
rect 29733 11299 29791 11305
rect 1762 11228 1768 11280
rect 1820 11228 1826 11280
rect 12710 11228 12716 11280
rect 12768 11228 12774 11280
rect 14642 11228 14648 11280
rect 14700 11268 14706 11280
rect 15565 11271 15623 11277
rect 14700 11240 14964 11268
rect 14700 11228 14706 11240
rect 10965 11203 11023 11209
rect 10965 11169 10977 11203
rect 11011 11200 11023 11203
rect 13814 11200 13820 11212
rect 11011 11172 13820 11200
rect 11011 11169 11023 11172
rect 10965 11163 11023 11169
rect 13814 11160 13820 11172
rect 13872 11160 13878 11212
rect 14826 11160 14832 11212
rect 14884 11160 14890 11212
rect 14936 11209 14964 11240
rect 15565 11237 15577 11271
rect 15611 11268 15623 11271
rect 18782 11268 18788 11280
rect 15611 11240 18788 11268
rect 15611 11237 15623 11240
rect 15565 11231 15623 11237
rect 18782 11228 18788 11240
rect 18840 11228 18846 11280
rect 22189 11271 22247 11277
rect 22189 11268 22201 11271
rect 21744 11240 22201 11268
rect 21744 11212 21772 11240
rect 22189 11237 22201 11240
rect 22235 11237 22247 11271
rect 22189 11231 22247 11237
rect 23293 11271 23351 11277
rect 23293 11237 23305 11271
rect 23339 11268 23351 11271
rect 23382 11268 23388 11280
rect 23339 11240 23388 11268
rect 23339 11237 23351 11240
rect 23293 11231 23351 11237
rect 23382 11228 23388 11240
rect 23440 11228 23446 11280
rect 26329 11271 26387 11277
rect 26329 11237 26341 11271
rect 26375 11268 26387 11271
rect 26602 11268 26608 11280
rect 26375 11240 26608 11268
rect 26375 11237 26387 11240
rect 26329 11231 26387 11237
rect 26602 11228 26608 11240
rect 26660 11228 26666 11280
rect 28442 11228 28448 11280
rect 28500 11268 28506 11280
rect 28629 11271 28687 11277
rect 28629 11268 28641 11271
rect 28500 11240 28641 11268
rect 28500 11228 28506 11240
rect 28629 11237 28641 11240
rect 28675 11237 28687 11271
rect 28629 11231 28687 11237
rect 29089 11271 29147 11277
rect 29089 11237 29101 11271
rect 29135 11268 29147 11271
rect 29365 11271 29423 11277
rect 29365 11268 29377 11271
rect 29135 11240 29377 11268
rect 29135 11237 29147 11240
rect 29089 11231 29147 11237
rect 14921 11203 14979 11209
rect 14921 11169 14933 11203
rect 14967 11169 14979 11203
rect 14921 11163 14979 11169
rect 15470 11160 15476 11212
rect 15528 11200 15534 11212
rect 16025 11203 16083 11209
rect 16025 11200 16037 11203
rect 15528 11172 16037 11200
rect 15528 11160 15534 11172
rect 16025 11169 16037 11172
rect 16071 11169 16083 11203
rect 16025 11163 16083 11169
rect 16209 11203 16267 11209
rect 16209 11169 16221 11203
rect 16255 11200 16267 11203
rect 17034 11200 17040 11212
rect 16255 11172 17040 11200
rect 16255 11169 16267 11172
rect 16209 11163 16267 11169
rect 17034 11160 17040 11172
rect 17092 11160 17098 11212
rect 17405 11203 17463 11209
rect 17405 11169 17417 11203
rect 17451 11200 17463 11203
rect 17451 11172 18552 11200
rect 17451 11169 17463 11172
rect 17405 11163 17463 11169
rect 1578 11092 1584 11144
rect 1636 11132 1642 11144
rect 2317 11135 2375 11141
rect 2317 11132 2329 11135
rect 1636 11104 2329 11132
rect 1636 11092 1642 11104
rect 2317 11101 2329 11104
rect 2363 11101 2375 11135
rect 2317 11095 2375 11101
rect 12342 11092 12348 11144
rect 12400 11092 12406 11144
rect 12894 11092 12900 11144
rect 12952 11132 12958 11144
rect 12989 11135 13047 11141
rect 12989 11132 13001 11135
rect 12952 11104 13001 11132
rect 12952 11092 12958 11104
rect 12989 11101 13001 11104
rect 13035 11132 13047 11135
rect 14734 11132 14740 11144
rect 13035 11104 14740 11132
rect 13035 11101 13047 11104
rect 12989 11095 13047 11101
rect 14734 11092 14740 11104
rect 14792 11092 14798 11144
rect 17221 11135 17279 11141
rect 17221 11101 17233 11135
rect 17267 11132 17279 11135
rect 18322 11132 18328 11144
rect 17267 11104 18328 11132
rect 17267 11101 17279 11104
rect 17221 11095 17279 11101
rect 18322 11092 18328 11104
rect 18380 11092 18386 11144
rect 18414 11092 18420 11144
rect 18472 11092 18478 11144
rect 18524 11132 18552 11172
rect 18598 11160 18604 11212
rect 18656 11200 18662 11212
rect 18874 11200 18880 11212
rect 18656 11172 18880 11200
rect 18656 11160 18662 11172
rect 18874 11160 18880 11172
rect 18932 11160 18938 11212
rect 20441 11203 20499 11209
rect 20441 11169 20453 11203
rect 20487 11200 20499 11203
rect 21450 11200 21456 11212
rect 20487 11172 21456 11200
rect 20487 11169 20499 11172
rect 20441 11163 20499 11169
rect 21450 11160 21456 11172
rect 21508 11160 21514 11212
rect 21726 11160 21732 11212
rect 21784 11160 21790 11212
rect 23753 11203 23811 11209
rect 23753 11169 23765 11203
rect 23799 11200 23811 11203
rect 23842 11200 23848 11212
rect 23799 11172 23848 11200
rect 23799 11169 23811 11172
rect 23753 11163 23811 11169
rect 23842 11160 23848 11172
rect 23900 11160 23906 11212
rect 23937 11203 23995 11209
rect 23937 11169 23949 11203
rect 23983 11200 23995 11203
rect 24118 11200 24124 11212
rect 23983 11172 24124 11200
rect 23983 11169 23995 11172
rect 23937 11163 23995 11169
rect 24118 11160 24124 11172
rect 24176 11160 24182 11212
rect 24486 11160 24492 11212
rect 24544 11200 24550 11212
rect 24857 11203 24915 11209
rect 24857 11200 24869 11203
rect 24544 11172 24869 11200
rect 24544 11160 24550 11172
rect 24857 11169 24869 11172
rect 24903 11169 24915 11203
rect 24857 11163 24915 11169
rect 27157 11203 27215 11209
rect 27157 11169 27169 11203
rect 27203 11200 27215 11203
rect 29178 11200 29184 11212
rect 27203 11172 29184 11200
rect 27203 11169 27215 11172
rect 27157 11163 27215 11169
rect 29178 11160 29184 11172
rect 29236 11160 29242 11212
rect 19518 11132 19524 11144
rect 18524 11104 19524 11132
rect 19518 11092 19524 11104
rect 19576 11092 19582 11144
rect 23474 11092 23480 11144
rect 23532 11132 23538 11144
rect 24578 11132 24584 11144
rect 23532 11104 24584 11132
rect 23532 11092 23538 11104
rect 24578 11092 24584 11104
rect 24636 11092 24642 11144
rect 25958 11092 25964 11144
rect 26016 11092 26022 11144
rect 26881 11135 26939 11141
rect 26881 11101 26893 11135
rect 26927 11101 26939 11135
rect 26881 11095 26939 11101
rect 11238 11024 11244 11076
rect 11296 11024 11302 11076
rect 13541 11067 13599 11073
rect 12912 11036 13124 11064
rect 1762 10956 1768 11008
rect 1820 10996 1826 11008
rect 12912 10996 12940 11036
rect 1820 10968 12940 10996
rect 13096 10996 13124 11036
rect 13541 11033 13553 11067
rect 13587 11064 13599 11067
rect 15838 11064 15844 11076
rect 13587 11036 15844 11064
rect 13587 11033 13599 11036
rect 13541 11027 13599 11033
rect 15838 11024 15844 11036
rect 15896 11024 15902 11076
rect 15933 11067 15991 11073
rect 15933 11033 15945 11067
rect 15979 11064 15991 11067
rect 16574 11064 16580 11076
rect 15979 11036 16580 11064
rect 15979 11033 15991 11036
rect 15933 11027 15991 11033
rect 16574 11024 16580 11036
rect 16632 11024 16638 11076
rect 17129 11067 17187 11073
rect 17129 11033 17141 11067
rect 17175 11064 17187 11067
rect 17770 11064 17776 11076
rect 17175 11036 17776 11064
rect 17175 11033 17187 11036
rect 17129 11027 17187 11033
rect 17770 11024 17776 11036
rect 17828 11024 17834 11076
rect 18138 11024 18144 11076
rect 18196 11064 18202 11076
rect 19058 11064 19064 11076
rect 18196 11036 19064 11064
rect 18196 11024 18202 11036
rect 13998 10996 14004 11008
rect 13096 10968 14004 10996
rect 1820 10956 1826 10968
rect 13998 10956 14004 10968
rect 14056 10956 14062 11008
rect 15378 10956 15384 11008
rect 15436 10996 15442 11008
rect 16390 10996 16396 11008
rect 15436 10968 16396 10996
rect 15436 10956 15442 10968
rect 16390 10956 16396 10968
rect 16448 10956 16454 11008
rect 17862 10956 17868 11008
rect 17920 10996 17926 11008
rect 18340 11005 18368 11036
rect 19058 11024 19064 11036
rect 19116 11024 19122 11076
rect 19797 11067 19855 11073
rect 19797 11033 19809 11067
rect 19843 11064 19855 11067
rect 20806 11064 20812 11076
rect 19843 11036 20812 11064
rect 19843 11033 19855 11036
rect 19797 11027 19855 11033
rect 20806 11024 20812 11036
rect 20864 11024 20870 11076
rect 21174 11024 21180 11076
rect 21232 11024 21238 11076
rect 23661 11067 23719 11073
rect 22572 11036 22784 11064
rect 17957 10999 18015 11005
rect 17957 10996 17969 10999
rect 17920 10968 17969 10996
rect 17920 10956 17926 10968
rect 17957 10965 17969 10968
rect 18003 10965 18015 10999
rect 17957 10959 18015 10965
rect 18325 10999 18383 11005
rect 18325 10965 18337 10999
rect 18371 10965 18383 10999
rect 18325 10959 18383 10965
rect 18598 10956 18604 11008
rect 18656 10996 18662 11008
rect 19886 10996 19892 11008
rect 18656 10968 19892 10996
rect 18656 10956 18662 10968
rect 19886 10956 19892 10968
rect 19944 10996 19950 11008
rect 22572 10996 22600 11036
rect 19944 10968 22600 10996
rect 19944 10956 19950 10968
rect 22646 10956 22652 11008
rect 22704 10956 22710 11008
rect 22756 10996 22784 11036
rect 23661 11033 23673 11067
rect 23707 11064 23719 11067
rect 24210 11064 24216 11076
rect 23707 11036 24216 11064
rect 23707 11033 23719 11036
rect 23661 11027 23719 11033
rect 24210 11024 24216 11036
rect 24268 11024 24274 11076
rect 26896 11064 26924 11095
rect 28810 11064 28816 11076
rect 26896 11036 27016 11064
rect 28382 11036 28816 11064
rect 26988 11008 27016 11036
rect 28810 11024 28816 11036
rect 28868 11064 28874 11076
rect 29288 11064 29316 11240
rect 29365 11237 29377 11240
rect 29411 11268 29423 11271
rect 30006 11268 30012 11280
rect 29411 11240 30012 11268
rect 29411 11237 29423 11240
rect 29365 11231 29423 11237
rect 30006 11228 30012 11240
rect 30064 11228 30070 11280
rect 33336 11268 33364 11308
rect 33410 11296 33416 11348
rect 33468 11336 33474 11348
rect 34974 11336 34980 11348
rect 33468 11308 34980 11336
rect 33468 11296 33474 11308
rect 34974 11296 34980 11308
rect 35032 11296 35038 11348
rect 36170 11336 36176 11348
rect 35084 11308 36176 11336
rect 35084 11268 35112 11308
rect 36170 11296 36176 11308
rect 36228 11296 36234 11348
rect 38749 11339 38807 11345
rect 38749 11305 38761 11339
rect 38795 11336 38807 11339
rect 39298 11336 39304 11348
rect 38795 11308 39304 11336
rect 38795 11305 38807 11308
rect 38749 11299 38807 11305
rect 39298 11296 39304 11308
rect 39356 11296 39362 11348
rect 39482 11296 39488 11348
rect 39540 11336 39546 11348
rect 39577 11339 39635 11345
rect 39577 11336 39589 11339
rect 39540 11308 39589 11336
rect 39540 11296 39546 11308
rect 39577 11305 39589 11308
rect 39623 11305 39635 11339
rect 41598 11336 41604 11348
rect 39577 11299 39635 11305
rect 39684 11308 41604 11336
rect 38197 11271 38255 11277
rect 33336 11240 35112 11268
rect 35176 11240 35848 11268
rect 30285 11203 30343 11209
rect 30285 11169 30297 11203
rect 30331 11200 30343 11203
rect 31018 11200 31024 11212
rect 30331 11172 31024 11200
rect 30331 11169 30343 11172
rect 30285 11163 30343 11169
rect 31018 11160 31024 11172
rect 31076 11160 31082 11212
rect 31389 11203 31447 11209
rect 31389 11169 31401 11203
rect 31435 11200 31447 11203
rect 31938 11200 31944 11212
rect 31435 11172 31944 11200
rect 31435 11169 31447 11172
rect 31389 11163 31447 11169
rect 31938 11160 31944 11172
rect 31996 11200 32002 11212
rect 32122 11200 32128 11212
rect 31996 11172 32128 11200
rect 31996 11160 32002 11172
rect 32122 11160 32128 11172
rect 32180 11160 32186 11212
rect 32766 11160 32772 11212
rect 32824 11200 32830 11212
rect 32861 11203 32919 11209
rect 32861 11200 32873 11203
rect 32824 11172 32873 11200
rect 32824 11160 32830 11172
rect 32861 11169 32873 11172
rect 32907 11169 32919 11203
rect 32861 11163 32919 11169
rect 34054 11160 34060 11212
rect 34112 11160 34118 11212
rect 34146 11160 34152 11212
rect 34204 11200 34210 11212
rect 35176 11200 35204 11240
rect 34204 11172 35204 11200
rect 34204 11160 34210 11172
rect 35710 11160 35716 11212
rect 35768 11160 35774 11212
rect 35820 11200 35848 11240
rect 38197 11237 38209 11271
rect 38243 11268 38255 11271
rect 39684 11268 39712 11308
rect 41598 11296 41604 11308
rect 41656 11296 41662 11348
rect 38243 11240 39712 11268
rect 40773 11271 40831 11277
rect 38243 11237 38255 11240
rect 38197 11231 38255 11237
rect 40773 11237 40785 11271
rect 40819 11268 40831 11271
rect 40819 11240 45554 11268
rect 40819 11237 40831 11240
rect 40773 11231 40831 11237
rect 35820 11172 37780 11200
rect 29546 11092 29552 11144
rect 29604 11132 29610 11144
rect 31113 11135 31171 11141
rect 31113 11132 31125 11135
rect 29604 11104 31125 11132
rect 29604 11092 29610 11104
rect 31113 11101 31125 11104
rect 31159 11101 31171 11135
rect 31113 11095 31171 11101
rect 33321 11135 33379 11141
rect 33321 11101 33333 11135
rect 33367 11132 33379 11135
rect 33778 11132 33784 11144
rect 33367 11104 33784 11132
rect 33367 11101 33379 11104
rect 33321 11095 33379 11101
rect 33778 11092 33784 11104
rect 33836 11132 33842 11144
rect 37752 11141 37780 11172
rect 34701 11135 34759 11141
rect 34701 11132 34713 11135
rect 33836 11104 34713 11132
rect 33836 11092 33842 11104
rect 34701 11101 34713 11104
rect 34747 11101 34759 11135
rect 34701 11095 34759 11101
rect 37737 11135 37795 11141
rect 37737 11101 37749 11135
rect 37783 11101 37795 11135
rect 37737 11095 37795 11101
rect 38381 11135 38439 11141
rect 38381 11101 38393 11135
rect 38427 11101 38439 11135
rect 38381 11095 38439 11101
rect 28868 11036 29316 11064
rect 28868 11024 28874 11036
rect 29362 11024 29368 11076
rect 29420 11064 29426 11076
rect 30190 11064 30196 11076
rect 29420 11036 30196 11064
rect 29420 11024 29426 11036
rect 30190 11024 30196 11036
rect 30248 11024 30254 11076
rect 30742 11064 30748 11076
rect 30300 11036 30748 11064
rect 26142 10996 26148 11008
rect 22756 10968 26148 10996
rect 26142 10956 26148 10968
rect 26200 10956 26206 11008
rect 26970 10956 26976 11008
rect 27028 10956 27034 11008
rect 27798 10956 27804 11008
rect 27856 10996 27862 11008
rect 29730 10996 29736 11008
rect 27856 10968 29736 10996
rect 27856 10956 27862 10968
rect 29730 10956 29736 10968
rect 29788 10956 29794 11008
rect 30006 10956 30012 11008
rect 30064 10996 30070 11008
rect 30101 10999 30159 11005
rect 30101 10996 30113 10999
rect 30064 10968 30113 10996
rect 30064 10956 30070 10968
rect 30101 10965 30113 10968
rect 30147 10996 30159 10999
rect 30300 10996 30328 11036
rect 30742 11024 30748 11036
rect 30800 11024 30806 11076
rect 33226 11064 33232 11076
rect 32614 11036 33232 11064
rect 33226 11024 33232 11036
rect 33284 11024 33290 11076
rect 35989 11067 36047 11073
rect 35989 11033 36001 11067
rect 36035 11064 36047 11067
rect 36078 11064 36084 11076
rect 36035 11036 36084 11064
rect 36035 11033 36047 11036
rect 35989 11027 36047 11033
rect 36078 11024 36084 11036
rect 36136 11024 36142 11076
rect 36722 11024 36728 11076
rect 36780 11024 36786 11076
rect 37366 11024 37372 11076
rect 37424 11064 37430 11076
rect 38396 11064 38424 11095
rect 39482 11092 39488 11144
rect 39540 11132 39546 11144
rect 40129 11135 40187 11141
rect 40129 11132 40141 11135
rect 39540 11104 40141 11132
rect 39540 11092 39546 11104
rect 40129 11101 40141 11104
rect 40175 11101 40187 11135
rect 40129 11095 40187 11101
rect 40218 11092 40224 11144
rect 40276 11132 40282 11144
rect 40957 11135 41015 11141
rect 40957 11132 40969 11135
rect 40276 11104 40969 11132
rect 40276 11092 40282 11104
rect 40957 11101 40969 11104
rect 41003 11101 41015 11135
rect 45526 11132 45554 11240
rect 49142 11160 49148 11212
rect 49200 11160 49206 11212
rect 45649 11135 45707 11141
rect 45649 11132 45661 11135
rect 45526 11104 45661 11132
rect 40957 11095 41015 11101
rect 45649 11101 45661 11104
rect 45695 11101 45707 11135
rect 45649 11095 45707 11101
rect 47026 11092 47032 11144
rect 47084 11132 47090 11144
rect 47949 11135 48007 11141
rect 47949 11132 47961 11135
rect 47084 11104 47961 11132
rect 47084 11092 47090 11104
rect 47949 11101 47961 11104
rect 47995 11101 48007 11135
rect 47949 11095 48007 11101
rect 37424 11036 38424 11064
rect 40313 11067 40371 11073
rect 37424 11024 37430 11036
rect 40313 11033 40325 11067
rect 40359 11064 40371 11067
rect 45738 11064 45744 11076
rect 40359 11036 45744 11064
rect 40359 11033 40371 11036
rect 40313 11027 40371 11033
rect 45738 11024 45744 11036
rect 45796 11024 45802 11076
rect 45833 11067 45891 11073
rect 45833 11033 45845 11067
rect 45879 11064 45891 11067
rect 46934 11064 46940 11076
rect 45879 11036 46940 11064
rect 45879 11033 45891 11036
rect 45833 11027 45891 11033
rect 46934 11024 46940 11036
rect 46992 11024 46998 11076
rect 30147 10968 30328 10996
rect 30147 10965 30159 10968
rect 30101 10959 30159 10965
rect 30374 10956 30380 11008
rect 30432 10996 30438 11008
rect 32306 10996 32312 11008
rect 30432 10968 32312 10996
rect 30432 10956 30438 10968
rect 32306 10956 32312 10968
rect 32364 10956 32370 11008
rect 32950 10956 32956 11008
rect 33008 10996 33014 11008
rect 37458 10996 37464 11008
rect 33008 10968 37464 10996
rect 33008 10956 33014 10968
rect 37458 10956 37464 10968
rect 37516 10956 37522 11008
rect 1104 10906 49864 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 27950 10906
rect 28002 10854 28014 10906
rect 28066 10854 28078 10906
rect 28130 10854 28142 10906
rect 28194 10854 28206 10906
rect 28258 10854 37950 10906
rect 38002 10854 38014 10906
rect 38066 10854 38078 10906
rect 38130 10854 38142 10906
rect 38194 10854 38206 10906
rect 38258 10854 47950 10906
rect 48002 10854 48014 10906
rect 48066 10854 48078 10906
rect 48130 10854 48142 10906
rect 48194 10854 48206 10906
rect 48258 10854 49864 10906
rect 1104 10832 49864 10854
rect 1762 10752 1768 10804
rect 1820 10752 1826 10804
rect 1854 10752 1860 10804
rect 1912 10792 1918 10804
rect 1912 10764 6914 10792
rect 1912 10752 1918 10764
rect 1210 10684 1216 10736
rect 1268 10724 1274 10736
rect 6886 10724 6914 10764
rect 12342 10752 12348 10804
rect 12400 10792 12406 10804
rect 12621 10795 12679 10801
rect 12621 10792 12633 10795
rect 12400 10764 12633 10792
rect 12400 10752 12406 10764
rect 12621 10761 12633 10764
rect 12667 10761 12679 10795
rect 12621 10755 12679 10761
rect 12802 10752 12808 10804
rect 12860 10792 12866 10804
rect 13173 10795 13231 10801
rect 13173 10792 13185 10795
rect 12860 10764 13185 10792
rect 12860 10752 12866 10764
rect 13173 10761 13185 10764
rect 13219 10761 13231 10795
rect 13173 10755 13231 10761
rect 14182 10752 14188 10804
rect 14240 10792 14246 10804
rect 14369 10795 14427 10801
rect 14369 10792 14381 10795
rect 14240 10764 14381 10792
rect 14240 10752 14246 10764
rect 14369 10761 14381 10764
rect 14415 10761 14427 10795
rect 14369 10755 14427 10761
rect 15933 10795 15991 10801
rect 15933 10761 15945 10795
rect 15979 10792 15991 10795
rect 17129 10795 17187 10801
rect 17129 10792 17141 10795
rect 15979 10764 17141 10792
rect 15979 10761 15991 10764
rect 15933 10755 15991 10761
rect 17129 10761 17141 10764
rect 17175 10761 17187 10795
rect 17129 10755 17187 10761
rect 18046 10752 18052 10804
rect 18104 10792 18110 10804
rect 18785 10795 18843 10801
rect 18785 10792 18797 10795
rect 18104 10764 18797 10792
rect 18104 10752 18110 10764
rect 18785 10761 18797 10764
rect 18831 10792 18843 10795
rect 19521 10795 19579 10801
rect 18831 10764 19380 10792
rect 18831 10761 18843 10764
rect 18785 10755 18843 10761
rect 14550 10724 14556 10736
rect 1268 10696 2360 10724
rect 6886 10696 14556 10724
rect 1268 10684 1274 10696
rect 1302 10616 1308 10668
rect 1360 10656 1366 10668
rect 2332 10665 2360 10696
rect 14550 10684 14556 10696
rect 14608 10684 14614 10736
rect 14737 10727 14795 10733
rect 14737 10693 14749 10727
rect 14783 10724 14795 10727
rect 15746 10724 15752 10736
rect 14783 10696 15752 10724
rect 14783 10693 14795 10696
rect 14737 10687 14795 10693
rect 1581 10659 1639 10665
rect 1581 10656 1593 10659
rect 1360 10628 1593 10656
rect 1360 10616 1366 10628
rect 1581 10625 1593 10628
rect 1627 10625 1639 10659
rect 1581 10619 1639 10625
rect 2317 10659 2375 10665
rect 2317 10625 2329 10659
rect 2363 10656 2375 10659
rect 2869 10659 2927 10665
rect 2869 10656 2881 10659
rect 2363 10628 2881 10656
rect 2363 10625 2375 10628
rect 2317 10619 2375 10625
rect 2869 10625 2881 10628
rect 2915 10625 2927 10659
rect 2869 10619 2927 10625
rect 1596 10588 1624 10619
rect 13538 10616 13544 10668
rect 13596 10616 13602 10668
rect 13630 10616 13636 10668
rect 13688 10616 13694 10668
rect 13906 10616 13912 10668
rect 13964 10656 13970 10668
rect 14752 10656 14780 10687
rect 15746 10684 15752 10696
rect 15804 10684 15810 10736
rect 15838 10684 15844 10736
rect 15896 10724 15902 10736
rect 17497 10727 17555 10733
rect 17497 10724 17509 10727
rect 15896 10696 17509 10724
rect 15896 10684 15902 10696
rect 17497 10693 17509 10696
rect 17543 10693 17555 10727
rect 17497 10687 17555 10693
rect 17586 10684 17592 10736
rect 17644 10684 17650 10736
rect 18156 10696 18828 10724
rect 13964 10628 14780 10656
rect 14829 10659 14887 10665
rect 13964 10616 13970 10628
rect 14829 10625 14841 10659
rect 14875 10656 14887 10659
rect 16482 10656 16488 10668
rect 14875 10628 16488 10656
rect 14875 10625 14887 10628
rect 14829 10619 14887 10625
rect 16482 10616 16488 10628
rect 16540 10616 16546 10668
rect 16853 10659 16911 10665
rect 16853 10625 16865 10659
rect 16899 10656 16911 10659
rect 17604 10656 17632 10684
rect 18156 10656 18184 10696
rect 16899 10628 18184 10656
rect 16899 10625 16911 10628
rect 16853 10619 16911 10625
rect 18230 10616 18236 10668
rect 18288 10656 18294 10668
rect 18288 10628 18644 10656
rect 18288 10616 18294 10628
rect 3053 10591 3111 10597
rect 3053 10588 3065 10591
rect 1596 10560 3065 10588
rect 3053 10557 3065 10560
rect 3099 10557 3111 10591
rect 3053 10551 3111 10557
rect 12897 10591 12955 10597
rect 12897 10557 12909 10591
rect 12943 10588 12955 10591
rect 13648 10588 13676 10616
rect 12943 10560 13676 10588
rect 13817 10591 13875 10597
rect 12943 10557 12955 10560
rect 12897 10551 12955 10557
rect 13817 10557 13829 10591
rect 13863 10588 13875 10591
rect 14366 10588 14372 10600
rect 13863 10560 14372 10588
rect 13863 10557 13875 10560
rect 13817 10551 13875 10557
rect 14366 10548 14372 10560
rect 14424 10548 14430 10600
rect 14918 10548 14924 10600
rect 14976 10548 14982 10600
rect 16022 10548 16028 10600
rect 16080 10548 16086 10600
rect 16114 10548 16120 10600
rect 16172 10548 16178 10600
rect 16574 10548 16580 10600
rect 16632 10588 16638 10600
rect 17589 10591 17647 10597
rect 17589 10588 17601 10591
rect 16632 10560 17601 10588
rect 16632 10548 16638 10560
rect 17589 10557 17601 10560
rect 17635 10557 17647 10591
rect 17589 10551 17647 10557
rect 17681 10591 17739 10597
rect 17681 10557 17693 10591
rect 17727 10557 17739 10591
rect 18616 10588 18644 10628
rect 18690 10616 18696 10668
rect 18748 10616 18754 10668
rect 18800 10656 18828 10696
rect 19352 10656 19380 10764
rect 19521 10761 19533 10795
rect 19567 10792 19579 10795
rect 19702 10792 19708 10804
rect 19567 10764 19708 10792
rect 19567 10761 19579 10764
rect 19521 10755 19579 10761
rect 19702 10752 19708 10764
rect 19760 10752 19766 10804
rect 19886 10752 19892 10804
rect 19944 10752 19950 10804
rect 21085 10795 21143 10801
rect 21085 10761 21097 10795
rect 21131 10792 21143 10795
rect 22646 10792 22652 10804
rect 21131 10764 22652 10792
rect 21131 10761 21143 10764
rect 21085 10755 21143 10761
rect 22646 10752 22652 10764
rect 22704 10752 22710 10804
rect 23658 10752 23664 10804
rect 23716 10792 23722 10804
rect 24213 10795 24271 10801
rect 24213 10792 24225 10795
rect 23716 10764 24225 10792
rect 23716 10752 23722 10764
rect 24213 10761 24225 10764
rect 24259 10761 24271 10795
rect 24213 10755 24271 10761
rect 26142 10752 26148 10804
rect 26200 10792 26206 10804
rect 27617 10795 27675 10801
rect 27617 10792 27629 10795
rect 26200 10764 27629 10792
rect 26200 10752 26206 10764
rect 27617 10761 27629 10764
rect 27663 10761 27675 10795
rect 27617 10755 27675 10761
rect 28537 10795 28595 10801
rect 28537 10761 28549 10795
rect 28583 10792 28595 10795
rect 28902 10792 28908 10804
rect 28583 10764 28908 10792
rect 28583 10761 28595 10764
rect 28537 10755 28595 10761
rect 21177 10727 21235 10733
rect 21177 10693 21189 10727
rect 21223 10724 21235 10727
rect 22278 10724 22284 10736
rect 21223 10696 22284 10724
rect 21223 10693 21235 10696
rect 21177 10687 21235 10693
rect 22278 10684 22284 10696
rect 22336 10684 22342 10736
rect 27632 10724 27660 10755
rect 28828 10733 28856 10764
rect 28902 10752 28908 10764
rect 28960 10752 28966 10804
rect 29730 10752 29736 10804
rect 29788 10792 29794 10804
rect 29788 10764 30880 10792
rect 29788 10752 29794 10764
rect 28813 10727 28871 10733
rect 23584 10696 26372 10724
rect 27632 10696 28028 10724
rect 21450 10656 21456 10668
rect 18800 10628 19104 10656
rect 19352 10628 21456 10656
rect 18877 10591 18935 10597
rect 18877 10588 18889 10591
rect 17681 10551 17739 10557
rect 17788 10560 18552 10588
rect 18616 10560 18889 10588
rect 2501 10523 2559 10529
rect 2501 10489 2513 10523
rect 2547 10520 2559 10523
rect 2547 10492 6914 10520
rect 2547 10489 2559 10492
rect 2501 10483 2559 10489
rect 6886 10452 6914 10492
rect 15010 10480 15016 10532
rect 15068 10520 15074 10532
rect 17696 10520 17724 10551
rect 15068 10492 17724 10520
rect 15068 10480 15074 10492
rect 14274 10452 14280 10464
rect 6886 10424 14280 10452
rect 14274 10412 14280 10424
rect 14332 10412 14338 10464
rect 15562 10412 15568 10464
rect 15620 10412 15626 10464
rect 16390 10412 16396 10464
rect 16448 10452 16454 10464
rect 17788 10452 17816 10560
rect 16448 10424 17816 10452
rect 18325 10455 18383 10461
rect 16448 10412 16454 10424
rect 18325 10421 18337 10455
rect 18371 10452 18383 10455
rect 18414 10452 18420 10464
rect 18371 10424 18420 10452
rect 18371 10421 18383 10424
rect 18325 10415 18383 10421
rect 18414 10412 18420 10424
rect 18472 10412 18478 10464
rect 18524 10452 18552 10560
rect 18877 10557 18889 10560
rect 18923 10557 18935 10591
rect 19076 10588 19104 10628
rect 21450 10616 21456 10628
rect 21508 10616 21514 10668
rect 23382 10616 23388 10668
rect 23440 10616 23446 10668
rect 19981 10591 20039 10597
rect 19981 10588 19993 10591
rect 19076 10560 19993 10588
rect 18877 10551 18935 10557
rect 19981 10557 19993 10560
rect 20027 10557 20039 10591
rect 19981 10551 20039 10557
rect 20165 10591 20223 10597
rect 20165 10557 20177 10591
rect 20211 10588 20223 10591
rect 20806 10588 20812 10600
rect 20211 10560 20812 10588
rect 20211 10557 20223 10560
rect 20165 10551 20223 10557
rect 20806 10548 20812 10560
rect 20864 10548 20870 10600
rect 21361 10591 21419 10597
rect 21361 10557 21373 10591
rect 21407 10557 21419 10591
rect 21361 10551 21419 10557
rect 20717 10455 20775 10461
rect 20717 10452 20729 10455
rect 18524 10424 20729 10452
rect 20717 10421 20729 10424
rect 20763 10421 20775 10455
rect 21376 10452 21404 10551
rect 21542 10548 21548 10600
rect 21600 10588 21606 10600
rect 22002 10588 22008 10600
rect 21600 10560 22008 10588
rect 21600 10548 21606 10560
rect 22002 10548 22008 10560
rect 22060 10548 22066 10600
rect 22281 10591 22339 10597
rect 22281 10588 22293 10591
rect 22112 10560 22293 10588
rect 21818 10480 21824 10532
rect 21876 10520 21882 10532
rect 22112 10520 22140 10560
rect 22281 10557 22293 10560
rect 22327 10557 22339 10591
rect 22281 10551 22339 10557
rect 22830 10548 22836 10600
rect 22888 10588 22894 10600
rect 23584 10588 23612 10696
rect 26344 10665 26372 10696
rect 24581 10659 24639 10665
rect 24581 10625 24593 10659
rect 24627 10656 24639 10659
rect 25409 10659 25467 10665
rect 25409 10656 25421 10659
rect 24627 10628 25421 10656
rect 24627 10625 24639 10628
rect 24581 10619 24639 10625
rect 25409 10625 25421 10628
rect 25455 10625 25467 10659
rect 25409 10619 25467 10625
rect 26329 10659 26387 10665
rect 26329 10625 26341 10659
rect 26375 10656 26387 10659
rect 27430 10656 27436 10668
rect 26375 10628 27436 10656
rect 26375 10625 26387 10628
rect 26329 10619 26387 10625
rect 27430 10616 27436 10628
rect 27488 10656 27494 10668
rect 27525 10659 27583 10665
rect 27525 10656 27537 10659
rect 27488 10628 27537 10656
rect 27488 10616 27494 10628
rect 27525 10625 27537 10628
rect 27571 10625 27583 10659
rect 27525 10619 27583 10625
rect 22888 10560 23612 10588
rect 22888 10548 22894 10560
rect 23934 10548 23940 10600
rect 23992 10588 23998 10600
rect 24673 10591 24731 10597
rect 24673 10588 24685 10591
rect 23992 10560 24685 10588
rect 23992 10548 23998 10560
rect 24673 10557 24685 10560
rect 24719 10557 24731 10591
rect 24673 10551 24731 10557
rect 21876 10492 22140 10520
rect 24688 10520 24716 10551
rect 24854 10548 24860 10600
rect 24912 10588 24918 10600
rect 26602 10588 26608 10600
rect 24912 10560 26608 10588
rect 24912 10548 24918 10560
rect 26602 10548 26608 10560
rect 26660 10548 26666 10600
rect 27798 10548 27804 10600
rect 27856 10548 27862 10600
rect 28000 10588 28028 10696
rect 28813 10693 28825 10727
rect 28859 10724 28871 10727
rect 28859 10696 28893 10724
rect 28859 10693 28871 10696
rect 28813 10687 28871 10693
rect 29546 10684 29552 10736
rect 29604 10684 29610 10736
rect 30282 10684 30288 10736
rect 30340 10724 30346 10736
rect 30852 10724 30880 10764
rect 31110 10752 31116 10804
rect 31168 10792 31174 10804
rect 31389 10795 31447 10801
rect 31389 10792 31401 10795
rect 31168 10764 31401 10792
rect 31168 10752 31174 10764
rect 31389 10761 31401 10764
rect 31435 10761 31447 10795
rect 31389 10755 31447 10761
rect 32309 10795 32367 10801
rect 32309 10761 32321 10795
rect 32355 10792 32367 10795
rect 32950 10792 32956 10804
rect 32355 10764 32956 10792
rect 32355 10761 32367 10764
rect 32309 10755 32367 10761
rect 32950 10752 32956 10764
rect 33008 10752 33014 10804
rect 33318 10752 33324 10804
rect 33376 10752 33382 10804
rect 35066 10792 35072 10804
rect 33796 10764 35072 10792
rect 31754 10724 31760 10736
rect 30340 10696 30788 10724
rect 30852 10696 31760 10724
rect 30340 10684 30346 10696
rect 29730 10616 29736 10668
rect 29788 10656 29794 10668
rect 30561 10659 30619 10665
rect 30561 10656 30573 10659
rect 29788 10628 30573 10656
rect 29788 10616 29794 10628
rect 30561 10625 30573 10628
rect 30607 10625 30619 10659
rect 30561 10619 30619 10625
rect 29086 10588 29092 10600
rect 28000 10560 29092 10588
rect 29086 10548 29092 10560
rect 29144 10588 29150 10600
rect 30374 10588 30380 10600
rect 29144 10560 30380 10588
rect 29144 10548 29150 10560
rect 30374 10548 30380 10560
rect 30432 10548 30438 10600
rect 30466 10548 30472 10600
rect 30524 10588 30530 10600
rect 30760 10597 30788 10696
rect 31754 10684 31760 10696
rect 31812 10724 31818 10736
rect 32214 10724 32220 10736
rect 31812 10696 32220 10724
rect 31812 10684 31818 10696
rect 32214 10684 32220 10696
rect 32272 10684 32278 10736
rect 32398 10684 32404 10736
rect 32456 10724 32462 10736
rect 32456 10696 32904 10724
rect 32456 10684 32462 10696
rect 32674 10616 32680 10668
rect 32732 10616 32738 10668
rect 32876 10597 32904 10696
rect 33796 10665 33824 10764
rect 35066 10752 35072 10764
rect 35124 10792 35130 10804
rect 35710 10792 35716 10804
rect 35124 10764 35716 10792
rect 35124 10752 35130 10764
rect 35710 10752 35716 10764
rect 35768 10752 35774 10804
rect 36081 10795 36139 10801
rect 36081 10761 36093 10795
rect 36127 10792 36139 10795
rect 36906 10792 36912 10804
rect 36127 10764 36912 10792
rect 36127 10761 36139 10764
rect 36081 10755 36139 10761
rect 36906 10752 36912 10764
rect 36964 10752 36970 10804
rect 35342 10684 35348 10736
rect 35400 10724 35406 10736
rect 35400 10696 36676 10724
rect 35400 10684 35406 10696
rect 33781 10659 33839 10665
rect 33781 10625 33793 10659
rect 33827 10625 33839 10659
rect 35526 10656 35532 10668
rect 35190 10628 35532 10656
rect 33781 10619 33839 10625
rect 35526 10616 35532 10628
rect 35584 10616 35590 10668
rect 35710 10616 35716 10668
rect 35768 10656 35774 10668
rect 36449 10659 36507 10665
rect 36449 10656 36461 10659
rect 35768 10628 36461 10656
rect 35768 10616 35774 10628
rect 36449 10625 36461 10628
rect 36495 10625 36507 10659
rect 36449 10619 36507 10625
rect 30653 10591 30711 10597
rect 30653 10588 30665 10591
rect 30524 10560 30665 10588
rect 30524 10548 30530 10560
rect 30653 10557 30665 10560
rect 30699 10557 30711 10591
rect 30653 10551 30711 10557
rect 30745 10591 30803 10597
rect 30745 10557 30757 10591
rect 30791 10557 30803 10591
rect 32769 10591 32827 10597
rect 32769 10588 32781 10591
rect 30745 10551 30803 10557
rect 31726 10560 32781 10588
rect 27157 10523 27215 10529
rect 24688 10492 27108 10520
rect 21876 10480 21882 10492
rect 22094 10452 22100 10464
rect 21376 10424 22100 10452
rect 20717 10415 20775 10421
rect 22094 10412 22100 10424
rect 22152 10412 22158 10464
rect 23658 10412 23664 10464
rect 23716 10452 23722 10464
rect 23753 10455 23811 10461
rect 23753 10452 23765 10455
rect 23716 10424 23765 10452
rect 23716 10412 23722 10424
rect 23753 10421 23765 10424
rect 23799 10421 23811 10455
rect 23753 10415 23811 10421
rect 25958 10412 25964 10464
rect 26016 10412 26022 10464
rect 26142 10412 26148 10464
rect 26200 10412 26206 10464
rect 26510 10412 26516 10464
rect 26568 10412 26574 10464
rect 26786 10412 26792 10464
rect 26844 10412 26850 10464
rect 27080 10452 27108 10492
rect 27157 10489 27169 10523
rect 27203 10520 27215 10523
rect 31726 10520 31754 10560
rect 32769 10557 32781 10560
rect 32815 10557 32827 10591
rect 32769 10551 32827 10557
rect 32861 10591 32919 10597
rect 32861 10557 32873 10591
rect 32907 10557 32919 10591
rect 32861 10551 32919 10557
rect 34057 10591 34115 10597
rect 34057 10557 34069 10591
rect 34103 10588 34115 10591
rect 34103 10560 35848 10588
rect 34103 10557 34115 10560
rect 34057 10551 34115 10557
rect 27203 10492 31754 10520
rect 27203 10489 27215 10492
rect 27157 10483 27215 10489
rect 32306 10480 32312 10532
rect 32364 10520 32370 10532
rect 32364 10492 33916 10520
rect 32364 10480 32370 10492
rect 30006 10452 30012 10464
rect 27080 10424 30012 10452
rect 30006 10412 30012 10424
rect 30064 10412 30070 10464
rect 30193 10455 30251 10461
rect 30193 10421 30205 10455
rect 30239 10452 30251 10455
rect 31294 10452 31300 10464
rect 30239 10424 31300 10452
rect 30239 10421 30251 10424
rect 30193 10415 30251 10421
rect 31294 10412 31300 10424
rect 31352 10412 31358 10464
rect 31938 10412 31944 10464
rect 31996 10412 32002 10464
rect 32214 10412 32220 10464
rect 32272 10452 32278 10464
rect 32858 10452 32864 10464
rect 32272 10424 32864 10452
rect 32272 10412 32278 10424
rect 32858 10412 32864 10424
rect 32916 10412 32922 10464
rect 33888 10452 33916 10492
rect 35158 10480 35164 10532
rect 35216 10520 35222 10532
rect 35529 10523 35587 10529
rect 35529 10520 35541 10523
rect 35216 10492 35541 10520
rect 35216 10480 35222 10492
rect 35529 10489 35541 10492
rect 35575 10489 35587 10523
rect 35820 10520 35848 10560
rect 35894 10548 35900 10600
rect 35952 10588 35958 10600
rect 36648 10597 36676 10696
rect 36722 10684 36728 10736
rect 36780 10724 36786 10736
rect 37277 10727 37335 10733
rect 37277 10724 37289 10727
rect 36780 10696 37289 10724
rect 36780 10684 36786 10696
rect 37277 10693 37289 10696
rect 37323 10693 37335 10727
rect 37277 10687 37335 10693
rect 49145 10727 49203 10733
rect 49145 10693 49157 10727
rect 49191 10724 49203 10727
rect 49234 10724 49240 10736
rect 49191 10696 49240 10724
rect 49191 10693 49203 10696
rect 49145 10687 49203 10693
rect 49234 10684 49240 10696
rect 49292 10684 49298 10736
rect 39758 10616 39764 10668
rect 39816 10656 39822 10668
rect 40221 10659 40279 10665
rect 40221 10656 40233 10659
rect 39816 10628 40233 10656
rect 39816 10616 39822 10628
rect 40221 10625 40233 10628
rect 40267 10625 40279 10659
rect 40221 10619 40279 10625
rect 46934 10616 46940 10668
rect 46992 10656 46998 10668
rect 47949 10659 48007 10665
rect 47949 10656 47961 10659
rect 46992 10628 47961 10656
rect 46992 10616 46998 10628
rect 47949 10625 47961 10628
rect 47995 10625 48007 10659
rect 47949 10619 48007 10625
rect 36541 10591 36599 10597
rect 36541 10588 36553 10591
rect 35952 10560 36553 10588
rect 35952 10548 35958 10560
rect 36541 10557 36553 10560
rect 36587 10557 36599 10591
rect 36541 10551 36599 10557
rect 36633 10591 36691 10597
rect 36633 10557 36645 10591
rect 36679 10557 36691 10591
rect 36633 10551 36691 10557
rect 39945 10523 40003 10529
rect 35820 10492 36676 10520
rect 35529 10483 35587 10489
rect 36648 10464 36676 10492
rect 39945 10489 39957 10523
rect 39991 10520 40003 10523
rect 46934 10520 46940 10532
rect 39991 10492 46940 10520
rect 39991 10489 40003 10492
rect 39945 10483 40003 10489
rect 46934 10480 46940 10492
rect 46992 10480 46998 10532
rect 35342 10452 35348 10464
rect 33888 10424 35348 10452
rect 35342 10412 35348 10424
rect 35400 10412 35406 10464
rect 36630 10412 36636 10464
rect 36688 10412 36694 10464
rect 1104 10362 49864 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 32950 10362
rect 33002 10310 33014 10362
rect 33066 10310 33078 10362
rect 33130 10310 33142 10362
rect 33194 10310 33206 10362
rect 33258 10310 42950 10362
rect 43002 10310 43014 10362
rect 43066 10310 43078 10362
rect 43130 10310 43142 10362
rect 43194 10310 43206 10362
rect 43258 10310 49864 10362
rect 1104 10288 49864 10310
rect 12713 10251 12771 10257
rect 12713 10217 12725 10251
rect 12759 10248 12771 10251
rect 16022 10248 16028 10260
rect 12759 10220 16028 10248
rect 12759 10217 12771 10220
rect 12713 10211 12771 10217
rect 16022 10208 16028 10220
rect 16080 10208 16086 10260
rect 16206 10208 16212 10260
rect 16264 10248 16270 10260
rect 16393 10251 16451 10257
rect 16393 10248 16405 10251
rect 16264 10220 16405 10248
rect 16264 10208 16270 10220
rect 16393 10217 16405 10220
rect 16439 10248 16451 10251
rect 18046 10248 18052 10260
rect 16439 10220 18052 10248
rect 16439 10217 16451 10220
rect 16393 10211 16451 10217
rect 18046 10208 18052 10220
rect 18104 10208 18110 10260
rect 18141 10251 18199 10257
rect 18141 10217 18153 10251
rect 18187 10248 18199 10251
rect 18322 10248 18328 10260
rect 18187 10220 18328 10248
rect 18187 10217 18199 10220
rect 18141 10211 18199 10217
rect 18322 10208 18328 10220
rect 18380 10208 18386 10260
rect 18432 10220 21588 10248
rect 13906 10140 13912 10192
rect 13964 10140 13970 10192
rect 17954 10180 17960 10192
rect 15580 10152 17960 10180
rect 1854 10072 1860 10124
rect 1912 10072 1918 10124
rect 13265 10115 13323 10121
rect 13265 10112 13277 10115
rect 13096 10084 13277 10112
rect 1302 10004 1308 10056
rect 1360 10044 1366 10056
rect 1581 10047 1639 10053
rect 1581 10044 1593 10047
rect 1360 10016 1593 10044
rect 1360 10004 1366 10016
rect 1581 10013 1593 10016
rect 1627 10013 1639 10047
rect 1581 10007 1639 10013
rect 13096 9976 13124 10084
rect 13265 10081 13277 10084
rect 13311 10081 13323 10115
rect 15580 10112 15608 10152
rect 17954 10140 17960 10152
rect 18012 10140 18018 10192
rect 13265 10075 13323 10081
rect 13740 10084 15608 10112
rect 16577 10115 16635 10121
rect 13173 10047 13231 10053
rect 13173 10013 13185 10047
rect 13219 10044 13231 10047
rect 13740 10044 13768 10084
rect 16577 10081 16589 10115
rect 16623 10112 16635 10115
rect 16850 10112 16856 10124
rect 16623 10084 16856 10112
rect 16623 10081 16635 10084
rect 16577 10075 16635 10081
rect 16850 10072 16856 10084
rect 16908 10072 16914 10124
rect 17402 10072 17408 10124
rect 17460 10072 17466 10124
rect 17494 10072 17500 10124
rect 17552 10112 17558 10124
rect 18230 10112 18236 10124
rect 17552 10084 18236 10112
rect 17552 10072 17558 10084
rect 18230 10072 18236 10084
rect 18288 10072 18294 10124
rect 13219 10016 13768 10044
rect 13219 10013 13231 10016
rect 13173 10007 13231 10013
rect 13814 10004 13820 10056
rect 13872 10044 13878 10056
rect 14277 10047 14335 10053
rect 14277 10044 14289 10047
rect 13872 10016 14289 10044
rect 13872 10004 13878 10016
rect 14277 10013 14289 10016
rect 14323 10013 14335 10047
rect 14277 10007 14335 10013
rect 16666 10004 16672 10056
rect 16724 10044 16730 10056
rect 18432 10044 18460 10220
rect 21560 10180 21588 10220
rect 21634 10208 21640 10260
rect 21692 10248 21698 10260
rect 22830 10248 22836 10260
rect 21692 10220 22836 10248
rect 21692 10208 21698 10220
rect 22830 10208 22836 10220
rect 22888 10208 22894 10260
rect 23750 10208 23756 10260
rect 23808 10248 23814 10260
rect 26329 10251 26387 10257
rect 26329 10248 26341 10251
rect 23808 10220 26341 10248
rect 23808 10208 23814 10220
rect 26329 10217 26341 10220
rect 26375 10217 26387 10251
rect 26329 10211 26387 10217
rect 32122 10208 32128 10260
rect 32180 10208 32186 10260
rect 32585 10251 32643 10257
rect 32585 10217 32597 10251
rect 32631 10248 32643 10251
rect 34422 10248 34428 10260
rect 32631 10220 34428 10248
rect 32631 10217 32643 10220
rect 32585 10211 32643 10217
rect 34422 10208 34428 10220
rect 34480 10208 34486 10260
rect 35158 10248 35164 10260
rect 34532 10220 35164 10248
rect 21560 10152 21864 10180
rect 18506 10072 18512 10124
rect 18564 10112 18570 10124
rect 18601 10115 18659 10121
rect 18601 10112 18613 10115
rect 18564 10084 18613 10112
rect 18564 10072 18570 10084
rect 18601 10081 18613 10084
rect 18647 10081 18659 10115
rect 18601 10075 18659 10081
rect 18785 10115 18843 10121
rect 18785 10081 18797 10115
rect 18831 10081 18843 10115
rect 18785 10075 18843 10081
rect 19521 10115 19579 10121
rect 19521 10081 19533 10115
rect 19567 10112 19579 10115
rect 19610 10112 19616 10124
rect 19567 10084 19616 10112
rect 19567 10081 19579 10084
rect 19521 10075 19579 10081
rect 16724 10016 18460 10044
rect 18800 10044 18828 10075
rect 19610 10072 19616 10084
rect 19668 10072 19674 10124
rect 19702 10072 19708 10124
rect 19760 10112 19766 10124
rect 20257 10115 20315 10121
rect 20257 10112 20269 10115
rect 19760 10084 20269 10112
rect 19760 10072 19766 10084
rect 20257 10081 20269 10084
rect 20303 10112 20315 10115
rect 21542 10112 21548 10124
rect 20303 10084 21548 10112
rect 20303 10081 20315 10084
rect 20257 10075 20315 10081
rect 21542 10072 21548 10084
rect 21600 10072 21606 10124
rect 19794 10044 19800 10056
rect 18800 10016 19800 10044
rect 16724 10004 16730 10016
rect 19794 10004 19800 10016
rect 19852 10004 19858 10056
rect 21836 10044 21864 10152
rect 23382 10140 23388 10192
rect 23440 10180 23446 10192
rect 23842 10180 23848 10192
rect 23440 10152 23848 10180
rect 23440 10140 23446 10152
rect 23842 10140 23848 10152
rect 23900 10140 23906 10192
rect 26510 10140 26516 10192
rect 26568 10180 26574 10192
rect 26697 10183 26755 10189
rect 26697 10180 26709 10183
rect 26568 10152 26709 10180
rect 26568 10140 26574 10152
rect 26697 10149 26709 10152
rect 26743 10180 26755 10183
rect 28721 10183 28779 10189
rect 26743 10152 27108 10180
rect 26743 10149 26755 10152
rect 26697 10143 26755 10149
rect 22002 10072 22008 10124
rect 22060 10112 22066 10124
rect 23201 10115 23259 10121
rect 23201 10112 23213 10115
rect 22060 10084 23213 10112
rect 22060 10072 22066 10084
rect 23201 10081 23213 10084
rect 23247 10081 23259 10115
rect 23201 10075 23259 10081
rect 23753 10115 23811 10121
rect 23753 10081 23765 10115
rect 23799 10112 23811 10115
rect 24118 10112 24124 10124
rect 23799 10084 24124 10112
rect 23799 10081 23811 10084
rect 23753 10075 23811 10081
rect 24118 10072 24124 10084
rect 24176 10072 24182 10124
rect 24581 10115 24639 10121
rect 24581 10081 24593 10115
rect 24627 10112 24639 10115
rect 27080 10112 27108 10152
rect 28721 10149 28733 10183
rect 28767 10180 28779 10183
rect 29086 10180 29092 10192
rect 28767 10152 29092 10180
rect 28767 10149 28779 10152
rect 28721 10143 28779 10149
rect 29086 10140 29092 10152
rect 29144 10180 29150 10192
rect 30282 10180 30288 10192
rect 29144 10152 30288 10180
rect 29144 10140 29150 10152
rect 30282 10140 30288 10152
rect 30340 10140 30346 10192
rect 33042 10140 33048 10192
rect 33100 10180 33106 10192
rect 34532 10180 34560 10220
rect 35158 10208 35164 10220
rect 35216 10208 35222 10260
rect 35342 10208 35348 10260
rect 35400 10248 35406 10260
rect 35400 10220 36400 10248
rect 35400 10208 35406 10220
rect 33100 10152 34560 10180
rect 33100 10140 33106 10152
rect 28810 10112 28816 10124
rect 24627 10084 27016 10112
rect 27080 10084 28816 10112
rect 24627 10081 24639 10084
rect 24581 10075 24639 10081
rect 26988 10056 27016 10084
rect 22465 10047 22523 10053
rect 21836 10016 22094 10044
rect 14553 9979 14611 9985
rect 14553 9976 14565 9979
rect 13096 9948 14565 9976
rect 14553 9945 14565 9948
rect 14599 9976 14611 9979
rect 14826 9976 14832 9988
rect 14599 9948 14832 9976
rect 14599 9945 14611 9948
rect 14553 9939 14611 9945
rect 14826 9936 14832 9948
rect 14884 9936 14890 9988
rect 15286 9936 15292 9988
rect 15344 9936 15350 9988
rect 15838 9936 15844 9988
rect 15896 9976 15902 9988
rect 16206 9976 16212 9988
rect 15896 9948 16212 9976
rect 15896 9936 15902 9948
rect 16206 9936 16212 9948
rect 16264 9976 16270 9988
rect 20533 9979 20591 9985
rect 16264 9948 18552 9976
rect 16264 9936 16270 9948
rect 12434 9868 12440 9920
rect 12492 9908 12498 9920
rect 13078 9908 13084 9920
rect 12492 9880 13084 9908
rect 12492 9868 12498 9880
rect 13078 9868 13084 9880
rect 13136 9868 13142 9920
rect 13906 9868 13912 9920
rect 13964 9908 13970 9920
rect 14458 9908 14464 9920
rect 13964 9880 14464 9908
rect 13964 9868 13970 9880
rect 14458 9868 14464 9880
rect 14516 9908 14522 9920
rect 16025 9911 16083 9917
rect 16025 9908 16037 9911
rect 14516 9880 16037 9908
rect 14516 9868 14522 9880
rect 16025 9877 16037 9880
rect 16071 9908 16083 9911
rect 16114 9908 16120 9920
rect 16071 9880 16120 9908
rect 16071 9877 16083 9880
rect 16025 9871 16083 9877
rect 16114 9868 16120 9880
rect 16172 9868 16178 9920
rect 16942 9868 16948 9920
rect 17000 9868 17006 9920
rect 17310 9868 17316 9920
rect 17368 9868 17374 9920
rect 18524 9917 18552 9948
rect 20533 9945 20545 9979
rect 20579 9976 20591 9979
rect 20806 9976 20812 9988
rect 20579 9948 20812 9976
rect 20579 9945 20591 9948
rect 20533 9939 20591 9945
rect 20806 9936 20812 9948
rect 20864 9936 20870 9988
rect 21174 9936 21180 9988
rect 21232 9936 21238 9988
rect 22066 9976 22094 10016
rect 22465 10013 22477 10047
rect 22511 10044 22523 10047
rect 22554 10044 22560 10056
rect 22511 10016 22560 10044
rect 22511 10013 22523 10016
rect 22465 10007 22523 10013
rect 22554 10004 22560 10016
rect 22612 10004 22618 10056
rect 25958 10004 25964 10056
rect 26016 10044 26022 10056
rect 26510 10044 26516 10056
rect 26016 10016 26516 10044
rect 26016 10004 26022 10016
rect 26510 10004 26516 10016
rect 26568 10004 26574 10056
rect 26970 10004 26976 10056
rect 27028 10004 27034 10056
rect 28368 10030 28396 10084
rect 28810 10072 28816 10084
rect 28868 10112 28874 10124
rect 28997 10115 29055 10121
rect 28997 10112 29009 10115
rect 28868 10084 29009 10112
rect 28868 10072 28874 10084
rect 28997 10081 29009 10084
rect 29043 10081 29055 10115
rect 28997 10075 29055 10081
rect 29362 10072 29368 10124
rect 29420 10072 29426 10124
rect 29733 10115 29791 10121
rect 29733 10081 29745 10115
rect 29779 10112 29791 10115
rect 32674 10112 32680 10124
rect 29779 10084 32680 10112
rect 29779 10081 29791 10084
rect 29733 10075 29791 10081
rect 32674 10072 32680 10084
rect 32732 10072 32738 10124
rect 33226 10072 33232 10124
rect 33284 10072 33290 10124
rect 34054 10072 34060 10124
rect 34112 10112 34118 10124
rect 34885 10115 34943 10121
rect 34885 10112 34897 10115
rect 34112 10084 34897 10112
rect 34112 10072 34118 10084
rect 34885 10081 34897 10084
rect 34931 10081 34943 10115
rect 34885 10075 34943 10081
rect 35161 10115 35219 10121
rect 35161 10081 35173 10115
rect 35207 10112 35219 10115
rect 35250 10112 35256 10124
rect 35207 10084 35256 10112
rect 35207 10081 35219 10084
rect 35161 10075 35219 10081
rect 35250 10072 35256 10084
rect 35308 10072 35314 10124
rect 30374 10004 30380 10056
rect 30432 10004 30438 10056
rect 31754 10004 31760 10056
rect 31812 10004 31818 10056
rect 36372 10044 36400 10220
rect 36630 10208 36636 10260
rect 36688 10208 36694 10260
rect 36722 10208 36728 10260
rect 36780 10248 36786 10260
rect 36909 10251 36967 10257
rect 36909 10248 36921 10251
rect 36780 10220 36921 10248
rect 36780 10208 36786 10220
rect 36909 10217 36921 10220
rect 36955 10217 36967 10251
rect 36909 10211 36967 10217
rect 49142 10072 49148 10124
rect 49200 10072 49206 10124
rect 38289 10047 38347 10053
rect 38289 10044 38301 10047
rect 36372 10016 38301 10044
rect 38289 10013 38301 10016
rect 38335 10044 38347 10047
rect 38749 10047 38807 10053
rect 38749 10044 38761 10047
rect 38335 10016 38761 10044
rect 38335 10013 38347 10016
rect 38289 10007 38347 10013
rect 38749 10013 38761 10016
rect 38795 10013 38807 10047
rect 40589 10047 40647 10053
rect 40589 10044 40601 10047
rect 38749 10007 38807 10013
rect 40144 10016 40601 10044
rect 22066 9948 24808 9976
rect 18509 9911 18567 9917
rect 18509 9877 18521 9911
rect 18555 9908 18567 9911
rect 21542 9908 21548 9920
rect 18555 9880 21548 9908
rect 18555 9877 18567 9880
rect 18509 9871 18567 9877
rect 21542 9868 21548 9880
rect 21600 9868 21606 9920
rect 21818 9868 21824 9920
rect 21876 9908 21882 9920
rect 22005 9911 22063 9917
rect 22005 9908 22017 9911
rect 21876 9880 22017 9908
rect 21876 9868 21882 9880
rect 22005 9877 22017 9880
rect 22051 9877 22063 9911
rect 22005 9871 22063 9877
rect 23934 9868 23940 9920
rect 23992 9908 23998 9920
rect 24029 9911 24087 9917
rect 24029 9908 24041 9911
rect 23992 9880 24041 9908
rect 23992 9868 23998 9880
rect 24029 9877 24041 9880
rect 24075 9877 24087 9911
rect 24780 9908 24808 9948
rect 24854 9936 24860 9988
rect 24912 9936 24918 9988
rect 26326 9936 26332 9988
rect 26384 9976 26390 9988
rect 27249 9979 27307 9985
rect 27249 9976 27261 9979
rect 26384 9948 27261 9976
rect 26384 9936 26390 9948
rect 27249 9945 27261 9948
rect 27295 9945 27307 9979
rect 30098 9976 30104 9988
rect 27249 9939 27307 9945
rect 28920 9948 30104 9976
rect 26142 9908 26148 9920
rect 24780 9880 26148 9908
rect 24029 9871 24087 9877
rect 26142 9868 26148 9880
rect 26200 9868 26206 9920
rect 27264 9908 27292 9939
rect 28920 9908 28948 9948
rect 30098 9936 30104 9948
rect 30156 9936 30162 9988
rect 30650 9936 30656 9988
rect 30708 9936 30714 9988
rect 32953 9979 33011 9985
rect 32953 9976 32965 9979
rect 31956 9948 32965 9976
rect 27264 9880 28948 9908
rect 28994 9868 29000 9920
rect 29052 9908 29058 9920
rect 31956 9908 31984 9948
rect 32953 9945 32965 9948
rect 32999 9945 33011 9979
rect 32953 9939 33011 9945
rect 33134 9936 33140 9988
rect 33192 9976 33198 9988
rect 33781 9979 33839 9985
rect 33781 9976 33793 9979
rect 33192 9948 33793 9976
rect 33192 9936 33198 9948
rect 33781 9945 33793 9948
rect 33827 9945 33839 9979
rect 36722 9976 36728 9988
rect 36386 9948 36728 9976
rect 33781 9939 33839 9945
rect 29052 9880 31984 9908
rect 29052 9868 29058 9880
rect 32674 9868 32680 9920
rect 32732 9908 32738 9920
rect 33045 9911 33103 9917
rect 33045 9908 33057 9911
rect 32732 9880 33057 9908
rect 32732 9868 32738 9880
rect 33045 9877 33057 9880
rect 33091 9877 33103 9911
rect 33045 9871 33103 9877
rect 35802 9868 35808 9920
rect 35860 9908 35866 9920
rect 36464 9908 36492 9948
rect 36722 9936 36728 9948
rect 36780 9936 36786 9988
rect 38562 9936 38568 9988
rect 38620 9976 38626 9988
rect 40144 9985 40172 10016
rect 40589 10013 40601 10016
rect 40635 10013 40647 10047
rect 40589 10007 40647 10013
rect 41598 10004 41604 10056
rect 41656 10044 41662 10056
rect 44361 10047 44419 10053
rect 44361 10044 44373 10047
rect 41656 10016 44373 10044
rect 41656 10004 41662 10016
rect 44361 10013 44373 10016
rect 44407 10013 44419 10047
rect 44361 10007 44419 10013
rect 45738 10004 45744 10056
rect 45796 10044 45802 10056
rect 46109 10047 46167 10053
rect 46109 10044 46121 10047
rect 45796 10016 46121 10044
rect 45796 10004 45802 10016
rect 46109 10013 46121 10016
rect 46155 10013 46167 10047
rect 46109 10007 46167 10013
rect 46290 10004 46296 10056
rect 46348 10044 46354 10056
rect 47949 10047 48007 10053
rect 47949 10044 47961 10047
rect 46348 10016 47961 10044
rect 46348 10004 46354 10016
rect 47949 10013 47961 10016
rect 47995 10013 48007 10047
rect 47949 10007 48007 10013
rect 40129 9979 40187 9985
rect 40129 9976 40141 9979
rect 38620 9948 40141 9976
rect 38620 9936 38626 9948
rect 40129 9945 40141 9948
rect 40175 9945 40187 9979
rect 40129 9939 40187 9945
rect 40313 9979 40371 9985
rect 40313 9945 40325 9979
rect 40359 9976 40371 9979
rect 44545 9979 44603 9985
rect 40359 9948 42932 9976
rect 40359 9945 40371 9948
rect 40313 9939 40371 9945
rect 35860 9880 36492 9908
rect 35860 9868 35866 9880
rect 38378 9868 38384 9920
rect 38436 9868 38442 9920
rect 42904 9908 42932 9948
rect 44545 9945 44557 9979
rect 44591 9976 44603 9979
rect 46014 9976 46020 9988
rect 44591 9948 46020 9976
rect 44591 9945 44603 9948
rect 44545 9939 44603 9945
rect 46014 9936 46020 9948
rect 46072 9936 46078 9988
rect 47302 9936 47308 9988
rect 47360 9936 47366 9988
rect 45830 9908 45836 9920
rect 42904 9880 45836 9908
rect 45830 9868 45836 9880
rect 45888 9868 45894 9920
rect 1104 9818 49864 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 27950 9818
rect 28002 9766 28014 9818
rect 28066 9766 28078 9818
rect 28130 9766 28142 9818
rect 28194 9766 28206 9818
rect 28258 9766 37950 9818
rect 38002 9766 38014 9818
rect 38066 9766 38078 9818
rect 38130 9766 38142 9818
rect 38194 9766 38206 9818
rect 38258 9766 47950 9818
rect 48002 9766 48014 9818
rect 48066 9766 48078 9818
rect 48130 9766 48142 9818
rect 48194 9766 48206 9818
rect 48258 9766 49864 9818
rect 1104 9744 49864 9766
rect 1302 9664 1308 9716
rect 1360 9704 1366 9716
rect 2133 9707 2191 9713
rect 2133 9704 2145 9707
rect 1360 9676 2145 9704
rect 1360 9664 1366 9676
rect 2133 9673 2145 9676
rect 2179 9673 2191 9707
rect 2133 9667 2191 9673
rect 16574 9664 16580 9716
rect 16632 9704 16638 9716
rect 17310 9704 17316 9716
rect 16632 9676 17316 9704
rect 16632 9664 16638 9676
rect 17310 9664 17316 9676
rect 17368 9664 17374 9716
rect 20898 9664 20904 9716
rect 20956 9704 20962 9716
rect 21085 9707 21143 9713
rect 21085 9704 21097 9707
rect 20956 9676 21097 9704
rect 20956 9664 20962 9676
rect 21085 9673 21097 9676
rect 21131 9673 21143 9707
rect 21085 9667 21143 9673
rect 21174 9664 21180 9716
rect 21232 9704 21238 9716
rect 21726 9704 21732 9716
rect 21232 9676 21732 9704
rect 21232 9664 21238 9676
rect 21726 9664 21732 9676
rect 21784 9664 21790 9716
rect 22278 9664 22284 9716
rect 22336 9664 22342 9716
rect 31478 9704 31484 9716
rect 23676 9676 25084 9704
rect 12526 9596 12532 9648
rect 12584 9596 12590 9648
rect 12618 9596 12624 9648
rect 12676 9596 12682 9648
rect 12710 9596 12716 9648
rect 12768 9596 12774 9648
rect 15286 9636 15292 9648
rect 14858 9608 15292 9636
rect 15286 9596 15292 9608
rect 15344 9596 15350 9648
rect 15381 9639 15439 9645
rect 15381 9605 15393 9639
rect 15427 9636 15439 9639
rect 17218 9636 17224 9648
rect 15427 9608 17224 9636
rect 15427 9605 15439 9608
rect 15381 9599 15439 9605
rect 17218 9596 17224 9608
rect 17276 9596 17282 9648
rect 17402 9596 17408 9648
rect 17460 9636 17466 9648
rect 17460 9608 17618 9636
rect 17460 9596 17466 9608
rect 18874 9596 18880 9648
rect 18932 9596 18938 9648
rect 19518 9596 19524 9648
rect 19576 9636 19582 9648
rect 19613 9639 19671 9645
rect 19613 9636 19625 9639
rect 19576 9608 19625 9636
rect 19576 9596 19582 9608
rect 19613 9605 19625 9608
rect 19659 9605 19671 9639
rect 19613 9599 19671 9605
rect 21450 9596 21456 9648
rect 21508 9636 21514 9648
rect 21545 9639 21603 9645
rect 21545 9636 21557 9639
rect 21508 9608 21557 9636
rect 21508 9596 21514 9608
rect 21545 9605 21557 9608
rect 21591 9636 21603 9639
rect 22741 9639 22799 9645
rect 22741 9636 22753 9639
rect 21591 9608 22753 9636
rect 21591 9605 21603 9608
rect 21545 9599 21603 9605
rect 22741 9605 22753 9608
rect 22787 9636 22799 9639
rect 23676 9636 23704 9676
rect 22787 9608 23704 9636
rect 22787 9605 22799 9608
rect 22741 9599 22799 9605
rect 23750 9596 23756 9648
rect 23808 9596 23814 9648
rect 25056 9636 25084 9676
rect 28184 9676 29132 9704
rect 25590 9636 25596 9648
rect 25056 9608 25596 9636
rect 25590 9596 25596 9608
rect 25648 9596 25654 9648
rect 25958 9636 25964 9648
rect 25700 9608 25964 9636
rect 1302 9528 1308 9580
rect 1360 9568 1366 9580
rect 1581 9571 1639 9577
rect 1581 9568 1593 9571
rect 1360 9540 1593 9568
rect 1360 9528 1366 9540
rect 1581 9537 1593 9540
rect 1627 9568 1639 9571
rect 2317 9571 2375 9577
rect 2317 9568 2329 9571
rect 1627 9540 2329 9568
rect 1627 9537 1639 9540
rect 1581 9531 1639 9537
rect 2317 9537 2329 9540
rect 2363 9537 2375 9571
rect 2317 9531 2375 9537
rect 12728 9509 12756 9596
rect 16117 9571 16175 9577
rect 16117 9537 16129 9571
rect 16163 9568 16175 9571
rect 16206 9568 16212 9580
rect 16163 9540 16212 9568
rect 16163 9537 16175 9540
rect 16117 9531 16175 9537
rect 16206 9528 16212 9540
rect 16264 9528 16270 9580
rect 16482 9528 16488 9580
rect 16540 9528 16546 9580
rect 21082 9568 21088 9580
rect 20746 9540 21088 9568
rect 21082 9528 21088 9540
rect 21140 9528 21146 9580
rect 22646 9528 22652 9580
rect 22704 9528 22710 9580
rect 23474 9528 23480 9580
rect 23532 9528 23538 9580
rect 25314 9568 25320 9580
rect 24886 9554 25320 9568
rect 24872 9540 25320 9554
rect 12713 9503 12771 9509
rect 12713 9469 12725 9503
rect 12759 9469 12771 9503
rect 12713 9463 12771 9469
rect 13357 9503 13415 9509
rect 13357 9469 13369 9503
rect 13403 9469 13415 9503
rect 13357 9463 13415 9469
rect 1762 9392 1768 9444
rect 1820 9392 1826 9444
rect 12161 9367 12219 9373
rect 12161 9333 12173 9367
rect 12207 9364 12219 9367
rect 12802 9364 12808 9376
rect 12207 9336 12808 9364
rect 12207 9333 12219 9336
rect 12161 9327 12219 9333
rect 12802 9324 12808 9336
rect 12860 9324 12866 9376
rect 13372 9364 13400 9463
rect 13630 9460 13636 9512
rect 13688 9460 13694 9512
rect 14182 9460 14188 9512
rect 14240 9500 14246 9512
rect 16666 9500 16672 9512
rect 14240 9472 16672 9500
rect 14240 9460 14246 9472
rect 16666 9460 16672 9472
rect 16724 9460 16730 9512
rect 16758 9460 16764 9512
rect 16816 9500 16822 9512
rect 16853 9503 16911 9509
rect 16853 9500 16865 9503
rect 16816 9472 16865 9500
rect 16816 9460 16822 9472
rect 16853 9469 16865 9472
rect 16899 9469 16911 9503
rect 16853 9463 16911 9469
rect 17129 9503 17187 9509
rect 17129 9469 17141 9503
rect 17175 9500 17187 9503
rect 18598 9500 18604 9512
rect 17175 9472 18604 9500
rect 17175 9469 17187 9472
rect 17129 9463 17187 9469
rect 14918 9392 14924 9444
rect 14976 9432 14982 9444
rect 15841 9435 15899 9441
rect 15841 9432 15853 9435
rect 14976 9404 15853 9432
rect 14976 9392 14982 9404
rect 15841 9401 15853 9404
rect 15887 9432 15899 9435
rect 16574 9432 16580 9444
rect 15887 9404 16580 9432
rect 15887 9401 15899 9404
rect 15841 9395 15899 9401
rect 16574 9392 16580 9404
rect 16632 9392 16638 9444
rect 13814 9364 13820 9376
rect 13372 9336 13820 9364
rect 13814 9324 13820 9336
rect 13872 9324 13878 9376
rect 15286 9324 15292 9376
rect 15344 9364 15350 9376
rect 15657 9367 15715 9373
rect 15657 9364 15669 9367
rect 15344 9336 15669 9364
rect 15344 9324 15350 9336
rect 15657 9333 15669 9336
rect 15703 9364 15715 9367
rect 16209 9367 16267 9373
rect 16209 9364 16221 9367
rect 15703 9336 16221 9364
rect 15703 9333 15715 9336
rect 15657 9327 15715 9333
rect 16209 9333 16221 9336
rect 16255 9333 16267 9367
rect 16868 9364 16896 9463
rect 18598 9460 18604 9472
rect 18656 9460 18662 9512
rect 19337 9503 19395 9509
rect 19337 9469 19349 9503
rect 19383 9469 19395 9503
rect 19337 9463 19395 9469
rect 22925 9503 22983 9509
rect 22925 9469 22937 9503
rect 22971 9500 22983 9503
rect 22971 9472 23612 9500
rect 22971 9469 22983 9472
rect 22925 9463 22983 9469
rect 19352 9364 19380 9463
rect 22554 9392 22560 9444
rect 22612 9432 22618 9444
rect 22940 9432 22968 9463
rect 22612 9404 22968 9432
rect 22612 9392 22618 9404
rect 16868 9336 19380 9364
rect 16209 9327 16267 9333
rect 21082 9324 21088 9376
rect 21140 9364 21146 9376
rect 21361 9367 21419 9373
rect 21361 9364 21373 9367
rect 21140 9336 21373 9364
rect 21140 9324 21146 9336
rect 21361 9333 21373 9336
rect 21407 9364 21419 9367
rect 21726 9364 21732 9376
rect 21407 9336 21732 9364
rect 21407 9333 21419 9336
rect 21361 9327 21419 9333
rect 21726 9324 21732 9336
rect 21784 9364 21790 9376
rect 21913 9367 21971 9373
rect 21913 9364 21925 9367
rect 21784 9336 21925 9364
rect 21784 9324 21790 9336
rect 21913 9333 21925 9336
rect 21959 9364 21971 9367
rect 23382 9364 23388 9376
rect 21959 9336 23388 9364
rect 21959 9333 21971 9336
rect 21913 9327 21971 9333
rect 23382 9324 23388 9336
rect 23440 9324 23446 9376
rect 23584 9364 23612 9472
rect 23842 9460 23848 9512
rect 23900 9500 23906 9512
rect 24872 9500 24900 9540
rect 25314 9528 25320 9540
rect 25372 9568 25378 9580
rect 25700 9568 25728 9608
rect 25958 9596 25964 9608
rect 26016 9596 26022 9648
rect 27801 9639 27859 9645
rect 27801 9605 27813 9639
rect 27847 9636 27859 9639
rect 28184 9636 28212 9676
rect 27847 9608 28212 9636
rect 27847 9605 27859 9608
rect 27801 9599 27859 9605
rect 28810 9596 28816 9648
rect 28868 9596 28874 9648
rect 29104 9636 29132 9676
rect 30392 9676 31484 9704
rect 30392 9636 30420 9676
rect 31478 9664 31484 9676
rect 31536 9664 31542 9716
rect 31754 9664 31760 9716
rect 31812 9704 31818 9716
rect 31849 9707 31907 9713
rect 31849 9704 31861 9707
rect 31812 9676 31861 9704
rect 31812 9664 31818 9676
rect 31849 9673 31861 9676
rect 31895 9704 31907 9707
rect 32309 9707 32367 9713
rect 32309 9704 32321 9707
rect 31895 9676 32321 9704
rect 31895 9673 31907 9676
rect 31849 9667 31907 9673
rect 32309 9673 32321 9676
rect 32355 9704 32367 9707
rect 32674 9704 32680 9716
rect 32355 9676 32680 9704
rect 32355 9673 32367 9676
rect 32309 9667 32367 9673
rect 32674 9664 32680 9676
rect 32732 9704 32738 9716
rect 33318 9704 33324 9716
rect 32732 9676 33324 9704
rect 32732 9664 32738 9676
rect 33318 9664 33324 9676
rect 33376 9664 33382 9716
rect 35802 9664 35808 9716
rect 35860 9704 35866 9716
rect 35897 9707 35955 9713
rect 35897 9704 35909 9707
rect 35860 9676 35909 9704
rect 35860 9664 35866 9676
rect 35897 9673 35909 9676
rect 35943 9704 35955 9707
rect 35943 9676 36032 9704
rect 35943 9673 35955 9676
rect 35897 9667 35955 9673
rect 29104 9608 30420 9636
rect 30558 9596 30564 9648
rect 30616 9596 30622 9648
rect 31294 9596 31300 9648
rect 31352 9636 31358 9648
rect 32953 9639 33011 9645
rect 32953 9636 32965 9639
rect 31352 9608 32965 9636
rect 31352 9596 31358 9608
rect 32953 9605 32965 9608
rect 32999 9605 33011 9639
rect 34054 9636 34060 9648
rect 32953 9599 33011 9605
rect 33888 9608 34060 9636
rect 25372 9540 25728 9568
rect 25372 9528 25378 9540
rect 25774 9528 25780 9580
rect 25832 9568 25838 9580
rect 26053 9571 26111 9577
rect 26053 9568 26065 9571
rect 25832 9540 26065 9568
rect 25832 9528 25838 9540
rect 26053 9537 26065 9540
rect 26099 9537 26111 9571
rect 26053 9531 26111 9537
rect 26142 9528 26148 9580
rect 26200 9528 26206 9580
rect 33888 9577 33916 9608
rect 34054 9596 34060 9608
rect 34112 9596 34118 9648
rect 34146 9596 34152 9648
rect 34204 9596 34210 9648
rect 35526 9636 35532 9648
rect 35374 9608 35532 9636
rect 35526 9596 35532 9608
rect 35584 9636 35590 9648
rect 36004 9636 36032 9676
rect 38378 9664 38384 9716
rect 38436 9704 38442 9716
rect 47026 9704 47032 9716
rect 38436 9676 47032 9704
rect 38436 9664 38442 9676
rect 47026 9664 47032 9676
rect 47084 9664 47090 9716
rect 35584 9608 36032 9636
rect 49145 9639 49203 9645
rect 35584 9596 35590 9608
rect 49145 9605 49157 9639
rect 49191 9636 49203 9639
rect 49326 9636 49332 9648
rect 49191 9608 49332 9636
rect 49191 9605 49203 9608
rect 49145 9599 49203 9605
rect 49326 9596 49332 9608
rect 49384 9596 49390 9648
rect 33873 9571 33931 9577
rect 31220 9540 33180 9568
rect 23900 9472 24900 9500
rect 23900 9460 23906 9472
rect 26326 9460 26332 9512
rect 26384 9460 26390 9512
rect 26970 9460 26976 9512
rect 27028 9500 27034 9512
rect 27525 9503 27583 9509
rect 27525 9500 27537 9503
rect 27028 9472 27537 9500
rect 27028 9460 27034 9472
rect 27525 9469 27537 9472
rect 27571 9500 27583 9503
rect 28810 9500 28816 9512
rect 27571 9472 28816 9500
rect 27571 9469 27583 9472
rect 27525 9463 27583 9469
rect 28810 9460 28816 9472
rect 28868 9500 28874 9512
rect 29546 9500 29552 9512
rect 28868 9472 29552 9500
rect 28868 9460 28874 9472
rect 29546 9460 29552 9472
rect 29604 9500 29610 9512
rect 29733 9503 29791 9509
rect 29733 9500 29745 9503
rect 29604 9472 29745 9500
rect 29604 9460 29610 9472
rect 29733 9469 29745 9472
rect 29779 9469 29791 9503
rect 30009 9503 30067 9509
rect 30009 9500 30021 9503
rect 29733 9463 29791 9469
rect 29840 9472 30021 9500
rect 29178 9392 29184 9444
rect 29236 9432 29242 9444
rect 29273 9435 29331 9441
rect 29273 9432 29285 9435
rect 29236 9404 29285 9432
rect 29236 9392 29242 9404
rect 29273 9401 29285 9404
rect 29319 9401 29331 9435
rect 29273 9395 29331 9401
rect 29638 9392 29644 9444
rect 29696 9432 29702 9444
rect 29840 9432 29868 9472
rect 30009 9469 30021 9472
rect 30055 9469 30067 9503
rect 30009 9463 30067 9469
rect 30650 9460 30656 9512
rect 30708 9500 30714 9512
rect 31220 9500 31248 9540
rect 30708 9472 31248 9500
rect 30708 9460 30714 9472
rect 31294 9460 31300 9512
rect 31352 9500 31358 9512
rect 33152 9509 33180 9540
rect 33873 9537 33885 9571
rect 33919 9537 33931 9571
rect 33873 9531 33931 9537
rect 33045 9503 33103 9509
rect 33045 9500 33057 9503
rect 31352 9472 33057 9500
rect 31352 9460 31358 9472
rect 33045 9469 33057 9472
rect 33091 9469 33103 9503
rect 33045 9463 33103 9469
rect 33137 9503 33195 9509
rect 33137 9469 33149 9503
rect 33183 9469 33195 9503
rect 33137 9463 33195 9469
rect 31662 9432 31668 9444
rect 29696 9404 29868 9432
rect 31128 9404 31668 9432
rect 29696 9392 29702 9404
rect 25225 9367 25283 9373
rect 25225 9364 25237 9367
rect 23584 9336 25237 9364
rect 25225 9333 25237 9336
rect 25271 9333 25283 9367
rect 25225 9327 25283 9333
rect 25682 9324 25688 9376
rect 25740 9324 25746 9376
rect 30374 9324 30380 9376
rect 30432 9364 30438 9376
rect 31128 9364 31156 9404
rect 31662 9392 31668 9404
rect 31720 9432 31726 9444
rect 33888 9432 33916 9531
rect 43346 9528 43352 9580
rect 43404 9568 43410 9580
rect 47949 9571 48007 9577
rect 47949 9568 47961 9571
rect 43404 9540 47961 9568
rect 43404 9528 43410 9540
rect 47949 9537 47961 9540
rect 47995 9537 48007 9571
rect 47949 9531 48007 9537
rect 31720 9404 33916 9432
rect 31720 9392 31726 9404
rect 35250 9392 35256 9444
rect 35308 9432 35314 9444
rect 35621 9435 35679 9441
rect 35621 9432 35633 9435
rect 35308 9404 35633 9432
rect 35308 9392 35314 9404
rect 35621 9401 35633 9404
rect 35667 9401 35679 9435
rect 35621 9395 35679 9401
rect 30432 9336 31156 9364
rect 32585 9367 32643 9373
rect 30432 9324 30438 9336
rect 32585 9333 32597 9367
rect 32631 9364 32643 9367
rect 35526 9364 35532 9376
rect 32631 9336 35532 9364
rect 32631 9333 32643 9336
rect 32585 9327 32643 9333
rect 35526 9324 35532 9336
rect 35584 9324 35590 9376
rect 1104 9274 49864 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 32950 9274
rect 33002 9222 33014 9274
rect 33066 9222 33078 9274
rect 33130 9222 33142 9274
rect 33194 9222 33206 9274
rect 33258 9222 42950 9274
rect 43002 9222 43014 9274
rect 43066 9222 43078 9274
rect 43130 9222 43142 9274
rect 43194 9222 43206 9274
rect 43258 9222 49864 9274
rect 1104 9200 49864 9222
rect 1765 9163 1823 9169
rect 1765 9129 1777 9163
rect 1811 9160 1823 9163
rect 14182 9160 14188 9172
rect 1811 9132 14188 9160
rect 1811 9129 1823 9132
rect 1765 9123 1823 9129
rect 14182 9120 14188 9132
rect 14240 9120 14246 9172
rect 14277 9163 14335 9169
rect 14277 9129 14289 9163
rect 14323 9160 14335 9163
rect 17862 9160 17868 9172
rect 14323 9132 17868 9160
rect 14323 9129 14335 9132
rect 14277 9123 14335 9129
rect 17862 9120 17868 9132
rect 17920 9120 17926 9172
rect 19518 9120 19524 9172
rect 19576 9160 19582 9172
rect 21177 9163 21235 9169
rect 21177 9160 21189 9163
rect 19576 9132 21189 9160
rect 19576 9120 19582 9132
rect 21177 9129 21189 9132
rect 21223 9129 21235 9163
rect 21177 9123 21235 9129
rect 24394 9120 24400 9172
rect 24452 9120 24458 9172
rect 24673 9163 24731 9169
rect 24673 9129 24685 9163
rect 24719 9160 24731 9163
rect 25314 9160 25320 9172
rect 24719 9132 25320 9160
rect 24719 9129 24731 9132
rect 24673 9123 24731 9129
rect 25314 9120 25320 9132
rect 25372 9120 25378 9172
rect 25590 9120 25596 9172
rect 25648 9160 25654 9172
rect 26142 9160 26148 9172
rect 25648 9132 26148 9160
rect 25648 9120 25654 9132
rect 26142 9120 26148 9132
rect 26200 9120 26206 9172
rect 28169 9163 28227 9169
rect 28169 9129 28181 9163
rect 28215 9160 28227 9163
rect 28994 9160 29000 9172
rect 28215 9132 29000 9160
rect 28215 9129 28227 9132
rect 28169 9123 28227 9129
rect 28994 9120 29000 9132
rect 29052 9120 29058 9172
rect 29638 9120 29644 9172
rect 29696 9160 29702 9172
rect 32493 9163 32551 9169
rect 32493 9160 32505 9163
rect 29696 9132 32505 9160
rect 29696 9120 29702 9132
rect 32493 9129 32505 9132
rect 32539 9129 32551 9163
rect 32493 9123 32551 9129
rect 32674 9120 32680 9172
rect 32732 9160 32738 9172
rect 32769 9163 32827 9169
rect 32769 9160 32781 9163
rect 32732 9132 32781 9160
rect 32732 9120 32738 9132
rect 32769 9129 32781 9132
rect 32815 9129 32827 9163
rect 32769 9123 32827 9129
rect 33321 9163 33379 9169
rect 33321 9129 33333 9163
rect 33367 9160 33379 9163
rect 35894 9160 35900 9172
rect 33367 9132 35900 9160
rect 33367 9129 33379 9132
rect 33321 9123 33379 9129
rect 35894 9120 35900 9132
rect 35952 9120 35958 9172
rect 36541 9163 36599 9169
rect 36541 9129 36553 9163
rect 36587 9160 36599 9163
rect 43622 9160 43628 9172
rect 36587 9132 43628 9160
rect 36587 9129 36599 9132
rect 36541 9123 36599 9129
rect 43622 9120 43628 9132
rect 43680 9120 43686 9172
rect 2314 9052 2320 9104
rect 2372 9092 2378 9104
rect 11146 9092 11152 9104
rect 2372 9064 11152 9092
rect 2372 9052 2378 9064
rect 11146 9052 11152 9064
rect 11204 9052 11210 9104
rect 13814 9052 13820 9104
rect 13872 9092 13878 9104
rect 13872 9064 16436 9092
rect 13872 9052 13878 9064
rect 2869 9027 2927 9033
rect 2869 9024 2881 9027
rect 2332 8996 2881 9024
rect 1210 8916 1216 8968
rect 1268 8956 1274 8968
rect 2332 8965 2360 8996
rect 2869 8993 2881 8996
rect 2915 8993 2927 9027
rect 2869 8987 2927 8993
rect 13630 8984 13636 9036
rect 13688 9024 13694 9036
rect 15378 9024 15384 9036
rect 13688 8996 15384 9024
rect 13688 8984 13694 8996
rect 15378 8984 15384 8996
rect 15436 9024 15442 9036
rect 16408 9033 16436 9064
rect 25682 9052 25688 9104
rect 25740 9092 25746 9104
rect 30466 9092 30472 9104
rect 25740 9064 30472 9092
rect 25740 9052 25746 9064
rect 30466 9052 30472 9064
rect 30524 9052 30530 9104
rect 32306 9052 32312 9104
rect 32364 9092 32370 9104
rect 35710 9092 35716 9104
rect 32364 9064 35716 9092
rect 32364 9052 32370 9064
rect 35710 9052 35716 9064
rect 35768 9052 35774 9104
rect 15749 9027 15807 9033
rect 15749 9024 15761 9027
rect 15436 8996 15761 9024
rect 15436 8984 15442 8996
rect 15749 8993 15761 8996
rect 15795 8993 15807 9027
rect 15749 8987 15807 8993
rect 16393 9027 16451 9033
rect 16393 8993 16405 9027
rect 16439 9024 16451 9027
rect 16758 9024 16764 9036
rect 16439 8996 16764 9024
rect 16439 8993 16451 8996
rect 16393 8987 16451 8993
rect 16758 8984 16764 8996
rect 16816 8984 16822 9036
rect 17034 8984 17040 9036
rect 17092 9024 17098 9036
rect 18141 9027 18199 9033
rect 18141 9024 18153 9027
rect 17092 8996 18153 9024
rect 17092 8984 17098 8996
rect 18141 8993 18153 8996
rect 18187 8993 18199 9027
rect 18141 8987 18199 8993
rect 18690 8984 18696 9036
rect 18748 8984 18754 9036
rect 19429 9027 19487 9033
rect 19429 8993 19441 9027
rect 19475 9024 19487 9027
rect 19702 9024 19708 9036
rect 19475 8996 19708 9024
rect 19475 8993 19487 8996
rect 19429 8987 19487 8993
rect 19702 8984 19708 8996
rect 19760 8984 19766 9036
rect 22002 8984 22008 9036
rect 22060 9024 22066 9036
rect 22281 9027 22339 9033
rect 22281 9024 22293 9027
rect 22060 8996 22293 9024
rect 22060 8984 22066 8996
rect 22281 8993 22293 8996
rect 22327 8993 22339 9027
rect 22281 8987 22339 8993
rect 22554 8984 22560 9036
rect 22612 8984 22618 9036
rect 22646 8984 22652 9036
rect 22704 9024 22710 9036
rect 24854 9024 24860 9036
rect 22704 8996 24860 9024
rect 22704 8984 22710 8996
rect 24854 8984 24860 8996
rect 24912 8984 24918 9036
rect 28813 9027 28871 9033
rect 28813 8993 28825 9027
rect 28859 9024 28871 9027
rect 29638 9024 29644 9036
rect 28859 8996 29644 9024
rect 28859 8993 28871 8996
rect 28813 8987 28871 8993
rect 29638 8984 29644 8996
rect 29696 8984 29702 9036
rect 30374 8984 30380 9036
rect 30432 9024 30438 9036
rect 30745 9027 30803 9033
rect 30745 9024 30757 9027
rect 30432 8996 30757 9024
rect 30432 8984 30438 8996
rect 30745 8993 30757 8996
rect 30791 8993 30803 9027
rect 30745 8987 30803 8993
rect 32582 8984 32588 9036
rect 32640 9024 32646 9036
rect 33965 9027 34023 9033
rect 32640 8996 33088 9024
rect 32640 8984 32646 8996
rect 2317 8959 2375 8965
rect 2317 8956 2329 8959
rect 1268 8928 2329 8956
rect 1268 8916 1274 8928
rect 2317 8925 2329 8928
rect 2363 8925 2375 8959
rect 3053 8959 3111 8965
rect 3053 8956 3065 8959
rect 2317 8919 2375 8925
rect 2424 8928 3065 8956
rect 1302 8848 1308 8900
rect 1360 8888 1366 8900
rect 1673 8891 1731 8897
rect 1673 8888 1685 8891
rect 1360 8860 1685 8888
rect 1360 8848 1366 8860
rect 1673 8857 1685 8860
rect 1719 8888 1731 8891
rect 2424 8888 2452 8928
rect 3053 8925 3065 8928
rect 3099 8925 3111 8959
rect 3053 8919 3111 8925
rect 11330 8916 11336 8968
rect 11388 8956 11394 8968
rect 14461 8959 14519 8965
rect 14461 8956 14473 8959
rect 11388 8928 14473 8956
rect 11388 8916 11394 8928
rect 14461 8925 14473 8928
rect 14507 8925 14519 8959
rect 14461 8919 14519 8925
rect 14921 8959 14979 8965
rect 14921 8925 14933 8959
rect 14967 8956 14979 8959
rect 15286 8956 15292 8968
rect 14967 8928 15292 8956
rect 14967 8925 14979 8928
rect 14921 8919 14979 8925
rect 15286 8916 15292 8928
rect 15344 8916 15350 8968
rect 15562 8916 15568 8968
rect 15620 8916 15626 8968
rect 15654 8916 15660 8968
rect 15712 8916 15718 8968
rect 32674 8956 32680 8968
rect 32154 8928 32680 8956
rect 32674 8916 32680 8928
rect 32732 8916 32738 8968
rect 33060 8965 33088 8996
rect 33965 8993 33977 9027
rect 34011 8993 34023 9027
rect 33965 8987 34023 8993
rect 33045 8959 33103 8965
rect 33045 8925 33057 8959
rect 33091 8956 33103 8959
rect 33689 8959 33747 8965
rect 33689 8956 33701 8959
rect 33091 8928 33701 8956
rect 33091 8925 33103 8928
rect 33045 8919 33103 8925
rect 33689 8925 33701 8928
rect 33735 8956 33747 8959
rect 33870 8956 33876 8968
rect 33735 8928 33876 8956
rect 33735 8925 33747 8928
rect 33689 8919 33747 8925
rect 33870 8916 33876 8928
rect 33928 8916 33934 8968
rect 33980 8956 34008 8987
rect 34054 8984 34060 9036
rect 34112 9024 34118 9036
rect 35437 9027 35495 9033
rect 35437 9024 35449 9027
rect 34112 8996 35449 9024
rect 34112 8984 34118 8996
rect 35437 8993 35449 8996
rect 35483 8993 35495 9027
rect 35437 8987 35495 8993
rect 35526 8984 35532 9036
rect 35584 9024 35590 9036
rect 49145 9027 49203 9033
rect 35584 8996 37872 9024
rect 35584 8984 35590 8996
rect 34146 8956 34152 8968
rect 33980 8928 34152 8956
rect 15102 8888 15108 8900
rect 1719 8860 2452 8888
rect 2516 8860 15108 8888
rect 1719 8857 1731 8860
rect 1673 8851 1731 8857
rect 2516 8829 2544 8860
rect 15102 8848 15108 8860
rect 15160 8848 15166 8900
rect 16574 8888 16580 8900
rect 15212 8860 16580 8888
rect 15212 8829 15240 8860
rect 16574 8848 16580 8860
rect 16632 8848 16638 8900
rect 16669 8891 16727 8897
rect 16669 8857 16681 8891
rect 16715 8857 16727 8891
rect 16669 8851 16727 8857
rect 2501 8823 2559 8829
rect 2501 8789 2513 8823
rect 2547 8789 2559 8823
rect 2501 8783 2559 8789
rect 15197 8823 15255 8829
rect 15197 8789 15209 8823
rect 15243 8789 15255 8823
rect 16684 8820 16712 8851
rect 17218 8848 17224 8900
rect 17276 8848 17282 8900
rect 19705 8891 19763 8897
rect 19705 8857 19717 8891
rect 19751 8888 19763 8891
rect 19794 8888 19800 8900
rect 19751 8860 19800 8888
rect 19751 8857 19763 8860
rect 19705 8851 19763 8857
rect 19794 8848 19800 8860
rect 19852 8848 19858 8900
rect 21082 8888 21088 8900
rect 20930 8860 21088 8888
rect 21082 8848 21088 8860
rect 21140 8848 21146 8900
rect 22094 8848 22100 8900
rect 22152 8888 22158 8900
rect 23842 8888 23848 8900
rect 22152 8860 22876 8888
rect 23782 8860 23848 8888
rect 22152 8848 22158 8860
rect 17586 8820 17592 8832
rect 16684 8792 17592 8820
rect 15197 8783 15255 8789
rect 17586 8780 17592 8792
rect 17644 8780 17650 8832
rect 21637 8823 21695 8829
rect 21637 8789 21649 8823
rect 21683 8820 21695 8823
rect 22370 8820 22376 8832
rect 21683 8792 22376 8820
rect 21683 8789 21695 8792
rect 21637 8783 21695 8789
rect 22370 8780 22376 8792
rect 22428 8780 22434 8832
rect 22848 8820 22876 8860
rect 23842 8848 23848 8860
rect 23900 8848 23906 8900
rect 28537 8891 28595 8897
rect 28537 8857 28549 8891
rect 28583 8888 28595 8891
rect 29733 8891 29791 8897
rect 29733 8888 29745 8891
rect 28583 8860 29745 8888
rect 28583 8857 28595 8860
rect 28537 8851 28595 8857
rect 29733 8857 29745 8860
rect 29779 8857 29791 8891
rect 29733 8851 29791 8857
rect 31018 8848 31024 8900
rect 31076 8848 31082 8900
rect 32582 8848 32588 8900
rect 32640 8888 32646 8900
rect 33980 8888 34008 8928
rect 34146 8916 34152 8928
rect 34204 8916 34210 8968
rect 34514 8916 34520 8968
rect 34572 8956 34578 8968
rect 37844 8965 37872 8996
rect 49145 8993 49157 9027
rect 49191 9024 49203 9027
rect 49234 9024 49240 9036
rect 49191 8996 49240 9024
rect 49191 8993 49203 8996
rect 49145 8987 49203 8993
rect 49234 8984 49240 8996
rect 49292 8984 49298 9036
rect 36725 8959 36783 8965
rect 36725 8956 36737 8959
rect 34572 8928 36737 8956
rect 34572 8916 34578 8928
rect 36725 8925 36737 8928
rect 36771 8925 36783 8959
rect 36725 8919 36783 8925
rect 37829 8959 37887 8965
rect 37829 8925 37841 8959
rect 37875 8925 37887 8959
rect 39853 8959 39911 8965
rect 39853 8956 39865 8959
rect 37829 8919 37887 8925
rect 39316 8928 39865 8956
rect 32640 8860 34008 8888
rect 32640 8848 32646 8860
rect 34974 8848 34980 8900
rect 35032 8888 35038 8900
rect 35345 8891 35403 8897
rect 35345 8888 35357 8891
rect 35032 8860 35357 8888
rect 35032 8848 35038 8860
rect 35345 8857 35357 8860
rect 35391 8857 35403 8891
rect 35345 8851 35403 8857
rect 35802 8848 35808 8900
rect 35860 8888 35866 8900
rect 39316 8897 39344 8928
rect 39853 8925 39865 8928
rect 39899 8925 39911 8959
rect 39853 8919 39911 8925
rect 43714 8916 43720 8968
rect 43772 8956 43778 8968
rect 47949 8959 48007 8965
rect 47949 8956 47961 8959
rect 43772 8928 47961 8956
rect 43772 8916 43778 8928
rect 47949 8925 47961 8928
rect 47995 8925 48007 8959
rect 47949 8919 48007 8925
rect 39301 8891 39359 8897
rect 39301 8888 39313 8891
rect 35860 8860 39313 8888
rect 35860 8848 35866 8860
rect 39301 8857 39313 8860
rect 39347 8857 39359 8891
rect 39301 8851 39359 8857
rect 39485 8891 39543 8897
rect 39485 8857 39497 8891
rect 39531 8888 39543 8891
rect 47486 8888 47492 8900
rect 39531 8860 47492 8888
rect 39531 8857 39543 8860
rect 39485 8851 39543 8857
rect 47486 8848 47492 8860
rect 47544 8848 47550 8900
rect 24029 8823 24087 8829
rect 24029 8820 24041 8823
rect 22848 8792 24041 8820
rect 24029 8789 24041 8792
rect 24075 8789 24087 8823
rect 24029 8783 24087 8789
rect 24854 8780 24860 8832
rect 24912 8780 24918 8832
rect 25682 8780 25688 8832
rect 25740 8780 25746 8832
rect 27798 8780 27804 8832
rect 27856 8820 27862 8832
rect 28626 8820 28632 8832
rect 27856 8792 28632 8820
rect 27856 8780 27862 8792
rect 28626 8780 28632 8792
rect 28684 8780 28690 8832
rect 30285 8823 30343 8829
rect 30285 8789 30297 8823
rect 30331 8820 30343 8823
rect 30374 8820 30380 8832
rect 30331 8792 30380 8820
rect 30331 8789 30343 8792
rect 30285 8783 30343 8789
rect 30374 8780 30380 8792
rect 30432 8820 30438 8832
rect 30558 8820 30564 8832
rect 30432 8792 30564 8820
rect 30432 8780 30438 8792
rect 30558 8780 30564 8792
rect 30616 8820 30622 8832
rect 31386 8820 31392 8832
rect 30616 8792 31392 8820
rect 30616 8780 30622 8792
rect 31386 8780 31392 8792
rect 31444 8780 31450 8832
rect 33778 8780 33784 8832
rect 33836 8780 33842 8832
rect 34882 8780 34888 8832
rect 34940 8780 34946 8832
rect 35250 8780 35256 8832
rect 35308 8780 35314 8832
rect 37645 8823 37703 8829
rect 37645 8789 37657 8823
rect 37691 8820 37703 8823
rect 39574 8820 39580 8832
rect 37691 8792 39580 8820
rect 37691 8789 37703 8792
rect 37645 8783 37703 8789
rect 39574 8780 39580 8792
rect 39632 8780 39638 8832
rect 1104 8730 49864 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 27950 8730
rect 28002 8678 28014 8730
rect 28066 8678 28078 8730
rect 28130 8678 28142 8730
rect 28194 8678 28206 8730
rect 28258 8678 37950 8730
rect 38002 8678 38014 8730
rect 38066 8678 38078 8730
rect 38130 8678 38142 8730
rect 38194 8678 38206 8730
rect 38258 8678 47950 8730
rect 48002 8678 48014 8730
rect 48066 8678 48078 8730
rect 48130 8678 48142 8730
rect 48194 8678 48206 8730
rect 48258 8678 49864 8730
rect 1104 8656 49864 8678
rect 15378 8576 15384 8628
rect 15436 8576 15442 8628
rect 16666 8576 16672 8628
rect 16724 8616 16730 8628
rect 17218 8616 17224 8628
rect 16724 8588 17224 8616
rect 16724 8576 16730 8588
rect 17218 8576 17224 8588
rect 17276 8616 17282 8628
rect 17276 8588 18552 8616
rect 17276 8576 17282 8588
rect 13814 8548 13820 8560
rect 13648 8520 13820 8548
rect 13648 8489 13676 8520
rect 13814 8508 13820 8520
rect 13872 8508 13878 8560
rect 13906 8508 13912 8560
rect 13964 8508 13970 8560
rect 15286 8548 15292 8560
rect 15134 8520 15292 8548
rect 15286 8508 15292 8520
rect 15344 8548 15350 8560
rect 15746 8548 15752 8560
rect 15344 8520 15752 8548
rect 15344 8508 15350 8520
rect 15746 8508 15752 8520
rect 15804 8508 15810 8560
rect 17034 8508 17040 8560
rect 17092 8548 17098 8560
rect 17129 8551 17187 8557
rect 17129 8548 17141 8551
rect 17092 8520 17141 8548
rect 17092 8508 17098 8520
rect 17129 8517 17141 8520
rect 17175 8517 17187 8551
rect 17328 8548 17356 8588
rect 17402 8548 17408 8560
rect 17328 8520 17408 8548
rect 17129 8511 17187 8517
rect 17402 8508 17408 8520
rect 17460 8548 17466 8560
rect 18524 8548 18552 8588
rect 18598 8576 18604 8628
rect 18656 8576 18662 8628
rect 19978 8576 19984 8628
rect 20036 8616 20042 8628
rect 21453 8619 21511 8625
rect 21453 8616 21465 8619
rect 20036 8588 21465 8616
rect 20036 8576 20042 8588
rect 21453 8585 21465 8588
rect 21499 8585 21511 8619
rect 21453 8579 21511 8585
rect 22094 8576 22100 8628
rect 22152 8576 22158 8628
rect 23842 8576 23848 8628
rect 23900 8616 23906 8628
rect 24029 8619 24087 8625
rect 24029 8616 24041 8619
rect 23900 8588 24041 8616
rect 23900 8576 23906 8588
rect 24029 8585 24041 8588
rect 24075 8585 24087 8619
rect 24029 8579 24087 8585
rect 30561 8619 30619 8625
rect 30561 8585 30573 8619
rect 30607 8616 30619 8619
rect 30650 8616 30656 8628
rect 30607 8588 30656 8616
rect 30607 8585 30619 8588
rect 30561 8579 30619 8585
rect 30650 8576 30656 8588
rect 30708 8576 30714 8628
rect 31018 8576 31024 8628
rect 31076 8616 31082 8628
rect 34054 8616 34060 8628
rect 31076 8588 34060 8616
rect 31076 8576 31082 8588
rect 34054 8576 34060 8588
rect 34112 8576 34118 8628
rect 34425 8619 34483 8625
rect 34425 8585 34437 8619
rect 34471 8616 34483 8619
rect 35618 8616 35624 8628
rect 34471 8588 35624 8616
rect 34471 8585 34483 8588
rect 34425 8579 34483 8585
rect 35618 8576 35624 8588
rect 35676 8576 35682 8628
rect 37461 8619 37519 8625
rect 37461 8585 37473 8619
rect 37507 8616 37519 8619
rect 40218 8616 40224 8628
rect 37507 8588 40224 8616
rect 37507 8585 37519 8588
rect 37461 8579 37519 8585
rect 40218 8576 40224 8588
rect 40276 8576 40282 8628
rect 40405 8619 40463 8625
rect 40405 8585 40417 8619
rect 40451 8616 40463 8619
rect 47670 8616 47676 8628
rect 40451 8588 47676 8616
rect 40451 8585 40463 8588
rect 40405 8579 40463 8585
rect 47670 8576 47676 8588
rect 47728 8576 47734 8628
rect 22112 8548 22140 8576
rect 22281 8551 22339 8557
rect 22281 8548 22293 8551
rect 17460 8520 17618 8548
rect 18524 8520 20470 8548
rect 22112 8520 22293 8548
rect 17460 8508 17466 8520
rect 22281 8517 22293 8520
rect 22327 8517 22339 8551
rect 23860 8548 23888 8576
rect 23506 8520 23888 8548
rect 22281 8511 22339 8517
rect 29086 8508 29092 8560
rect 29144 8508 29150 8560
rect 32582 8548 32588 8560
rect 31588 8520 32588 8548
rect 1857 8483 1915 8489
rect 1857 8449 1869 8483
rect 1903 8480 1915 8483
rect 13633 8483 13691 8489
rect 1903 8452 6914 8480
rect 1903 8449 1915 8452
rect 1857 8443 1915 8449
rect 1394 8372 1400 8424
rect 1452 8412 1458 8424
rect 1581 8415 1639 8421
rect 1581 8412 1593 8415
rect 1452 8384 1593 8412
rect 1452 8372 1458 8384
rect 1581 8381 1593 8384
rect 1627 8381 1639 8415
rect 6886 8412 6914 8452
rect 13633 8449 13645 8483
rect 13679 8449 13691 8483
rect 13633 8443 13691 8449
rect 16758 8440 16764 8492
rect 16816 8480 16822 8492
rect 16853 8483 16911 8489
rect 16853 8480 16865 8483
rect 16816 8452 16865 8480
rect 16816 8440 16822 8452
rect 16853 8449 16865 8452
rect 16899 8449 16911 8483
rect 16853 8443 16911 8449
rect 19702 8440 19708 8492
rect 19760 8440 19766 8492
rect 21082 8440 21088 8492
rect 21140 8440 21146 8492
rect 22002 8440 22008 8492
rect 22060 8440 22066 8492
rect 30374 8480 30380 8492
rect 30222 8452 30380 8480
rect 30374 8440 30380 8452
rect 30432 8480 30438 8492
rect 30650 8480 30656 8492
rect 30432 8452 30656 8480
rect 30432 8440 30438 8452
rect 30650 8440 30656 8452
rect 30708 8440 30714 8492
rect 30926 8440 30932 8492
rect 30984 8480 30990 8492
rect 31389 8483 31447 8489
rect 31389 8480 31401 8483
rect 30984 8452 31401 8480
rect 30984 8440 30990 8452
rect 31389 8449 31401 8452
rect 31435 8449 31447 8483
rect 31389 8443 31447 8449
rect 6886 8384 16896 8412
rect 1581 8375 1639 8381
rect 16868 8356 16896 8384
rect 17770 8372 17776 8424
rect 17828 8412 17834 8424
rect 19061 8415 19119 8421
rect 19061 8412 19073 8415
rect 17828 8384 19073 8412
rect 17828 8372 17834 8384
rect 19061 8381 19073 8384
rect 19107 8381 19119 8415
rect 19061 8375 19119 8381
rect 19981 8415 20039 8421
rect 19981 8381 19993 8415
rect 20027 8412 20039 8415
rect 20027 8384 22094 8412
rect 20027 8381 20039 8384
rect 19981 8375 20039 8381
rect 15746 8304 15752 8356
rect 15804 8344 15810 8356
rect 16666 8344 16672 8356
rect 15804 8316 16672 8344
rect 15804 8304 15810 8316
rect 16666 8304 16672 8316
rect 16724 8304 16730 8356
rect 16850 8304 16856 8356
rect 16908 8304 16914 8356
rect 6914 8236 6920 8288
rect 6972 8276 6978 8288
rect 15194 8276 15200 8288
rect 6972 8248 15200 8276
rect 6972 8236 6978 8248
rect 15194 8236 15200 8248
rect 15252 8236 15258 8288
rect 22066 8276 22094 8384
rect 28810 8372 28816 8424
rect 28868 8372 28874 8424
rect 31478 8372 31484 8424
rect 31536 8372 31542 8424
rect 31588 8421 31616 8520
rect 32582 8508 32588 8520
rect 32640 8508 32646 8560
rect 32674 8508 32680 8560
rect 32732 8548 32738 8560
rect 32732 8520 33074 8548
rect 32732 8508 32738 8520
rect 34882 8508 34888 8560
rect 34940 8548 34946 8560
rect 34940 8520 39160 8548
rect 34940 8508 34946 8520
rect 31662 8440 31668 8492
rect 31720 8480 31726 8492
rect 32309 8483 32367 8489
rect 32309 8480 32321 8483
rect 31720 8452 32321 8480
rect 31720 8440 31726 8452
rect 32309 8449 32321 8452
rect 32355 8449 32367 8483
rect 32309 8443 32367 8449
rect 34422 8440 34428 8492
rect 34480 8480 34486 8492
rect 39132 8489 39160 8520
rect 39574 8508 39580 8560
rect 39632 8548 39638 8560
rect 44177 8551 44235 8557
rect 44177 8548 44189 8551
rect 39632 8520 44189 8548
rect 39632 8508 39638 8520
rect 44177 8517 44189 8520
rect 44223 8517 44235 8551
rect 44177 8511 44235 8517
rect 49142 8508 49148 8560
rect 49200 8508 49206 8560
rect 37645 8483 37703 8489
rect 37645 8480 37657 8483
rect 34480 8452 37657 8480
rect 34480 8440 34486 8452
rect 37645 8449 37657 8452
rect 37691 8449 37703 8483
rect 37645 8443 37703 8449
rect 39117 8483 39175 8489
rect 39117 8449 39129 8483
rect 39163 8449 39175 8483
rect 39117 8443 39175 8449
rect 40313 8483 40371 8489
rect 40313 8449 40325 8483
rect 40359 8480 40371 8483
rect 40773 8483 40831 8489
rect 40773 8480 40785 8483
rect 40359 8452 40785 8480
rect 40359 8449 40371 8452
rect 40313 8443 40371 8449
rect 40773 8449 40785 8452
rect 40819 8449 40831 8483
rect 40773 8443 40831 8449
rect 31573 8415 31631 8421
rect 31573 8381 31585 8415
rect 31619 8381 31631 8415
rect 31573 8375 31631 8381
rect 32214 8372 32220 8424
rect 32272 8412 32278 8424
rect 32585 8415 32643 8421
rect 32585 8412 32597 8415
rect 32272 8384 32597 8412
rect 32272 8372 32278 8384
rect 32585 8381 32597 8384
rect 32631 8412 32643 8415
rect 32674 8412 32680 8424
rect 32631 8384 32680 8412
rect 32631 8381 32643 8384
rect 32585 8375 32643 8381
rect 32674 8372 32680 8384
rect 32732 8372 32738 8424
rect 33042 8372 33048 8424
rect 33100 8412 33106 8424
rect 38746 8412 38752 8424
rect 33100 8384 38752 8412
rect 33100 8372 33106 8384
rect 38746 8372 38752 8384
rect 38804 8372 38810 8424
rect 40328 8412 40356 8443
rect 45830 8440 45836 8492
rect 45888 8440 45894 8492
rect 46014 8440 46020 8492
rect 46072 8480 46078 8492
rect 47949 8483 48007 8489
rect 47949 8480 47961 8483
rect 46072 8452 47961 8480
rect 46072 8440 46078 8452
rect 47949 8449 47961 8452
rect 47995 8449 48007 8483
rect 47949 8443 48007 8449
rect 38856 8384 40356 8412
rect 23753 8347 23811 8353
rect 23753 8344 23765 8347
rect 23308 8316 23765 8344
rect 22646 8276 22652 8288
rect 22066 8248 22652 8276
rect 22646 8236 22652 8248
rect 22704 8276 22710 8288
rect 23308 8276 23336 8316
rect 23753 8313 23765 8316
rect 23799 8313 23811 8347
rect 23753 8307 23811 8313
rect 31021 8347 31079 8353
rect 31021 8313 31033 8347
rect 31067 8344 31079 8347
rect 32306 8344 32312 8356
rect 31067 8316 32312 8344
rect 31067 8313 31079 8316
rect 31021 8307 31079 8313
rect 32306 8304 32312 8316
rect 32364 8304 32370 8356
rect 33594 8304 33600 8356
rect 33652 8344 33658 8356
rect 36262 8344 36268 8356
rect 33652 8316 36268 8344
rect 33652 8304 33658 8316
rect 36262 8304 36268 8316
rect 36320 8344 36326 8356
rect 38856 8344 38884 8384
rect 46842 8372 46848 8424
rect 46900 8372 46906 8424
rect 36320 8316 38884 8344
rect 38933 8347 38991 8353
rect 36320 8304 36326 8316
rect 38933 8313 38945 8347
rect 38979 8344 38991 8347
rect 40126 8344 40132 8356
rect 38979 8316 40132 8344
rect 38979 8313 38991 8316
rect 38933 8307 38991 8313
rect 40126 8304 40132 8316
rect 40184 8304 40190 8356
rect 44361 8347 44419 8353
rect 44361 8313 44373 8347
rect 44407 8344 44419 8347
rect 47854 8344 47860 8356
rect 44407 8316 47860 8344
rect 44407 8313 44419 8316
rect 44361 8307 44419 8313
rect 47854 8304 47860 8316
rect 47912 8304 47918 8356
rect 22704 8248 23336 8276
rect 22704 8236 22710 8248
rect 27154 8236 27160 8288
rect 27212 8276 27218 8288
rect 33962 8276 33968 8288
rect 27212 8248 33968 8276
rect 27212 8236 27218 8248
rect 33962 8236 33968 8248
rect 34020 8236 34026 8288
rect 1104 8186 49864 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 32950 8186
rect 33002 8134 33014 8186
rect 33066 8134 33078 8186
rect 33130 8134 33142 8186
rect 33194 8134 33206 8186
rect 33258 8134 42950 8186
rect 43002 8134 43014 8186
rect 43066 8134 43078 8186
rect 43130 8134 43142 8186
rect 43194 8134 43206 8186
rect 43258 8134 49864 8186
rect 1104 8112 49864 8134
rect 1394 8032 1400 8084
rect 1452 8072 1458 8084
rect 2133 8075 2191 8081
rect 2133 8072 2145 8075
rect 1452 8044 2145 8072
rect 1452 8032 1458 8044
rect 2133 8041 2145 8044
rect 2179 8041 2191 8075
rect 2133 8035 2191 8041
rect 15565 8075 15623 8081
rect 15565 8041 15577 8075
rect 15611 8072 15623 8075
rect 18874 8072 18880 8084
rect 15611 8044 18880 8072
rect 15611 8041 15623 8044
rect 15565 8035 15623 8041
rect 18874 8032 18880 8044
rect 18932 8032 18938 8084
rect 19794 8032 19800 8084
rect 19852 8072 19858 8084
rect 21177 8075 21235 8081
rect 21177 8072 21189 8075
rect 19852 8044 21189 8072
rect 19852 8032 19858 8044
rect 21177 8041 21189 8044
rect 21223 8041 21235 8075
rect 21177 8035 21235 8041
rect 21910 8032 21916 8084
rect 21968 8072 21974 8084
rect 22005 8075 22063 8081
rect 22005 8072 22017 8075
rect 21968 8044 22017 8072
rect 21968 8032 21974 8044
rect 22005 8041 22017 8044
rect 22051 8041 22063 8075
rect 22005 8035 22063 8041
rect 31021 8075 31079 8081
rect 31021 8041 31033 8075
rect 31067 8072 31079 8075
rect 31067 8044 33548 8072
rect 31067 8041 31079 8044
rect 31021 8035 31079 8041
rect 17034 7964 17040 8016
rect 17092 8004 17098 8016
rect 17865 8007 17923 8013
rect 17092 7976 17264 8004
rect 17092 7964 17098 7976
rect 13998 7936 14004 7948
rect 6886 7908 14004 7936
rect 1302 7828 1308 7880
rect 1360 7868 1366 7880
rect 1581 7871 1639 7877
rect 1581 7868 1593 7871
rect 1360 7840 1593 7868
rect 1360 7828 1366 7840
rect 1581 7837 1593 7840
rect 1627 7868 1639 7871
rect 2317 7871 2375 7877
rect 2317 7868 2329 7871
rect 1627 7840 2329 7868
rect 1627 7837 1639 7840
rect 1581 7831 1639 7837
rect 2317 7837 2329 7840
rect 2363 7837 2375 7871
rect 2317 7831 2375 7837
rect 2406 7828 2412 7880
rect 2464 7868 2470 7880
rect 6886 7868 6914 7908
rect 13998 7896 14004 7908
rect 14056 7896 14062 7948
rect 16942 7896 16948 7948
rect 17000 7936 17006 7948
rect 17236 7945 17264 7976
rect 17865 7973 17877 8007
rect 17911 8004 17923 8007
rect 19242 8004 19248 8016
rect 17911 7976 19248 8004
rect 17911 7973 17923 7976
rect 17865 7967 17923 7973
rect 19242 7964 19248 7976
rect 19300 7964 19306 8016
rect 24854 7964 24860 8016
rect 24912 8004 24918 8016
rect 32766 8004 32772 8016
rect 24912 7976 32772 8004
rect 24912 7964 24918 7976
rect 32766 7964 32772 7976
rect 32824 7964 32830 8016
rect 33410 8004 33416 8016
rect 32876 7976 33416 8004
rect 17129 7939 17187 7945
rect 17129 7936 17141 7939
rect 17000 7908 17141 7936
rect 17000 7896 17006 7908
rect 17129 7905 17141 7908
rect 17175 7905 17187 7939
rect 17129 7899 17187 7905
rect 17221 7939 17279 7945
rect 17221 7905 17233 7939
rect 17267 7905 17279 7939
rect 17221 7899 17279 7905
rect 18509 7939 18567 7945
rect 18509 7905 18521 7939
rect 18555 7936 18567 7939
rect 18598 7936 18604 7948
rect 18555 7908 18604 7936
rect 18555 7905 18567 7908
rect 18509 7899 18567 7905
rect 18598 7896 18604 7908
rect 18656 7896 18662 7948
rect 19429 7939 19487 7945
rect 19429 7905 19441 7939
rect 19475 7936 19487 7939
rect 19702 7936 19708 7948
rect 19475 7908 19708 7936
rect 19475 7905 19487 7908
rect 19429 7899 19487 7905
rect 19702 7896 19708 7908
rect 19760 7896 19766 7948
rect 22649 7939 22707 7945
rect 22649 7905 22661 7939
rect 22695 7936 22707 7939
rect 23658 7936 23664 7948
rect 22695 7908 23664 7936
rect 22695 7905 22707 7908
rect 22649 7899 22707 7905
rect 23658 7896 23664 7908
rect 23716 7896 23722 7948
rect 29730 7896 29736 7948
rect 29788 7896 29794 7948
rect 30558 7896 30564 7948
rect 30616 7936 30622 7948
rect 31478 7936 31484 7948
rect 30616 7908 31484 7936
rect 30616 7896 30622 7908
rect 31478 7896 31484 7908
rect 31536 7896 31542 7948
rect 31665 7939 31723 7945
rect 31665 7905 31677 7939
rect 31711 7936 31723 7939
rect 32214 7936 32220 7948
rect 31711 7908 32220 7936
rect 31711 7905 31723 7908
rect 31665 7899 31723 7905
rect 32214 7896 32220 7908
rect 32272 7896 32278 7948
rect 32876 7936 32904 7976
rect 33410 7964 33416 7976
rect 33468 7964 33474 8016
rect 33520 8004 33548 8044
rect 33962 8032 33968 8084
rect 34020 8072 34026 8084
rect 37553 8075 37611 8081
rect 37553 8072 37565 8075
rect 34020 8044 37565 8072
rect 34020 8032 34026 8044
rect 37553 8041 37565 8044
rect 37599 8041 37611 8075
rect 37553 8035 37611 8041
rect 35250 8004 35256 8016
rect 33520 7976 35256 8004
rect 35250 7964 35256 7976
rect 35308 7964 35314 8016
rect 32416 7908 32904 7936
rect 32953 7939 33011 7945
rect 2464 7840 6914 7868
rect 2464 7828 2470 7840
rect 12802 7828 12808 7880
rect 12860 7868 12866 7880
rect 15749 7871 15807 7877
rect 15749 7868 15761 7871
rect 12860 7840 15761 7868
rect 12860 7828 12866 7840
rect 15749 7837 15761 7840
rect 15795 7837 15807 7871
rect 15749 7831 15807 7837
rect 17037 7871 17095 7877
rect 17037 7837 17049 7871
rect 17083 7868 17095 7871
rect 18414 7868 18420 7880
rect 17083 7840 18420 7868
rect 17083 7837 17095 7840
rect 17037 7831 17095 7837
rect 18414 7828 18420 7840
rect 18472 7828 18478 7880
rect 22370 7828 22376 7880
rect 22428 7828 22434 7880
rect 32416 7868 32444 7908
rect 32953 7905 32965 7939
rect 32999 7936 33011 7939
rect 34790 7936 34796 7948
rect 32999 7908 34796 7936
rect 32999 7905 33011 7908
rect 32953 7899 33011 7905
rect 34790 7896 34796 7908
rect 34848 7896 34854 7948
rect 37568 7868 37596 8035
rect 49145 7939 49203 7945
rect 49145 7905 49157 7939
rect 49191 7936 49203 7939
rect 49234 7936 49240 7948
rect 49191 7908 49240 7936
rect 49191 7905 49203 7908
rect 49145 7899 49203 7905
rect 49234 7896 49240 7908
rect 49292 7896 49298 7948
rect 38013 7871 38071 7877
rect 38013 7868 38025 7871
rect 31726 7840 32444 7868
rect 32508 7840 35664 7868
rect 37568 7840 38025 7868
rect 14182 7800 14188 7812
rect 1780 7772 14188 7800
rect 1780 7741 1808 7772
rect 14182 7760 14188 7772
rect 14240 7760 14246 7812
rect 18233 7803 18291 7809
rect 18233 7800 18245 7803
rect 16684 7772 18245 7800
rect 16684 7741 16712 7772
rect 18233 7769 18245 7772
rect 18279 7769 18291 7803
rect 18233 7763 18291 7769
rect 18506 7760 18512 7812
rect 18564 7800 18570 7812
rect 18969 7803 19027 7809
rect 18969 7800 18981 7803
rect 18564 7772 18981 7800
rect 18564 7760 18570 7772
rect 18969 7769 18981 7772
rect 19015 7769 19027 7803
rect 18969 7763 19027 7769
rect 19705 7803 19763 7809
rect 19705 7769 19717 7803
rect 19751 7800 19763 7803
rect 19978 7800 19984 7812
rect 19751 7772 19984 7800
rect 19751 7769 19763 7772
rect 19705 7763 19763 7769
rect 19978 7760 19984 7772
rect 20036 7760 20042 7812
rect 21082 7800 21088 7812
rect 20930 7772 21088 7800
rect 21082 7760 21088 7772
rect 21140 7800 21146 7812
rect 30377 7803 30435 7809
rect 21140 7772 21496 7800
rect 21140 7760 21146 7772
rect 21468 7744 21496 7772
rect 30377 7769 30389 7803
rect 30423 7800 30435 7803
rect 31481 7803 31539 7809
rect 31481 7800 31493 7803
rect 30423 7772 31493 7800
rect 30423 7769 30435 7772
rect 30377 7763 30435 7769
rect 31481 7769 31493 7772
rect 31527 7800 31539 7803
rect 31726 7800 31754 7840
rect 31527 7772 31754 7800
rect 31527 7769 31539 7772
rect 31481 7763 31539 7769
rect 1765 7735 1823 7741
rect 1765 7701 1777 7735
rect 1811 7701 1823 7735
rect 1765 7695 1823 7701
rect 16669 7735 16727 7741
rect 16669 7701 16681 7735
rect 16715 7701 16727 7735
rect 16669 7695 16727 7701
rect 18325 7735 18383 7741
rect 18325 7701 18337 7735
rect 18371 7732 18383 7735
rect 18782 7732 18788 7744
rect 18371 7704 18788 7732
rect 18371 7701 18383 7704
rect 18325 7695 18383 7701
rect 18782 7692 18788 7704
rect 18840 7692 18846 7744
rect 21450 7692 21456 7744
rect 21508 7732 21514 7744
rect 21637 7735 21695 7741
rect 21637 7732 21649 7735
rect 21508 7704 21649 7732
rect 21508 7692 21514 7704
rect 21637 7701 21649 7704
rect 21683 7701 21695 7735
rect 21637 7695 21695 7701
rect 22278 7692 22284 7744
rect 22336 7732 22342 7744
rect 22465 7735 22523 7741
rect 22465 7732 22477 7735
rect 22336 7704 22477 7732
rect 22336 7692 22342 7704
rect 22465 7701 22477 7704
rect 22511 7732 22523 7735
rect 23017 7735 23075 7741
rect 23017 7732 23029 7735
rect 22511 7704 23029 7732
rect 22511 7701 22523 7704
rect 22465 7695 22523 7701
rect 23017 7701 23029 7704
rect 23063 7732 23075 7735
rect 25682 7732 25688 7744
rect 23063 7704 25688 7732
rect 23063 7701 23075 7704
rect 23017 7695 23075 7701
rect 25682 7692 25688 7704
rect 25740 7692 25746 7744
rect 30650 7692 30656 7744
rect 30708 7692 30714 7744
rect 31386 7692 31392 7744
rect 31444 7692 31450 7744
rect 32309 7735 32367 7741
rect 32309 7701 32321 7735
rect 32355 7732 32367 7735
rect 32508 7732 32536 7840
rect 32677 7803 32735 7809
rect 32677 7769 32689 7803
rect 32723 7800 32735 7803
rect 32858 7800 32864 7812
rect 32723 7772 32864 7800
rect 32723 7769 32735 7772
rect 32677 7763 32735 7769
rect 32858 7760 32864 7772
rect 32916 7760 32922 7812
rect 35636 7800 35664 7840
rect 38013 7837 38025 7840
rect 38059 7837 38071 7871
rect 39022 7868 39028 7880
rect 38013 7831 38071 7837
rect 38120 7840 39028 7868
rect 38120 7800 38148 7840
rect 39022 7828 39028 7840
rect 39080 7828 39086 7880
rect 46934 7828 46940 7880
rect 46992 7868 46998 7880
rect 47949 7871 48007 7877
rect 47949 7868 47961 7871
rect 46992 7840 47961 7868
rect 46992 7828 46998 7840
rect 47949 7837 47961 7840
rect 47995 7837 48007 7871
rect 47949 7831 48007 7837
rect 35636 7772 38148 7800
rect 38746 7760 38752 7812
rect 38804 7760 38810 7812
rect 38933 7803 38991 7809
rect 38933 7769 38945 7803
rect 38979 7800 38991 7803
rect 40034 7800 40040 7812
rect 38979 7772 40040 7800
rect 38979 7769 38991 7772
rect 38933 7763 38991 7769
rect 40034 7760 40040 7772
rect 40092 7760 40098 7812
rect 32355 7704 32536 7732
rect 32355 7701 32367 7704
rect 32309 7695 32367 7701
rect 32766 7692 32772 7744
rect 32824 7692 32830 7744
rect 38105 7735 38163 7741
rect 38105 7701 38117 7735
rect 38151 7732 38163 7735
rect 38654 7732 38660 7744
rect 38151 7704 38660 7732
rect 38151 7701 38163 7704
rect 38105 7695 38163 7701
rect 38654 7692 38660 7704
rect 38712 7692 38718 7744
rect 38764 7732 38792 7760
rect 39209 7735 39267 7741
rect 39209 7732 39221 7735
rect 38764 7704 39221 7732
rect 39209 7701 39221 7704
rect 39255 7701 39267 7735
rect 39209 7695 39267 7701
rect 1104 7642 49864 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 27950 7642
rect 28002 7590 28014 7642
rect 28066 7590 28078 7642
rect 28130 7590 28142 7642
rect 28194 7590 28206 7642
rect 28258 7590 37950 7642
rect 38002 7590 38014 7642
rect 38066 7590 38078 7642
rect 38130 7590 38142 7642
rect 38194 7590 38206 7642
rect 38258 7590 47950 7642
rect 48002 7590 48014 7642
rect 48066 7590 48078 7642
rect 48130 7590 48142 7642
rect 48194 7590 48206 7642
rect 48258 7590 49864 7642
rect 1104 7568 49864 7590
rect 17402 7488 17408 7540
rect 17460 7528 17466 7540
rect 18233 7531 18291 7537
rect 18233 7528 18245 7531
rect 17460 7500 18245 7528
rect 17460 7488 17466 7500
rect 18233 7497 18245 7500
rect 18279 7528 18291 7531
rect 18693 7531 18751 7537
rect 18693 7528 18705 7531
rect 18279 7500 18705 7528
rect 18279 7497 18291 7500
rect 18233 7491 18291 7497
rect 18693 7497 18705 7500
rect 18739 7497 18751 7531
rect 18693 7491 18751 7497
rect 20530 7488 20536 7540
rect 20588 7528 20594 7540
rect 22005 7531 22063 7537
rect 22005 7528 22017 7531
rect 20588 7500 22017 7528
rect 20588 7488 20594 7500
rect 22005 7497 22017 7500
rect 22051 7497 22063 7531
rect 22005 7491 22063 7497
rect 22462 7488 22468 7540
rect 22520 7528 22526 7540
rect 23017 7531 23075 7537
rect 23017 7528 23029 7531
rect 22520 7500 23029 7528
rect 22520 7488 22526 7500
rect 23017 7497 23029 7500
rect 23063 7497 23075 7531
rect 23017 7491 23075 7497
rect 28534 7488 28540 7540
rect 28592 7528 28598 7540
rect 28592 7500 30696 7528
rect 28592 7488 28598 7500
rect 17310 7420 17316 7472
rect 17368 7460 17374 7472
rect 21361 7463 21419 7469
rect 21361 7460 21373 7463
rect 17368 7432 21373 7460
rect 17368 7420 17374 7432
rect 21361 7429 21373 7432
rect 21407 7460 21419 7463
rect 22373 7463 22431 7469
rect 22373 7460 22385 7463
rect 21407 7432 22385 7460
rect 21407 7429 21419 7432
rect 21361 7423 21419 7429
rect 22373 7429 22385 7432
rect 22419 7460 22431 7463
rect 30558 7460 30564 7472
rect 22419 7432 30564 7460
rect 22419 7429 22431 7432
rect 22373 7423 22431 7429
rect 30558 7420 30564 7432
rect 30616 7420 30622 7472
rect 30668 7460 30696 7500
rect 30926 7488 30932 7540
rect 30984 7488 30990 7540
rect 31386 7488 31392 7540
rect 31444 7528 31450 7540
rect 32309 7531 32367 7537
rect 32309 7528 32321 7531
rect 31444 7500 32321 7528
rect 31444 7488 31450 7500
rect 32309 7497 32321 7500
rect 32355 7497 32367 7531
rect 32309 7491 32367 7497
rect 38654 7488 38660 7540
rect 38712 7528 38718 7540
rect 46934 7528 46940 7540
rect 38712 7500 46940 7528
rect 38712 7488 38718 7500
rect 46934 7488 46940 7500
rect 46992 7488 46998 7540
rect 37369 7463 37427 7469
rect 37369 7460 37381 7463
rect 30668 7432 37381 7460
rect 37369 7429 37381 7432
rect 37415 7460 37427 7463
rect 37829 7463 37887 7469
rect 37829 7460 37841 7463
rect 37415 7432 37841 7460
rect 37415 7429 37427 7432
rect 37369 7423 37427 7429
rect 37829 7429 37841 7432
rect 37875 7429 37887 7463
rect 37829 7423 37887 7429
rect 40126 7420 40132 7472
rect 40184 7460 40190 7472
rect 44913 7463 44971 7469
rect 44913 7460 44925 7463
rect 40184 7432 44925 7460
rect 40184 7420 40190 7432
rect 44913 7429 44925 7432
rect 44959 7429 44971 7463
rect 44913 7423 44971 7429
rect 49145 7463 49203 7469
rect 49145 7429 49157 7463
rect 49191 7460 49203 7463
rect 49326 7460 49332 7472
rect 49191 7432 49332 7460
rect 49191 7429 49203 7432
rect 49145 7423 49203 7429
rect 49326 7420 49332 7432
rect 49384 7420 49390 7472
rect 1302 7352 1308 7404
rect 1360 7392 1366 7404
rect 1581 7395 1639 7401
rect 1581 7392 1593 7395
rect 1360 7364 1593 7392
rect 1360 7352 1366 7364
rect 1581 7361 1593 7364
rect 1627 7392 1639 7395
rect 2133 7395 2191 7401
rect 2133 7392 2145 7395
rect 1627 7364 2145 7392
rect 1627 7361 1639 7364
rect 1581 7355 1639 7361
rect 2133 7361 2145 7364
rect 2179 7361 2191 7395
rect 2133 7355 2191 7361
rect 34330 7352 34336 7404
rect 34388 7392 34394 7404
rect 38565 7395 38623 7401
rect 38565 7392 38577 7395
rect 34388 7364 38577 7392
rect 34388 7352 34394 7364
rect 38565 7361 38577 7364
rect 38611 7392 38623 7395
rect 39025 7395 39083 7401
rect 39025 7392 39037 7395
rect 38611 7364 39037 7392
rect 38611 7361 38623 7364
rect 38565 7355 38623 7361
rect 39025 7361 39037 7364
rect 39071 7361 39083 7395
rect 39025 7355 39083 7361
rect 47026 7352 47032 7404
rect 47084 7392 47090 7404
rect 47949 7395 48007 7401
rect 47949 7392 47961 7395
rect 47084 7364 47961 7392
rect 47084 7352 47090 7364
rect 47949 7361 47961 7364
rect 47995 7361 48007 7395
rect 47949 7355 48007 7361
rect 22646 7284 22652 7336
rect 22704 7284 22710 7336
rect 1765 7259 1823 7265
rect 1765 7225 1777 7259
rect 1811 7256 1823 7259
rect 19150 7256 19156 7268
rect 1811 7228 19156 7256
rect 1811 7225 1823 7228
rect 1765 7219 1823 7225
rect 19150 7216 19156 7228
rect 19208 7216 19214 7268
rect 38749 7259 38807 7265
rect 38749 7225 38761 7259
rect 38795 7256 38807 7259
rect 45097 7259 45155 7265
rect 38795 7228 42104 7256
rect 38795 7225 38807 7228
rect 38749 7219 38807 7225
rect 21269 7191 21327 7197
rect 21269 7157 21281 7191
rect 21315 7188 21327 7191
rect 21450 7188 21456 7200
rect 21315 7160 21456 7188
rect 21315 7157 21327 7160
rect 21269 7151 21327 7157
rect 21450 7148 21456 7160
rect 21508 7188 21514 7200
rect 21637 7191 21695 7197
rect 21637 7188 21649 7191
rect 21508 7160 21649 7188
rect 21508 7148 21514 7160
rect 21637 7157 21649 7160
rect 21683 7188 21695 7191
rect 22462 7188 22468 7200
rect 21683 7160 22468 7188
rect 21683 7157 21695 7160
rect 21637 7151 21695 7157
rect 22462 7148 22468 7160
rect 22520 7148 22526 7200
rect 32766 7148 32772 7200
rect 32824 7188 32830 7200
rect 32861 7191 32919 7197
rect 32861 7188 32873 7191
rect 32824 7160 32873 7188
rect 32824 7148 32830 7160
rect 32861 7157 32873 7160
rect 32907 7188 32919 7191
rect 37366 7188 37372 7200
rect 32907 7160 37372 7188
rect 32907 7157 32919 7160
rect 32861 7151 32919 7157
rect 37366 7148 37372 7160
rect 37424 7148 37430 7200
rect 37918 7148 37924 7200
rect 37976 7148 37982 7200
rect 42076 7188 42104 7228
rect 45097 7225 45109 7259
rect 45143 7256 45155 7259
rect 47762 7256 47768 7268
rect 45143 7228 47768 7256
rect 45143 7225 45155 7228
rect 45097 7219 45155 7225
rect 47762 7216 47768 7228
rect 47820 7216 47826 7268
rect 45830 7188 45836 7200
rect 42076 7160 45836 7188
rect 45830 7148 45836 7160
rect 45888 7148 45894 7200
rect 1104 7098 49864 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 32950 7098
rect 33002 7046 33014 7098
rect 33066 7046 33078 7098
rect 33130 7046 33142 7098
rect 33194 7046 33206 7098
rect 33258 7046 42950 7098
rect 43002 7046 43014 7098
rect 43066 7046 43078 7098
rect 43130 7046 43142 7098
rect 43194 7046 43206 7098
rect 43258 7046 49864 7098
rect 1104 7024 49864 7046
rect 37918 6876 37924 6928
rect 37976 6916 37982 6928
rect 47026 6916 47032 6928
rect 37976 6888 47032 6916
rect 37976 6876 37982 6888
rect 47026 6876 47032 6888
rect 47084 6876 47090 6928
rect 33778 6808 33784 6860
rect 33836 6848 33842 6860
rect 40126 6848 40132 6860
rect 33836 6820 40132 6848
rect 33836 6808 33842 6820
rect 40126 6808 40132 6820
rect 40184 6808 40190 6860
rect 49142 6808 49148 6860
rect 49200 6808 49206 6860
rect 1302 6740 1308 6792
rect 1360 6780 1366 6792
rect 2501 6783 2559 6789
rect 2501 6780 2513 6783
rect 1360 6752 2513 6780
rect 1360 6740 1366 6752
rect 2501 6749 2513 6752
rect 2547 6780 2559 6783
rect 2777 6783 2835 6789
rect 2777 6780 2789 6783
rect 2547 6752 2789 6780
rect 2547 6749 2559 6752
rect 2501 6743 2559 6749
rect 2777 6749 2789 6752
rect 2823 6749 2835 6783
rect 2777 6743 2835 6749
rect 16574 6740 16580 6792
rect 16632 6780 16638 6792
rect 17865 6783 17923 6789
rect 17865 6780 17877 6783
rect 16632 6752 17877 6780
rect 16632 6740 16638 6752
rect 17865 6749 17877 6752
rect 17911 6749 17923 6783
rect 17865 6743 17923 6749
rect 19242 6740 19248 6792
rect 19300 6780 19306 6792
rect 19797 6783 19855 6789
rect 19797 6780 19809 6783
rect 19300 6752 19809 6780
rect 19300 6740 19306 6752
rect 19797 6749 19809 6752
rect 19843 6749 19855 6783
rect 19797 6743 19855 6749
rect 40034 6740 40040 6792
rect 40092 6780 40098 6792
rect 46109 6783 46167 6789
rect 46109 6780 46121 6783
rect 40092 6752 46121 6780
rect 40092 6740 40098 6752
rect 46109 6749 46121 6752
rect 46155 6749 46167 6783
rect 46109 6743 46167 6749
rect 47854 6740 47860 6792
rect 47912 6780 47918 6792
rect 47949 6783 48007 6789
rect 47949 6780 47961 6783
rect 47912 6752 47961 6780
rect 47912 6740 47918 6752
rect 47949 6749 47961 6752
rect 47995 6749 48007 6783
rect 47949 6743 48007 6749
rect 1210 6672 1216 6724
rect 1268 6712 1274 6724
rect 1673 6715 1731 6721
rect 1673 6712 1685 6715
rect 1268 6684 1685 6712
rect 1268 6672 1274 6684
rect 1673 6681 1685 6684
rect 1719 6681 1731 6715
rect 1673 6675 1731 6681
rect 1857 6715 1915 6721
rect 1857 6681 1869 6715
rect 1903 6712 1915 6715
rect 27798 6712 27804 6724
rect 1903 6684 27804 6712
rect 1903 6681 1915 6684
rect 1857 6675 1915 6681
rect 27798 6672 27804 6684
rect 27856 6672 27862 6724
rect 47305 6715 47363 6721
rect 47305 6681 47317 6715
rect 47351 6712 47363 6715
rect 48866 6712 48872 6724
rect 47351 6684 48872 6712
rect 47351 6681 47363 6684
rect 47305 6675 47363 6681
rect 48866 6672 48872 6684
rect 48924 6672 48930 6724
rect 2314 6604 2320 6656
rect 2372 6604 2378 6656
rect 17681 6647 17739 6653
rect 17681 6613 17693 6647
rect 17727 6644 17739 6647
rect 19150 6644 19156 6656
rect 17727 6616 19156 6644
rect 17727 6613 17739 6616
rect 17681 6607 17739 6613
rect 19150 6604 19156 6616
rect 19208 6604 19214 6656
rect 19613 6647 19671 6653
rect 19613 6613 19625 6647
rect 19659 6644 19671 6647
rect 21910 6644 21916 6656
rect 19659 6616 21916 6644
rect 19659 6613 19671 6616
rect 19613 6607 19671 6613
rect 21910 6604 21916 6616
rect 21968 6604 21974 6656
rect 1104 6554 49864 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 27950 6554
rect 28002 6502 28014 6554
rect 28066 6502 28078 6554
rect 28130 6502 28142 6554
rect 28194 6502 28206 6554
rect 28258 6502 37950 6554
rect 38002 6502 38014 6554
rect 38066 6502 38078 6554
rect 38130 6502 38142 6554
rect 38194 6502 38206 6554
rect 38258 6502 47950 6554
rect 48002 6502 48014 6554
rect 48066 6502 48078 6554
rect 48130 6502 48142 6554
rect 48194 6502 48206 6554
rect 48258 6502 49864 6554
rect 1104 6480 49864 6502
rect 1210 6400 1216 6452
rect 1268 6440 1274 6452
rect 2133 6443 2191 6449
rect 2133 6440 2145 6443
rect 1268 6412 2145 6440
rect 1268 6400 1274 6412
rect 2133 6409 2145 6412
rect 2179 6409 2191 6443
rect 2133 6403 2191 6409
rect 40218 6332 40224 6384
rect 40276 6372 40282 6384
rect 43993 6375 44051 6381
rect 43993 6372 44005 6375
rect 40276 6344 44005 6372
rect 40276 6332 40282 6344
rect 43993 6341 44005 6344
rect 44039 6341 44051 6375
rect 43993 6335 44051 6341
rect 49145 6375 49203 6381
rect 49145 6341 49157 6375
rect 49191 6372 49203 6375
rect 49234 6372 49240 6384
rect 49191 6344 49240 6372
rect 49191 6341 49203 6344
rect 49145 6335 49203 6341
rect 49234 6332 49240 6344
rect 49292 6332 49298 6384
rect 1302 6264 1308 6316
rect 1360 6304 1366 6316
rect 1581 6307 1639 6313
rect 1581 6304 1593 6307
rect 1360 6276 1593 6304
rect 1360 6264 1366 6276
rect 1581 6273 1593 6276
rect 1627 6304 1639 6307
rect 2317 6307 2375 6313
rect 2317 6304 2329 6307
rect 1627 6276 2329 6304
rect 1627 6273 1639 6276
rect 1581 6267 1639 6273
rect 2317 6273 2329 6276
rect 2363 6273 2375 6307
rect 2317 6267 2375 6273
rect 17862 6264 17868 6316
rect 17920 6304 17926 6316
rect 18049 6307 18107 6313
rect 18049 6304 18061 6307
rect 17920 6276 18061 6304
rect 17920 6264 17926 6276
rect 18049 6273 18061 6276
rect 18095 6273 18107 6307
rect 18049 6267 18107 6273
rect 37553 6307 37611 6313
rect 37553 6273 37565 6307
rect 37599 6273 37611 6307
rect 37553 6267 37611 6273
rect 18233 6239 18291 6245
rect 18233 6205 18245 6239
rect 18279 6236 18291 6239
rect 18322 6236 18328 6248
rect 18279 6208 18328 6236
rect 18279 6205 18291 6208
rect 18233 6199 18291 6205
rect 18322 6196 18328 6208
rect 18380 6196 18386 6248
rect 25682 6196 25688 6248
rect 25740 6236 25746 6248
rect 36446 6236 36452 6248
rect 25740 6208 36452 6236
rect 25740 6196 25746 6208
rect 36446 6196 36452 6208
rect 36504 6196 36510 6248
rect 1765 6171 1823 6177
rect 1765 6137 1777 6171
rect 1811 6168 1823 6171
rect 14090 6168 14096 6180
rect 1811 6140 14096 6168
rect 1811 6137 1823 6140
rect 1765 6131 1823 6137
rect 14090 6128 14096 6140
rect 14148 6128 14154 6180
rect 22554 6168 22560 6180
rect 17236 6140 22560 6168
rect 7834 6060 7840 6112
rect 7892 6100 7898 6112
rect 17236 6100 17264 6140
rect 22554 6128 22560 6140
rect 22612 6128 22618 6180
rect 28350 6128 28356 6180
rect 28408 6168 28414 6180
rect 37274 6168 37280 6180
rect 28408 6140 37280 6168
rect 28408 6128 28414 6140
rect 37274 6128 37280 6140
rect 37332 6128 37338 6180
rect 37568 6168 37596 6267
rect 47486 6264 47492 6316
rect 47544 6304 47550 6316
rect 47949 6307 48007 6313
rect 47949 6304 47961 6307
rect 47544 6276 47961 6304
rect 47544 6264 47550 6276
rect 47949 6273 47961 6276
rect 47995 6273 48007 6307
rect 47949 6267 48007 6273
rect 38013 6171 38071 6177
rect 38013 6168 38025 6171
rect 37568 6140 38025 6168
rect 7892 6072 17264 6100
rect 18693 6103 18751 6109
rect 7892 6060 7898 6072
rect 18693 6069 18705 6103
rect 18739 6100 18751 6103
rect 19610 6100 19616 6112
rect 18739 6072 19616 6100
rect 18739 6069 18751 6072
rect 18693 6063 18751 6069
rect 19610 6060 19616 6072
rect 19668 6060 19674 6112
rect 30742 6060 30748 6112
rect 30800 6100 30806 6112
rect 37568 6100 37596 6140
rect 38013 6137 38025 6140
rect 38059 6137 38071 6171
rect 38013 6131 38071 6137
rect 44177 6171 44235 6177
rect 44177 6137 44189 6171
rect 44223 6168 44235 6171
rect 47118 6168 47124 6180
rect 44223 6140 47124 6168
rect 44223 6137 44235 6140
rect 44177 6131 44235 6137
rect 47118 6128 47124 6140
rect 47176 6128 47182 6180
rect 30800 6072 37596 6100
rect 30800 6060 30806 6072
rect 37642 6060 37648 6112
rect 37700 6060 37706 6112
rect 1104 6010 49864 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 32950 6010
rect 33002 5958 33014 6010
rect 33066 5958 33078 6010
rect 33130 5958 33142 6010
rect 33194 5958 33206 6010
rect 33258 5958 42950 6010
rect 43002 5958 43014 6010
rect 43066 5958 43078 6010
rect 43130 5958 43142 6010
rect 43194 5958 43206 6010
rect 43258 5958 49864 6010
rect 1104 5936 49864 5958
rect 2501 5899 2559 5905
rect 2501 5865 2513 5899
rect 2547 5896 2559 5899
rect 6914 5896 6920 5908
rect 2547 5868 6920 5896
rect 2547 5865 2559 5868
rect 2501 5859 2559 5865
rect 6914 5856 6920 5868
rect 6972 5856 6978 5908
rect 37642 5856 37648 5908
rect 37700 5896 37706 5908
rect 47302 5896 47308 5908
rect 37700 5868 47308 5896
rect 37700 5856 37706 5868
rect 47302 5856 47308 5868
rect 47360 5856 47366 5908
rect 27430 5788 27436 5840
rect 27488 5828 27494 5840
rect 35802 5828 35808 5840
rect 27488 5800 35808 5828
rect 27488 5788 27494 5800
rect 35802 5788 35808 5800
rect 35860 5788 35866 5840
rect 3053 5763 3111 5769
rect 3053 5760 3065 5763
rect 1596 5732 3065 5760
rect 1302 5652 1308 5704
rect 1360 5692 1366 5704
rect 1596 5701 1624 5732
rect 3053 5729 3065 5732
rect 3099 5729 3111 5763
rect 3053 5723 3111 5729
rect 49145 5763 49203 5769
rect 49145 5729 49157 5763
rect 49191 5760 49203 5763
rect 49418 5760 49424 5772
rect 49191 5732 49424 5760
rect 49191 5729 49203 5732
rect 49145 5723 49203 5729
rect 49418 5720 49424 5732
rect 49476 5720 49482 5772
rect 1581 5695 1639 5701
rect 1581 5692 1593 5695
rect 1360 5664 1593 5692
rect 1360 5652 1366 5664
rect 1581 5661 1593 5664
rect 1627 5661 1639 5695
rect 1581 5655 1639 5661
rect 2317 5695 2375 5701
rect 2317 5661 2329 5695
rect 2363 5692 2375 5695
rect 2774 5692 2780 5704
rect 2363 5664 2780 5692
rect 2363 5661 2375 5664
rect 2317 5655 2375 5661
rect 2774 5652 2780 5664
rect 2832 5692 2838 5704
rect 2869 5695 2927 5701
rect 2869 5692 2881 5695
rect 2832 5664 2881 5692
rect 2832 5652 2838 5664
rect 2869 5661 2881 5664
rect 2915 5661 2927 5695
rect 2869 5655 2927 5661
rect 19334 5652 19340 5704
rect 19392 5692 19398 5704
rect 23934 5692 23940 5704
rect 19392 5664 23940 5692
rect 19392 5652 19398 5664
rect 23934 5652 23940 5664
rect 23992 5652 23998 5704
rect 27338 5652 27344 5704
rect 27396 5692 27402 5704
rect 32766 5692 32772 5704
rect 27396 5664 32772 5692
rect 27396 5652 27402 5664
rect 32766 5652 32772 5664
rect 32824 5652 32830 5704
rect 43714 5652 43720 5704
rect 43772 5652 43778 5704
rect 47670 5652 47676 5704
rect 47728 5692 47734 5704
rect 47949 5695 48007 5701
rect 47949 5692 47961 5695
rect 47728 5664 47961 5692
rect 47728 5652 47734 5664
rect 47949 5661 47961 5664
rect 47995 5661 48007 5695
rect 47949 5655 48007 5661
rect 43901 5627 43959 5633
rect 1780 5596 6914 5624
rect 1780 5565 1808 5596
rect 1765 5559 1823 5565
rect 1765 5525 1777 5559
rect 1811 5525 1823 5559
rect 6886 5556 6914 5596
rect 43901 5593 43913 5627
rect 43947 5624 43959 5627
rect 45738 5624 45744 5636
rect 43947 5596 45744 5624
rect 43947 5593 43959 5596
rect 43901 5587 43959 5593
rect 45738 5584 45744 5596
rect 45796 5584 45802 5636
rect 17678 5556 17684 5568
rect 6886 5528 17684 5556
rect 1765 5519 1823 5525
rect 17678 5516 17684 5528
rect 17736 5516 17742 5568
rect 1104 5466 49864 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 27950 5466
rect 28002 5414 28014 5466
rect 28066 5414 28078 5466
rect 28130 5414 28142 5466
rect 28194 5414 28206 5466
rect 28258 5414 37950 5466
rect 38002 5414 38014 5466
rect 38066 5414 38078 5466
rect 38130 5414 38142 5466
rect 38194 5414 38206 5466
rect 38258 5414 47950 5466
rect 48002 5414 48014 5466
rect 48066 5414 48078 5466
rect 48130 5414 48142 5466
rect 48194 5414 48206 5466
rect 48258 5414 49864 5466
rect 1104 5392 49864 5414
rect 31478 5244 31484 5296
rect 31536 5284 31542 5296
rect 38473 5287 38531 5293
rect 38473 5284 38485 5287
rect 31536 5256 38485 5284
rect 31536 5244 31542 5256
rect 38473 5253 38485 5256
rect 38519 5284 38531 5287
rect 38933 5287 38991 5293
rect 38933 5284 38945 5287
rect 38519 5256 38945 5284
rect 38519 5253 38531 5256
rect 38473 5247 38531 5253
rect 38933 5253 38945 5256
rect 38979 5253 38991 5287
rect 38933 5247 38991 5253
rect 49142 5244 49148 5296
rect 49200 5244 49206 5296
rect 18874 5176 18880 5228
rect 18932 5176 18938 5228
rect 37366 5176 37372 5228
rect 37424 5216 37430 5228
rect 37737 5219 37795 5225
rect 37737 5216 37749 5219
rect 37424 5188 37749 5216
rect 37424 5176 37430 5188
rect 37737 5185 37749 5188
rect 37783 5185 37795 5219
rect 37737 5179 37795 5185
rect 45830 5176 45836 5228
rect 45888 5176 45894 5228
rect 47762 5176 47768 5228
rect 47820 5216 47826 5228
rect 47949 5219 48007 5225
rect 47949 5216 47961 5219
rect 47820 5188 47961 5216
rect 47820 5176 47826 5188
rect 47949 5185 47961 5188
rect 47995 5185 48007 5219
rect 47949 5179 48007 5185
rect 1302 5108 1308 5160
rect 1360 5148 1366 5160
rect 1581 5151 1639 5157
rect 1581 5148 1593 5151
rect 1360 5120 1593 5148
rect 1360 5108 1366 5120
rect 1581 5117 1593 5120
rect 1627 5117 1639 5151
rect 1581 5111 1639 5117
rect 1857 5151 1915 5157
rect 1857 5117 1869 5151
rect 1903 5148 1915 5151
rect 11790 5148 11796 5160
rect 1903 5120 11796 5148
rect 1903 5117 1915 5120
rect 1857 5111 1915 5117
rect 11790 5108 11796 5120
rect 11848 5108 11854 5160
rect 19058 5108 19064 5160
rect 19116 5108 19122 5160
rect 46845 5151 46903 5157
rect 46845 5117 46857 5151
rect 46891 5148 46903 5151
rect 48314 5148 48320 5160
rect 46891 5120 48320 5148
rect 46891 5117 46903 5120
rect 46845 5111 46903 5117
rect 48314 5108 48320 5120
rect 48372 5108 48378 5160
rect 38657 5083 38715 5089
rect 38657 5049 38669 5083
rect 38703 5080 38715 5083
rect 40402 5080 40408 5092
rect 38703 5052 40408 5080
rect 38703 5049 38715 5052
rect 38657 5043 38715 5049
rect 40402 5040 40408 5052
rect 40460 5040 40466 5092
rect 1854 4972 1860 5024
rect 1912 5012 1918 5024
rect 12434 5012 12440 5024
rect 1912 4984 12440 5012
rect 1912 4972 1918 4984
rect 12434 4972 12440 4984
rect 12492 4972 12498 5024
rect 19521 5015 19579 5021
rect 19521 4981 19533 5015
rect 19567 5012 19579 5015
rect 20806 5012 20812 5024
rect 19567 4984 20812 5012
rect 19567 4981 19579 4984
rect 19521 4975 19579 4981
rect 20806 4972 20812 4984
rect 20864 4972 20870 5024
rect 37826 4972 37832 5024
rect 37884 4972 37890 5024
rect 1104 4922 49864 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 32950 4922
rect 33002 4870 33014 4922
rect 33066 4870 33078 4922
rect 33130 4870 33142 4922
rect 33194 4870 33206 4922
rect 33258 4870 42950 4922
rect 43002 4870 43014 4922
rect 43066 4870 43078 4922
rect 43130 4870 43142 4922
rect 43194 4870 43206 4922
rect 43258 4870 49864 4922
rect 1104 4848 49864 4870
rect 1302 4768 1308 4820
rect 1360 4808 1366 4820
rect 2133 4811 2191 4817
rect 2133 4808 2145 4811
rect 1360 4780 2145 4808
rect 1360 4768 1366 4780
rect 2133 4777 2145 4780
rect 2179 4777 2191 4811
rect 2133 4771 2191 4777
rect 35802 4768 35808 4820
rect 35860 4808 35866 4820
rect 36817 4811 36875 4817
rect 36817 4808 36829 4811
rect 35860 4780 36829 4808
rect 35860 4768 35866 4780
rect 36817 4777 36829 4780
rect 36863 4777 36875 4811
rect 36817 4771 36875 4777
rect 11698 4700 11704 4752
rect 11756 4740 11762 4752
rect 20990 4740 20996 4752
rect 11756 4712 20996 4740
rect 11756 4700 11762 4712
rect 20990 4700 20996 4712
rect 21048 4740 21054 4752
rect 21048 4712 25636 4740
rect 21048 4700 21054 4712
rect 19150 4632 19156 4684
rect 19208 4672 19214 4684
rect 20441 4675 20499 4681
rect 20441 4672 20453 4675
rect 19208 4644 20453 4672
rect 19208 4632 19214 4644
rect 20441 4641 20453 4644
rect 20487 4641 20499 4675
rect 20441 4635 20499 4641
rect 21910 4632 21916 4684
rect 21968 4632 21974 4684
rect 22922 4672 22928 4684
rect 22020 4644 22928 4672
rect 1302 4564 1308 4616
rect 1360 4604 1366 4616
rect 1581 4607 1639 4613
rect 1581 4604 1593 4607
rect 1360 4576 1593 4604
rect 1360 4564 1366 4576
rect 1581 4573 1593 4576
rect 1627 4604 1639 4607
rect 2317 4607 2375 4613
rect 2317 4604 2329 4607
rect 1627 4576 2329 4604
rect 1627 4573 1639 4576
rect 1581 4567 1639 4573
rect 2317 4573 2329 4576
rect 2363 4573 2375 4607
rect 2317 4567 2375 4573
rect 19518 4564 19524 4616
rect 19576 4604 19582 4616
rect 20625 4607 20683 4613
rect 20625 4604 20637 4607
rect 19576 4576 20637 4604
rect 19576 4564 19582 4576
rect 20625 4573 20637 4576
rect 20671 4604 20683 4607
rect 22020 4604 22048 4644
rect 22922 4632 22928 4644
rect 22980 4632 22986 4684
rect 23198 4632 23204 4684
rect 23256 4672 23262 4684
rect 25608 4681 25636 4712
rect 25317 4675 25375 4681
rect 25317 4672 25329 4675
rect 23256 4644 25329 4672
rect 23256 4632 23262 4644
rect 25317 4641 25329 4644
rect 25363 4641 25375 4675
rect 25317 4635 25375 4641
rect 25593 4675 25651 4681
rect 25593 4641 25605 4675
rect 25639 4641 25651 4675
rect 25593 4635 25651 4641
rect 20671 4576 22048 4604
rect 20671 4573 20683 4576
rect 20625 4567 20683 4573
rect 22094 4564 22100 4616
rect 22152 4564 22158 4616
rect 23084 4607 23142 4613
rect 23084 4604 23096 4607
rect 22480 4576 23096 4604
rect 1780 4508 6914 4536
rect 1780 4477 1808 4508
rect 1765 4471 1823 4477
rect 1765 4437 1777 4471
rect 1811 4437 1823 4471
rect 6886 4468 6914 4508
rect 19058 4496 19064 4548
rect 19116 4536 19122 4548
rect 22480 4536 22508 4576
rect 23084 4573 23096 4576
rect 23130 4604 23142 4607
rect 24026 4604 24032 4616
rect 23130 4576 24032 4604
rect 23130 4573 23142 4576
rect 23084 4567 23142 4573
rect 24026 4564 24032 4576
rect 24084 4564 24090 4616
rect 25133 4607 25191 4613
rect 25133 4573 25145 4607
rect 25179 4573 25191 4607
rect 36832 4604 36860 4771
rect 40126 4768 40132 4820
rect 40184 4808 40190 4820
rect 46661 4811 46719 4817
rect 46661 4808 46673 4811
rect 40184 4780 46673 4808
rect 40184 4768 40190 4780
rect 46661 4777 46673 4780
rect 46707 4777 46719 4811
rect 46661 4771 46719 4777
rect 37826 4700 37832 4752
rect 37884 4740 37890 4752
rect 47210 4740 47216 4752
rect 37884 4712 47216 4740
rect 37884 4700 37890 4712
rect 47210 4700 47216 4712
rect 47268 4700 47274 4752
rect 36998 4632 37004 4684
rect 37056 4672 37062 4684
rect 47489 4675 47547 4681
rect 47489 4672 47501 4675
rect 37056 4644 47501 4672
rect 37056 4632 37062 4644
rect 47489 4641 47501 4644
rect 47535 4641 47547 4675
rect 47489 4635 47547 4641
rect 49145 4675 49203 4681
rect 49145 4641 49157 4675
rect 49191 4672 49203 4675
rect 49418 4672 49424 4684
rect 49191 4644 49424 4672
rect 49191 4641 49203 4644
rect 49145 4635 49203 4641
rect 49418 4632 49424 4644
rect 49476 4632 49482 4684
rect 37277 4607 37335 4613
rect 37277 4604 37289 4607
rect 36832 4576 37289 4604
rect 25133 4567 25191 4573
rect 37277 4573 37289 4576
rect 37323 4573 37335 4607
rect 38473 4607 38531 4613
rect 38473 4604 38485 4607
rect 37277 4567 37335 4573
rect 38028 4576 38485 4604
rect 19116 4508 22508 4536
rect 22557 4539 22615 4545
rect 19116 4496 19122 4508
rect 22557 4505 22569 4539
rect 22603 4536 22615 4539
rect 24578 4536 24584 4548
rect 22603 4508 24584 4536
rect 22603 4505 22615 4508
rect 22557 4499 22615 4505
rect 24578 4496 24584 4508
rect 24636 4496 24642 4548
rect 19334 4468 19340 4480
rect 6886 4440 19340 4468
rect 1765 4431 1823 4437
rect 19334 4428 19340 4440
rect 19392 4428 19398 4480
rect 21085 4471 21143 4477
rect 21085 4437 21097 4471
rect 21131 4468 21143 4471
rect 21450 4468 21456 4480
rect 21131 4440 21456 4468
rect 21131 4437 21143 4440
rect 21085 4431 21143 4437
rect 21450 4428 21456 4440
rect 21508 4428 21514 4480
rect 23155 4471 23213 4477
rect 23155 4437 23167 4471
rect 23201 4468 23213 4471
rect 24394 4468 24400 4480
rect 23201 4440 24400 4468
rect 23201 4437 23213 4440
rect 23155 4431 23213 4437
rect 24394 4428 24400 4440
rect 24452 4428 24458 4480
rect 25148 4468 25176 4567
rect 32766 4496 32772 4548
rect 32824 4536 32830 4548
rect 38028 4545 38056 4576
rect 38473 4573 38485 4576
rect 38519 4573 38531 4607
rect 38473 4567 38531 4573
rect 46934 4564 46940 4616
rect 46992 4604 46998 4616
rect 47949 4607 48007 4613
rect 47949 4604 47961 4607
rect 46992 4576 47961 4604
rect 46992 4564 46998 4576
rect 47949 4573 47961 4576
rect 47995 4573 48007 4607
rect 47949 4567 48007 4573
rect 38013 4539 38071 4545
rect 38013 4536 38025 4539
rect 32824 4508 38025 4536
rect 32824 4496 32830 4508
rect 38013 4505 38025 4508
rect 38059 4505 38071 4539
rect 38013 4499 38071 4505
rect 38197 4539 38255 4545
rect 38197 4505 38209 4539
rect 38243 4536 38255 4539
rect 39758 4536 39764 4548
rect 38243 4508 39764 4536
rect 38243 4505 38255 4508
rect 38197 4499 38255 4505
rect 39758 4496 39764 4508
rect 39816 4496 39822 4548
rect 46569 4539 46627 4545
rect 46569 4505 46581 4539
rect 46615 4505 46627 4539
rect 46569 4499 46627 4505
rect 47305 4539 47363 4545
rect 47305 4505 47317 4539
rect 47351 4536 47363 4539
rect 47670 4536 47676 4548
rect 47351 4508 47676 4536
rect 47351 4505 47363 4508
rect 47305 4499 47363 4505
rect 32858 4468 32864 4480
rect 25148 4440 32864 4468
rect 32858 4428 32864 4440
rect 32916 4428 32922 4480
rect 37366 4428 37372 4480
rect 37424 4428 37430 4480
rect 46201 4471 46259 4477
rect 46201 4437 46213 4471
rect 46247 4468 46259 4471
rect 46584 4468 46612 4499
rect 47670 4496 47676 4508
rect 47728 4496 47734 4548
rect 49786 4468 49792 4480
rect 46247 4440 49792 4468
rect 46247 4437 46259 4440
rect 46201 4431 46259 4437
rect 49786 4428 49792 4440
rect 49844 4428 49850 4480
rect 1104 4378 49864 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 27950 4378
rect 28002 4326 28014 4378
rect 28066 4326 28078 4378
rect 28130 4326 28142 4378
rect 28194 4326 28206 4378
rect 28258 4326 37950 4378
rect 38002 4326 38014 4378
rect 38066 4326 38078 4378
rect 38130 4326 38142 4378
rect 38194 4326 38206 4378
rect 38258 4326 47950 4378
rect 48002 4326 48014 4378
rect 48066 4326 48078 4378
rect 48130 4326 48142 4378
rect 48194 4326 48206 4378
rect 48258 4326 49864 4378
rect 1104 4304 49864 4326
rect 37366 4224 37372 4276
rect 37424 4264 37430 4276
rect 45646 4264 45652 4276
rect 37424 4236 45652 4264
rect 37424 4224 37430 4236
rect 45646 4224 45652 4236
rect 45704 4224 45710 4276
rect 1394 4156 1400 4208
rect 1452 4196 1458 4208
rect 1673 4199 1731 4205
rect 1673 4196 1685 4199
rect 1452 4168 1685 4196
rect 1452 4156 1458 4168
rect 1673 4165 1685 4168
rect 1719 4196 1731 4199
rect 1719 4168 2728 4196
rect 1719 4165 1731 4168
rect 1673 4159 1731 4165
rect 1302 4088 1308 4140
rect 1360 4128 1366 4140
rect 2317 4131 2375 4137
rect 2317 4128 2329 4131
rect 1360 4100 2329 4128
rect 1360 4088 1366 4100
rect 2317 4097 2329 4100
rect 2363 4128 2375 4131
rect 2498 4128 2504 4140
rect 2363 4100 2504 4128
rect 2363 4097 2375 4100
rect 2317 4091 2375 4097
rect 2498 4088 2504 4100
rect 2556 4088 2562 4140
rect 2700 4128 2728 4168
rect 22094 4156 22100 4208
rect 22152 4196 22158 4208
rect 27341 4199 27399 4205
rect 27341 4196 27353 4199
rect 22152 4168 23336 4196
rect 22152 4156 22158 4168
rect 3053 4131 3111 4137
rect 3053 4128 3065 4131
rect 2700 4100 3065 4128
rect 3053 4097 3065 4100
rect 3099 4097 3111 4131
rect 3053 4091 3111 4097
rect 22348 4130 22406 4136
rect 22348 4096 22360 4130
rect 22394 4127 22406 4130
rect 22394 4099 22462 4127
rect 22394 4096 22406 4099
rect 22348 4090 22406 4096
rect 14918 4060 14924 4072
rect 2516 4032 14924 4060
rect 2516 4001 2544 4032
rect 14918 4020 14924 4032
rect 14976 4020 14982 4072
rect 2501 3995 2559 4001
rect 2501 3961 2513 3995
rect 2547 3961 2559 3995
rect 2501 3955 2559 3961
rect 2608 3964 4384 3992
rect 1765 3927 1823 3933
rect 1765 3893 1777 3927
rect 1811 3924 1823 3927
rect 2608 3924 2636 3964
rect 1811 3896 2636 3924
rect 1811 3893 1823 3896
rect 1765 3887 1823 3893
rect 2682 3884 2688 3936
rect 2740 3924 2746 3936
rect 2869 3927 2927 3933
rect 2869 3924 2881 3927
rect 2740 3896 2881 3924
rect 2740 3884 2746 3896
rect 2869 3893 2881 3896
rect 2915 3893 2927 3927
rect 4356 3924 4384 3964
rect 17954 3952 17960 4004
rect 18012 3992 18018 4004
rect 18322 3992 18328 4004
rect 18012 3964 18328 3992
rect 18012 3952 18018 3964
rect 18322 3952 18328 3964
rect 18380 3992 18386 4004
rect 22434 3992 22462 4099
rect 22922 4088 22928 4140
rect 22980 4137 22986 4140
rect 22980 4131 23018 4137
rect 23006 4097 23018 4131
rect 22980 4091 23018 4097
rect 23063 4131 23121 4137
rect 23063 4097 23075 4131
rect 23109 4128 23121 4131
rect 23198 4128 23204 4140
rect 23109 4100 23204 4128
rect 23109 4097 23121 4100
rect 23063 4091 23121 4097
rect 22980 4088 23003 4091
rect 23198 4088 23204 4100
rect 23256 4088 23262 4140
rect 23308 4128 23336 4168
rect 27172 4168 27353 4196
rect 23604 4131 23662 4137
rect 23604 4128 23616 4131
rect 23308 4100 23616 4128
rect 23604 4097 23616 4100
rect 23650 4097 23662 4131
rect 27172 4128 27200 4168
rect 27341 4165 27353 4168
rect 27387 4165 27399 4199
rect 27341 4159 27399 4165
rect 23604 4091 23662 4097
rect 27080 4100 27200 4128
rect 22975 4060 23003 4088
rect 23474 4060 23480 4072
rect 22975 4032 23480 4060
rect 23474 4020 23480 4032
rect 23532 4020 23538 4072
rect 24210 4020 24216 4072
rect 24268 4020 24274 4072
rect 24394 4020 24400 4072
rect 24452 4020 24458 4072
rect 25406 4020 25412 4072
rect 25464 4020 25470 4072
rect 23707 3995 23765 4001
rect 18380 3964 22968 3992
rect 18380 3952 18386 3964
rect 7834 3924 7840 3936
rect 4356 3896 7840 3924
rect 2869 3887 2927 3893
rect 7834 3884 7840 3896
rect 7892 3884 7898 3936
rect 22419 3927 22477 3933
rect 22419 3893 22431 3927
rect 22465 3924 22477 3927
rect 22830 3924 22836 3936
rect 22465 3896 22836 3924
rect 22465 3893 22477 3896
rect 22419 3887 22477 3893
rect 22830 3884 22836 3896
rect 22888 3884 22894 3936
rect 22940 3924 22968 3964
rect 23707 3961 23719 3995
rect 23753 3992 23765 3995
rect 27080 3992 27108 4100
rect 37274 4088 37280 4140
rect 37332 4128 37338 4140
rect 39206 4128 39212 4140
rect 37332 4100 39212 4128
rect 37332 4088 37338 4100
rect 39206 4088 39212 4100
rect 39264 4088 39270 4140
rect 45830 4088 45836 4140
rect 45888 4088 45894 4140
rect 47026 4088 47032 4140
rect 47084 4128 47090 4140
rect 47949 4131 48007 4137
rect 47949 4128 47961 4131
rect 47084 4100 47961 4128
rect 47084 4088 47090 4100
rect 47949 4097 47961 4100
rect 47995 4097 48007 4131
rect 47949 4091 48007 4097
rect 49145 4131 49203 4137
rect 49145 4097 49157 4131
rect 49191 4128 49203 4131
rect 49326 4128 49332 4140
rect 49191 4100 49332 4128
rect 49191 4097 49203 4100
rect 49145 4091 49203 4097
rect 49326 4088 49332 4100
rect 49384 4088 49390 4140
rect 27157 4063 27215 4069
rect 27157 4029 27169 4063
rect 27203 4060 27215 4063
rect 27203 4032 27568 4060
rect 27203 4029 27215 4032
rect 27157 4023 27215 4029
rect 23753 3964 27108 3992
rect 27540 3992 27568 4032
rect 27614 4020 27620 4072
rect 27672 4020 27678 4072
rect 46658 4020 46664 4072
rect 46716 4020 46722 4072
rect 34422 3992 34428 4004
rect 27540 3964 34428 3992
rect 23753 3961 23765 3964
rect 23707 3955 23765 3961
rect 34422 3952 34428 3964
rect 34480 3952 34486 4004
rect 27798 3924 27804 3936
rect 22940 3896 27804 3924
rect 27798 3884 27804 3896
rect 27856 3884 27862 3936
rect 47670 3884 47676 3936
rect 47728 3884 47734 3936
rect 1104 3834 49864 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 32950 3834
rect 33002 3782 33014 3834
rect 33066 3782 33078 3834
rect 33130 3782 33142 3834
rect 33194 3782 33206 3834
rect 33258 3782 42950 3834
rect 43002 3782 43014 3834
rect 43066 3782 43078 3834
rect 43130 3782 43142 3834
rect 43194 3782 43206 3834
rect 43258 3782 49864 3834
rect 1104 3760 49864 3782
rect 23845 3723 23903 3729
rect 23845 3689 23857 3723
rect 23891 3720 23903 3723
rect 25958 3720 25964 3732
rect 23891 3692 25964 3720
rect 23891 3689 23903 3692
rect 23845 3683 23903 3689
rect 25958 3680 25964 3692
rect 26016 3680 26022 3732
rect 26050 3680 26056 3732
rect 26108 3720 26114 3732
rect 27614 3720 27620 3732
rect 26108 3692 27620 3720
rect 26108 3680 26114 3692
rect 27614 3680 27620 3692
rect 27672 3680 27678 3732
rect 22554 3612 22560 3664
rect 22612 3652 22618 3664
rect 23017 3655 23075 3661
rect 23017 3652 23029 3655
rect 22612 3624 23029 3652
rect 22612 3612 22618 3624
rect 23017 3621 23029 3624
rect 23063 3621 23075 3655
rect 23017 3615 23075 3621
rect 24026 3612 24032 3664
rect 24084 3612 24090 3664
rect 24118 3612 24124 3664
rect 24176 3652 24182 3664
rect 24176 3624 25084 3652
rect 24176 3612 24182 3624
rect 1854 3544 1860 3596
rect 1912 3544 1918 3596
rect 7466 3544 7472 3596
rect 7524 3584 7530 3596
rect 7524 3556 22784 3584
rect 7524 3544 7530 3556
rect 1302 3476 1308 3528
rect 1360 3516 1366 3528
rect 1581 3519 1639 3525
rect 1581 3516 1593 3519
rect 1360 3488 1593 3516
rect 1360 3476 1366 3488
rect 1581 3485 1593 3488
rect 1627 3485 1639 3519
rect 1581 3479 1639 3485
rect 3326 3476 3332 3528
rect 3384 3516 3390 3528
rect 11698 3516 11704 3528
rect 3384 3488 11704 3516
rect 3384 3476 3390 3488
rect 11698 3476 11704 3488
rect 11756 3476 11762 3528
rect 16485 3519 16543 3525
rect 16485 3485 16497 3519
rect 16531 3516 16543 3519
rect 17954 3516 17960 3528
rect 16531 3488 17960 3516
rect 16531 3485 16543 3488
rect 16485 3479 16543 3485
rect 17954 3476 17960 3488
rect 18012 3476 18018 3528
rect 20990 3476 20996 3528
rect 21048 3476 21054 3528
rect 21174 3408 21180 3460
rect 21232 3448 21238 3460
rect 21269 3451 21327 3457
rect 21269 3448 21281 3451
rect 21232 3420 21281 3448
rect 21232 3408 21238 3420
rect 21269 3417 21281 3420
rect 21315 3417 21327 3451
rect 22554 3448 22560 3460
rect 22494 3420 22560 3448
rect 21269 3411 21327 3417
rect 22554 3408 22560 3420
rect 22612 3408 22618 3460
rect 22756 3448 22784 3556
rect 22830 3544 22836 3596
rect 22888 3584 22894 3596
rect 25056 3593 25084 3624
rect 40402 3612 40408 3664
rect 40460 3652 40466 3664
rect 40460 3624 46152 3652
rect 40460 3612 40466 3624
rect 24765 3587 24823 3593
rect 24765 3584 24777 3587
rect 22888 3556 24777 3584
rect 22888 3544 22894 3556
rect 24765 3553 24777 3556
rect 24811 3553 24823 3587
rect 24765 3547 24823 3553
rect 25041 3587 25099 3593
rect 25041 3553 25053 3587
rect 25087 3553 25099 3587
rect 25041 3547 25099 3553
rect 36633 3587 36691 3593
rect 36633 3553 36645 3587
rect 36679 3584 36691 3587
rect 45830 3584 45836 3596
rect 36679 3556 45836 3584
rect 36679 3553 36691 3556
rect 36633 3547 36691 3553
rect 45830 3544 45836 3556
rect 45888 3544 45894 3596
rect 23566 3476 23572 3528
rect 23624 3476 23630 3528
rect 24581 3519 24639 3525
rect 24581 3485 24593 3519
rect 24627 3485 24639 3519
rect 24581 3479 24639 3485
rect 24118 3448 24124 3460
rect 22756 3420 24124 3448
rect 24118 3408 24124 3420
rect 24176 3408 24182 3460
rect 12802 3340 12808 3392
rect 12860 3380 12866 3392
rect 16577 3383 16635 3389
rect 16577 3380 16589 3383
rect 12860 3352 16589 3380
rect 12860 3340 12866 3352
rect 16577 3349 16589 3352
rect 16623 3349 16635 3383
rect 16577 3343 16635 3349
rect 22741 3383 22799 3389
rect 22741 3349 22753 3383
rect 22787 3380 22799 3383
rect 23382 3380 23388 3392
rect 22787 3352 23388 3380
rect 22787 3349 22799 3352
rect 22741 3343 22799 3349
rect 23382 3340 23388 3352
rect 23440 3340 23446 3392
rect 24596 3380 24624 3479
rect 36446 3476 36452 3528
rect 36504 3516 36510 3528
rect 36909 3519 36967 3525
rect 36909 3516 36921 3519
rect 36504 3488 36921 3516
rect 36504 3476 36510 3488
rect 36909 3485 36921 3488
rect 36955 3485 36967 3519
rect 45554 3516 45560 3528
rect 36909 3479 36967 3485
rect 45480 3488 45560 3516
rect 45480 3457 45508 3488
rect 45554 3476 45560 3488
rect 45612 3476 45618 3528
rect 46124 3525 46152 3624
rect 49142 3544 49148 3596
rect 49200 3544 49206 3596
rect 46109 3519 46167 3525
rect 46109 3485 46121 3519
rect 46155 3485 46167 3519
rect 46109 3479 46167 3485
rect 47118 3476 47124 3528
rect 47176 3516 47182 3528
rect 47949 3519 48007 3525
rect 47949 3516 47961 3519
rect 47176 3488 47961 3516
rect 47176 3476 47182 3488
rect 47949 3485 47961 3488
rect 47995 3485 48007 3519
rect 47949 3479 48007 3485
rect 45097 3451 45155 3457
rect 45097 3417 45109 3451
rect 45143 3448 45155 3451
rect 45465 3451 45523 3457
rect 45465 3448 45477 3451
rect 45143 3420 45477 3448
rect 45143 3417 45155 3420
rect 45097 3411 45155 3417
rect 45465 3417 45477 3420
rect 45511 3417 45523 3451
rect 45465 3411 45523 3417
rect 47305 3451 47363 3457
rect 47305 3417 47317 3451
rect 47351 3448 47363 3451
rect 48682 3448 48688 3460
rect 47351 3420 48688 3448
rect 47351 3417 47363 3420
rect 47305 3411 47363 3417
rect 48682 3408 48688 3420
rect 48740 3408 48746 3460
rect 27522 3380 27528 3392
rect 24596 3352 27528 3380
rect 27522 3340 27528 3352
rect 27580 3340 27586 3392
rect 35434 3340 35440 3392
rect 35492 3380 35498 3392
rect 45557 3383 45615 3389
rect 45557 3380 45569 3383
rect 35492 3352 45569 3380
rect 35492 3340 35498 3352
rect 45557 3349 45569 3352
rect 45603 3349 45615 3383
rect 45557 3343 45615 3349
rect 1104 3290 49864 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 27950 3290
rect 28002 3238 28014 3290
rect 28066 3238 28078 3290
rect 28130 3238 28142 3290
rect 28194 3238 28206 3290
rect 28258 3238 37950 3290
rect 38002 3238 38014 3290
rect 38066 3238 38078 3290
rect 38130 3238 38142 3290
rect 38194 3238 38206 3290
rect 38258 3238 47950 3290
rect 48002 3238 48014 3290
rect 48066 3238 48078 3290
rect 48130 3238 48142 3290
rect 48194 3238 48206 3290
rect 48258 3238 49864 3290
rect 1104 3216 49864 3238
rect 1302 3136 1308 3188
rect 1360 3176 1366 3188
rect 2133 3179 2191 3185
rect 2133 3176 2145 3179
rect 1360 3148 2145 3176
rect 1360 3136 1366 3148
rect 2133 3145 2145 3148
rect 2179 3145 2191 3179
rect 2133 3139 2191 3145
rect 16301 3179 16359 3185
rect 16301 3145 16313 3179
rect 16347 3176 16359 3179
rect 21174 3176 21180 3188
rect 16347 3148 21180 3176
rect 16347 3145 16359 3148
rect 16301 3139 16359 3145
rect 21174 3136 21180 3148
rect 21232 3136 21238 3188
rect 21269 3179 21327 3185
rect 21269 3145 21281 3179
rect 21315 3176 21327 3179
rect 23198 3176 23204 3188
rect 21315 3148 23204 3176
rect 21315 3145 21327 3148
rect 21269 3139 21327 3145
rect 23198 3136 23204 3148
rect 23256 3136 23262 3188
rect 23566 3176 23572 3188
rect 23308 3148 23572 3176
rect 16666 3108 16672 3120
rect 16054 3080 16672 3108
rect 16666 3068 16672 3080
rect 16724 3068 16730 3120
rect 19058 3108 19064 3120
rect 17604 3080 19064 3108
rect 1302 3000 1308 3052
rect 1360 3040 1366 3052
rect 1581 3043 1639 3049
rect 1581 3040 1593 3043
rect 1360 3012 1593 3040
rect 1360 3000 1366 3012
rect 1581 3009 1593 3012
rect 1627 3040 1639 3043
rect 2501 3043 2559 3049
rect 2501 3040 2513 3043
rect 1627 3012 2513 3040
rect 1627 3009 1639 3012
rect 1581 3003 1639 3009
rect 2501 3009 2513 3012
rect 2547 3009 2559 3043
rect 2501 3003 2559 3009
rect 13814 3000 13820 3052
rect 13872 3040 13878 3052
rect 17604 3049 17632 3080
rect 19058 3068 19064 3080
rect 19116 3068 19122 3120
rect 22094 3108 22100 3120
rect 20180 3080 22100 3108
rect 20180 3049 20208 3080
rect 22094 3068 22100 3080
rect 22152 3108 22158 3120
rect 22646 3108 22652 3120
rect 22152 3080 22652 3108
rect 22152 3068 22158 3080
rect 22646 3068 22652 3080
rect 22704 3068 22710 3120
rect 14553 3043 14611 3049
rect 14553 3040 14565 3043
rect 13872 3012 14565 3040
rect 13872 3000 13878 3012
rect 14553 3009 14565 3012
rect 14599 3009 14611 3043
rect 14553 3003 14611 3009
rect 17589 3043 17647 3049
rect 17589 3009 17601 3043
rect 17635 3009 17647 3043
rect 17589 3003 17647 3009
rect 18325 3043 18383 3049
rect 18325 3009 18337 3043
rect 18371 3009 18383 3043
rect 18325 3003 18383 3009
rect 20165 3043 20223 3049
rect 20165 3009 20177 3043
rect 20211 3009 20223 3043
rect 20165 3003 20223 3009
rect 11054 2932 11060 2984
rect 11112 2972 11118 2984
rect 14829 2975 14887 2981
rect 14829 2972 14841 2975
rect 11112 2944 14841 2972
rect 11112 2932 11118 2944
rect 14829 2941 14841 2944
rect 14875 2941 14887 2975
rect 14829 2935 14887 2941
rect 1765 2907 1823 2913
rect 1765 2873 1777 2907
rect 1811 2904 1823 2907
rect 2406 2904 2412 2916
rect 1811 2876 2412 2904
rect 1811 2873 1823 2876
rect 1765 2867 1823 2873
rect 2406 2864 2412 2876
rect 2464 2864 2470 2916
rect 15838 2864 15844 2916
rect 15896 2904 15902 2916
rect 17405 2907 17463 2913
rect 17405 2904 17417 2907
rect 15896 2876 17417 2904
rect 15896 2864 15902 2876
rect 17405 2873 17417 2876
rect 17451 2873 17463 2907
rect 18340 2904 18368 3003
rect 20806 3000 20812 3052
rect 20864 3000 20870 3052
rect 21450 3000 21456 3052
rect 21508 3000 21514 3052
rect 23308 3049 23336 3148
rect 23566 3136 23572 3148
rect 23624 3176 23630 3188
rect 37734 3176 37740 3188
rect 23624 3148 37740 3176
rect 23624 3136 23630 3148
rect 23382 3068 23388 3120
rect 23440 3108 23446 3120
rect 24489 3111 24547 3117
rect 24489 3108 24501 3111
rect 23440 3080 24501 3108
rect 23440 3068 23446 3080
rect 24489 3077 24501 3080
rect 24535 3077 24547 3111
rect 26878 3108 26884 3120
rect 25714 3080 26884 3108
rect 24489 3071 24547 3077
rect 26878 3068 26884 3080
rect 26936 3068 26942 3120
rect 22189 3043 22247 3049
rect 22189 3009 22201 3043
rect 22235 3040 22247 3043
rect 23293 3043 23351 3049
rect 23293 3040 23305 3043
rect 22235 3012 23305 3040
rect 22235 3009 22247 3012
rect 22189 3003 22247 3009
rect 23293 3009 23305 3012
rect 23339 3009 23351 3043
rect 26605 3043 26663 3049
rect 26605 3040 26617 3043
rect 23293 3003 23351 3009
rect 25700 3012 26617 3040
rect 18414 2932 18420 2984
rect 18472 2972 18478 2984
rect 18601 2975 18659 2981
rect 18601 2972 18613 2975
rect 18472 2944 18613 2972
rect 18472 2932 18478 2944
rect 18601 2941 18613 2944
rect 18647 2941 18659 2975
rect 18601 2935 18659 2941
rect 20990 2932 20996 2984
rect 21048 2972 21054 2984
rect 22002 2972 22008 2984
rect 21048 2944 22008 2972
rect 21048 2932 21054 2944
rect 22002 2932 22008 2944
rect 22060 2972 22066 2984
rect 24213 2975 24271 2981
rect 24213 2972 24225 2975
rect 22060 2944 24225 2972
rect 22060 2932 22066 2944
rect 24213 2941 24225 2944
rect 24259 2941 24271 2975
rect 24213 2935 24271 2941
rect 24578 2932 24584 2984
rect 24636 2972 24642 2984
rect 25700 2972 25728 3012
rect 26605 3009 26617 3012
rect 26651 3009 26663 3043
rect 27448 3038 27476 3148
rect 37734 3136 37740 3148
rect 37792 3136 37798 3188
rect 27706 3068 27712 3120
rect 27764 3108 27770 3120
rect 29638 3108 29644 3120
rect 27764 3080 29644 3108
rect 27764 3068 27770 3080
rect 29638 3068 29644 3080
rect 29696 3068 29702 3120
rect 49145 3111 49203 3117
rect 49145 3077 49157 3111
rect 49191 3108 49203 3111
rect 49234 3108 49240 3120
rect 49191 3080 49240 3108
rect 49191 3077 49203 3080
rect 49145 3071 49203 3077
rect 49234 3068 49240 3080
rect 49292 3068 49298 3120
rect 27525 3043 27583 3049
rect 27525 3038 27537 3043
rect 27448 3010 27537 3038
rect 26605 3003 26663 3009
rect 27525 3009 27537 3010
rect 27571 3009 27583 3043
rect 27525 3003 27583 3009
rect 28810 3000 28816 3052
rect 28868 3040 28874 3052
rect 28905 3043 28963 3049
rect 28905 3040 28917 3043
rect 28868 3012 28917 3040
rect 28868 3000 28874 3012
rect 28905 3009 28917 3012
rect 28951 3009 28963 3043
rect 28905 3003 28963 3009
rect 39758 3000 39764 3052
rect 39816 3040 39822 3052
rect 43993 3043 44051 3049
rect 43993 3040 44005 3043
rect 39816 3012 44005 3040
rect 39816 3000 39822 3012
rect 43993 3009 44005 3012
rect 44039 3009 44051 3043
rect 43993 3003 44051 3009
rect 45738 3000 45744 3052
rect 45796 3040 45802 3052
rect 45833 3043 45891 3049
rect 45833 3040 45845 3043
rect 45796 3012 45845 3040
rect 45796 3000 45802 3012
rect 45833 3009 45845 3012
rect 45879 3009 45891 3043
rect 45833 3003 45891 3009
rect 47302 3000 47308 3052
rect 47360 3040 47366 3052
rect 47949 3043 48007 3049
rect 47949 3040 47961 3043
rect 47360 3012 47961 3040
rect 47360 3000 47366 3012
rect 47949 3009 47961 3012
rect 47995 3009 48007 3043
rect 47949 3003 48007 3009
rect 24636 2944 25728 2972
rect 24636 2932 24642 2944
rect 25958 2932 25964 2984
rect 26016 2972 26022 2984
rect 29181 2975 29239 2981
rect 29181 2972 29193 2975
rect 26016 2944 29193 2972
rect 26016 2932 26022 2944
rect 29181 2941 29193 2944
rect 29227 2941 29239 2975
rect 29181 2935 29239 2941
rect 29638 2932 29644 2984
rect 29696 2972 29702 2984
rect 30650 2972 30656 2984
rect 29696 2944 30656 2972
rect 29696 2932 29702 2944
rect 30650 2932 30656 2944
rect 30708 2972 30714 2984
rect 31021 2975 31079 2981
rect 31021 2972 31033 2975
rect 30708 2944 31033 2972
rect 30708 2932 30714 2944
rect 31021 2941 31033 2944
rect 31067 2941 31079 2975
rect 31021 2935 31079 2941
rect 45189 2975 45247 2981
rect 45189 2941 45201 2975
rect 45235 2972 45247 2975
rect 46750 2972 46756 2984
rect 45235 2944 46756 2972
rect 45235 2941 45247 2944
rect 45189 2935 45247 2941
rect 46750 2932 46756 2944
rect 46808 2932 46814 2984
rect 46842 2932 46848 2984
rect 46900 2932 46906 2984
rect 19981 2907 20039 2913
rect 19981 2904 19993 2907
rect 18340 2876 19993 2904
rect 17405 2867 17463 2873
rect 19981 2873 19993 2876
rect 20027 2873 20039 2907
rect 19981 2867 20039 2873
rect 20625 2907 20683 2913
rect 20625 2873 20637 2907
rect 20671 2904 20683 2907
rect 22370 2904 22376 2916
rect 20671 2876 22376 2904
rect 20671 2873 20683 2876
rect 20625 2867 20683 2873
rect 22370 2864 22376 2876
rect 22428 2864 22434 2916
rect 22646 2864 22652 2916
rect 22704 2864 22710 2916
rect 23198 2864 23204 2916
rect 23256 2904 23262 2916
rect 23256 2876 23888 2904
rect 23256 2864 23262 2876
rect 2314 2796 2320 2848
rect 2372 2796 2378 2848
rect 2774 2796 2780 2848
rect 2832 2796 2838 2848
rect 21174 2796 21180 2848
rect 21232 2836 21238 2848
rect 22281 2839 22339 2845
rect 22281 2836 22293 2839
rect 21232 2808 22293 2836
rect 21232 2796 21238 2808
rect 22281 2805 22293 2808
rect 22327 2805 22339 2839
rect 22281 2799 22339 2805
rect 23382 2796 23388 2848
rect 23440 2796 23446 2848
rect 23474 2796 23480 2848
rect 23532 2836 23538 2848
rect 23753 2839 23811 2845
rect 23753 2836 23765 2839
rect 23532 2808 23765 2836
rect 23532 2796 23538 2808
rect 23753 2805 23765 2808
rect 23799 2805 23811 2839
rect 23860 2836 23888 2876
rect 26878 2864 26884 2916
rect 26936 2904 26942 2916
rect 27706 2904 27712 2916
rect 26936 2876 27712 2904
rect 26936 2864 26942 2876
rect 27706 2864 27712 2876
rect 27764 2864 27770 2916
rect 38286 2904 38292 2916
rect 27816 2876 29040 2904
rect 24578 2836 24584 2848
rect 23860 2808 24584 2836
rect 23753 2799 23811 2805
rect 24578 2796 24584 2808
rect 24636 2796 24642 2848
rect 26421 2839 26479 2845
rect 26421 2805 26433 2839
rect 26467 2836 26479 2839
rect 27154 2836 27160 2848
rect 26467 2808 27160 2836
rect 26467 2805 26479 2808
rect 26421 2799 26479 2805
rect 27154 2796 27160 2808
rect 27212 2796 27218 2848
rect 27816 2845 27844 2876
rect 27801 2839 27859 2845
rect 27801 2805 27813 2839
rect 27847 2805 27859 2839
rect 27801 2799 27859 2805
rect 27890 2796 27896 2848
rect 27948 2836 27954 2848
rect 27985 2839 28043 2845
rect 27985 2836 27997 2839
rect 27948 2808 27997 2836
rect 27948 2796 27954 2808
rect 27985 2805 27997 2808
rect 28031 2805 28043 2839
rect 29012 2836 29040 2876
rect 30668 2876 38292 2904
rect 30668 2845 30696 2876
rect 38286 2864 38292 2876
rect 38344 2864 38350 2916
rect 30653 2839 30711 2845
rect 30653 2836 30665 2839
rect 29012 2808 30665 2836
rect 27985 2799 28043 2805
rect 30653 2805 30665 2808
rect 30699 2805 30711 2839
rect 30653 2799 30711 2805
rect 1104 2746 49864 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 32950 2746
rect 33002 2694 33014 2746
rect 33066 2694 33078 2746
rect 33130 2694 33142 2746
rect 33194 2694 33206 2746
rect 33258 2694 42950 2746
rect 43002 2694 43014 2746
rect 43066 2694 43078 2746
rect 43130 2694 43142 2746
rect 43194 2694 43206 2746
rect 43258 2694 49864 2746
rect 1104 2672 49864 2694
rect 3053 2635 3111 2641
rect 3053 2601 3065 2635
rect 3099 2632 3111 2635
rect 9677 2635 9735 2641
rect 3099 2604 6914 2632
rect 3099 2601 3111 2604
rect 3053 2595 3111 2601
rect 1765 2567 1823 2573
rect 1765 2533 1777 2567
rect 1811 2564 1823 2567
rect 4338 2564 4344 2576
rect 1811 2536 4344 2564
rect 1811 2533 1823 2536
rect 1765 2527 1823 2533
rect 4338 2524 4344 2536
rect 4396 2524 4402 2576
rect 6886 2564 6914 2604
rect 9677 2601 9689 2635
rect 9723 2632 9735 2635
rect 11054 2632 11060 2644
rect 9723 2604 11060 2632
rect 9723 2601 9735 2604
rect 9677 2595 9735 2601
rect 11054 2592 11060 2604
rect 11112 2592 11118 2644
rect 13538 2632 13544 2644
rect 11164 2604 13544 2632
rect 11164 2564 11192 2604
rect 13538 2592 13544 2604
rect 13596 2592 13602 2644
rect 22278 2632 22284 2644
rect 16546 2604 22284 2632
rect 16546 2564 16574 2604
rect 22278 2592 22284 2604
rect 22336 2592 22342 2644
rect 26329 2635 26387 2641
rect 26329 2601 26341 2635
rect 26375 2632 26387 2635
rect 26878 2632 26884 2644
rect 26375 2604 26884 2632
rect 26375 2601 26387 2604
rect 26329 2595 26387 2601
rect 26878 2592 26884 2604
rect 26936 2592 26942 2644
rect 27522 2592 27528 2644
rect 27580 2632 27586 2644
rect 28997 2635 29055 2641
rect 28997 2632 29009 2635
rect 27580 2604 29009 2632
rect 27580 2592 27586 2604
rect 28997 2601 29009 2604
rect 29043 2601 29055 2635
rect 28997 2595 29055 2601
rect 32858 2592 32864 2644
rect 32916 2632 32922 2644
rect 32953 2635 33011 2641
rect 32953 2632 32965 2635
rect 32916 2604 32965 2632
rect 32916 2592 32922 2604
rect 32953 2601 32965 2604
rect 32999 2601 33011 2635
rect 32953 2595 33011 2601
rect 34422 2592 34428 2644
rect 34480 2632 34486 2644
rect 35069 2635 35127 2641
rect 35069 2632 35081 2635
rect 34480 2604 35081 2632
rect 34480 2592 34486 2604
rect 35069 2601 35081 2604
rect 35115 2601 35127 2635
rect 35069 2595 35127 2601
rect 18693 2567 18751 2573
rect 18693 2564 18705 2567
rect 6886 2536 11192 2564
rect 11624 2536 16574 2564
rect 17236 2536 18705 2564
rect 2593 2499 2651 2505
rect 2593 2465 2605 2499
rect 2639 2496 2651 2499
rect 11624 2496 11652 2536
rect 2639 2468 11652 2496
rect 2639 2465 2651 2468
rect 2593 2459 2651 2465
rect 11698 2456 11704 2508
rect 11756 2496 11762 2508
rect 12253 2499 12311 2505
rect 12253 2496 12265 2499
rect 11756 2468 12265 2496
rect 11756 2456 11762 2468
rect 12253 2465 12265 2468
rect 12299 2465 12311 2499
rect 12253 2459 12311 2465
rect 13814 2456 13820 2508
rect 13872 2496 13878 2508
rect 14737 2499 14795 2505
rect 14737 2496 14749 2499
rect 13872 2468 14749 2496
rect 13872 2456 13878 2468
rect 14737 2465 14749 2468
rect 14783 2465 14795 2499
rect 14737 2459 14795 2465
rect 1302 2388 1308 2440
rect 1360 2428 1366 2440
rect 1581 2431 1639 2437
rect 1581 2428 1593 2431
rect 1360 2400 1593 2428
rect 1360 2388 1366 2400
rect 1581 2397 1593 2400
rect 1627 2428 1639 2431
rect 2774 2428 2780 2440
rect 1627 2400 2780 2428
rect 1627 2397 1639 2400
rect 1581 2391 1639 2397
rect 2774 2388 2780 2400
rect 2832 2388 2838 2440
rect 3237 2431 3295 2437
rect 3237 2397 3249 2431
rect 3283 2397 3295 2431
rect 3237 2391 3295 2397
rect 1210 2320 1216 2372
rect 1268 2360 1274 2372
rect 2314 2360 2320 2372
rect 1268 2332 2320 2360
rect 1268 2320 1274 2332
rect 2314 2320 2320 2332
rect 2372 2360 2378 2372
rect 2409 2363 2467 2369
rect 2409 2360 2421 2363
rect 2372 2332 2421 2360
rect 2372 2320 2378 2332
rect 2409 2329 2421 2332
rect 2455 2329 2467 2363
rect 2409 2323 2467 2329
rect 1302 2252 1308 2304
rect 1360 2292 1366 2304
rect 3252 2292 3280 2391
rect 9674 2388 9680 2440
rect 9732 2428 9738 2440
rect 9861 2431 9919 2437
rect 9861 2428 9873 2431
rect 9732 2400 9873 2428
rect 9732 2388 9738 2400
rect 9861 2397 9873 2400
rect 9907 2428 9919 2431
rect 10137 2431 10195 2437
rect 10137 2428 10149 2431
rect 9907 2400 10149 2428
rect 9907 2397 9919 2400
rect 9861 2391 9919 2397
rect 10137 2397 10149 2400
rect 10183 2397 10195 2431
rect 10137 2391 10195 2397
rect 11977 2431 12035 2437
rect 11977 2397 11989 2431
rect 12023 2428 12035 2431
rect 12802 2428 12808 2440
rect 12023 2400 12808 2428
rect 12023 2397 12035 2400
rect 11977 2391 12035 2397
rect 12802 2388 12808 2400
rect 12860 2388 12866 2440
rect 14461 2431 14519 2437
rect 14461 2397 14473 2431
rect 14507 2428 14519 2431
rect 15838 2428 15844 2440
rect 14507 2400 15844 2428
rect 14507 2397 14519 2400
rect 14461 2391 14519 2397
rect 15838 2388 15844 2400
rect 15896 2388 15902 2440
rect 17037 2431 17095 2437
rect 17037 2397 17049 2431
rect 17083 2428 17095 2431
rect 17236 2428 17264 2536
rect 18693 2533 18705 2536
rect 18739 2533 18751 2567
rect 18693 2527 18751 2533
rect 19429 2567 19487 2573
rect 19429 2533 19441 2567
rect 19475 2564 19487 2567
rect 19475 2536 20116 2564
rect 19475 2533 19487 2536
rect 19429 2527 19487 2533
rect 17313 2499 17371 2505
rect 17313 2465 17325 2499
rect 17359 2465 17371 2499
rect 17313 2459 17371 2465
rect 17083 2400 17264 2428
rect 17083 2397 17095 2400
rect 17037 2391 17095 2397
rect 4338 2320 4344 2372
rect 4396 2360 4402 2372
rect 4396 2332 6914 2360
rect 4396 2320 4402 2332
rect 3513 2295 3571 2301
rect 3513 2292 3525 2295
rect 1360 2264 3525 2292
rect 1360 2252 1366 2264
rect 3513 2261 3525 2264
rect 3559 2261 3571 2295
rect 6886 2292 6914 2332
rect 15930 2320 15936 2372
rect 15988 2360 15994 2372
rect 17328 2360 17356 2459
rect 18877 2431 18935 2437
rect 18877 2397 18889 2431
rect 18923 2428 18935 2431
rect 19518 2428 19524 2440
rect 18923 2400 19524 2428
rect 18923 2397 18935 2400
rect 18877 2391 18935 2397
rect 19518 2388 19524 2400
rect 19576 2388 19582 2440
rect 19610 2388 19616 2440
rect 19668 2388 19674 2440
rect 20088 2437 20116 2536
rect 24210 2524 24216 2576
rect 24268 2564 24274 2576
rect 30837 2567 30895 2573
rect 30837 2564 30849 2567
rect 24268 2536 30849 2564
rect 24268 2524 24274 2536
rect 30837 2533 30849 2536
rect 30883 2533 30895 2567
rect 30837 2527 30895 2533
rect 35894 2524 35900 2576
rect 35952 2564 35958 2576
rect 35952 2536 43852 2564
rect 35952 2524 35958 2536
rect 20162 2456 20168 2508
rect 20220 2496 20226 2508
rect 20533 2499 20591 2505
rect 20533 2496 20545 2499
rect 20220 2468 20545 2496
rect 20220 2456 20226 2468
rect 20533 2465 20545 2468
rect 20579 2465 20591 2499
rect 20533 2459 20591 2465
rect 22278 2456 22284 2508
rect 22336 2496 22342 2508
rect 22833 2499 22891 2505
rect 22833 2496 22845 2499
rect 22336 2468 22845 2496
rect 22336 2456 22342 2468
rect 22833 2465 22845 2468
rect 22879 2465 22891 2499
rect 22833 2459 22891 2465
rect 24394 2456 24400 2508
rect 24452 2496 24458 2508
rect 25041 2499 25099 2505
rect 25041 2496 25053 2499
rect 24452 2468 25053 2496
rect 24452 2456 24458 2468
rect 25041 2465 25053 2468
rect 25087 2465 25099 2499
rect 25041 2459 25099 2465
rect 26510 2456 26516 2508
rect 26568 2496 26574 2508
rect 27617 2499 27675 2505
rect 27617 2496 27629 2499
rect 26568 2468 27629 2496
rect 26568 2456 26574 2468
rect 27617 2465 27629 2468
rect 27663 2465 27675 2499
rect 27617 2459 27675 2465
rect 37734 2456 37740 2508
rect 37792 2456 37798 2508
rect 41322 2456 41328 2508
rect 41380 2496 41386 2508
rect 43824 2505 43852 2536
rect 41417 2499 41475 2505
rect 41417 2496 41429 2499
rect 41380 2468 41429 2496
rect 41380 2456 41386 2468
rect 41417 2465 41429 2468
rect 41463 2465 41475 2499
rect 41417 2459 41475 2465
rect 43809 2499 43867 2505
rect 43809 2465 43821 2499
rect 43855 2465 43867 2499
rect 43809 2459 43867 2465
rect 49142 2456 49148 2508
rect 49200 2456 49206 2508
rect 20073 2431 20131 2437
rect 20073 2397 20085 2431
rect 20119 2397 20131 2431
rect 20073 2391 20131 2397
rect 22370 2388 22376 2440
rect 22428 2388 22434 2440
rect 24578 2388 24584 2440
rect 24636 2388 24642 2440
rect 27154 2388 27160 2440
rect 27212 2388 27218 2440
rect 28994 2388 29000 2440
rect 29052 2428 29058 2440
rect 29181 2431 29239 2437
rect 29181 2428 29193 2431
rect 29052 2400 29193 2428
rect 29052 2388 29058 2400
rect 29181 2397 29193 2400
rect 29227 2428 29239 2431
rect 29549 2431 29607 2437
rect 29549 2428 29561 2431
rect 29227 2400 29561 2428
rect 29227 2397 29239 2400
rect 29181 2391 29239 2397
rect 29549 2397 29561 2400
rect 29595 2397 29607 2431
rect 29549 2391 29607 2397
rect 30742 2388 30748 2440
rect 30800 2428 30806 2440
rect 31021 2431 31079 2437
rect 31021 2428 31033 2431
rect 30800 2400 31033 2428
rect 30800 2388 30806 2400
rect 31021 2397 31033 2400
rect 31067 2428 31079 2431
rect 31297 2431 31355 2437
rect 31297 2428 31309 2431
rect 31067 2400 31309 2428
rect 31067 2397 31079 2400
rect 31021 2391 31079 2397
rect 31297 2397 31309 2400
rect 31343 2397 31355 2431
rect 31297 2391 31355 2397
rect 33134 2388 33140 2440
rect 33192 2428 33198 2440
rect 33413 2431 33471 2437
rect 33413 2428 33425 2431
rect 33192 2400 33425 2428
rect 33192 2388 33198 2400
rect 33413 2397 33425 2400
rect 33459 2397 33471 2431
rect 33413 2391 33471 2397
rect 34974 2388 34980 2440
rect 35032 2428 35038 2440
rect 35253 2431 35311 2437
rect 35253 2428 35265 2431
rect 35032 2400 35265 2428
rect 35032 2388 35038 2400
rect 35253 2397 35265 2400
rect 35299 2428 35311 2431
rect 35529 2431 35587 2437
rect 35529 2428 35541 2431
rect 35299 2400 35541 2428
rect 35299 2397 35311 2400
rect 35253 2391 35311 2397
rect 35529 2397 35541 2400
rect 35575 2397 35587 2431
rect 37461 2431 37519 2437
rect 37461 2428 37473 2431
rect 35529 2391 35587 2397
rect 37108 2400 37473 2428
rect 15988 2332 17356 2360
rect 15988 2320 15994 2332
rect 37108 2304 37136 2400
rect 37461 2397 37473 2400
rect 37507 2397 37519 2431
rect 37461 2391 37519 2397
rect 38286 2388 38292 2440
rect 38344 2428 38350 2440
rect 40681 2431 40739 2437
rect 40681 2428 40693 2431
rect 38344 2400 40693 2428
rect 38344 2388 38350 2400
rect 40681 2397 40693 2400
rect 40727 2397 40739 2431
rect 43533 2431 43591 2437
rect 43533 2428 43545 2431
rect 40681 2391 40739 2397
rect 43456 2400 43545 2428
rect 43456 2304 43484 2400
rect 43533 2397 43545 2400
rect 43579 2397 43591 2431
rect 43533 2391 43591 2397
rect 45646 2388 45652 2440
rect 45704 2428 45710 2440
rect 45833 2431 45891 2437
rect 45833 2428 45845 2431
rect 45704 2400 45845 2428
rect 45704 2388 45710 2400
rect 45833 2397 45845 2400
rect 45879 2397 45891 2431
rect 45833 2391 45891 2397
rect 47210 2388 47216 2440
rect 47268 2428 47274 2440
rect 47949 2431 48007 2437
rect 47949 2428 47961 2431
rect 47268 2400 47961 2428
rect 47268 2388 47274 2400
rect 47949 2397 47961 2400
rect 47995 2397 48007 2431
rect 47949 2391 48007 2397
rect 47029 2363 47087 2369
rect 47029 2329 47041 2363
rect 47075 2360 47087 2363
rect 48498 2360 48504 2372
rect 47075 2332 48504 2360
rect 47075 2329 47087 2332
rect 47029 2323 47087 2329
rect 48498 2320 48504 2332
rect 48556 2320 48562 2372
rect 12710 2292 12716 2304
rect 6886 2264 12716 2292
rect 3513 2255 3571 2261
rect 12710 2252 12716 2264
rect 12768 2252 12774 2304
rect 37090 2252 37096 2304
rect 37148 2252 37154 2304
rect 43257 2295 43315 2301
rect 43257 2261 43269 2295
rect 43303 2292 43315 2295
rect 43438 2292 43444 2304
rect 43303 2264 43444 2292
rect 43303 2261 43315 2264
rect 43257 2255 43315 2261
rect 43438 2252 43444 2264
rect 43496 2252 43502 2304
rect 1104 2202 49864 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 27950 2202
rect 28002 2150 28014 2202
rect 28066 2150 28078 2202
rect 28130 2150 28142 2202
rect 28194 2150 28206 2202
rect 28258 2150 37950 2202
rect 38002 2150 38014 2202
rect 38066 2150 38078 2202
rect 38130 2150 38142 2202
rect 38194 2150 38206 2202
rect 38258 2150 47950 2202
rect 48002 2150 48014 2202
rect 48066 2150 48078 2202
rect 48130 2150 48142 2202
rect 48194 2150 48206 2202
rect 48258 2150 49864 2202
rect 1104 2128 49864 2150
<< via1 >>
rect 30656 26324 30708 26376
rect 40132 26324 40184 26376
rect 3424 25032 3476 25084
rect 10048 25032 10100 25084
rect 29368 25032 29420 25084
rect 40408 25032 40460 25084
rect 31300 24964 31352 25016
rect 42800 24964 42852 25016
rect 4068 24896 4120 24948
rect 8852 24896 8904 24948
rect 29644 24896 29696 24948
rect 44272 24896 44324 24948
rect 25596 24828 25648 24880
rect 48320 24828 48372 24880
rect 25872 24760 25924 24812
rect 35440 24760 35492 24812
rect 37924 24760 37976 24812
rect 40500 24760 40552 24812
rect 16028 24692 16080 24744
rect 24584 24692 24636 24744
rect 27988 24692 28040 24744
rect 29184 24692 29236 24744
rect 34796 24692 34848 24744
rect 38660 24692 38712 24744
rect 17868 24624 17920 24676
rect 23296 24624 23348 24676
rect 23388 24624 23440 24676
rect 26700 24624 26752 24676
rect 29092 24624 29144 24676
rect 3884 24556 3936 24608
rect 6644 24556 6696 24608
rect 17040 24556 17092 24608
rect 24308 24556 24360 24608
rect 24768 24556 24820 24608
rect 30564 24556 30616 24608
rect 31852 24624 31904 24676
rect 40040 24624 40092 24676
rect 32312 24556 32364 24608
rect 34060 24556 34112 24608
rect 39672 24556 39724 24608
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 32950 24454 33002 24506
rect 33014 24454 33066 24506
rect 33078 24454 33130 24506
rect 33142 24454 33194 24506
rect 33206 24454 33258 24506
rect 42950 24454 43002 24506
rect 43014 24454 43066 24506
rect 43078 24454 43130 24506
rect 43142 24454 43194 24506
rect 43206 24454 43258 24506
rect 2780 24352 2832 24404
rect 6184 24352 6236 24404
rect 7748 24352 7800 24404
rect 20720 24352 20772 24404
rect 3516 24216 3568 24268
rect 6736 24284 6788 24336
rect 2320 24148 2372 24200
rect 10140 24284 10192 24336
rect 8668 24216 8720 24268
rect 11888 24284 11940 24336
rect 2136 24080 2188 24132
rect 7380 24191 7432 24200
rect 7380 24157 7389 24191
rect 7389 24157 7423 24191
rect 7423 24157 7432 24191
rect 7380 24148 7432 24157
rect 5540 24012 5592 24064
rect 7472 24012 7524 24064
rect 9128 24055 9180 24064
rect 9128 24021 9137 24055
rect 9137 24021 9171 24055
rect 9171 24021 9180 24055
rect 9128 24012 9180 24021
rect 10876 24080 10928 24132
rect 14924 24284 14976 24336
rect 13820 24216 13872 24268
rect 17684 24216 17736 24268
rect 19616 24284 19668 24336
rect 20996 24284 21048 24336
rect 24032 24284 24084 24336
rect 24584 24395 24636 24404
rect 24584 24361 24593 24395
rect 24593 24361 24627 24395
rect 24627 24361 24636 24395
rect 24584 24352 24636 24361
rect 25964 24395 26016 24404
rect 25964 24361 25973 24395
rect 25973 24361 26007 24395
rect 26007 24361 26016 24395
rect 25964 24352 26016 24361
rect 29920 24352 29972 24404
rect 27252 24284 27304 24336
rect 28632 24284 28684 24336
rect 31484 24284 31536 24336
rect 32312 24395 32364 24404
rect 32312 24361 32321 24395
rect 32321 24361 32355 24395
rect 32355 24361 32364 24395
rect 32312 24352 32364 24361
rect 32404 24352 32456 24404
rect 13728 24148 13780 24200
rect 14372 24148 14424 24200
rect 12624 24080 12676 24132
rect 19340 24148 19392 24200
rect 20904 24259 20956 24268
rect 20904 24225 20913 24259
rect 20913 24225 20947 24259
rect 20947 24225 20956 24259
rect 20904 24216 20956 24225
rect 18420 24080 18472 24132
rect 9772 24012 9824 24064
rect 11704 24055 11756 24064
rect 11704 24021 11713 24055
rect 11713 24021 11747 24055
rect 11747 24021 11756 24055
rect 11704 24012 11756 24021
rect 11796 24012 11848 24064
rect 18512 24012 18564 24064
rect 19432 24055 19484 24064
rect 19432 24021 19441 24055
rect 19441 24021 19475 24055
rect 19475 24021 19484 24055
rect 19432 24012 19484 24021
rect 20536 24148 20588 24200
rect 21272 24148 21324 24200
rect 25044 24148 25096 24200
rect 20444 24080 20496 24132
rect 27344 24216 27396 24268
rect 25872 24191 25924 24200
rect 25872 24157 25881 24191
rect 25881 24157 25915 24191
rect 25915 24157 25924 24191
rect 25872 24148 25924 24157
rect 26056 24148 26108 24200
rect 27160 24080 27212 24132
rect 30104 24148 30156 24200
rect 30564 24191 30616 24200
rect 30564 24157 30573 24191
rect 30573 24157 30607 24191
rect 30607 24157 30616 24191
rect 30564 24148 30616 24157
rect 31116 24148 31168 24200
rect 31484 24148 31536 24200
rect 32128 24148 32180 24200
rect 34428 24284 34480 24336
rect 34060 24259 34112 24268
rect 34060 24225 34069 24259
rect 34069 24225 34103 24259
rect 34103 24225 34112 24259
rect 34060 24216 34112 24225
rect 35348 24216 35400 24268
rect 35532 24259 35584 24268
rect 35532 24225 35541 24259
rect 35541 24225 35575 24259
rect 35575 24225 35584 24259
rect 35532 24216 35584 24225
rect 30748 24080 30800 24132
rect 31944 24080 31996 24132
rect 36084 24148 36136 24200
rect 40316 24352 40368 24404
rect 40500 24352 40552 24404
rect 40868 24352 40920 24404
rect 39120 24284 39172 24336
rect 37372 24216 37424 24268
rect 37924 24259 37976 24268
rect 37924 24225 37933 24259
rect 37933 24225 37967 24259
rect 37967 24225 37976 24259
rect 37924 24216 37976 24225
rect 38292 24216 38344 24268
rect 34152 24080 34204 24132
rect 22560 24012 22612 24064
rect 24676 24012 24728 24064
rect 24952 24055 25004 24064
rect 24952 24021 24961 24055
rect 24961 24021 24995 24055
rect 24995 24021 25004 24055
rect 24952 24012 25004 24021
rect 26148 24012 26200 24064
rect 26240 24012 26292 24064
rect 26424 24012 26476 24064
rect 27344 24055 27396 24064
rect 27344 24021 27353 24055
rect 27353 24021 27387 24055
rect 27387 24021 27396 24055
rect 27344 24012 27396 24021
rect 28632 24012 28684 24064
rect 30380 24055 30432 24064
rect 30380 24021 30389 24055
rect 30389 24021 30423 24055
rect 30423 24021 30432 24055
rect 30380 24012 30432 24021
rect 30932 24012 30984 24064
rect 31116 24012 31168 24064
rect 32956 24055 33008 24064
rect 32956 24021 32965 24055
rect 32965 24021 32999 24055
rect 32999 24021 33008 24055
rect 32956 24012 33008 24021
rect 37740 24080 37792 24132
rect 38936 24191 38988 24200
rect 38936 24157 38945 24191
rect 38945 24157 38979 24191
rect 38979 24157 38988 24191
rect 38936 24148 38988 24157
rect 40132 24148 40184 24200
rect 40684 24259 40736 24268
rect 40684 24225 40693 24259
rect 40693 24225 40727 24259
rect 40727 24225 40736 24259
rect 40684 24216 40736 24225
rect 40960 24259 41012 24268
rect 40960 24225 40969 24259
rect 40969 24225 41003 24259
rect 41003 24225 41012 24259
rect 40960 24216 41012 24225
rect 47492 24216 47544 24268
rect 48228 24216 48280 24268
rect 41328 24148 41380 24200
rect 42156 24148 42208 24200
rect 44640 24148 44692 24200
rect 44732 24148 44784 24200
rect 45284 24191 45336 24200
rect 45284 24157 45293 24191
rect 45293 24157 45327 24191
rect 45327 24157 45336 24191
rect 45284 24148 45336 24157
rect 45560 24148 45612 24200
rect 47308 24148 47360 24200
rect 48780 24191 48832 24200
rect 48780 24157 48789 24191
rect 48789 24157 48823 24191
rect 48823 24157 48832 24191
rect 48780 24148 48832 24157
rect 41788 24080 41840 24132
rect 42248 24080 42300 24132
rect 46020 24080 46072 24132
rect 46756 24123 46808 24132
rect 46756 24089 46765 24123
rect 46765 24089 46799 24123
rect 46799 24089 46808 24123
rect 46756 24080 46808 24089
rect 35256 24055 35308 24064
rect 35256 24021 35265 24055
rect 35265 24021 35299 24055
rect 35299 24021 35308 24055
rect 35256 24012 35308 24021
rect 35440 24012 35492 24064
rect 35992 24012 36044 24064
rect 36176 24012 36228 24064
rect 37648 24012 37700 24064
rect 40500 24012 40552 24064
rect 41972 24055 42024 24064
rect 41972 24021 41981 24055
rect 41981 24021 42015 24055
rect 42015 24021 42024 24055
rect 41972 24012 42024 24021
rect 42156 24055 42208 24064
rect 42156 24021 42165 24055
rect 42165 24021 42199 24055
rect 42199 24021 42208 24055
rect 42156 24012 42208 24021
rect 43996 24012 44048 24064
rect 46112 24055 46164 24064
rect 46112 24021 46121 24055
rect 46121 24021 46155 24055
rect 46155 24021 46164 24055
rect 46112 24012 46164 24021
rect 46204 24012 46256 24064
rect 46940 24012 46992 24064
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 27950 23910 28002 23962
rect 28014 23910 28066 23962
rect 28078 23910 28130 23962
rect 28142 23910 28194 23962
rect 28206 23910 28258 23962
rect 37950 23910 38002 23962
rect 38014 23910 38066 23962
rect 38078 23910 38130 23962
rect 38142 23910 38194 23962
rect 38206 23910 38258 23962
rect 47950 23910 48002 23962
rect 48014 23910 48066 23962
rect 48078 23910 48130 23962
rect 48142 23910 48194 23962
rect 48206 23910 48258 23962
rect 2136 23851 2188 23860
rect 2136 23817 2145 23851
rect 2145 23817 2179 23851
rect 2179 23817 2188 23851
rect 2136 23808 2188 23817
rect 4160 23740 4212 23792
rect 3700 23672 3752 23724
rect 4712 23715 4764 23724
rect 4712 23681 4721 23715
rect 4721 23681 4755 23715
rect 4755 23681 4764 23715
rect 4712 23672 4764 23681
rect 5448 23647 5500 23656
rect 5448 23613 5457 23647
rect 5457 23613 5491 23647
rect 5491 23613 5500 23647
rect 5448 23604 5500 23613
rect 7748 23672 7800 23724
rect 11796 23808 11848 23860
rect 17040 23808 17092 23860
rect 9312 23740 9364 23792
rect 10692 23783 10744 23792
rect 10692 23749 10701 23783
rect 10701 23749 10735 23783
rect 10735 23749 10744 23783
rect 10692 23740 10744 23749
rect 10876 23740 10928 23792
rect 12348 23740 12400 23792
rect 12440 23672 12492 23724
rect 4068 23536 4120 23588
rect 6736 23536 6788 23588
rect 8392 23604 8444 23656
rect 14188 23740 14240 23792
rect 14464 23740 14516 23792
rect 16120 23783 16172 23792
rect 16120 23749 16129 23783
rect 16129 23749 16163 23783
rect 16163 23749 16172 23783
rect 16120 23740 16172 23749
rect 20996 23808 21048 23860
rect 21272 23851 21324 23860
rect 21272 23817 21281 23851
rect 21281 23817 21315 23851
rect 21315 23817 21324 23851
rect 21272 23808 21324 23817
rect 18328 23740 18380 23792
rect 10324 23536 10376 23588
rect 20168 23672 20220 23724
rect 17960 23604 18012 23656
rect 4804 23468 4856 23520
rect 12348 23468 12400 23520
rect 15384 23468 15436 23520
rect 19064 23647 19116 23656
rect 19064 23613 19073 23647
rect 19073 23613 19107 23647
rect 19107 23613 19116 23647
rect 19064 23604 19116 23613
rect 22100 23604 22152 23656
rect 23296 23851 23348 23860
rect 23296 23817 23305 23851
rect 23305 23817 23339 23851
rect 23339 23817 23348 23851
rect 23296 23808 23348 23817
rect 23848 23740 23900 23792
rect 23940 23740 23992 23792
rect 24952 23808 25004 23860
rect 26148 23808 26200 23860
rect 26516 23808 26568 23860
rect 25412 23740 25464 23792
rect 26424 23740 26476 23792
rect 26976 23740 27028 23792
rect 20168 23536 20220 23588
rect 20352 23468 20404 23520
rect 20536 23511 20588 23520
rect 20536 23477 20545 23511
rect 20545 23477 20579 23511
rect 20579 23477 20588 23511
rect 20536 23468 20588 23477
rect 20720 23536 20772 23588
rect 22008 23536 22060 23588
rect 23756 23604 23808 23656
rect 24492 23536 24544 23588
rect 21088 23468 21140 23520
rect 24584 23468 24636 23520
rect 24860 23647 24912 23656
rect 24860 23613 24869 23647
rect 24869 23613 24903 23647
rect 24903 23613 24912 23647
rect 24860 23604 24912 23613
rect 26516 23468 26568 23520
rect 26608 23511 26660 23520
rect 26608 23477 26617 23511
rect 26617 23477 26651 23511
rect 26651 23477 26660 23511
rect 26608 23468 26660 23477
rect 26700 23468 26752 23520
rect 27988 23715 28040 23724
rect 27988 23681 27997 23715
rect 27997 23681 28031 23715
rect 28031 23681 28040 23715
rect 27988 23672 28040 23681
rect 31576 23808 31628 23860
rect 31668 23808 31720 23860
rect 32956 23808 33008 23860
rect 29460 23740 29512 23792
rect 30748 23740 30800 23792
rect 34428 23740 34480 23792
rect 29184 23672 29236 23724
rect 32680 23715 32732 23724
rect 32680 23681 32689 23715
rect 32689 23681 32723 23715
rect 32723 23681 32732 23715
rect 32680 23672 32732 23681
rect 27804 23604 27856 23656
rect 29736 23536 29788 23588
rect 27620 23468 27672 23520
rect 27712 23468 27764 23520
rect 29184 23468 29236 23520
rect 30656 23604 30708 23656
rect 32588 23604 32640 23656
rect 31576 23536 31628 23588
rect 31392 23468 31444 23520
rect 31760 23511 31812 23520
rect 31760 23477 31769 23511
rect 31769 23477 31803 23511
rect 31803 23477 31812 23511
rect 31760 23468 31812 23477
rect 33600 23647 33652 23656
rect 33600 23613 33609 23647
rect 33609 23613 33643 23647
rect 33643 23613 33652 23647
rect 33600 23604 33652 23613
rect 34336 23604 34388 23656
rect 44180 23808 44232 23860
rect 45284 23808 45336 23860
rect 35348 23740 35400 23792
rect 37556 23740 37608 23792
rect 37740 23740 37792 23792
rect 38384 23740 38436 23792
rect 35808 23672 35860 23724
rect 37464 23672 37516 23724
rect 40040 23672 40092 23724
rect 40132 23672 40184 23724
rect 40592 23672 40644 23724
rect 40776 23740 40828 23792
rect 42432 23740 42484 23792
rect 46848 23783 46900 23792
rect 46848 23749 46857 23783
rect 46857 23749 46891 23783
rect 46891 23749 46900 23783
rect 46848 23740 46900 23749
rect 42156 23672 42208 23724
rect 42800 23672 42852 23724
rect 44272 23672 44324 23724
rect 45376 23715 45428 23724
rect 45376 23681 45385 23715
rect 45385 23681 45419 23715
rect 45419 23681 45428 23715
rect 45376 23672 45428 23681
rect 36360 23647 36412 23656
rect 36360 23613 36369 23647
rect 36369 23613 36403 23647
rect 36403 23613 36412 23647
rect 36360 23604 36412 23613
rect 36452 23647 36504 23656
rect 36452 23613 36461 23647
rect 36461 23613 36495 23647
rect 36495 23613 36504 23647
rect 36452 23604 36504 23613
rect 39304 23647 39356 23656
rect 39304 23613 39313 23647
rect 39313 23613 39347 23647
rect 39347 23613 39356 23647
rect 39304 23604 39356 23613
rect 39396 23647 39448 23656
rect 39396 23613 39405 23647
rect 39405 23613 39439 23647
rect 39439 23613 39448 23647
rect 39396 23604 39448 23613
rect 40408 23604 40460 23656
rect 41788 23647 41840 23656
rect 41788 23613 41797 23647
rect 41797 23613 41831 23647
rect 41831 23613 41840 23647
rect 41788 23604 41840 23613
rect 42616 23647 42668 23656
rect 42616 23613 42625 23647
rect 42625 23613 42659 23647
rect 42659 23613 42668 23647
rect 42616 23604 42668 23613
rect 43904 23647 43956 23656
rect 43904 23613 43913 23647
rect 43913 23613 43947 23647
rect 43947 23613 43956 23647
rect 43904 23604 43956 23613
rect 46756 23672 46808 23724
rect 47860 23672 47912 23724
rect 48596 23672 48648 23724
rect 46480 23604 46532 23656
rect 48412 23604 48464 23656
rect 37648 23536 37700 23588
rect 38476 23579 38528 23588
rect 38476 23545 38485 23579
rect 38485 23545 38519 23579
rect 38519 23545 38528 23579
rect 38476 23536 38528 23545
rect 34980 23468 35032 23520
rect 35900 23511 35952 23520
rect 35900 23477 35909 23511
rect 35909 23477 35943 23511
rect 35943 23477 35952 23511
rect 35900 23468 35952 23477
rect 37280 23468 37332 23520
rect 38384 23468 38436 23520
rect 38660 23468 38712 23520
rect 41604 23468 41656 23520
rect 42432 23536 42484 23588
rect 45192 23579 45244 23588
rect 45192 23545 45201 23579
rect 45201 23545 45235 23579
rect 45235 23545 45244 23579
rect 45192 23536 45244 23545
rect 42248 23468 42300 23520
rect 45376 23468 45428 23520
rect 47124 23468 47176 23520
rect 49148 23468 49200 23520
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 32950 23366 33002 23418
rect 33014 23366 33066 23418
rect 33078 23366 33130 23418
rect 33142 23366 33194 23418
rect 33206 23366 33258 23418
rect 42950 23366 43002 23418
rect 43014 23366 43066 23418
rect 43078 23366 43130 23418
rect 43142 23366 43194 23418
rect 43206 23366 43258 23418
rect 2872 23264 2924 23316
rect 4344 23264 4396 23316
rect 4712 23307 4764 23316
rect 4712 23273 4721 23307
rect 4721 23273 4755 23307
rect 4755 23273 4764 23307
rect 4712 23264 4764 23273
rect 14188 23307 14240 23316
rect 14188 23273 14197 23307
rect 14197 23273 14231 23307
rect 14231 23273 14240 23307
rect 14188 23264 14240 23273
rect 1584 23128 1636 23180
rect 4436 23128 4488 23180
rect 6092 23171 6144 23180
rect 6092 23137 6101 23171
rect 6101 23137 6135 23171
rect 6135 23137 6144 23171
rect 6092 23128 6144 23137
rect 7840 23171 7892 23180
rect 7840 23137 7849 23171
rect 7849 23137 7883 23171
rect 7883 23137 7892 23171
rect 7840 23128 7892 23137
rect 15844 23196 15896 23248
rect 11244 23171 11296 23180
rect 11244 23137 11253 23171
rect 11253 23137 11287 23171
rect 11287 23137 11296 23171
rect 11244 23128 11296 23137
rect 13360 23171 13412 23180
rect 13360 23137 13369 23171
rect 13369 23137 13403 23171
rect 13403 23137 13412 23171
rect 13360 23128 13412 23137
rect 2780 23035 2832 23044
rect 2780 23001 2789 23035
rect 2789 23001 2823 23035
rect 2823 23001 2832 23035
rect 2780 22992 2832 23001
rect 3608 22924 3660 22976
rect 4528 23060 4580 23112
rect 5080 23060 5132 23112
rect 5540 23060 5592 23112
rect 9128 23060 9180 23112
rect 12348 23060 12400 23112
rect 13912 23060 13964 23112
rect 7748 22992 7800 23044
rect 6920 22924 6972 22976
rect 7012 22924 7064 22976
rect 14648 22967 14700 22976
rect 14648 22933 14657 22967
rect 14657 22933 14691 22967
rect 14691 22933 14700 22967
rect 14648 22924 14700 22933
rect 15752 23171 15804 23180
rect 15752 23137 15761 23171
rect 15761 23137 15795 23171
rect 15795 23137 15804 23171
rect 15752 23128 15804 23137
rect 17960 23264 18012 23316
rect 22836 23264 22888 23316
rect 19340 23171 19392 23180
rect 17040 23060 17092 23112
rect 19340 23137 19349 23171
rect 19349 23137 19383 23171
rect 19383 23137 19392 23171
rect 19340 23128 19392 23137
rect 20168 23128 20220 23180
rect 19248 23060 19300 23112
rect 20352 23171 20404 23180
rect 20352 23137 20361 23171
rect 20361 23137 20395 23171
rect 20395 23137 20404 23171
rect 20352 23128 20404 23137
rect 22008 23196 22060 23248
rect 22100 23239 22152 23248
rect 22100 23205 22109 23239
rect 22109 23205 22143 23239
rect 22143 23205 22152 23239
rect 22100 23196 22152 23205
rect 23756 23264 23808 23316
rect 24032 23264 24084 23316
rect 25228 23307 25280 23316
rect 25228 23273 25237 23307
rect 25237 23273 25271 23307
rect 25271 23273 25280 23307
rect 25228 23264 25280 23273
rect 25412 23264 25464 23316
rect 27988 23264 28040 23316
rect 29736 23307 29788 23316
rect 29736 23273 29745 23307
rect 29745 23273 29779 23307
rect 29779 23273 29788 23307
rect 29736 23264 29788 23273
rect 24584 23196 24636 23248
rect 25504 23196 25556 23248
rect 27528 23196 27580 23248
rect 17316 22992 17368 23044
rect 17408 23035 17460 23044
rect 17408 23001 17417 23035
rect 17417 23001 17451 23035
rect 17451 23001 17460 23035
rect 17408 22992 17460 23001
rect 19708 23035 19760 23044
rect 19708 23001 19717 23035
rect 19717 23001 19751 23035
rect 19751 23001 19760 23035
rect 19708 22992 19760 23001
rect 20720 22992 20772 23044
rect 21088 22992 21140 23044
rect 22008 23060 22060 23112
rect 26608 23128 26660 23180
rect 26700 23128 26752 23180
rect 29276 23196 29328 23248
rect 32128 23264 32180 23316
rect 33968 23264 34020 23316
rect 35072 23264 35124 23316
rect 37280 23264 37332 23316
rect 37556 23264 37608 23316
rect 40040 23307 40092 23316
rect 40040 23273 40049 23307
rect 40049 23273 40083 23307
rect 40083 23273 40092 23307
rect 40040 23264 40092 23273
rect 40224 23264 40276 23316
rect 40868 23264 40920 23316
rect 29460 23128 29512 23180
rect 30196 23171 30248 23180
rect 30196 23137 30205 23171
rect 30205 23137 30239 23171
rect 30239 23137 30248 23171
rect 30196 23128 30248 23137
rect 24400 23060 24452 23112
rect 17500 22924 17552 22976
rect 18880 22967 18932 22976
rect 18880 22933 18889 22967
rect 18889 22933 18923 22967
rect 18923 22933 18932 22967
rect 18880 22924 18932 22933
rect 20536 22924 20588 22976
rect 22284 22924 22336 22976
rect 25320 23060 25372 23112
rect 25688 23103 25740 23112
rect 25688 23069 25697 23103
rect 25697 23069 25731 23103
rect 25731 23069 25740 23103
rect 25688 23060 25740 23069
rect 27620 23060 27672 23112
rect 28540 23060 28592 23112
rect 24676 23035 24728 23044
rect 24676 23001 24685 23035
rect 24685 23001 24719 23035
rect 24719 23001 24728 23035
rect 24676 22992 24728 23001
rect 26424 22992 26476 23044
rect 24492 22924 24544 22976
rect 25136 22924 25188 22976
rect 28448 22992 28500 23044
rect 31392 23171 31444 23180
rect 31392 23137 31401 23171
rect 31401 23137 31435 23171
rect 31435 23137 31444 23171
rect 31392 23128 31444 23137
rect 34980 23196 35032 23248
rect 31760 23128 31812 23180
rect 33692 23128 33744 23180
rect 35072 23171 35124 23180
rect 35072 23137 35081 23171
rect 35081 23137 35115 23171
rect 35115 23137 35124 23171
rect 35072 23128 35124 23137
rect 39212 23196 39264 23248
rect 42800 23264 42852 23316
rect 44640 23264 44692 23316
rect 45468 23264 45520 23316
rect 47768 23264 47820 23316
rect 43904 23196 43956 23248
rect 37280 23171 37332 23180
rect 37280 23137 37289 23171
rect 37289 23137 37323 23171
rect 37323 23137 37332 23171
rect 37280 23128 37332 23137
rect 28264 22967 28316 22976
rect 28264 22933 28273 22967
rect 28273 22933 28307 22967
rect 28307 22933 28316 22967
rect 28264 22924 28316 22933
rect 29460 22924 29512 22976
rect 30104 22967 30156 22976
rect 30104 22933 30113 22967
rect 30113 22933 30147 22967
rect 30147 22933 30156 22967
rect 30104 22924 30156 22933
rect 31944 22992 31996 23044
rect 31024 22924 31076 22976
rect 31116 22924 31168 22976
rect 38844 23128 38896 23180
rect 41420 23128 41472 23180
rect 47676 23239 47728 23248
rect 47676 23205 47685 23239
rect 47685 23205 47719 23239
rect 47719 23205 47728 23239
rect 47676 23196 47728 23205
rect 46480 23171 46532 23180
rect 46480 23137 46489 23171
rect 46489 23137 46523 23171
rect 46523 23137 46532 23171
rect 46480 23128 46532 23137
rect 42892 23060 42944 23112
rect 43996 23060 44048 23112
rect 44088 23060 44140 23112
rect 49240 23128 49292 23180
rect 47860 23103 47912 23112
rect 47860 23069 47869 23103
rect 47869 23069 47903 23103
rect 47903 23069 47912 23103
rect 47860 23060 47912 23069
rect 48320 23103 48372 23112
rect 48320 23069 48329 23103
rect 48329 23069 48363 23103
rect 48363 23069 48372 23103
rect 48320 23060 48372 23069
rect 49332 23060 49384 23112
rect 33600 22992 33652 23044
rect 34428 22992 34480 23044
rect 35808 22992 35860 23044
rect 37832 22992 37884 23044
rect 33784 22924 33836 22976
rect 33876 22924 33928 22976
rect 34796 22924 34848 22976
rect 34980 22924 35032 22976
rect 35256 22924 35308 22976
rect 38844 22924 38896 22976
rect 39580 22967 39632 22976
rect 39580 22933 39589 22967
rect 39589 22933 39623 22967
rect 39623 22933 39632 22967
rect 39580 22924 39632 22933
rect 40408 22967 40460 22976
rect 40408 22933 40417 22967
rect 40417 22933 40451 22967
rect 40451 22933 40460 22967
rect 40408 22924 40460 22933
rect 41236 22992 41288 23044
rect 42064 22992 42116 23044
rect 43536 23035 43588 23044
rect 43536 23001 43545 23035
rect 43545 23001 43579 23035
rect 43579 23001 43588 23035
rect 43536 22992 43588 23001
rect 42156 22924 42208 22976
rect 42616 22924 42668 22976
rect 43996 22924 44048 22976
rect 48596 22992 48648 23044
rect 48504 22967 48556 22976
rect 48504 22933 48513 22967
rect 48513 22933 48547 22967
rect 48547 22933 48556 22967
rect 48504 22924 48556 22933
rect 49240 22967 49292 22976
rect 49240 22933 49249 22967
rect 49249 22933 49283 22967
rect 49283 22933 49292 22967
rect 49240 22924 49292 22933
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 27950 22822 28002 22874
rect 28014 22822 28066 22874
rect 28078 22822 28130 22874
rect 28142 22822 28194 22874
rect 28206 22822 28258 22874
rect 37950 22822 38002 22874
rect 38014 22822 38066 22874
rect 38078 22822 38130 22874
rect 38142 22822 38194 22874
rect 38206 22822 38258 22874
rect 47950 22822 48002 22874
rect 48014 22822 48066 22874
rect 48078 22822 48130 22874
rect 48142 22822 48194 22874
rect 48206 22822 48258 22874
rect 4068 22720 4120 22772
rect 5540 22720 5592 22772
rect 11060 22720 11112 22772
rect 12256 22763 12308 22772
rect 12256 22729 12265 22763
rect 12265 22729 12299 22763
rect 12299 22729 12308 22763
rect 12256 22720 12308 22729
rect 12716 22720 12768 22772
rect 13544 22720 13596 22772
rect 17408 22720 17460 22772
rect 20444 22720 20496 22772
rect 15292 22652 15344 22704
rect 2872 22516 2924 22568
rect 4804 22627 4856 22636
rect 4804 22593 4813 22627
rect 4813 22593 4847 22627
rect 4847 22593 4856 22627
rect 4804 22584 4856 22593
rect 4988 22516 5040 22568
rect 7472 22627 7524 22636
rect 7472 22593 7481 22627
rect 7481 22593 7515 22627
rect 7515 22593 7524 22627
rect 7472 22584 7524 22593
rect 7656 22516 7708 22568
rect 4160 22491 4212 22500
rect 4160 22457 4169 22491
rect 4169 22457 4203 22491
rect 4203 22457 4212 22491
rect 4160 22448 4212 22457
rect 9128 22448 9180 22500
rect 11704 22584 11756 22636
rect 12716 22584 12768 22636
rect 14648 22584 14700 22636
rect 16672 22584 16724 22636
rect 17040 22652 17092 22704
rect 18788 22652 18840 22704
rect 21088 22652 21140 22704
rect 22284 22695 22336 22704
rect 22284 22661 22293 22695
rect 22293 22661 22327 22695
rect 22327 22661 22336 22695
rect 22284 22652 22336 22661
rect 24216 22720 24268 22772
rect 24308 22720 24360 22772
rect 24860 22720 24912 22772
rect 27804 22720 27856 22772
rect 25044 22652 25096 22704
rect 25136 22695 25188 22704
rect 25136 22661 25145 22695
rect 25145 22661 25179 22695
rect 25179 22661 25188 22695
rect 25136 22652 25188 22661
rect 26424 22652 26476 22704
rect 27528 22652 27580 22704
rect 28356 22652 28408 22704
rect 30748 22763 30800 22772
rect 30748 22729 30757 22763
rect 30757 22729 30791 22763
rect 30791 22729 30800 22763
rect 30748 22720 30800 22729
rect 31208 22720 31260 22772
rect 31392 22720 31444 22772
rect 31484 22763 31536 22772
rect 31484 22729 31493 22763
rect 31493 22729 31527 22763
rect 31527 22729 31536 22763
rect 31484 22720 31536 22729
rect 31576 22652 31628 22704
rect 18236 22584 18288 22636
rect 19340 22584 19392 22636
rect 10232 22559 10284 22568
rect 10232 22525 10241 22559
rect 10241 22525 10275 22559
rect 10275 22525 10284 22559
rect 10232 22516 10284 22525
rect 7104 22380 7156 22432
rect 8668 22380 8720 22432
rect 12256 22516 12308 22568
rect 12532 22516 12584 22568
rect 13544 22516 13596 22568
rect 14464 22516 14516 22568
rect 15108 22516 15160 22568
rect 16764 22516 16816 22568
rect 18604 22516 18656 22568
rect 14188 22380 14240 22432
rect 18696 22448 18748 22500
rect 20720 22448 20772 22500
rect 21180 22491 21232 22500
rect 21180 22457 21189 22491
rect 21189 22457 21223 22491
rect 21223 22457 21232 22491
rect 21180 22448 21232 22457
rect 20352 22380 20404 22432
rect 24860 22627 24912 22636
rect 24860 22593 24869 22627
rect 24869 22593 24903 22627
rect 24903 22593 24912 22627
rect 24860 22584 24912 22593
rect 27344 22627 27396 22636
rect 27344 22593 27353 22627
rect 27353 22593 27387 22627
rect 27387 22593 27396 22627
rect 27344 22584 27396 22593
rect 27804 22584 27856 22636
rect 29460 22584 29512 22636
rect 30656 22627 30708 22636
rect 30656 22593 30665 22627
rect 30665 22593 30699 22627
rect 30699 22593 30708 22627
rect 30656 22584 30708 22593
rect 35992 22720 36044 22772
rect 36084 22763 36136 22772
rect 36084 22729 36093 22763
rect 36093 22729 36127 22763
rect 36127 22729 36136 22763
rect 36084 22720 36136 22729
rect 38568 22720 38620 22772
rect 41236 22720 41288 22772
rect 33876 22652 33928 22704
rect 33968 22695 34020 22704
rect 33968 22661 33977 22695
rect 33977 22661 34011 22695
rect 34011 22661 34020 22695
rect 33968 22652 34020 22661
rect 34428 22652 34480 22704
rect 21548 22516 21600 22568
rect 23480 22516 23532 22568
rect 24492 22516 24544 22568
rect 27528 22516 27580 22568
rect 28356 22559 28408 22568
rect 28356 22525 28365 22559
rect 28365 22525 28399 22559
rect 28399 22525 28408 22559
rect 28356 22516 28408 22525
rect 28448 22516 28500 22568
rect 33692 22627 33744 22636
rect 33692 22593 33701 22627
rect 33701 22593 33735 22627
rect 33735 22593 33744 22627
rect 33692 22584 33744 22593
rect 35992 22584 36044 22636
rect 36820 22584 36872 22636
rect 24584 22448 24636 22500
rect 27160 22491 27212 22500
rect 27160 22457 27169 22491
rect 27169 22457 27203 22491
rect 27203 22457 27212 22491
rect 27160 22448 27212 22457
rect 29368 22448 29420 22500
rect 22468 22380 22520 22432
rect 26608 22423 26660 22432
rect 26608 22389 26617 22423
rect 26617 22389 26651 22423
rect 26651 22389 26660 22423
rect 26608 22380 26660 22389
rect 28908 22380 28960 22432
rect 29920 22380 29972 22432
rect 31852 22380 31904 22432
rect 32864 22380 32916 22432
rect 33600 22380 33652 22432
rect 34336 22516 34388 22568
rect 37832 22652 37884 22704
rect 39580 22652 39632 22704
rect 41972 22720 42024 22772
rect 42248 22720 42300 22772
rect 42892 22720 42944 22772
rect 44548 22763 44600 22772
rect 44548 22729 44557 22763
rect 44557 22729 44591 22763
rect 44591 22729 44600 22763
rect 44548 22720 44600 22729
rect 47308 22720 47360 22772
rect 47860 22720 47912 22772
rect 48412 22720 48464 22772
rect 37280 22584 37332 22636
rect 39488 22584 39540 22636
rect 40040 22627 40092 22636
rect 40040 22593 40049 22627
rect 40049 22593 40083 22627
rect 40083 22593 40092 22627
rect 40040 22584 40092 22593
rect 41420 22652 41472 22704
rect 41696 22627 41748 22636
rect 41696 22593 41705 22627
rect 41705 22593 41739 22627
rect 41739 22593 41748 22627
rect 41696 22584 41748 22593
rect 42064 22652 42116 22704
rect 43720 22652 43772 22704
rect 42248 22584 42300 22636
rect 42800 22627 42852 22636
rect 42800 22593 42809 22627
rect 42809 22593 42843 22627
rect 42843 22593 42852 22627
rect 42800 22584 42852 22593
rect 37740 22559 37792 22568
rect 37740 22525 37749 22559
rect 37749 22525 37783 22559
rect 37783 22525 37792 22559
rect 37740 22516 37792 22525
rect 37832 22516 37884 22568
rect 37464 22448 37516 22500
rect 40132 22559 40184 22568
rect 40132 22525 40141 22559
rect 40141 22525 40175 22559
rect 40175 22525 40184 22559
rect 40132 22516 40184 22525
rect 40868 22516 40920 22568
rect 43352 22516 43404 22568
rect 46664 22584 46716 22636
rect 47584 22584 47636 22636
rect 49056 22627 49108 22636
rect 49056 22593 49065 22627
rect 49065 22593 49099 22627
rect 49099 22593 49108 22627
rect 49056 22584 49108 22593
rect 35348 22380 35400 22432
rect 35532 22380 35584 22432
rect 37740 22380 37792 22432
rect 39488 22380 39540 22432
rect 39672 22423 39724 22432
rect 39672 22389 39681 22423
rect 39681 22389 39715 22423
rect 39715 22389 39724 22423
rect 39672 22380 39724 22389
rect 39856 22380 39908 22432
rect 40960 22380 41012 22432
rect 41512 22423 41564 22432
rect 41512 22389 41521 22423
rect 41521 22389 41555 22423
rect 41555 22389 41564 22423
rect 41512 22380 41564 22389
rect 42156 22423 42208 22432
rect 42156 22389 42165 22423
rect 42165 22389 42199 22423
rect 42199 22389 42208 22423
rect 42156 22380 42208 22389
rect 42616 22491 42668 22500
rect 42616 22457 42625 22491
rect 42625 22457 42659 22491
rect 42659 22457 42668 22491
rect 42616 22448 42668 22457
rect 44180 22448 44232 22500
rect 42800 22380 42852 22432
rect 43904 22423 43956 22432
rect 43904 22389 43913 22423
rect 43913 22389 43947 22423
rect 43947 22389 43956 22423
rect 43904 22380 43956 22389
rect 48596 22380 48648 22432
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 32950 22278 33002 22330
rect 33014 22278 33066 22330
rect 33078 22278 33130 22330
rect 33142 22278 33194 22330
rect 33206 22278 33258 22330
rect 42950 22278 43002 22330
rect 43014 22278 43066 22330
rect 43078 22278 43130 22330
rect 43142 22278 43194 22330
rect 43206 22278 43258 22330
rect 2228 22176 2280 22228
rect 4896 22176 4948 22228
rect 6920 22176 6972 22228
rect 8392 22219 8444 22228
rect 8392 22185 8401 22219
rect 8401 22185 8435 22219
rect 8435 22185 8444 22219
rect 8392 22176 8444 22185
rect 12348 22219 12400 22228
rect 12348 22185 12357 22219
rect 12357 22185 12391 22219
rect 12391 22185 12400 22219
rect 12348 22176 12400 22185
rect 3976 22108 4028 22160
rect 1308 22040 1360 22092
rect 3884 22040 3936 22092
rect 11152 22108 11204 22160
rect 4068 22015 4120 22024
rect 4068 21981 4077 22015
rect 4077 21981 4111 22015
rect 4111 21981 4120 22015
rect 4068 21972 4120 21981
rect 6460 21972 6512 22024
rect 9128 22015 9180 22024
rect 9128 21981 9137 22015
rect 9137 21981 9171 22015
rect 9171 21981 9180 22015
rect 9128 21972 9180 21981
rect 10048 22083 10100 22092
rect 10048 22049 10057 22083
rect 10057 22049 10091 22083
rect 10091 22049 10100 22083
rect 10048 22040 10100 22049
rect 11060 22083 11112 22092
rect 11060 22049 11069 22083
rect 11069 22049 11103 22083
rect 11103 22049 11112 22083
rect 11060 22040 11112 22049
rect 16764 22176 16816 22228
rect 17040 22176 17092 22228
rect 18604 22176 18656 22228
rect 18696 22176 18748 22228
rect 22192 22176 22244 22228
rect 23756 22176 23808 22228
rect 24400 22176 24452 22228
rect 27804 22176 27856 22228
rect 28356 22176 28408 22228
rect 29000 22176 29052 22228
rect 29368 22176 29420 22228
rect 29460 22176 29512 22228
rect 31576 22176 31628 22228
rect 32588 22219 32640 22228
rect 32588 22185 32597 22219
rect 32597 22185 32631 22219
rect 32631 22185 32640 22219
rect 32588 22176 32640 22185
rect 33324 22176 33376 22228
rect 37188 22176 37240 22228
rect 37556 22219 37608 22228
rect 37556 22185 37586 22219
rect 37586 22185 37608 22219
rect 37556 22176 37608 22185
rect 40040 22176 40092 22228
rect 41696 22176 41748 22228
rect 42708 22176 42760 22228
rect 43352 22176 43404 22228
rect 43720 22219 43772 22228
rect 43720 22185 43729 22219
rect 43729 22185 43763 22219
rect 43763 22185 43772 22219
rect 43720 22176 43772 22185
rect 49332 22176 49384 22228
rect 17224 22108 17276 22160
rect 13728 22040 13780 22092
rect 16120 22040 16172 22092
rect 16488 22040 16540 22092
rect 18972 22108 19024 22160
rect 21456 22108 21508 22160
rect 11152 21904 11204 21956
rect 11336 22015 11388 22024
rect 11336 21981 11345 22015
rect 11345 21981 11379 22015
rect 11379 21981 11388 22015
rect 11336 21972 11388 21981
rect 12532 22015 12584 22024
rect 12532 21981 12541 22015
rect 12541 21981 12575 22015
rect 12575 21981 12584 22015
rect 12532 21972 12584 21981
rect 15200 22015 15252 22024
rect 15200 21981 15209 22015
rect 15209 21981 15243 22015
rect 15243 21981 15252 22015
rect 15200 21972 15252 21981
rect 12716 21904 12768 21956
rect 14740 21904 14792 21956
rect 16764 21904 16816 21956
rect 9680 21836 9732 21888
rect 9864 21836 9916 21888
rect 16488 21836 16540 21888
rect 20720 22040 20772 22092
rect 21088 22083 21140 22092
rect 21088 22049 21097 22083
rect 21097 22049 21131 22083
rect 21131 22049 21140 22083
rect 21088 22040 21140 22049
rect 23204 22083 23256 22092
rect 23204 22049 23213 22083
rect 23213 22049 23247 22083
rect 23247 22049 23256 22083
rect 23204 22040 23256 22049
rect 23572 22040 23624 22092
rect 24584 22040 24636 22092
rect 25136 22083 25188 22092
rect 25136 22049 25145 22083
rect 25145 22049 25179 22083
rect 25179 22049 25188 22083
rect 25136 22040 25188 22049
rect 26424 22040 26476 22092
rect 26608 22108 26660 22160
rect 27068 22108 27120 22160
rect 27252 22040 27304 22092
rect 17684 21972 17736 22024
rect 18236 21972 18288 22024
rect 19432 22015 19484 22024
rect 19432 21981 19441 22015
rect 19441 21981 19475 22015
rect 19475 21981 19484 22015
rect 19432 21972 19484 21981
rect 21916 21972 21968 22024
rect 23756 21972 23808 22024
rect 24952 21972 25004 22024
rect 25320 21972 25372 22024
rect 28540 22040 28592 22092
rect 28908 22083 28960 22092
rect 28908 22049 28917 22083
rect 28917 22049 28951 22083
rect 28951 22049 28960 22083
rect 28908 22040 28960 22049
rect 30380 22040 30432 22092
rect 31208 22040 31260 22092
rect 32312 22040 32364 22092
rect 34336 22108 34388 22160
rect 34428 22151 34480 22160
rect 34428 22117 34437 22151
rect 34437 22117 34471 22151
rect 34471 22117 34480 22151
rect 34428 22108 34480 22117
rect 35716 22108 35768 22160
rect 38844 22108 38896 22160
rect 34152 22083 34204 22092
rect 34152 22049 34161 22083
rect 34161 22049 34195 22083
rect 34195 22049 34204 22083
rect 34152 22040 34204 22049
rect 30564 21972 30616 22024
rect 33048 21972 33100 22024
rect 35072 22040 35124 22092
rect 35624 22040 35676 22092
rect 34428 21972 34480 22024
rect 36084 21972 36136 22024
rect 36636 21972 36688 22024
rect 37280 22083 37332 22092
rect 37280 22049 37289 22083
rect 37289 22049 37323 22083
rect 37323 22049 37332 22083
rect 37280 22040 37332 22049
rect 37648 22040 37700 22092
rect 38292 22040 38344 22092
rect 40776 22108 40828 22160
rect 42432 22151 42484 22160
rect 42432 22117 42441 22151
rect 42441 22117 42475 22151
rect 42475 22117 42484 22151
rect 42432 22108 42484 22117
rect 41604 22040 41656 22092
rect 42064 22040 42116 22092
rect 49240 22040 49292 22092
rect 24768 21904 24820 21956
rect 21916 21879 21968 21888
rect 21916 21845 21925 21879
rect 21925 21845 21959 21879
rect 21959 21845 21968 21879
rect 21916 21836 21968 21845
rect 22652 21879 22704 21888
rect 22652 21845 22661 21879
rect 22661 21845 22695 21879
rect 22695 21845 22704 21879
rect 22652 21836 22704 21845
rect 23572 21836 23624 21888
rect 23848 21836 23900 21888
rect 24860 21836 24912 21888
rect 25780 21904 25832 21956
rect 26148 21904 26200 21956
rect 29828 21904 29880 21956
rect 30748 21904 30800 21956
rect 31392 21904 31444 21956
rect 31576 21904 31628 21956
rect 25044 21879 25096 21888
rect 25044 21845 25053 21879
rect 25053 21845 25087 21879
rect 25087 21845 25096 21879
rect 25044 21836 25096 21845
rect 25964 21879 26016 21888
rect 25964 21845 25973 21879
rect 25973 21845 26007 21879
rect 26007 21845 26016 21879
rect 25964 21836 26016 21845
rect 26516 21836 26568 21888
rect 27436 21836 27488 21888
rect 27620 21836 27672 21888
rect 31852 21836 31904 21888
rect 32680 21836 32732 21888
rect 33416 21879 33468 21888
rect 33416 21845 33425 21879
rect 33425 21845 33459 21879
rect 33459 21845 33468 21879
rect 33416 21836 33468 21845
rect 33508 21879 33560 21888
rect 33508 21845 33517 21879
rect 33517 21845 33551 21879
rect 33551 21845 33560 21879
rect 33508 21836 33560 21845
rect 36360 21904 36412 21956
rect 35164 21836 35216 21888
rect 35532 21836 35584 21888
rect 36176 21836 36228 21888
rect 37280 21904 37332 21956
rect 38844 21904 38896 21956
rect 39580 21947 39632 21956
rect 39580 21913 39589 21947
rect 39589 21913 39623 21947
rect 39623 21913 39632 21947
rect 39580 21904 39632 21913
rect 41420 21904 41472 21956
rect 38568 21836 38620 21888
rect 40040 21879 40092 21888
rect 40040 21845 40049 21879
rect 40049 21845 40083 21879
rect 40083 21845 40092 21879
rect 40040 21836 40092 21845
rect 40684 21836 40736 21888
rect 41788 21904 41840 21956
rect 41972 21972 42024 22024
rect 46572 21972 46624 22024
rect 47860 21972 47912 22024
rect 48780 21972 48832 22024
rect 45376 21904 45428 21956
rect 49148 21947 49200 21956
rect 49148 21913 49157 21947
rect 49157 21913 49191 21947
rect 49191 21913 49200 21947
rect 49148 21904 49200 21913
rect 47676 21836 47728 21888
rect 47768 21879 47820 21888
rect 47768 21845 47777 21879
rect 47777 21845 47811 21879
rect 47811 21845 47820 21879
rect 47768 21836 47820 21845
rect 48412 21879 48464 21888
rect 48412 21845 48421 21879
rect 48421 21845 48455 21879
rect 48455 21845 48464 21879
rect 48412 21836 48464 21845
rect 48504 21836 48556 21888
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 27950 21734 28002 21786
rect 28014 21734 28066 21786
rect 28078 21734 28130 21786
rect 28142 21734 28194 21786
rect 28206 21734 28258 21786
rect 37950 21734 38002 21786
rect 38014 21734 38066 21786
rect 38078 21734 38130 21786
rect 38142 21734 38194 21786
rect 38206 21734 38258 21786
rect 47950 21734 48002 21786
rect 48014 21734 48066 21786
rect 48078 21734 48130 21786
rect 48142 21734 48194 21786
rect 48206 21734 48258 21786
rect 4068 21632 4120 21684
rect 4344 21607 4396 21616
rect 4344 21573 4353 21607
rect 4353 21573 4387 21607
rect 4387 21573 4396 21607
rect 4344 21564 4396 21573
rect 9772 21632 9824 21684
rect 12624 21632 12676 21684
rect 13912 21675 13964 21684
rect 13912 21641 13921 21675
rect 13921 21641 13955 21675
rect 13955 21641 13964 21675
rect 13912 21632 13964 21641
rect 10048 21564 10100 21616
rect 3332 21428 3384 21480
rect 3608 21539 3660 21548
rect 3608 21505 3617 21539
rect 3617 21505 3651 21539
rect 3651 21505 3660 21539
rect 3608 21496 3660 21505
rect 5908 21539 5960 21548
rect 5908 21505 5917 21539
rect 5917 21505 5951 21539
rect 5951 21505 5960 21539
rect 5908 21496 5960 21505
rect 5264 21428 5316 21480
rect 8576 21539 8628 21548
rect 8576 21505 8585 21539
rect 8585 21505 8619 21539
rect 8619 21505 8628 21539
rect 8576 21496 8628 21505
rect 6736 21428 6788 21480
rect 8852 21471 8904 21480
rect 8852 21437 8861 21471
rect 8861 21437 8895 21471
rect 8895 21437 8904 21471
rect 8852 21428 8904 21437
rect 11980 21496 12032 21548
rect 12808 21539 12860 21548
rect 12808 21505 12817 21539
rect 12817 21505 12851 21539
rect 12851 21505 12860 21539
rect 12808 21496 12860 21505
rect 14004 21496 14056 21548
rect 13452 21428 13504 21480
rect 14280 21496 14332 21548
rect 17040 21632 17092 21684
rect 14832 21607 14884 21616
rect 14832 21573 14841 21607
rect 14841 21573 14875 21607
rect 14875 21573 14884 21607
rect 14832 21564 14884 21573
rect 16764 21607 16816 21616
rect 16764 21573 16773 21607
rect 16773 21573 16807 21607
rect 16807 21573 16816 21607
rect 16764 21564 16816 21573
rect 17684 21632 17736 21684
rect 17868 21675 17920 21684
rect 17868 21641 17877 21675
rect 17877 21641 17911 21675
rect 17911 21641 17920 21675
rect 17868 21632 17920 21641
rect 18328 21496 18380 21548
rect 16120 21428 16172 21480
rect 20536 21632 20588 21684
rect 21916 21632 21968 21684
rect 22284 21632 22336 21684
rect 20720 21564 20772 21616
rect 18604 21471 18656 21480
rect 18604 21437 18613 21471
rect 18613 21437 18647 21471
rect 18647 21437 18656 21471
rect 18604 21428 18656 21437
rect 18880 21471 18932 21480
rect 18880 21437 18889 21471
rect 18889 21437 18923 21471
rect 18923 21437 18932 21471
rect 18880 21428 18932 21437
rect 27804 21632 27856 21684
rect 32404 21632 32456 21684
rect 33416 21632 33468 21684
rect 22744 21607 22796 21616
rect 22744 21573 22753 21607
rect 22753 21573 22787 21607
rect 22787 21573 22796 21607
rect 22744 21564 22796 21573
rect 23204 21564 23256 21616
rect 25044 21564 25096 21616
rect 26976 21564 27028 21616
rect 25872 21496 25924 21548
rect 26884 21496 26936 21548
rect 22468 21471 22520 21480
rect 22468 21437 22477 21471
rect 22477 21437 22511 21471
rect 22511 21437 22520 21471
rect 22468 21428 22520 21437
rect 5632 21360 5684 21412
rect 8576 21360 8628 21412
rect 4344 21292 4396 21344
rect 8760 21292 8812 21344
rect 9956 21292 10008 21344
rect 11888 21292 11940 21344
rect 16304 21335 16356 21344
rect 16304 21301 16313 21335
rect 16313 21301 16347 21335
rect 16347 21301 16356 21335
rect 16304 21292 16356 21301
rect 18696 21292 18748 21344
rect 22284 21360 22336 21412
rect 24768 21403 24820 21412
rect 24768 21369 24777 21403
rect 24777 21369 24811 21403
rect 24811 21369 24820 21403
rect 24768 21360 24820 21369
rect 25228 21471 25280 21480
rect 25228 21437 25237 21471
rect 25237 21437 25271 21471
rect 25271 21437 25280 21471
rect 25228 21428 25280 21437
rect 25320 21428 25372 21480
rect 27436 21564 27488 21616
rect 27712 21564 27764 21616
rect 29828 21564 29880 21616
rect 31208 21607 31260 21616
rect 31208 21573 31217 21607
rect 31217 21573 31251 21607
rect 31251 21573 31260 21607
rect 31208 21564 31260 21573
rect 31576 21564 31628 21616
rect 32864 21564 32916 21616
rect 34888 21675 34940 21684
rect 34888 21641 34897 21675
rect 34897 21641 34931 21675
rect 34931 21641 34940 21675
rect 34888 21632 34940 21641
rect 35072 21632 35124 21684
rect 35900 21632 35952 21684
rect 40040 21632 40092 21684
rect 40132 21632 40184 21684
rect 40408 21632 40460 21684
rect 36452 21564 36504 21616
rect 36636 21564 36688 21616
rect 38384 21564 38436 21616
rect 38844 21564 38896 21616
rect 39856 21564 39908 21616
rect 28724 21539 28776 21548
rect 28724 21505 28733 21539
rect 28733 21505 28767 21539
rect 28767 21505 28776 21539
rect 28724 21496 28776 21505
rect 28816 21539 28868 21548
rect 28816 21505 28825 21539
rect 28825 21505 28859 21539
rect 28859 21505 28868 21539
rect 28816 21496 28868 21505
rect 28908 21471 28960 21480
rect 28908 21437 28917 21471
rect 28917 21437 28951 21471
rect 28951 21437 28960 21471
rect 28908 21428 28960 21437
rect 29276 21428 29328 21480
rect 29092 21360 29144 21412
rect 29920 21360 29972 21412
rect 20352 21335 20404 21344
rect 20352 21301 20361 21335
rect 20361 21301 20395 21335
rect 20395 21301 20404 21335
rect 20352 21292 20404 21301
rect 20720 21335 20772 21344
rect 20720 21301 20729 21335
rect 20729 21301 20763 21335
rect 20763 21301 20772 21335
rect 21916 21335 21968 21344
rect 20720 21292 20772 21301
rect 21916 21301 21925 21335
rect 21925 21301 21959 21335
rect 21959 21301 21968 21335
rect 21916 21292 21968 21301
rect 23204 21292 23256 21344
rect 25412 21292 25464 21344
rect 25872 21335 25924 21344
rect 25872 21301 25881 21335
rect 25881 21301 25915 21335
rect 25915 21301 25924 21335
rect 25872 21292 25924 21301
rect 26148 21292 26200 21344
rect 26332 21292 26384 21344
rect 29552 21335 29604 21344
rect 29552 21301 29561 21335
rect 29561 21301 29595 21335
rect 29595 21301 29604 21335
rect 29552 21292 29604 21301
rect 30656 21292 30708 21344
rect 33600 21539 33652 21548
rect 33600 21505 33609 21539
rect 33609 21505 33643 21539
rect 33643 21505 33652 21539
rect 33600 21496 33652 21505
rect 33692 21539 33744 21548
rect 33692 21505 33701 21539
rect 33701 21505 33735 21539
rect 33735 21505 33744 21539
rect 33692 21496 33744 21505
rect 34796 21539 34848 21548
rect 34796 21505 34805 21539
rect 34805 21505 34839 21539
rect 34839 21505 34848 21539
rect 34796 21496 34848 21505
rect 31576 21428 31628 21480
rect 33416 21428 33468 21480
rect 36728 21496 36780 21548
rect 36176 21471 36228 21480
rect 36176 21437 36185 21471
rect 36185 21437 36219 21471
rect 36219 21437 36228 21471
rect 36176 21428 36228 21437
rect 36636 21428 36688 21480
rect 37740 21428 37792 21480
rect 38292 21471 38344 21480
rect 36360 21360 36412 21412
rect 37464 21360 37516 21412
rect 38292 21437 38301 21471
rect 38301 21437 38335 21471
rect 38335 21437 38344 21471
rect 38292 21428 38344 21437
rect 38384 21428 38436 21480
rect 41236 21564 41288 21616
rect 41788 21564 41840 21616
rect 42248 21632 42300 21684
rect 42892 21632 42944 21684
rect 43996 21632 44048 21684
rect 47492 21632 47544 21684
rect 48780 21675 48832 21684
rect 48780 21641 48789 21675
rect 48789 21641 48823 21675
rect 48823 21641 48832 21675
rect 48780 21632 48832 21641
rect 49056 21632 49108 21684
rect 47768 21564 47820 21616
rect 40868 21496 40920 21548
rect 47860 21496 47912 21548
rect 49056 21539 49108 21548
rect 49056 21505 49065 21539
rect 49065 21505 49099 21539
rect 49099 21505 49108 21539
rect 49056 21496 49108 21505
rect 40776 21471 40828 21480
rect 40776 21437 40785 21471
rect 40785 21437 40819 21471
rect 40819 21437 40828 21471
rect 40776 21428 40828 21437
rect 40040 21360 40092 21412
rect 40500 21360 40552 21412
rect 32680 21292 32732 21344
rect 34336 21292 34388 21344
rect 34520 21292 34572 21344
rect 37280 21292 37332 21344
rect 39764 21335 39816 21344
rect 39764 21301 39773 21335
rect 39773 21301 39807 21335
rect 39807 21301 39816 21335
rect 39764 21292 39816 21301
rect 39856 21292 39908 21344
rect 41420 21403 41472 21412
rect 41420 21369 41429 21403
rect 41429 21369 41463 21403
rect 41463 21369 41472 21403
rect 41420 21360 41472 21369
rect 41788 21428 41840 21480
rect 42892 21428 42944 21480
rect 46204 21360 46256 21412
rect 49240 21335 49292 21344
rect 49240 21301 49249 21335
rect 49249 21301 49283 21335
rect 49283 21301 49292 21335
rect 49240 21292 49292 21301
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 32950 21190 33002 21242
rect 33014 21190 33066 21242
rect 33078 21190 33130 21242
rect 33142 21190 33194 21242
rect 33206 21190 33258 21242
rect 42950 21190 43002 21242
rect 43014 21190 43066 21242
rect 43078 21190 43130 21242
rect 43142 21190 43194 21242
rect 43206 21190 43258 21242
rect 4252 20952 4304 21004
rect 5540 20952 5592 21004
rect 4344 20884 4396 20936
rect 2780 20859 2832 20868
rect 2780 20825 2789 20859
rect 2789 20825 2823 20859
rect 2823 20825 2832 20859
rect 2780 20816 2832 20825
rect 7748 21088 7800 21140
rect 6460 21020 6512 21072
rect 12440 21088 12492 21140
rect 12992 21088 13044 21140
rect 16580 21088 16632 21140
rect 18972 21088 19024 21140
rect 19156 21088 19208 21140
rect 20720 21088 20772 21140
rect 21272 21088 21324 21140
rect 21548 21088 21600 21140
rect 22652 21088 22704 21140
rect 22836 21088 22888 21140
rect 24676 21088 24728 21140
rect 26700 21131 26752 21140
rect 26700 21097 26709 21131
rect 26709 21097 26743 21131
rect 26743 21097 26752 21131
rect 26700 21088 26752 21097
rect 27160 21088 27212 21140
rect 27804 21088 27856 21140
rect 30104 21088 30156 21140
rect 30380 21088 30432 21140
rect 31392 21088 31444 21140
rect 10508 21020 10560 21072
rect 11796 20952 11848 21004
rect 9864 20927 9916 20936
rect 9864 20893 9873 20927
rect 9873 20893 9907 20927
rect 9907 20893 9916 20927
rect 9864 20884 9916 20893
rect 11244 20884 11296 20936
rect 11336 20927 11388 20936
rect 11336 20893 11345 20927
rect 11345 20893 11379 20927
rect 11379 20893 11388 20927
rect 11336 20884 11388 20893
rect 12808 21020 12860 21072
rect 13728 21020 13780 21072
rect 13636 20952 13688 21004
rect 23848 21020 23900 21072
rect 20444 20952 20496 21004
rect 12072 20816 12124 20868
rect 12808 20859 12860 20868
rect 12808 20825 12817 20859
rect 12817 20825 12851 20859
rect 12851 20825 12860 20859
rect 12808 20816 12860 20825
rect 11060 20748 11112 20800
rect 12440 20791 12492 20800
rect 12440 20757 12449 20791
rect 12449 20757 12483 20791
rect 12483 20757 12492 20791
rect 12440 20748 12492 20757
rect 12992 20748 13044 20800
rect 14280 20927 14332 20936
rect 14280 20893 14289 20927
rect 14289 20893 14323 20927
rect 14323 20893 14332 20927
rect 14280 20884 14332 20893
rect 17040 20884 17092 20936
rect 21088 20884 21140 20936
rect 21180 20927 21232 20936
rect 21180 20893 21189 20927
rect 21189 20893 21223 20927
rect 21223 20893 21232 20927
rect 21180 20884 21232 20893
rect 25596 20952 25648 21004
rect 29552 21020 29604 21072
rect 24124 20884 24176 20936
rect 25780 20884 25832 20936
rect 28724 20952 28776 21004
rect 30472 21020 30524 21072
rect 30840 21063 30892 21072
rect 30840 21029 30849 21063
rect 30849 21029 30883 21063
rect 30883 21029 30892 21063
rect 30840 21020 30892 21029
rect 34520 21088 34572 21140
rect 30196 20995 30248 21004
rect 27344 20884 27396 20936
rect 28632 20884 28684 20936
rect 28816 20884 28868 20936
rect 30196 20961 30205 20995
rect 30205 20961 30239 20995
rect 30239 20961 30248 20995
rect 30196 20952 30248 20961
rect 34336 21020 34388 21072
rect 39948 21088 40000 21140
rect 40224 21088 40276 21140
rect 40316 21088 40368 21140
rect 41052 21088 41104 21140
rect 39120 21020 39172 21072
rect 34060 20952 34112 21004
rect 35716 20952 35768 21004
rect 35808 20952 35860 21004
rect 37004 20952 37056 21004
rect 37280 20952 37332 21004
rect 38292 20952 38344 21004
rect 39764 21020 39816 21072
rect 42156 21020 42208 21072
rect 30288 20884 30340 20936
rect 30564 20884 30616 20936
rect 14556 20859 14608 20868
rect 14556 20825 14565 20859
rect 14565 20825 14599 20859
rect 14599 20825 14608 20859
rect 14556 20816 14608 20825
rect 16764 20816 16816 20868
rect 19156 20816 19208 20868
rect 21548 20816 21600 20868
rect 21916 20816 21968 20868
rect 14832 20748 14884 20800
rect 17776 20748 17828 20800
rect 18788 20748 18840 20800
rect 25964 20816 26016 20868
rect 26792 20816 26844 20868
rect 27160 20816 27212 20868
rect 29276 20816 29328 20868
rect 30104 20816 30156 20868
rect 24032 20748 24084 20800
rect 28632 20748 28684 20800
rect 28724 20791 28776 20800
rect 28724 20757 28733 20791
rect 28733 20757 28767 20791
rect 28767 20757 28776 20791
rect 28724 20748 28776 20757
rect 28816 20791 28868 20800
rect 28816 20757 28825 20791
rect 28825 20757 28859 20791
rect 28859 20757 28868 20791
rect 28816 20748 28868 20757
rect 29368 20748 29420 20800
rect 29552 20748 29604 20800
rect 29736 20791 29788 20800
rect 29736 20757 29745 20791
rect 29745 20757 29779 20791
rect 29779 20757 29788 20791
rect 29736 20748 29788 20757
rect 32312 20884 32364 20936
rect 37648 20927 37700 20936
rect 37648 20893 37657 20927
rect 37657 20893 37691 20927
rect 37691 20893 37700 20927
rect 37648 20884 37700 20893
rect 48412 20884 48464 20936
rect 49056 20927 49108 20936
rect 49056 20893 49065 20927
rect 49065 20893 49099 20927
rect 49099 20893 49108 20927
rect 49056 20884 49108 20893
rect 31392 20816 31444 20868
rect 32772 20816 32824 20868
rect 32864 20816 32916 20868
rect 33232 20816 33284 20868
rect 35072 20816 35124 20868
rect 35256 20816 35308 20868
rect 35808 20816 35860 20868
rect 38660 20816 38712 20868
rect 34244 20791 34296 20800
rect 34244 20757 34253 20791
rect 34253 20757 34287 20791
rect 34287 20757 34296 20791
rect 34244 20748 34296 20757
rect 34704 20748 34756 20800
rect 36176 20748 36228 20800
rect 36636 20791 36688 20800
rect 36636 20757 36645 20791
rect 36645 20757 36679 20791
rect 36679 20757 36688 20791
rect 36636 20748 36688 20757
rect 38292 20748 38344 20800
rect 41420 20816 41472 20868
rect 42156 20816 42208 20868
rect 48964 20748 49016 20800
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 27950 20646 28002 20698
rect 28014 20646 28066 20698
rect 28078 20646 28130 20698
rect 28142 20646 28194 20698
rect 28206 20646 28258 20698
rect 37950 20646 38002 20698
rect 38014 20646 38066 20698
rect 38078 20646 38130 20698
rect 38142 20646 38194 20698
rect 38206 20646 38258 20698
rect 47950 20646 48002 20698
rect 48014 20646 48066 20698
rect 48078 20646 48130 20698
rect 48142 20646 48194 20698
rect 48206 20646 48258 20698
rect 5264 20587 5316 20596
rect 5264 20553 5273 20587
rect 5273 20553 5307 20587
rect 5307 20553 5316 20587
rect 5264 20544 5316 20553
rect 9680 20587 9732 20596
rect 9680 20553 9689 20587
rect 9689 20553 9723 20587
rect 9723 20553 9732 20587
rect 9680 20544 9732 20553
rect 10324 20587 10376 20596
rect 10324 20553 10333 20587
rect 10333 20553 10367 20587
rect 10367 20553 10376 20587
rect 10324 20544 10376 20553
rect 1952 20408 2004 20460
rect 2872 20340 2924 20392
rect 3884 20383 3936 20392
rect 3884 20349 3893 20383
rect 3893 20349 3927 20383
rect 3927 20349 3936 20383
rect 3884 20340 3936 20349
rect 8392 20476 8444 20528
rect 11888 20544 11940 20596
rect 10600 20476 10652 20528
rect 13360 20544 13412 20596
rect 13636 20544 13688 20596
rect 14924 20587 14976 20596
rect 14924 20553 14933 20587
rect 14933 20553 14967 20587
rect 14967 20553 14976 20587
rect 14924 20544 14976 20553
rect 15108 20544 15160 20596
rect 15384 20544 15436 20596
rect 15844 20544 15896 20596
rect 16028 20587 16080 20596
rect 16028 20553 16037 20587
rect 16037 20553 16071 20587
rect 16071 20553 16080 20587
rect 16028 20544 16080 20553
rect 4160 20340 4212 20392
rect 6644 20340 6696 20392
rect 11428 20408 11480 20460
rect 10416 20340 10468 20392
rect 10968 20383 11020 20392
rect 10968 20349 10977 20383
rect 10977 20349 11011 20383
rect 11011 20349 11020 20383
rect 10968 20340 11020 20349
rect 11888 20408 11940 20460
rect 12716 20519 12768 20528
rect 12716 20485 12725 20519
rect 12725 20485 12759 20519
rect 12759 20485 12768 20519
rect 12716 20476 12768 20485
rect 13268 20519 13320 20528
rect 13268 20485 13277 20519
rect 13277 20485 13311 20519
rect 13311 20485 13320 20519
rect 18880 20544 18932 20596
rect 19156 20587 19208 20596
rect 19156 20553 19165 20587
rect 19165 20553 19199 20587
rect 19199 20553 19208 20587
rect 19156 20544 19208 20553
rect 13268 20476 13320 20485
rect 14924 20408 14976 20460
rect 10876 20272 10928 20324
rect 1768 20204 1820 20256
rect 4804 20204 4856 20256
rect 4988 20204 5040 20256
rect 10048 20204 10100 20256
rect 14832 20340 14884 20392
rect 19340 20476 19392 20528
rect 15936 20408 15988 20460
rect 19156 20408 19208 20460
rect 20260 20544 20312 20596
rect 22468 20544 22520 20596
rect 22744 20544 22796 20596
rect 22836 20544 22888 20596
rect 19984 20519 20036 20528
rect 19984 20485 19993 20519
rect 19993 20485 20027 20519
rect 20027 20485 20036 20519
rect 19984 20476 20036 20485
rect 21272 20476 21324 20528
rect 21548 20408 21600 20460
rect 15476 20340 15528 20392
rect 16212 20383 16264 20392
rect 16212 20349 16221 20383
rect 16221 20349 16255 20383
rect 16255 20349 16264 20383
rect 16212 20340 16264 20349
rect 16764 20383 16816 20392
rect 16764 20349 16773 20383
rect 16773 20349 16807 20383
rect 16807 20349 16816 20383
rect 16764 20340 16816 20349
rect 17040 20383 17092 20392
rect 17040 20349 17049 20383
rect 17049 20349 17083 20383
rect 17083 20349 17092 20383
rect 17040 20340 17092 20349
rect 17684 20340 17736 20392
rect 18052 20340 18104 20392
rect 18788 20340 18840 20392
rect 18972 20340 19024 20392
rect 21456 20383 21508 20392
rect 21456 20349 21465 20383
rect 21465 20349 21499 20383
rect 21499 20349 21508 20383
rect 21456 20340 21508 20349
rect 22468 20383 22520 20392
rect 22468 20349 22477 20383
rect 22477 20349 22511 20383
rect 22511 20349 22520 20383
rect 22468 20340 22520 20349
rect 23388 20451 23440 20460
rect 23388 20417 23397 20451
rect 23397 20417 23431 20451
rect 23431 20417 23440 20451
rect 23388 20408 23440 20417
rect 23480 20408 23532 20460
rect 25688 20544 25740 20596
rect 24676 20476 24728 20528
rect 25504 20476 25556 20528
rect 26884 20476 26936 20528
rect 16856 20272 16908 20324
rect 13268 20204 13320 20256
rect 13544 20204 13596 20256
rect 13820 20204 13872 20256
rect 15752 20204 15804 20256
rect 22192 20272 22244 20324
rect 23756 20340 23808 20392
rect 24492 20340 24544 20392
rect 25780 20340 25832 20392
rect 26700 20408 26752 20460
rect 32312 20544 32364 20596
rect 28264 20476 28316 20528
rect 29828 20519 29880 20528
rect 29828 20485 29837 20519
rect 29837 20485 29871 20519
rect 29871 20485 29880 20519
rect 29828 20476 29880 20485
rect 30012 20476 30064 20528
rect 31116 20519 31168 20528
rect 31116 20485 31125 20519
rect 31125 20485 31159 20519
rect 31159 20485 31168 20519
rect 31116 20476 31168 20485
rect 27160 20340 27212 20392
rect 27528 20383 27580 20392
rect 27528 20349 27537 20383
rect 27537 20349 27571 20383
rect 27571 20349 27580 20383
rect 27528 20340 27580 20349
rect 27620 20340 27672 20392
rect 30840 20408 30892 20460
rect 31668 20476 31720 20528
rect 31392 20408 31444 20460
rect 33232 20476 33284 20528
rect 34060 20587 34112 20596
rect 34060 20553 34069 20587
rect 34069 20553 34103 20587
rect 34103 20553 34112 20587
rect 34060 20544 34112 20553
rect 34704 20544 34756 20596
rect 34428 20476 34480 20528
rect 34612 20476 34664 20528
rect 29000 20383 29052 20392
rect 29000 20349 29009 20383
rect 29009 20349 29043 20383
rect 29043 20349 29052 20383
rect 29000 20340 29052 20349
rect 25412 20272 25464 20324
rect 29276 20340 29328 20392
rect 31208 20383 31260 20392
rect 31208 20349 31217 20383
rect 31217 20349 31251 20383
rect 31251 20349 31260 20383
rect 31208 20340 31260 20349
rect 32312 20383 32364 20392
rect 32312 20349 32321 20383
rect 32321 20349 32355 20383
rect 32355 20349 32364 20383
rect 32312 20340 32364 20349
rect 18788 20204 18840 20256
rect 22008 20247 22060 20256
rect 22008 20213 22017 20247
rect 22017 20213 22051 20247
rect 22051 20213 22060 20247
rect 22008 20204 22060 20213
rect 25504 20204 25556 20256
rect 26608 20247 26660 20256
rect 26608 20213 26617 20247
rect 26617 20213 26651 20247
rect 26651 20213 26660 20247
rect 26608 20204 26660 20213
rect 29000 20204 29052 20256
rect 30564 20204 30616 20256
rect 31024 20204 31076 20256
rect 31852 20315 31904 20324
rect 31852 20281 31861 20315
rect 31861 20281 31895 20315
rect 31895 20281 31904 20315
rect 31852 20272 31904 20281
rect 37372 20476 37424 20528
rect 38292 20476 38344 20528
rect 38660 20476 38712 20528
rect 40592 20544 40644 20596
rect 37188 20408 37240 20460
rect 35256 20340 35308 20392
rect 35532 20340 35584 20392
rect 35072 20272 35124 20324
rect 35256 20204 35308 20256
rect 35808 20247 35860 20256
rect 35808 20213 35817 20247
rect 35817 20213 35851 20247
rect 35851 20213 35860 20247
rect 35808 20204 35860 20213
rect 36636 20340 36688 20392
rect 37556 20340 37608 20392
rect 37740 20383 37792 20392
rect 37740 20349 37749 20383
rect 37749 20349 37783 20383
rect 37783 20349 37792 20383
rect 37740 20340 37792 20349
rect 38568 20340 38620 20392
rect 40500 20383 40552 20392
rect 40500 20349 40509 20383
rect 40509 20349 40543 20383
rect 40543 20349 40552 20383
rect 40500 20340 40552 20349
rect 39028 20272 39080 20324
rect 41328 20272 41380 20324
rect 48780 20408 48832 20460
rect 49056 20451 49108 20460
rect 49056 20417 49065 20451
rect 49065 20417 49099 20451
rect 49099 20417 49108 20451
rect 49056 20408 49108 20417
rect 38660 20204 38712 20256
rect 39212 20204 39264 20256
rect 39948 20247 40000 20256
rect 39948 20213 39957 20247
rect 39957 20213 39991 20247
rect 39991 20213 40000 20247
rect 39948 20204 40000 20213
rect 48412 20247 48464 20256
rect 48412 20213 48421 20247
rect 48421 20213 48455 20247
rect 48455 20213 48464 20247
rect 48412 20204 48464 20213
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 32950 20102 33002 20154
rect 33014 20102 33066 20154
rect 33078 20102 33130 20154
rect 33142 20102 33194 20154
rect 33206 20102 33258 20154
rect 42950 20102 43002 20154
rect 43014 20102 43066 20154
rect 43078 20102 43130 20154
rect 43142 20102 43194 20154
rect 43206 20102 43258 20154
rect 1768 19839 1820 19848
rect 1768 19805 1777 19839
rect 1777 19805 1811 19839
rect 1811 19805 1820 19839
rect 1768 19796 1820 19805
rect 7012 20000 7064 20052
rect 9956 20043 10008 20052
rect 9956 20009 9965 20043
rect 9965 20009 9999 20043
rect 9999 20009 10008 20043
rect 9956 20000 10008 20009
rect 4804 19932 4856 19984
rect 4896 19907 4948 19916
rect 4896 19873 4905 19907
rect 4905 19873 4939 19907
rect 4939 19873 4948 19907
rect 4896 19864 4948 19873
rect 6184 19864 6236 19916
rect 2780 19771 2832 19780
rect 2780 19737 2789 19771
rect 2789 19737 2823 19771
rect 2823 19737 2832 19771
rect 2780 19728 2832 19737
rect 9772 19796 9824 19848
rect 10600 19796 10652 19848
rect 7104 19728 7156 19780
rect 7840 19728 7892 19780
rect 10048 19728 10100 19780
rect 10508 19660 10560 19712
rect 10876 19932 10928 19984
rect 13912 19932 13964 19984
rect 14372 20000 14424 20052
rect 14924 20000 14976 20052
rect 18052 20000 18104 20052
rect 18328 20000 18380 20052
rect 20536 20000 20588 20052
rect 14280 19864 14332 19916
rect 14096 19796 14148 19848
rect 15568 19864 15620 19916
rect 18880 19932 18932 19984
rect 19064 19864 19116 19916
rect 19340 19907 19392 19916
rect 19340 19873 19349 19907
rect 19349 19873 19383 19907
rect 19383 19873 19392 19907
rect 19340 19864 19392 19873
rect 21180 19864 21232 19916
rect 21364 19864 21416 19916
rect 22468 20000 22520 20052
rect 26792 20043 26844 20052
rect 26792 20009 26801 20043
rect 26801 20009 26835 20043
rect 26835 20009 26844 20043
rect 26792 20000 26844 20009
rect 28356 20000 28408 20052
rect 29460 20000 29512 20052
rect 23388 19932 23440 19984
rect 23664 19864 23716 19916
rect 24124 19932 24176 19984
rect 24676 19932 24728 19984
rect 26424 19932 26476 19984
rect 30380 20000 30432 20052
rect 33508 20000 33560 20052
rect 34612 20000 34664 20052
rect 35808 20000 35860 20052
rect 23940 19864 23992 19916
rect 25412 19864 25464 19916
rect 26056 19864 26108 19916
rect 26148 19907 26200 19916
rect 26148 19873 26157 19907
rect 26157 19873 26191 19907
rect 26191 19873 26200 19907
rect 26148 19864 26200 19873
rect 27160 19864 27212 19916
rect 12164 19728 12216 19780
rect 12256 19771 12308 19780
rect 12256 19737 12265 19771
rect 12265 19737 12299 19771
rect 12299 19737 12308 19771
rect 12256 19728 12308 19737
rect 13544 19728 13596 19780
rect 13912 19728 13964 19780
rect 14556 19728 14608 19780
rect 17408 19796 17460 19848
rect 18512 19839 18564 19848
rect 18512 19805 18521 19839
rect 18521 19805 18555 19839
rect 18555 19805 18564 19839
rect 18512 19796 18564 19805
rect 15016 19771 15068 19780
rect 15016 19737 15025 19771
rect 15025 19737 15059 19771
rect 15059 19737 15068 19771
rect 15016 19728 15068 19737
rect 17040 19728 17092 19780
rect 19616 19728 19668 19780
rect 20168 19728 20220 19780
rect 16396 19660 16448 19712
rect 17224 19703 17276 19712
rect 17224 19669 17233 19703
rect 17233 19669 17267 19703
rect 17267 19669 17276 19703
rect 17224 19660 17276 19669
rect 17500 19660 17552 19712
rect 22376 19796 22428 19848
rect 29000 19907 29052 19916
rect 21548 19728 21600 19780
rect 21088 19660 21140 19712
rect 21180 19660 21232 19712
rect 24032 19728 24084 19780
rect 25228 19728 25280 19780
rect 25872 19728 25924 19780
rect 29000 19873 29009 19907
rect 29009 19873 29043 19907
rect 29043 19873 29052 19907
rect 29000 19864 29052 19873
rect 29460 19864 29512 19916
rect 30380 19864 30432 19916
rect 31300 19864 31352 19916
rect 31484 19907 31536 19916
rect 31484 19873 31493 19907
rect 31493 19873 31527 19907
rect 31527 19873 31536 19907
rect 31484 19864 31536 19873
rect 31944 19932 31996 19984
rect 33508 19864 33560 19916
rect 28908 19796 28960 19848
rect 22928 19703 22980 19712
rect 22928 19669 22937 19703
rect 22937 19669 22971 19703
rect 22971 19669 22980 19703
rect 22928 19660 22980 19669
rect 25964 19703 26016 19712
rect 25964 19669 25973 19703
rect 25973 19669 26007 19703
rect 26007 19669 26016 19703
rect 25964 19660 26016 19669
rect 26056 19703 26108 19712
rect 26056 19669 26065 19703
rect 26065 19669 26099 19703
rect 26099 19669 26108 19703
rect 26056 19660 26108 19669
rect 26884 19660 26936 19712
rect 27620 19660 27672 19712
rect 28724 19660 28776 19712
rect 28908 19660 28960 19712
rect 29736 19703 29788 19712
rect 29736 19669 29745 19703
rect 29745 19669 29779 19703
rect 29779 19669 29788 19703
rect 29736 19660 29788 19669
rect 30012 19728 30064 19780
rect 31116 19796 31168 19848
rect 31852 19796 31904 19848
rect 34980 19796 35032 19848
rect 35532 19907 35584 19916
rect 35532 19873 35541 19907
rect 35541 19873 35575 19907
rect 35575 19873 35584 19907
rect 35532 19864 35584 19873
rect 36176 19864 36228 19916
rect 37280 20000 37332 20052
rect 48596 20000 48648 20052
rect 48780 20043 48832 20052
rect 48780 20009 48789 20043
rect 48789 20009 48823 20043
rect 48823 20009 48832 20043
rect 48780 20000 48832 20009
rect 37096 19932 37148 19984
rect 38200 19932 38252 19984
rect 39764 19932 39816 19984
rect 41236 19975 41288 19984
rect 37372 19864 37424 19916
rect 37648 19864 37700 19916
rect 38752 19864 38804 19916
rect 39488 19864 39540 19916
rect 41236 19941 41245 19975
rect 41245 19941 41279 19975
rect 41279 19941 41288 19975
rect 41236 19932 41288 19941
rect 40592 19907 40644 19916
rect 40592 19873 40601 19907
rect 40601 19873 40635 19907
rect 40635 19873 40644 19907
rect 40592 19864 40644 19873
rect 41052 19907 41104 19916
rect 41052 19873 41061 19907
rect 41061 19873 41095 19907
rect 41095 19873 41104 19907
rect 41052 19864 41104 19873
rect 43904 19796 43956 19848
rect 32220 19728 32272 19780
rect 33784 19771 33836 19780
rect 33784 19737 33793 19771
rect 33793 19737 33827 19771
rect 33827 19737 33836 19771
rect 33784 19728 33836 19737
rect 30840 19660 30892 19712
rect 31668 19660 31720 19712
rect 32128 19703 32180 19712
rect 32128 19669 32137 19703
rect 32137 19669 32171 19703
rect 32171 19669 32180 19703
rect 32128 19660 32180 19669
rect 32404 19660 32456 19712
rect 32772 19660 32824 19712
rect 35072 19728 35124 19780
rect 35440 19728 35492 19780
rect 35624 19728 35676 19780
rect 34336 19660 34388 19712
rect 35808 19660 35860 19712
rect 40132 19728 40184 19780
rect 41052 19728 41104 19780
rect 49332 19728 49384 19780
rect 37832 19703 37884 19712
rect 37832 19669 37841 19703
rect 37841 19669 37875 19703
rect 37875 19669 37884 19703
rect 37832 19660 37884 19669
rect 38200 19703 38252 19712
rect 38200 19669 38209 19703
rect 38209 19669 38243 19703
rect 38243 19669 38252 19703
rect 38200 19660 38252 19669
rect 38660 19660 38712 19712
rect 39856 19660 39908 19712
rect 40040 19703 40092 19712
rect 40040 19669 40049 19703
rect 40049 19669 40083 19703
rect 40083 19669 40092 19703
rect 40040 19660 40092 19669
rect 45284 19660 45336 19712
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 27950 19558 28002 19610
rect 28014 19558 28066 19610
rect 28078 19558 28130 19610
rect 28142 19558 28194 19610
rect 28206 19558 28258 19610
rect 37950 19558 38002 19610
rect 38014 19558 38066 19610
rect 38078 19558 38130 19610
rect 38142 19558 38194 19610
rect 38206 19558 38258 19610
rect 47950 19558 48002 19610
rect 48014 19558 48066 19610
rect 48078 19558 48130 19610
rect 48142 19558 48194 19610
rect 48206 19558 48258 19610
rect 2872 19388 2924 19440
rect 9312 19456 9364 19508
rect 10048 19456 10100 19508
rect 13360 19456 13412 19508
rect 15016 19456 15068 19508
rect 16856 19499 16908 19508
rect 16856 19465 16865 19499
rect 16865 19465 16899 19499
rect 16899 19465 16908 19499
rect 16856 19456 16908 19465
rect 19340 19456 19392 19508
rect 19708 19456 19760 19508
rect 23848 19456 23900 19508
rect 4436 19431 4488 19440
rect 4436 19397 4445 19431
rect 4445 19397 4479 19431
rect 4479 19397 4488 19431
rect 4436 19388 4488 19397
rect 5356 19363 5408 19372
rect 5356 19329 5365 19363
rect 5365 19329 5399 19363
rect 5399 19329 5408 19363
rect 5356 19320 5408 19329
rect 12624 19388 12676 19440
rect 13544 19388 13596 19440
rect 16764 19388 16816 19440
rect 10876 19320 10928 19372
rect 11152 19363 11204 19372
rect 11152 19329 11161 19363
rect 11161 19329 11195 19363
rect 11195 19329 11204 19363
rect 11152 19320 11204 19329
rect 12072 19363 12124 19372
rect 12072 19329 12081 19363
rect 12081 19329 12115 19363
rect 12115 19329 12124 19363
rect 12072 19320 12124 19329
rect 12716 19363 12768 19372
rect 12716 19329 12725 19363
rect 12725 19329 12759 19363
rect 12759 19329 12768 19363
rect 12716 19320 12768 19329
rect 15384 19363 15436 19372
rect 9680 19295 9732 19304
rect 9680 19261 9689 19295
rect 9689 19261 9723 19295
rect 9723 19261 9732 19295
rect 9680 19252 9732 19261
rect 11336 19252 11388 19304
rect 9404 19184 9456 19236
rect 11244 19184 11296 19236
rect 15384 19329 15393 19363
rect 15393 19329 15427 19363
rect 15427 19329 15436 19363
rect 15384 19320 15436 19329
rect 18604 19388 18656 19440
rect 20536 19388 20588 19440
rect 21732 19388 21784 19440
rect 22744 19431 22796 19440
rect 22744 19397 22753 19431
rect 22753 19397 22787 19431
rect 22787 19397 22796 19431
rect 22744 19388 22796 19397
rect 24032 19388 24084 19440
rect 25780 19456 25832 19508
rect 25964 19456 26016 19508
rect 27344 19456 27396 19508
rect 27712 19456 27764 19508
rect 28448 19499 28500 19508
rect 28448 19465 28457 19499
rect 28457 19465 28491 19499
rect 28491 19465 28500 19499
rect 28448 19456 28500 19465
rect 24768 19388 24820 19440
rect 25228 19388 25280 19440
rect 15292 19252 15344 19304
rect 15752 19252 15804 19304
rect 16028 19184 16080 19236
rect 2320 19116 2372 19168
rect 8392 19116 8444 19168
rect 11888 19116 11940 19168
rect 16212 19159 16264 19168
rect 16212 19125 16221 19159
rect 16221 19125 16255 19159
rect 16255 19125 16264 19159
rect 16212 19116 16264 19125
rect 16764 19252 16816 19304
rect 20076 19363 20128 19372
rect 20076 19329 20085 19363
rect 20085 19329 20119 19363
rect 20119 19329 20128 19363
rect 20076 19320 20128 19329
rect 17408 19295 17460 19304
rect 17408 19261 17417 19295
rect 17417 19261 17451 19295
rect 17451 19261 17460 19295
rect 17408 19252 17460 19261
rect 20168 19252 20220 19304
rect 22928 19320 22980 19372
rect 23480 19363 23532 19372
rect 23480 19329 23489 19363
rect 23489 19329 23523 19363
rect 23523 19329 23532 19363
rect 23480 19320 23532 19329
rect 25504 19320 25556 19372
rect 25964 19320 26016 19372
rect 20444 19184 20496 19236
rect 25136 19252 25188 19304
rect 28264 19388 28316 19440
rect 28540 19388 28592 19440
rect 30012 19456 30064 19508
rect 30748 19456 30800 19508
rect 32864 19456 32916 19508
rect 26424 19295 26476 19346
rect 26424 19294 26433 19295
rect 26433 19294 26467 19295
rect 26467 19294 26476 19295
rect 28632 19320 28684 19372
rect 26608 19252 26660 19304
rect 28724 19252 28776 19304
rect 29184 19252 29236 19304
rect 32680 19431 32732 19440
rect 32680 19397 32689 19431
rect 32689 19397 32723 19431
rect 32723 19397 32732 19431
rect 32680 19388 32732 19397
rect 32772 19431 32824 19440
rect 32772 19397 32781 19431
rect 32781 19397 32815 19431
rect 32815 19397 32824 19431
rect 32772 19388 32824 19397
rect 33968 19499 34020 19508
rect 33968 19465 33977 19499
rect 33977 19465 34011 19499
rect 34011 19465 34020 19499
rect 33968 19456 34020 19465
rect 34428 19456 34480 19508
rect 35624 19456 35676 19508
rect 35900 19499 35952 19508
rect 35900 19465 35909 19499
rect 35909 19465 35943 19499
rect 35943 19465 35952 19499
rect 35900 19456 35952 19465
rect 37924 19456 37976 19508
rect 38384 19456 38436 19508
rect 40132 19499 40184 19508
rect 40132 19465 40141 19499
rect 40141 19465 40175 19499
rect 40175 19465 40184 19499
rect 40132 19456 40184 19465
rect 40408 19456 40460 19508
rect 49240 19456 49292 19508
rect 30380 19320 30432 19372
rect 32312 19320 32364 19372
rect 32588 19320 32640 19372
rect 34244 19320 34296 19372
rect 34612 19320 34664 19372
rect 36544 19388 36596 19440
rect 38476 19388 38528 19440
rect 39488 19388 39540 19440
rect 48412 19388 48464 19440
rect 36084 19320 36136 19372
rect 36268 19363 36320 19372
rect 36268 19329 36277 19363
rect 36277 19329 36311 19363
rect 36311 19329 36320 19363
rect 36268 19320 36320 19329
rect 36360 19363 36412 19372
rect 36360 19329 36369 19363
rect 36369 19329 36403 19363
rect 36403 19329 36412 19363
rect 36360 19320 36412 19329
rect 37740 19320 37792 19372
rect 40132 19320 40184 19372
rect 41236 19320 41288 19372
rect 45284 19320 45336 19372
rect 49148 19363 49200 19372
rect 49148 19329 49157 19363
rect 49157 19329 49191 19363
rect 49191 19329 49200 19363
rect 49148 19320 49200 19329
rect 19800 19116 19852 19168
rect 20536 19116 20588 19168
rect 21548 19116 21600 19168
rect 27804 19184 27856 19236
rect 28540 19184 28592 19236
rect 28632 19184 28684 19236
rect 31484 19252 31536 19304
rect 25228 19159 25280 19168
rect 25228 19125 25237 19159
rect 25237 19125 25271 19159
rect 25271 19125 25280 19159
rect 25228 19116 25280 19125
rect 25780 19159 25832 19168
rect 25780 19125 25789 19159
rect 25789 19125 25823 19159
rect 25823 19125 25832 19159
rect 25780 19116 25832 19125
rect 27252 19159 27304 19168
rect 27252 19125 27261 19159
rect 27261 19125 27295 19159
rect 27295 19125 27304 19159
rect 27252 19116 27304 19125
rect 27988 19116 28040 19168
rect 31116 19184 31168 19236
rect 35256 19252 35308 19304
rect 35900 19252 35952 19304
rect 38200 19295 38252 19304
rect 38200 19261 38209 19295
rect 38209 19261 38243 19295
rect 38243 19261 38252 19295
rect 38200 19252 38252 19261
rect 39212 19252 39264 19304
rect 41144 19295 41196 19304
rect 30380 19159 30432 19168
rect 30380 19125 30389 19159
rect 30389 19125 30423 19159
rect 30423 19125 30432 19159
rect 30380 19116 30432 19125
rect 32772 19116 32824 19168
rect 35900 19116 35952 19168
rect 36176 19116 36228 19168
rect 36360 19184 36412 19236
rect 36912 19227 36964 19236
rect 36912 19193 36921 19227
rect 36921 19193 36955 19227
rect 36955 19193 36964 19227
rect 36912 19184 36964 19193
rect 37372 19227 37424 19236
rect 37372 19193 37381 19227
rect 37381 19193 37415 19227
rect 37415 19193 37424 19227
rect 37372 19184 37424 19193
rect 37924 19184 37976 19236
rect 39488 19184 39540 19236
rect 40224 19184 40276 19236
rect 41144 19261 41153 19295
rect 41153 19261 41187 19295
rect 41187 19261 41196 19295
rect 41144 19252 41196 19261
rect 37464 19116 37516 19168
rect 38292 19116 38344 19168
rect 39764 19116 39816 19168
rect 41144 19116 41196 19168
rect 41604 19116 41656 19168
rect 49056 19116 49108 19168
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 32950 19014 33002 19066
rect 33014 19014 33066 19066
rect 33078 19014 33130 19066
rect 33142 19014 33194 19066
rect 33206 19014 33258 19066
rect 42950 19014 43002 19066
rect 43014 19014 43066 19066
rect 43078 19014 43130 19066
rect 43142 19014 43194 19066
rect 43206 19014 43258 19066
rect 3792 18776 3844 18828
rect 2780 18683 2832 18692
rect 2780 18649 2789 18683
rect 2789 18649 2823 18683
rect 2823 18649 2832 18683
rect 2780 18640 2832 18649
rect 8668 18776 8720 18828
rect 11060 18912 11112 18964
rect 11428 18912 11480 18964
rect 15108 18912 15160 18964
rect 10876 18887 10928 18896
rect 10876 18853 10885 18887
rect 10885 18853 10919 18887
rect 10919 18853 10928 18887
rect 10876 18844 10928 18853
rect 11888 18887 11940 18896
rect 11888 18853 11897 18887
rect 11897 18853 11931 18887
rect 11931 18853 11940 18887
rect 11888 18844 11940 18853
rect 10600 18776 10652 18828
rect 14096 18844 14148 18896
rect 13360 18776 13412 18828
rect 14280 18819 14332 18828
rect 14280 18785 14289 18819
rect 14289 18785 14323 18819
rect 14323 18785 14332 18819
rect 14280 18776 14332 18785
rect 15292 18776 15344 18828
rect 11520 18751 11572 18760
rect 11520 18717 11529 18751
rect 11529 18717 11563 18751
rect 11563 18717 11572 18751
rect 11520 18708 11572 18717
rect 11888 18708 11940 18760
rect 8300 18615 8352 18624
rect 8300 18581 8309 18615
rect 8309 18581 8343 18615
rect 8343 18581 8352 18615
rect 8300 18572 8352 18581
rect 9404 18683 9456 18692
rect 9404 18649 9413 18683
rect 9413 18649 9447 18683
rect 9447 18649 9456 18683
rect 9404 18640 9456 18649
rect 11704 18640 11756 18692
rect 12624 18708 12676 18760
rect 13268 18708 13320 18760
rect 13452 18708 13504 18760
rect 16028 18955 16080 18964
rect 16028 18921 16037 18955
rect 16037 18921 16071 18955
rect 16071 18921 16080 18955
rect 16028 18912 16080 18921
rect 16488 18912 16540 18964
rect 17040 18912 17092 18964
rect 19616 18912 19668 18964
rect 21088 18955 21140 18964
rect 21088 18921 21097 18955
rect 21097 18921 21131 18955
rect 21131 18921 21140 18955
rect 21088 18912 21140 18921
rect 15936 18844 15988 18896
rect 16304 18776 16356 18828
rect 17684 18844 17736 18896
rect 18696 18776 18748 18828
rect 18972 18776 19024 18828
rect 21364 18776 21416 18828
rect 21640 18819 21692 18828
rect 21640 18785 21649 18819
rect 21649 18785 21683 18819
rect 21683 18785 21692 18819
rect 21640 18776 21692 18785
rect 16672 18708 16724 18760
rect 17408 18751 17460 18760
rect 17408 18717 17417 18751
rect 17417 18717 17451 18751
rect 17451 18717 17460 18751
rect 17408 18708 17460 18717
rect 17776 18708 17828 18760
rect 13452 18572 13504 18624
rect 16948 18640 17000 18692
rect 15568 18572 15620 18624
rect 16764 18572 16816 18624
rect 19064 18708 19116 18760
rect 18880 18640 18932 18692
rect 19156 18572 19208 18624
rect 19340 18615 19392 18624
rect 19340 18581 19349 18615
rect 19349 18581 19383 18615
rect 19383 18581 19392 18615
rect 19340 18572 19392 18581
rect 25136 18912 25188 18964
rect 33048 18912 33100 18964
rect 33968 18912 34020 18964
rect 34336 18912 34388 18964
rect 34520 18955 34572 18964
rect 34520 18921 34529 18955
rect 34529 18921 34563 18955
rect 34563 18921 34572 18955
rect 34520 18912 34572 18921
rect 23664 18844 23716 18896
rect 22652 18776 22704 18828
rect 23296 18776 23348 18828
rect 25688 18776 25740 18828
rect 28356 18844 28408 18896
rect 28908 18844 28960 18896
rect 36912 18912 36964 18964
rect 38200 18912 38252 18964
rect 37464 18844 37516 18896
rect 38752 18844 38804 18896
rect 42708 18844 42760 18896
rect 27068 18776 27120 18828
rect 27344 18776 27396 18828
rect 29460 18776 29512 18828
rect 29644 18776 29696 18828
rect 30288 18819 30340 18828
rect 30288 18785 30297 18819
rect 30297 18785 30331 18819
rect 30331 18785 30340 18819
rect 30288 18776 30340 18785
rect 31944 18819 31996 18828
rect 31944 18785 31953 18819
rect 31953 18785 31987 18819
rect 31987 18785 31996 18819
rect 31944 18776 31996 18785
rect 27436 18708 27488 18760
rect 22284 18640 22336 18692
rect 21180 18572 21232 18624
rect 21456 18615 21508 18624
rect 21456 18581 21465 18615
rect 21465 18581 21499 18615
rect 21499 18581 21508 18615
rect 21456 18572 21508 18581
rect 21640 18572 21692 18624
rect 22376 18572 22428 18624
rect 24124 18640 24176 18692
rect 24768 18640 24820 18692
rect 25044 18683 25096 18692
rect 25044 18649 25053 18683
rect 25053 18649 25087 18683
rect 25087 18649 25096 18683
rect 25044 18640 25096 18649
rect 25228 18640 25280 18692
rect 27804 18640 27856 18692
rect 28448 18708 28500 18760
rect 29184 18751 29236 18760
rect 29184 18717 29193 18751
rect 29193 18717 29227 18751
rect 29227 18717 29236 18751
rect 29184 18708 29236 18717
rect 29920 18708 29972 18760
rect 29000 18640 29052 18692
rect 34152 18776 34204 18828
rect 35992 18776 36044 18828
rect 37556 18776 37608 18828
rect 32588 18708 32640 18760
rect 37004 18708 37056 18760
rect 35348 18640 35400 18692
rect 23940 18572 23992 18624
rect 24400 18572 24452 18624
rect 27988 18615 28040 18624
rect 27988 18581 27997 18615
rect 27997 18581 28031 18615
rect 28031 18581 28040 18615
rect 27988 18572 28040 18581
rect 28724 18572 28776 18624
rect 29920 18572 29972 18624
rect 30472 18572 30524 18624
rect 31668 18572 31720 18624
rect 31852 18615 31904 18624
rect 31852 18581 31861 18615
rect 31861 18581 31895 18615
rect 31895 18581 31904 18615
rect 31852 18572 31904 18581
rect 32036 18572 32088 18624
rect 32956 18572 33008 18624
rect 33140 18615 33192 18624
rect 33140 18581 33149 18615
rect 33149 18581 33183 18615
rect 33183 18581 33192 18615
rect 33140 18572 33192 18581
rect 33692 18572 33744 18624
rect 34152 18572 34204 18624
rect 34244 18615 34296 18624
rect 34244 18581 34253 18615
rect 34253 18581 34287 18615
rect 34287 18581 34296 18615
rect 34244 18572 34296 18581
rect 34704 18572 34756 18624
rect 38016 18615 38068 18624
rect 38016 18581 38025 18615
rect 38025 18581 38059 18615
rect 38059 18581 38068 18615
rect 38016 18572 38068 18581
rect 38568 18819 38620 18828
rect 38568 18785 38577 18819
rect 38577 18785 38611 18819
rect 38611 18785 38620 18819
rect 38568 18776 38620 18785
rect 38384 18708 38436 18760
rect 48780 18708 48832 18760
rect 49148 18708 49200 18760
rect 39764 18640 39816 18692
rect 41604 18640 41656 18692
rect 40500 18572 40552 18624
rect 40592 18572 40644 18624
rect 48412 18615 48464 18624
rect 48412 18581 48421 18615
rect 48421 18581 48455 18615
rect 48455 18581 48464 18615
rect 48412 18572 48464 18581
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 27950 18470 28002 18522
rect 28014 18470 28066 18522
rect 28078 18470 28130 18522
rect 28142 18470 28194 18522
rect 28206 18470 28258 18522
rect 37950 18470 38002 18522
rect 38014 18470 38066 18522
rect 38078 18470 38130 18522
rect 38142 18470 38194 18522
rect 38206 18470 38258 18522
rect 47950 18470 48002 18522
rect 48014 18470 48066 18522
rect 48078 18470 48130 18522
rect 48142 18470 48194 18522
rect 48206 18470 48258 18522
rect 5080 18368 5132 18420
rect 5632 18368 5684 18420
rect 9680 18368 9732 18420
rect 4988 18300 5040 18352
rect 2780 18207 2832 18216
rect 2780 18173 2789 18207
rect 2789 18173 2823 18207
rect 2823 18173 2832 18207
rect 2780 18164 2832 18173
rect 3700 18232 3752 18284
rect 11612 18300 11664 18352
rect 4160 18207 4212 18216
rect 4160 18173 4169 18207
rect 4169 18173 4203 18207
rect 4203 18173 4212 18207
rect 4160 18164 4212 18173
rect 11428 18232 11480 18284
rect 10232 18096 10284 18148
rect 10416 18139 10468 18148
rect 10416 18105 10425 18139
rect 10425 18105 10459 18139
rect 10459 18105 10468 18139
rect 10416 18096 10468 18105
rect 10324 18028 10376 18080
rect 11060 18164 11112 18216
rect 12716 18368 12768 18420
rect 13544 18368 13596 18420
rect 13636 18368 13688 18420
rect 15016 18411 15068 18420
rect 15016 18377 15025 18411
rect 15025 18377 15059 18411
rect 15059 18377 15068 18411
rect 15016 18368 15068 18377
rect 11888 18300 11940 18352
rect 13452 18300 13504 18352
rect 25780 18368 25832 18420
rect 27252 18368 27304 18420
rect 29000 18368 29052 18420
rect 29184 18368 29236 18420
rect 36176 18368 36228 18420
rect 39212 18368 39264 18420
rect 39764 18411 39816 18420
rect 39764 18377 39773 18411
rect 39773 18377 39807 18411
rect 39807 18377 39816 18411
rect 39764 18368 39816 18377
rect 40040 18368 40092 18420
rect 48780 18411 48832 18420
rect 48780 18377 48789 18411
rect 48789 18377 48823 18411
rect 48823 18377 48832 18411
rect 48780 18368 48832 18377
rect 14188 18232 14240 18284
rect 16672 18343 16724 18352
rect 16672 18309 16681 18343
rect 16681 18309 16715 18343
rect 16715 18309 16724 18343
rect 16672 18300 16724 18309
rect 10600 18096 10652 18148
rect 13360 18164 13412 18216
rect 13268 18096 13320 18148
rect 15292 18164 15344 18216
rect 16212 18164 16264 18216
rect 17776 18164 17828 18216
rect 12164 18028 12216 18080
rect 12348 18028 12400 18080
rect 15384 18096 15436 18148
rect 16120 18139 16172 18148
rect 16120 18105 16129 18139
rect 16129 18105 16163 18139
rect 16163 18105 16172 18139
rect 16120 18096 16172 18105
rect 19524 18232 19576 18284
rect 19892 18300 19944 18352
rect 21548 18300 21600 18352
rect 22836 18300 22888 18352
rect 23480 18300 23532 18352
rect 20904 18164 20956 18216
rect 22744 18207 22796 18216
rect 22744 18173 22753 18207
rect 22753 18173 22787 18207
rect 22787 18173 22796 18207
rect 22744 18164 22796 18173
rect 24676 18232 24728 18284
rect 27620 18300 27672 18352
rect 32128 18300 32180 18352
rect 32588 18300 32640 18352
rect 33140 18300 33192 18352
rect 34428 18300 34480 18352
rect 35716 18300 35768 18352
rect 25044 18275 25096 18284
rect 25044 18241 25053 18275
rect 25053 18241 25087 18275
rect 25087 18241 25096 18275
rect 25044 18232 25096 18241
rect 25136 18275 25188 18284
rect 25136 18241 25145 18275
rect 25145 18241 25179 18275
rect 25179 18241 25188 18275
rect 25136 18232 25188 18241
rect 27436 18232 27488 18284
rect 25320 18207 25372 18216
rect 25320 18173 25329 18207
rect 25329 18173 25363 18207
rect 25363 18173 25372 18207
rect 25320 18164 25372 18173
rect 19616 18096 19668 18148
rect 23756 18096 23808 18148
rect 26240 18164 26292 18216
rect 26424 18207 26476 18216
rect 26424 18173 26433 18207
rect 26433 18173 26467 18207
rect 26467 18173 26476 18207
rect 26424 18164 26476 18173
rect 27252 18164 27304 18216
rect 16580 18028 16632 18080
rect 18972 18071 19024 18080
rect 18972 18037 18981 18071
rect 18981 18037 19015 18071
rect 19015 18037 19024 18071
rect 18972 18028 19024 18037
rect 21916 18028 21968 18080
rect 22284 18028 22336 18080
rect 25504 18096 25556 18148
rect 25044 18028 25096 18080
rect 27160 18071 27212 18080
rect 27160 18037 27169 18071
rect 27169 18037 27203 18071
rect 27203 18037 27212 18071
rect 27160 18028 27212 18037
rect 27436 18028 27488 18080
rect 29736 18232 29788 18284
rect 32680 18275 32732 18284
rect 32680 18241 32689 18275
rect 32689 18241 32723 18275
rect 32723 18241 32732 18275
rect 32680 18232 32732 18241
rect 33048 18232 33100 18284
rect 35992 18232 36044 18284
rect 37372 18232 37424 18284
rect 37464 18232 37516 18284
rect 38384 18300 38436 18352
rect 40224 18300 40276 18352
rect 48412 18232 48464 18284
rect 49056 18275 49108 18284
rect 49056 18241 49065 18275
rect 49065 18241 49099 18275
rect 49099 18241 49108 18275
rect 49056 18232 49108 18241
rect 28816 18164 28868 18216
rect 29368 18096 29420 18148
rect 31392 18164 31444 18216
rect 30104 18139 30156 18148
rect 30104 18105 30113 18139
rect 30113 18105 30147 18139
rect 30147 18105 30156 18139
rect 30104 18096 30156 18105
rect 28540 18028 28592 18080
rect 33416 18164 33468 18216
rect 32496 18096 32548 18148
rect 33876 18207 33928 18216
rect 33876 18173 33885 18207
rect 33885 18173 33919 18207
rect 33919 18173 33928 18207
rect 33876 18164 33928 18173
rect 34336 18164 34388 18216
rect 35348 18207 35400 18216
rect 35348 18173 35357 18207
rect 35357 18173 35391 18207
rect 35391 18173 35400 18207
rect 35348 18164 35400 18173
rect 37832 18164 37884 18216
rect 38292 18207 38344 18216
rect 38292 18173 38301 18207
rect 38301 18173 38335 18207
rect 38335 18173 38344 18207
rect 38292 18164 38344 18173
rect 36268 18028 36320 18080
rect 36636 18096 36688 18148
rect 37280 18028 37332 18080
rect 48320 18028 48372 18080
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 32950 17926 33002 17978
rect 33014 17926 33066 17978
rect 33078 17926 33130 17978
rect 33142 17926 33194 17978
rect 33206 17926 33258 17978
rect 42950 17926 43002 17978
rect 43014 17926 43066 17978
rect 43078 17926 43130 17978
rect 43142 17926 43194 17978
rect 43206 17926 43258 17978
rect 11060 17824 11112 17876
rect 12256 17824 12308 17876
rect 12532 17824 12584 17876
rect 11980 17756 12032 17808
rect 1216 17688 1268 17740
rect 10600 17731 10652 17740
rect 10600 17697 10609 17731
rect 10609 17697 10643 17731
rect 10643 17697 10652 17731
rect 10600 17688 10652 17697
rect 8576 17620 8628 17672
rect 12256 17688 12308 17740
rect 12900 17688 12952 17740
rect 15016 17824 15068 17876
rect 15292 17824 15344 17876
rect 17224 17824 17276 17876
rect 17316 17824 17368 17876
rect 19616 17824 19668 17876
rect 16120 17756 16172 17808
rect 21732 17824 21784 17876
rect 24676 17824 24728 17876
rect 28908 17824 28960 17876
rect 29460 17824 29512 17876
rect 32588 17824 32640 17876
rect 34152 17824 34204 17876
rect 34888 17824 34940 17876
rect 34980 17824 35032 17876
rect 35164 17824 35216 17876
rect 13544 17688 13596 17740
rect 15200 17688 15252 17740
rect 16304 17688 16356 17740
rect 17684 17688 17736 17740
rect 18788 17731 18840 17740
rect 18788 17697 18797 17731
rect 18797 17697 18831 17731
rect 18831 17697 18840 17731
rect 18788 17688 18840 17697
rect 19892 17688 19944 17740
rect 20260 17731 20312 17740
rect 20260 17697 20269 17731
rect 20269 17697 20303 17731
rect 20303 17697 20312 17731
rect 20260 17688 20312 17697
rect 25596 17756 25648 17808
rect 26332 17799 26384 17808
rect 26332 17765 26341 17799
rect 26341 17765 26375 17799
rect 26375 17765 26384 17799
rect 26332 17756 26384 17765
rect 28540 17756 28592 17808
rect 30380 17756 30432 17808
rect 34612 17756 34664 17808
rect 13084 17663 13136 17672
rect 13084 17629 13093 17663
rect 13093 17629 13127 17663
rect 13127 17629 13136 17663
rect 13084 17620 13136 17629
rect 11520 17552 11572 17604
rect 12256 17484 12308 17536
rect 12900 17484 12952 17536
rect 13636 17484 13688 17536
rect 16212 17620 16264 17672
rect 18328 17620 18380 17672
rect 18972 17620 19024 17672
rect 20168 17620 20220 17672
rect 22192 17688 22244 17740
rect 23756 17731 23808 17740
rect 23756 17697 23765 17731
rect 23765 17697 23799 17731
rect 23799 17697 23808 17731
rect 23756 17688 23808 17697
rect 24032 17688 24084 17740
rect 25044 17731 25096 17740
rect 25044 17697 25053 17731
rect 25053 17697 25087 17731
rect 25087 17697 25096 17731
rect 25044 17688 25096 17697
rect 14648 17552 14700 17604
rect 15108 17552 15160 17604
rect 19708 17552 19760 17604
rect 19892 17552 19944 17604
rect 17500 17484 17552 17536
rect 18512 17484 18564 17536
rect 20352 17484 20404 17536
rect 20536 17595 20588 17604
rect 20536 17561 20545 17595
rect 20545 17561 20579 17595
rect 20579 17561 20588 17595
rect 20536 17552 20588 17561
rect 21548 17552 21600 17604
rect 20720 17484 20772 17536
rect 21180 17484 21232 17536
rect 21456 17484 21508 17536
rect 23940 17620 23992 17672
rect 28356 17688 28408 17740
rect 25596 17620 25648 17672
rect 24400 17552 24452 17604
rect 28908 17620 28960 17672
rect 30380 17620 30432 17672
rect 24768 17484 24820 17536
rect 24860 17484 24912 17536
rect 26608 17484 26660 17536
rect 27344 17595 27396 17604
rect 27344 17561 27353 17595
rect 27353 17561 27387 17595
rect 27387 17561 27396 17595
rect 27344 17552 27396 17561
rect 27620 17552 27672 17604
rect 30104 17552 30156 17604
rect 30932 17688 30984 17740
rect 30840 17620 30892 17672
rect 31944 17731 31996 17740
rect 31944 17697 31953 17731
rect 31953 17697 31987 17731
rect 31987 17697 31996 17731
rect 31944 17688 31996 17697
rect 33232 17731 33284 17740
rect 33232 17697 33241 17731
rect 33241 17697 33275 17731
rect 33275 17697 33284 17731
rect 33232 17688 33284 17697
rect 35164 17688 35216 17740
rect 48596 17824 48648 17876
rect 39856 17756 39908 17808
rect 40500 17799 40552 17808
rect 40500 17765 40509 17799
rect 40509 17765 40543 17799
rect 40543 17765 40552 17799
rect 40500 17756 40552 17765
rect 35716 17688 35768 17740
rect 36176 17688 36228 17740
rect 36544 17688 36596 17740
rect 38476 17731 38528 17740
rect 38476 17697 38485 17731
rect 38485 17697 38519 17731
rect 38519 17697 38528 17731
rect 38476 17688 38528 17697
rect 37464 17620 37516 17672
rect 32496 17552 32548 17604
rect 39948 17688 40000 17740
rect 41052 17731 41104 17740
rect 41052 17697 41061 17731
rect 41061 17697 41095 17731
rect 41095 17697 41104 17731
rect 41052 17688 41104 17697
rect 49056 17663 49108 17672
rect 49056 17629 49065 17663
rect 49065 17629 49099 17663
rect 49099 17629 49108 17663
rect 49056 17620 49108 17629
rect 28816 17527 28868 17536
rect 28816 17493 28825 17527
rect 28825 17493 28859 17527
rect 28859 17493 28868 17527
rect 28816 17484 28868 17493
rect 29644 17527 29696 17536
rect 29644 17493 29653 17527
rect 29653 17493 29687 17527
rect 29687 17493 29696 17527
rect 29644 17484 29696 17493
rect 30380 17484 30432 17536
rect 31208 17484 31260 17536
rect 31392 17484 31444 17536
rect 31484 17484 31536 17536
rect 32128 17484 32180 17536
rect 32680 17484 32732 17536
rect 33416 17484 33468 17536
rect 34888 17527 34940 17536
rect 34888 17493 34897 17527
rect 34897 17493 34931 17527
rect 34931 17493 34940 17527
rect 34888 17484 34940 17493
rect 35256 17484 35308 17536
rect 35440 17484 35492 17536
rect 35900 17484 35952 17536
rect 36176 17484 36228 17536
rect 36820 17484 36872 17536
rect 48412 17552 48464 17604
rect 48504 17552 48556 17604
rect 38384 17527 38436 17536
rect 38384 17493 38393 17527
rect 38393 17493 38427 17527
rect 38427 17493 38436 17527
rect 38384 17484 38436 17493
rect 49148 17484 49200 17536
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 27950 17382 28002 17434
rect 28014 17382 28066 17434
rect 28078 17382 28130 17434
rect 28142 17382 28194 17434
rect 28206 17382 28258 17434
rect 37950 17382 38002 17434
rect 38014 17382 38066 17434
rect 38078 17382 38130 17434
rect 38142 17382 38194 17434
rect 38206 17382 38258 17434
rect 47950 17382 48002 17434
rect 48014 17382 48066 17434
rect 48078 17382 48130 17434
rect 48142 17382 48194 17434
rect 48206 17382 48258 17434
rect 13452 17280 13504 17332
rect 14004 17280 14056 17332
rect 15568 17323 15620 17332
rect 15568 17289 15577 17323
rect 15577 17289 15611 17323
rect 15611 17289 15620 17323
rect 15568 17280 15620 17289
rect 16120 17280 16172 17332
rect 16488 17280 16540 17332
rect 18420 17280 18472 17332
rect 11796 17255 11848 17264
rect 11796 17221 11805 17255
rect 11805 17221 11839 17255
rect 11839 17221 11848 17255
rect 11796 17212 11848 17221
rect 13728 17212 13780 17264
rect 14280 17212 14332 17264
rect 15016 17212 15068 17264
rect 8300 17144 8352 17196
rect 9956 17144 10008 17196
rect 1308 17076 1360 17128
rect 10692 17076 10744 17128
rect 11980 17076 12032 17128
rect 14372 17144 14424 17196
rect 15108 17187 15160 17196
rect 15108 17153 15117 17187
rect 15117 17153 15151 17187
rect 15151 17153 15160 17187
rect 15108 17144 15160 17153
rect 15752 17144 15804 17196
rect 18328 17212 18380 17264
rect 16028 17076 16080 17128
rect 11060 17008 11112 17060
rect 18512 17144 18564 17196
rect 20260 17280 20312 17332
rect 20352 17280 20404 17332
rect 20536 17144 20588 17196
rect 17040 17076 17092 17128
rect 18604 17119 18656 17128
rect 18604 17085 18613 17119
rect 18613 17085 18647 17119
rect 18647 17085 18656 17119
rect 18604 17076 18656 17085
rect 20076 17076 20128 17128
rect 20904 17323 20956 17332
rect 20904 17289 20913 17323
rect 20913 17289 20947 17323
rect 20947 17289 20956 17323
rect 20904 17280 20956 17289
rect 20996 17280 21048 17332
rect 22192 17280 22244 17332
rect 23940 17280 23992 17332
rect 24952 17280 25004 17332
rect 24768 17212 24820 17264
rect 22652 17187 22704 17196
rect 22652 17153 22661 17187
rect 22661 17153 22695 17187
rect 22695 17153 22704 17187
rect 22652 17144 22704 17153
rect 24032 17144 24084 17196
rect 25228 17187 25280 17196
rect 25228 17153 25237 17187
rect 25237 17153 25271 17187
rect 25271 17153 25280 17187
rect 25228 17144 25280 17153
rect 25964 17255 26016 17264
rect 25964 17221 25973 17255
rect 25973 17221 26007 17255
rect 26007 17221 26016 17255
rect 25964 17212 26016 17221
rect 28540 17280 28592 17332
rect 32312 17280 32364 17332
rect 32404 17280 32456 17332
rect 33324 17280 33376 17332
rect 34888 17280 34940 17332
rect 27896 17212 27948 17264
rect 29276 17212 29328 17264
rect 27344 17144 27396 17196
rect 27528 17144 27580 17196
rect 9864 16983 9916 16992
rect 9864 16949 9873 16983
rect 9873 16949 9907 16983
rect 9907 16949 9916 16983
rect 9864 16940 9916 16949
rect 11704 16940 11756 16992
rect 12716 16983 12768 16992
rect 12716 16949 12725 16983
rect 12725 16949 12759 16983
rect 12759 16949 12768 16983
rect 12716 16940 12768 16949
rect 13084 16940 13136 16992
rect 17408 16940 17460 16992
rect 17500 16983 17552 16992
rect 17500 16949 17509 16983
rect 17509 16949 17543 16983
rect 17543 16949 17552 16983
rect 17500 16940 17552 16949
rect 22652 17008 22704 17060
rect 19892 16940 19944 16992
rect 21548 16940 21600 16992
rect 22560 16940 22612 16992
rect 23664 17076 23716 17128
rect 25136 17076 25188 17128
rect 27252 17076 27304 17128
rect 28080 17144 28132 17196
rect 29460 17144 29512 17196
rect 29644 17144 29696 17196
rect 28540 17076 28592 17128
rect 29184 17119 29236 17128
rect 29184 17085 29193 17119
rect 29193 17085 29227 17119
rect 29227 17085 29236 17119
rect 29184 17076 29236 17085
rect 29828 17076 29880 17128
rect 30380 17119 30432 17128
rect 30380 17085 30389 17119
rect 30389 17085 30423 17119
rect 30423 17085 30432 17119
rect 30380 17076 30432 17085
rect 25872 17008 25924 17060
rect 28816 17008 28868 17060
rect 30932 17144 30984 17196
rect 31208 17144 31260 17196
rect 32128 17144 32180 17196
rect 32496 17212 32548 17264
rect 32588 17255 32640 17264
rect 32588 17221 32597 17255
rect 32597 17221 32631 17255
rect 32631 17221 32640 17255
rect 32588 17212 32640 17221
rect 34152 17212 34204 17264
rect 34612 17255 34664 17264
rect 34612 17221 34621 17255
rect 34621 17221 34655 17255
rect 34655 17221 34664 17255
rect 34612 17212 34664 17221
rect 35348 17212 35400 17264
rect 35624 17212 35676 17264
rect 36452 17255 36504 17264
rect 36452 17221 36461 17255
rect 36461 17221 36495 17255
rect 36495 17221 36504 17255
rect 36452 17212 36504 17221
rect 37740 17212 37792 17264
rect 40132 17280 40184 17332
rect 40224 17280 40276 17332
rect 48320 17280 48372 17332
rect 48412 17323 48464 17332
rect 48412 17289 48421 17323
rect 48421 17289 48455 17323
rect 48455 17289 48464 17323
rect 48412 17280 48464 17289
rect 48596 17280 48648 17332
rect 41144 17212 41196 17264
rect 36084 17144 36136 17196
rect 30564 17076 30616 17128
rect 25964 16940 26016 16992
rect 26332 16940 26384 16992
rect 27804 16940 27856 16992
rect 30748 17008 30800 17060
rect 31668 17076 31720 17128
rect 33876 17076 33928 17128
rect 34888 17076 34940 17128
rect 36268 17144 36320 17196
rect 48780 17144 48832 17196
rect 49240 17144 49292 17196
rect 36544 17076 36596 17128
rect 36636 17119 36688 17128
rect 36636 17085 36645 17119
rect 36645 17085 36679 17119
rect 36679 17085 36688 17119
rect 36636 17076 36688 17085
rect 38292 17076 38344 17128
rect 38476 17119 38528 17128
rect 38476 17085 38485 17119
rect 38485 17085 38519 17119
rect 38519 17085 38528 17119
rect 38476 17076 38528 17085
rect 30932 16940 30984 16992
rect 33968 16940 34020 16992
rect 36544 16940 36596 16992
rect 37188 17008 37240 17060
rect 37740 17008 37792 17060
rect 40592 17076 40644 17128
rect 40408 17008 40460 17060
rect 41328 17008 41380 17060
rect 37648 16940 37700 16992
rect 38292 16940 38344 16992
rect 41052 16940 41104 16992
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 32950 16838 33002 16890
rect 33014 16838 33066 16890
rect 33078 16838 33130 16890
rect 33142 16838 33194 16890
rect 33206 16838 33258 16890
rect 42950 16838 43002 16890
rect 43014 16838 43066 16890
rect 43078 16838 43130 16890
rect 43142 16838 43194 16890
rect 43206 16838 43258 16890
rect 5356 16736 5408 16788
rect 11980 16736 12032 16788
rect 14280 16736 14332 16788
rect 14740 16736 14792 16788
rect 17224 16736 17276 16788
rect 18788 16736 18840 16788
rect 20996 16736 21048 16788
rect 4528 16600 4580 16652
rect 5448 16600 5500 16652
rect 8484 16600 8536 16652
rect 8576 16600 8628 16652
rect 10876 16600 10928 16652
rect 13912 16600 13964 16652
rect 15200 16668 15252 16720
rect 16948 16668 17000 16720
rect 18420 16668 18472 16720
rect 23940 16736 23992 16788
rect 27344 16779 27396 16788
rect 22744 16711 22796 16720
rect 22744 16677 22753 16711
rect 22753 16677 22787 16711
rect 22787 16677 22796 16711
rect 22744 16668 22796 16677
rect 27344 16745 27353 16779
rect 27353 16745 27387 16779
rect 27387 16745 27396 16779
rect 27344 16736 27396 16745
rect 28632 16779 28684 16788
rect 28632 16745 28641 16779
rect 28641 16745 28675 16779
rect 28675 16745 28684 16779
rect 28632 16736 28684 16745
rect 11060 16532 11112 16584
rect 11520 16532 11572 16584
rect 11704 16532 11756 16584
rect 13360 16532 13412 16584
rect 14188 16532 14240 16584
rect 16120 16643 16172 16652
rect 16120 16609 16129 16643
rect 16129 16609 16163 16643
rect 16163 16609 16172 16643
rect 16120 16600 16172 16609
rect 16304 16600 16356 16652
rect 18604 16600 18656 16652
rect 20352 16600 20404 16652
rect 1308 16464 1360 16516
rect 9588 16464 9640 16516
rect 10508 16464 10560 16516
rect 12624 16464 12676 16516
rect 16488 16532 16540 16584
rect 7840 16396 7892 16448
rect 11336 16396 11388 16448
rect 11520 16439 11572 16448
rect 11520 16405 11529 16439
rect 11529 16405 11563 16439
rect 11563 16405 11572 16439
rect 11520 16396 11572 16405
rect 12532 16396 12584 16448
rect 12992 16439 13044 16448
rect 12992 16405 13001 16439
rect 13001 16405 13035 16439
rect 13035 16405 13044 16439
rect 12992 16396 13044 16405
rect 13636 16396 13688 16448
rect 15016 16464 15068 16516
rect 15476 16464 15528 16516
rect 14740 16396 14792 16448
rect 14832 16396 14884 16448
rect 15660 16439 15712 16448
rect 15660 16405 15669 16439
rect 15669 16405 15703 16439
rect 15703 16405 15712 16439
rect 15660 16396 15712 16405
rect 17224 16396 17276 16448
rect 18880 16439 18932 16448
rect 18880 16405 18889 16439
rect 18889 16405 18923 16439
rect 18923 16405 18932 16439
rect 18880 16396 18932 16405
rect 18972 16396 19024 16448
rect 21272 16643 21324 16652
rect 21272 16609 21281 16643
rect 21281 16609 21315 16643
rect 21315 16609 21324 16643
rect 21272 16600 21324 16609
rect 25504 16668 25556 16720
rect 27620 16668 27672 16720
rect 24584 16600 24636 16652
rect 25596 16643 25648 16652
rect 25596 16609 25605 16643
rect 25605 16609 25639 16643
rect 25639 16609 25648 16643
rect 25596 16600 25648 16609
rect 25872 16643 25924 16652
rect 25872 16609 25881 16643
rect 25881 16609 25915 16643
rect 25915 16609 25924 16643
rect 25872 16600 25924 16609
rect 26608 16600 26660 16652
rect 26976 16532 27028 16584
rect 27528 16532 27580 16584
rect 29276 16643 29328 16652
rect 29276 16609 29285 16643
rect 29285 16609 29319 16643
rect 29319 16609 29328 16643
rect 29276 16600 29328 16609
rect 29460 16600 29512 16652
rect 31668 16600 31720 16652
rect 32496 16600 32548 16652
rect 28816 16532 28868 16584
rect 34152 16668 34204 16720
rect 34612 16736 34664 16788
rect 48504 16736 48556 16788
rect 48780 16779 48832 16788
rect 48780 16745 48789 16779
rect 48789 16745 48823 16779
rect 48823 16745 48832 16779
rect 48780 16736 48832 16745
rect 34428 16600 34480 16652
rect 35716 16643 35768 16652
rect 35716 16609 35725 16643
rect 35725 16609 35759 16643
rect 35759 16609 35768 16643
rect 35716 16600 35768 16609
rect 36268 16711 36320 16720
rect 36268 16677 36277 16711
rect 36277 16677 36311 16711
rect 36311 16677 36320 16711
rect 36268 16668 36320 16677
rect 36728 16643 36780 16652
rect 36728 16609 36737 16643
rect 36737 16609 36771 16643
rect 36771 16609 36780 16643
rect 36728 16600 36780 16609
rect 37004 16668 37056 16720
rect 37464 16668 37516 16720
rect 41236 16711 41288 16720
rect 20536 16396 20588 16448
rect 20812 16396 20864 16448
rect 22560 16464 22612 16516
rect 22836 16464 22888 16516
rect 24676 16507 24728 16516
rect 24676 16473 24685 16507
rect 24685 16473 24719 16507
rect 24719 16473 24728 16507
rect 24676 16464 24728 16473
rect 22652 16396 22704 16448
rect 23296 16439 23348 16448
rect 23296 16405 23305 16439
rect 23305 16405 23339 16439
rect 23339 16405 23348 16439
rect 23296 16396 23348 16405
rect 23388 16396 23440 16448
rect 24032 16396 24084 16448
rect 25964 16464 26016 16516
rect 27252 16464 27304 16516
rect 28264 16464 28316 16516
rect 29000 16464 29052 16516
rect 30196 16507 30248 16516
rect 30196 16473 30205 16507
rect 30205 16473 30239 16507
rect 30239 16473 30248 16507
rect 30196 16464 30248 16473
rect 25044 16396 25096 16448
rect 28080 16396 28132 16448
rect 30840 16396 30892 16448
rect 31852 16464 31904 16516
rect 31300 16439 31352 16448
rect 31300 16405 31309 16439
rect 31309 16405 31343 16439
rect 31343 16405 31352 16439
rect 31300 16396 31352 16405
rect 32128 16464 32180 16516
rect 32404 16464 32456 16516
rect 34520 16532 34572 16584
rect 34612 16532 34664 16584
rect 35900 16532 35952 16584
rect 40224 16600 40276 16652
rect 36912 16532 36964 16584
rect 37464 16532 37516 16584
rect 37740 16575 37792 16584
rect 37740 16541 37749 16575
rect 37749 16541 37783 16575
rect 37783 16541 37792 16575
rect 37740 16532 37792 16541
rect 41236 16677 41245 16711
rect 41245 16677 41279 16711
rect 41279 16677 41288 16711
rect 41236 16668 41288 16677
rect 41328 16668 41380 16720
rect 46112 16668 46164 16720
rect 40500 16643 40552 16652
rect 40500 16609 40509 16643
rect 40509 16609 40543 16643
rect 40543 16609 40552 16643
rect 40500 16600 40552 16609
rect 40592 16643 40644 16652
rect 40592 16609 40601 16643
rect 40601 16609 40635 16643
rect 40635 16609 40644 16643
rect 40592 16600 40644 16609
rect 41144 16600 41196 16652
rect 34060 16464 34112 16516
rect 36360 16464 36412 16516
rect 36452 16464 36504 16516
rect 37004 16464 37056 16516
rect 38292 16464 38344 16516
rect 39764 16464 39816 16516
rect 41604 16532 41656 16584
rect 49148 16532 49200 16584
rect 34520 16396 34572 16448
rect 34980 16396 35032 16448
rect 36544 16396 36596 16448
rect 36728 16396 36780 16448
rect 38384 16396 38436 16448
rect 38660 16396 38712 16448
rect 40040 16439 40092 16448
rect 40040 16405 40049 16439
rect 40049 16405 40083 16439
rect 40083 16405 40092 16439
rect 40040 16396 40092 16405
rect 41328 16396 41380 16448
rect 48780 16396 48832 16448
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 27950 16294 28002 16346
rect 28014 16294 28066 16346
rect 28078 16294 28130 16346
rect 28142 16294 28194 16346
rect 28206 16294 28258 16346
rect 37950 16294 38002 16346
rect 38014 16294 38066 16346
rect 38078 16294 38130 16346
rect 38142 16294 38194 16346
rect 38206 16294 38258 16346
rect 47950 16294 48002 16346
rect 48014 16294 48066 16346
rect 48078 16294 48130 16346
rect 48142 16294 48194 16346
rect 48206 16294 48258 16346
rect 8392 16192 8444 16244
rect 9312 16235 9364 16244
rect 9312 16201 9321 16235
rect 9321 16201 9355 16235
rect 9355 16201 9364 16235
rect 9312 16192 9364 16201
rect 10324 16192 10376 16244
rect 11520 16192 11572 16244
rect 14556 16192 14608 16244
rect 11152 16124 11204 16176
rect 11244 16124 11296 16176
rect 10784 16056 10836 16108
rect 10876 16056 10928 16108
rect 12440 16056 12492 16108
rect 1308 15988 1360 16040
rect 4160 15988 4212 16040
rect 8484 16031 8536 16040
rect 8484 15997 8493 16031
rect 8493 15997 8527 16031
rect 8527 15997 8536 16031
rect 8484 15988 8536 15997
rect 12992 16124 13044 16176
rect 14924 16192 14976 16244
rect 18328 16192 18380 16244
rect 19064 16192 19116 16244
rect 22008 16192 22060 16244
rect 24860 16192 24912 16244
rect 15936 16167 15988 16176
rect 15936 16133 15945 16167
rect 15945 16133 15979 16167
rect 15979 16133 15988 16167
rect 15936 16124 15988 16133
rect 17040 16056 17092 16108
rect 18420 16056 18472 16108
rect 11060 15988 11112 16040
rect 11980 15920 12032 15972
rect 12532 16031 12584 16040
rect 12532 15997 12541 16031
rect 12541 15997 12575 16031
rect 12575 15997 12584 16031
rect 12532 15988 12584 15997
rect 12900 15988 12952 16040
rect 14556 15988 14608 16040
rect 14832 16031 14884 16040
rect 14832 15997 14841 16031
rect 14841 15997 14875 16031
rect 14875 15997 14884 16031
rect 14832 15988 14884 15997
rect 15016 16031 15068 16040
rect 15016 15997 15025 16031
rect 15025 15997 15059 16031
rect 15059 15997 15068 16031
rect 15016 15988 15068 15997
rect 15200 15988 15252 16040
rect 13636 15920 13688 15972
rect 15844 16031 15896 16040
rect 15844 15997 15853 16031
rect 15853 15997 15887 16031
rect 15887 15997 15896 16031
rect 15844 15988 15896 15997
rect 15936 15988 15988 16040
rect 18880 16124 18932 16176
rect 20812 16124 20864 16176
rect 21548 16124 21600 16176
rect 23572 16124 23624 16176
rect 23664 16124 23716 16176
rect 26424 16192 26476 16244
rect 26884 16192 26936 16244
rect 18604 16056 18656 16108
rect 16488 15920 16540 15972
rect 16948 15920 17000 15972
rect 22744 15988 22796 16040
rect 26792 16124 26844 16176
rect 27620 16167 27672 16176
rect 27620 16133 27629 16167
rect 27629 16133 27663 16167
rect 27663 16133 27672 16167
rect 27620 16124 27672 16133
rect 30748 16192 30800 16244
rect 30932 16235 30984 16244
rect 30932 16201 30941 16235
rect 30941 16201 30975 16235
rect 30975 16201 30984 16235
rect 30932 16192 30984 16201
rect 31024 16235 31076 16244
rect 31024 16201 31033 16235
rect 31033 16201 31067 16235
rect 31067 16201 31076 16235
rect 31024 16192 31076 16201
rect 33968 16235 34020 16244
rect 33968 16201 33977 16235
rect 33977 16201 34011 16235
rect 34011 16201 34020 16235
rect 33968 16192 34020 16201
rect 34520 16192 34572 16244
rect 24584 16099 24636 16108
rect 24584 16065 24593 16099
rect 24593 16065 24627 16099
rect 24627 16065 24636 16099
rect 24584 16056 24636 16065
rect 25964 16056 26016 16108
rect 26608 16056 26660 16108
rect 28356 16099 28408 16108
rect 28356 16065 28365 16099
rect 28365 16065 28399 16099
rect 28399 16065 28408 16099
rect 28356 16056 28408 16065
rect 24124 15988 24176 16040
rect 26056 15988 26108 16040
rect 26240 15988 26292 16040
rect 27436 15988 27488 16040
rect 19064 15920 19116 15972
rect 9220 15852 9272 15904
rect 10232 15852 10284 15904
rect 11060 15852 11112 15904
rect 11888 15852 11940 15904
rect 15844 15852 15896 15904
rect 16672 15852 16724 15904
rect 16856 15895 16908 15904
rect 16856 15861 16865 15895
rect 16865 15861 16899 15895
rect 16899 15861 16908 15895
rect 16856 15852 16908 15861
rect 17132 15895 17184 15904
rect 17132 15861 17141 15895
rect 17141 15861 17175 15895
rect 17175 15861 17184 15895
rect 17132 15852 17184 15861
rect 20536 15852 20588 15904
rect 22836 15963 22888 15972
rect 22836 15929 22845 15963
rect 22845 15929 22879 15963
rect 22879 15929 22888 15963
rect 22836 15920 22888 15929
rect 24032 15920 24084 15972
rect 26424 15920 26476 15972
rect 28632 16031 28684 16040
rect 28632 15997 28641 16031
rect 28641 15997 28675 16031
rect 28675 15997 28684 16031
rect 28632 15988 28684 15997
rect 29092 15988 29144 16040
rect 29276 15988 29328 16040
rect 31484 16056 31536 16108
rect 33416 16124 33468 16176
rect 35164 16192 35216 16244
rect 36912 16192 36964 16244
rect 40040 16192 40092 16244
rect 33324 16056 33376 16108
rect 22284 15852 22336 15904
rect 25320 15852 25372 15904
rect 25964 15852 26016 15904
rect 26608 15895 26660 15904
rect 26608 15861 26617 15895
rect 26617 15861 26651 15895
rect 26651 15861 26660 15895
rect 26608 15852 26660 15861
rect 26700 15852 26752 15904
rect 29736 15852 29788 15904
rect 31852 15988 31904 16040
rect 32772 15988 32824 16040
rect 35440 16124 35492 16176
rect 37464 16124 37516 16176
rect 36452 16056 36504 16108
rect 38568 16124 38620 16176
rect 39764 16124 39816 16176
rect 41328 16124 41380 16176
rect 48688 16056 48740 16108
rect 49056 16099 49108 16108
rect 49056 16065 49065 16099
rect 49065 16065 49099 16099
rect 49099 16065 49108 16099
rect 49056 16056 49108 16065
rect 30840 15920 30892 15972
rect 32404 15920 32456 15972
rect 32588 15920 32640 15972
rect 34796 15988 34848 16040
rect 34888 15988 34940 16040
rect 36820 15988 36872 16040
rect 37280 15988 37332 16040
rect 40316 15988 40368 16040
rect 40592 15988 40644 16040
rect 41052 16031 41104 16040
rect 41052 15997 41061 16031
rect 41061 15997 41095 16031
rect 41095 15997 41104 16031
rect 41052 15988 41104 15997
rect 30564 15895 30616 15904
rect 30564 15861 30573 15895
rect 30573 15861 30607 15895
rect 30607 15861 30616 15895
rect 30564 15852 30616 15861
rect 31484 15852 31536 15904
rect 31668 15852 31720 15904
rect 33416 15852 33468 15904
rect 37740 15920 37792 15972
rect 49240 15963 49292 15972
rect 49240 15929 49249 15963
rect 49249 15929 49283 15963
rect 49283 15929 49292 15963
rect 49240 15920 49292 15929
rect 37372 15852 37424 15904
rect 41604 15895 41656 15904
rect 41604 15861 41613 15895
rect 41613 15861 41647 15895
rect 41647 15861 41656 15895
rect 41604 15852 41656 15861
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 32950 15750 33002 15802
rect 33014 15750 33066 15802
rect 33078 15750 33130 15802
rect 33142 15750 33194 15802
rect 33206 15750 33258 15802
rect 42950 15750 43002 15802
rect 43014 15750 43066 15802
rect 43078 15750 43130 15802
rect 43142 15750 43194 15802
rect 43206 15750 43258 15802
rect 10784 15648 10836 15700
rect 12072 15580 12124 15632
rect 14832 15648 14884 15700
rect 15476 15580 15528 15632
rect 1308 15512 1360 15564
rect 10600 15512 10652 15564
rect 12808 15512 12860 15564
rect 13452 15555 13504 15564
rect 13452 15521 13461 15555
rect 13461 15521 13495 15555
rect 13495 15521 13504 15555
rect 13452 15512 13504 15521
rect 10416 15444 10468 15496
rect 12716 15444 12768 15496
rect 14832 15555 14884 15564
rect 14832 15521 14841 15555
rect 14841 15521 14875 15555
rect 14875 15521 14884 15555
rect 14832 15512 14884 15521
rect 15384 15512 15436 15564
rect 15936 15580 15988 15632
rect 16580 15648 16632 15700
rect 17132 15648 17184 15700
rect 18512 15648 18564 15700
rect 19432 15648 19484 15700
rect 19892 15691 19944 15700
rect 19892 15657 19901 15691
rect 19901 15657 19935 15691
rect 19935 15657 19944 15691
rect 19892 15648 19944 15657
rect 15844 15444 15896 15496
rect 16948 15580 17000 15632
rect 16488 15512 16540 15564
rect 19156 15580 19208 15632
rect 21732 15648 21784 15700
rect 22468 15691 22520 15700
rect 22468 15657 22477 15691
rect 22477 15657 22511 15691
rect 22511 15657 22520 15691
rect 22468 15648 22520 15657
rect 23480 15648 23532 15700
rect 26608 15648 26660 15700
rect 26884 15648 26936 15700
rect 27344 15648 27396 15700
rect 32588 15648 32640 15700
rect 34152 15648 34204 15700
rect 36820 15648 36872 15700
rect 37004 15648 37056 15700
rect 37832 15648 37884 15700
rect 41604 15648 41656 15700
rect 48688 15648 48740 15700
rect 17316 15555 17368 15564
rect 17316 15521 17325 15555
rect 17325 15521 17359 15555
rect 17359 15521 17368 15555
rect 17316 15512 17368 15521
rect 6552 15351 6604 15360
rect 6552 15317 6561 15351
rect 6561 15317 6595 15351
rect 6595 15317 6604 15351
rect 6552 15308 6604 15317
rect 11704 15376 11756 15428
rect 11796 15308 11848 15360
rect 12532 15351 12584 15360
rect 12532 15317 12541 15351
rect 12541 15317 12575 15351
rect 12575 15317 12584 15351
rect 12532 15308 12584 15317
rect 13636 15376 13688 15428
rect 17868 15376 17920 15428
rect 19800 15444 19852 15496
rect 28816 15580 28868 15632
rect 21364 15512 21416 15564
rect 21088 15444 21140 15496
rect 21732 15512 21784 15564
rect 21916 15512 21968 15564
rect 23848 15512 23900 15564
rect 23940 15512 23992 15564
rect 25044 15512 25096 15564
rect 25320 15555 25372 15564
rect 25320 15521 25329 15555
rect 25329 15521 25363 15555
rect 25363 15521 25372 15555
rect 25320 15512 25372 15521
rect 26240 15512 26292 15564
rect 26516 15555 26568 15564
rect 26516 15521 26525 15555
rect 26525 15521 26559 15555
rect 26559 15521 26568 15555
rect 26516 15512 26568 15521
rect 26608 15512 26660 15564
rect 30748 15555 30800 15564
rect 30748 15521 30757 15555
rect 30757 15521 30791 15555
rect 30791 15521 30800 15555
rect 30748 15512 30800 15521
rect 31484 15512 31536 15564
rect 21548 15487 21600 15496
rect 21548 15453 21557 15487
rect 21557 15453 21591 15487
rect 21591 15453 21600 15487
rect 21548 15444 21600 15453
rect 27160 15444 27212 15496
rect 27804 15487 27856 15496
rect 27804 15453 27813 15487
rect 27813 15453 27847 15487
rect 27847 15453 27856 15487
rect 27804 15444 27856 15453
rect 30472 15487 30524 15496
rect 30472 15453 30481 15487
rect 30481 15453 30515 15487
rect 30515 15453 30524 15487
rect 30472 15444 30524 15453
rect 32220 15512 32272 15564
rect 33508 15512 33560 15564
rect 34152 15512 34204 15564
rect 36360 15512 36412 15564
rect 32680 15444 32732 15496
rect 34520 15444 34572 15496
rect 34888 15487 34940 15496
rect 34888 15453 34897 15487
rect 34897 15453 34931 15487
rect 34931 15453 34940 15487
rect 34888 15444 34940 15453
rect 37464 15444 37516 15496
rect 40316 15555 40368 15564
rect 40316 15521 40325 15555
rect 40325 15521 40359 15555
rect 40359 15521 40368 15555
rect 40316 15512 40368 15521
rect 49332 15487 49384 15496
rect 49332 15453 49341 15487
rect 49341 15453 49375 15487
rect 49375 15453 49384 15487
rect 49332 15444 49384 15453
rect 14464 15308 14516 15360
rect 15476 15308 15528 15360
rect 16028 15308 16080 15360
rect 20260 15351 20312 15360
rect 20260 15317 20269 15351
rect 20269 15317 20303 15351
rect 20303 15317 20312 15351
rect 20260 15308 20312 15317
rect 25596 15376 25648 15428
rect 26332 15419 26384 15428
rect 26332 15385 26341 15419
rect 26341 15385 26375 15419
rect 26375 15385 26384 15419
rect 26332 15376 26384 15385
rect 27344 15376 27396 15428
rect 27712 15376 27764 15428
rect 30380 15376 30432 15428
rect 26976 15351 27028 15360
rect 26976 15317 26985 15351
rect 26985 15317 27019 15351
rect 27019 15317 27028 15351
rect 26976 15308 27028 15317
rect 27436 15351 27488 15360
rect 27436 15317 27445 15351
rect 27445 15317 27479 15351
rect 27479 15317 27488 15351
rect 27436 15308 27488 15317
rect 29276 15351 29328 15360
rect 29276 15317 29285 15351
rect 29285 15317 29319 15351
rect 29319 15317 29328 15351
rect 29276 15308 29328 15317
rect 31116 15308 31168 15360
rect 31484 15308 31536 15360
rect 31668 15308 31720 15360
rect 32680 15351 32732 15360
rect 32680 15317 32689 15351
rect 32689 15317 32723 15351
rect 32723 15317 32732 15351
rect 32680 15308 32732 15317
rect 33876 15351 33928 15360
rect 33876 15317 33885 15351
rect 33885 15317 33919 15351
rect 33919 15317 33928 15351
rect 33876 15308 33928 15317
rect 36452 15376 36504 15428
rect 37372 15376 37424 15428
rect 36084 15308 36136 15360
rect 36544 15308 36596 15360
rect 37096 15351 37148 15360
rect 37096 15317 37105 15351
rect 37105 15317 37139 15351
rect 37139 15317 37148 15351
rect 37096 15308 37148 15317
rect 39764 15376 39816 15428
rect 41328 15376 41380 15428
rect 41052 15308 41104 15360
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 27950 15206 28002 15258
rect 28014 15206 28066 15258
rect 28078 15206 28130 15258
rect 28142 15206 28194 15258
rect 28206 15206 28258 15258
rect 37950 15206 38002 15258
rect 38014 15206 38066 15258
rect 38078 15206 38130 15258
rect 38142 15206 38194 15258
rect 38206 15206 38258 15258
rect 47950 15206 48002 15258
rect 48014 15206 48066 15258
rect 48078 15206 48130 15258
rect 48142 15206 48194 15258
rect 48206 15206 48258 15258
rect 9220 15104 9272 15156
rect 9588 15036 9640 15088
rect 11152 15079 11204 15088
rect 11152 15045 11161 15079
rect 11161 15045 11195 15079
rect 11195 15045 11204 15079
rect 11152 15036 11204 15045
rect 12348 15036 12400 15088
rect 12992 15104 13044 15156
rect 6552 14968 6604 15020
rect 1308 14900 1360 14952
rect 10048 14943 10100 14952
rect 10048 14909 10057 14943
rect 10057 14909 10091 14943
rect 10091 14909 10100 14943
rect 10048 14900 10100 14909
rect 11152 14900 11204 14952
rect 12348 14943 12400 14952
rect 12348 14909 12357 14943
rect 12357 14909 12391 14943
rect 12391 14909 12400 14943
rect 12348 14900 12400 14909
rect 11428 14832 11480 14884
rect 11980 14832 12032 14884
rect 12808 14832 12860 14884
rect 10968 14764 11020 14816
rect 11704 14764 11756 14816
rect 12992 14764 13044 14816
rect 13544 15036 13596 15088
rect 14556 15104 14608 15156
rect 14004 15036 14056 15088
rect 13912 14900 13964 14952
rect 15568 15147 15620 15156
rect 15568 15113 15577 15147
rect 15577 15113 15611 15147
rect 15611 15113 15620 15147
rect 15568 15104 15620 15113
rect 19432 15104 19484 15156
rect 19524 15147 19576 15156
rect 19524 15113 19533 15147
rect 19533 15113 19567 15147
rect 19567 15113 19576 15147
rect 19524 15104 19576 15113
rect 15660 15036 15712 15088
rect 16488 15036 16540 15088
rect 19984 15104 20036 15156
rect 21824 15147 21876 15156
rect 20812 15036 20864 15088
rect 17224 15011 17276 15020
rect 17224 14977 17233 15011
rect 17233 14977 17267 15011
rect 17267 14977 17276 15011
rect 17224 14968 17276 14977
rect 16120 14943 16172 14952
rect 16120 14909 16129 14943
rect 16129 14909 16163 14943
rect 16163 14909 16172 14943
rect 16120 14900 16172 14909
rect 16764 14900 16816 14952
rect 18604 14968 18656 15020
rect 19248 14968 19300 15020
rect 20904 14968 20956 15020
rect 21824 15113 21833 15147
rect 21833 15113 21867 15147
rect 21867 15113 21876 15147
rect 21824 15104 21876 15113
rect 22652 15104 22704 15156
rect 23480 15104 23532 15156
rect 23756 15104 23808 15156
rect 21272 15036 21324 15088
rect 25044 15036 25096 15088
rect 15936 14832 15988 14884
rect 16580 14832 16632 14884
rect 18880 14943 18932 14952
rect 18880 14909 18889 14943
rect 18889 14909 18923 14943
rect 18923 14909 18932 14943
rect 18880 14900 18932 14909
rect 20076 14943 20128 14952
rect 20076 14909 20085 14943
rect 20085 14909 20119 14943
rect 20119 14909 20128 14943
rect 20076 14900 20128 14909
rect 20536 14900 20588 14952
rect 23296 15011 23348 15020
rect 23296 14977 23305 15011
rect 23305 14977 23339 15011
rect 23339 14977 23348 15011
rect 23296 14968 23348 14977
rect 25412 14968 25464 15020
rect 25504 14968 25556 15020
rect 27068 14968 27120 15020
rect 17500 14832 17552 14884
rect 21732 14832 21784 14884
rect 15844 14764 15896 14816
rect 17408 14764 17460 14816
rect 19340 14764 19392 14816
rect 19616 14764 19668 14816
rect 19892 14764 19944 14816
rect 24584 14943 24636 14952
rect 24584 14909 24593 14943
rect 24593 14909 24627 14943
rect 24627 14909 24636 14943
rect 24584 14900 24636 14909
rect 24676 14943 24728 14952
rect 24676 14909 24685 14943
rect 24685 14909 24719 14943
rect 24719 14909 24728 14943
rect 24676 14900 24728 14909
rect 24768 14900 24820 14952
rect 24308 14832 24360 14884
rect 25044 14764 25096 14816
rect 25596 14807 25648 14816
rect 25596 14773 25605 14807
rect 25605 14773 25639 14807
rect 25639 14773 25648 14807
rect 25596 14764 25648 14773
rect 27528 15036 27580 15088
rect 28356 15036 28408 15088
rect 29276 15036 29328 15088
rect 29736 15147 29788 15156
rect 29736 15113 29745 15147
rect 29745 15113 29779 15147
rect 29779 15113 29788 15147
rect 29736 15104 29788 15113
rect 30288 15104 30340 15156
rect 30012 15036 30064 15088
rect 30196 15036 30248 15088
rect 27344 14900 27396 14952
rect 29828 14900 29880 14952
rect 26884 14764 26936 14816
rect 28448 14764 28500 14816
rect 29828 14764 29880 14816
rect 30656 15147 30708 15156
rect 30656 15113 30665 15147
rect 30665 15113 30699 15147
rect 30699 15113 30708 15147
rect 30656 15104 30708 15113
rect 30932 15104 30984 15156
rect 31300 15104 31352 15156
rect 31576 15104 31628 15156
rect 33876 15147 33928 15156
rect 33876 15113 33885 15147
rect 33885 15113 33919 15147
rect 33919 15113 33928 15147
rect 33876 15104 33928 15113
rect 34704 15147 34756 15156
rect 34704 15113 34713 15147
rect 34713 15113 34747 15147
rect 34747 15113 34756 15147
rect 34704 15104 34756 15113
rect 37280 15104 37332 15156
rect 31484 15036 31536 15088
rect 30932 14968 30984 15020
rect 37188 15036 37240 15088
rect 38568 15104 38620 15156
rect 40132 15147 40184 15156
rect 40132 15113 40141 15147
rect 40141 15113 40175 15147
rect 40175 15113 40184 15147
rect 40132 15104 40184 15113
rect 40316 15104 40368 15156
rect 35900 14968 35952 15020
rect 36176 14968 36228 15020
rect 36452 14968 36504 15020
rect 37832 15036 37884 15088
rect 48412 15036 48464 15088
rect 37464 15011 37516 15020
rect 37464 14977 37473 15011
rect 37473 14977 37507 15011
rect 37507 14977 37516 15011
rect 37464 14968 37516 14977
rect 39856 14968 39908 15020
rect 49056 15011 49108 15020
rect 49056 14977 49065 15011
rect 49065 14977 49099 15011
rect 49099 14977 49108 15011
rect 49056 14968 49108 14977
rect 30840 14900 30892 14952
rect 33876 14900 33928 14952
rect 33968 14943 34020 14952
rect 33968 14909 33977 14943
rect 33977 14909 34011 14943
rect 34011 14909 34020 14943
rect 33968 14900 34020 14909
rect 34060 14943 34112 14952
rect 34060 14909 34069 14943
rect 34069 14909 34103 14943
rect 34103 14909 34112 14943
rect 34060 14900 34112 14909
rect 34612 14900 34664 14952
rect 35348 14943 35400 14952
rect 35348 14909 35357 14943
rect 35357 14909 35391 14943
rect 35391 14909 35400 14943
rect 35348 14900 35400 14909
rect 36544 14943 36596 14952
rect 36544 14909 36553 14943
rect 36553 14909 36587 14943
rect 36587 14909 36596 14943
rect 36544 14900 36596 14909
rect 37004 14900 37056 14952
rect 38476 14900 38528 14952
rect 37280 14832 37332 14884
rect 38936 14900 38988 14952
rect 40316 14832 40368 14884
rect 32772 14764 32824 14816
rect 36728 14764 36780 14816
rect 37556 14764 37608 14816
rect 45836 14764 45888 14816
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 32950 14662 33002 14714
rect 33014 14662 33066 14714
rect 33078 14662 33130 14714
rect 33142 14662 33194 14714
rect 33206 14662 33258 14714
rect 42950 14662 43002 14714
rect 43014 14662 43066 14714
rect 43078 14662 43130 14714
rect 43142 14662 43194 14714
rect 43206 14662 43258 14714
rect 10416 14603 10468 14612
rect 10416 14569 10425 14603
rect 10425 14569 10459 14603
rect 10459 14569 10468 14603
rect 10416 14560 10468 14569
rect 11612 14560 11664 14612
rect 12624 14560 12676 14612
rect 13176 14560 13228 14612
rect 17132 14560 17184 14612
rect 17224 14560 17276 14612
rect 17868 14560 17920 14612
rect 18604 14560 18656 14612
rect 1308 14424 1360 14476
rect 13268 14492 13320 14544
rect 14464 14535 14516 14544
rect 14464 14501 14473 14535
rect 14473 14501 14507 14535
rect 14507 14501 14516 14535
rect 14464 14492 14516 14501
rect 14924 14492 14976 14544
rect 18880 14492 18932 14544
rect 12532 14424 12584 14476
rect 10324 14399 10376 14408
rect 10324 14365 10333 14399
rect 10333 14365 10367 14399
rect 10367 14365 10376 14399
rect 10324 14356 10376 14365
rect 10692 14356 10744 14408
rect 9588 14331 9640 14340
rect 9588 14297 9597 14331
rect 9597 14297 9631 14331
rect 9631 14297 9640 14331
rect 9588 14288 9640 14297
rect 12532 14288 12584 14340
rect 12808 14356 12860 14408
rect 14188 14399 14240 14408
rect 14188 14365 14197 14399
rect 14197 14365 14231 14399
rect 14231 14365 14240 14399
rect 14188 14356 14240 14365
rect 16120 14424 16172 14476
rect 17132 14424 17184 14476
rect 17592 14424 17644 14476
rect 19064 14560 19116 14612
rect 21088 14560 21140 14612
rect 21456 14560 21508 14612
rect 23204 14560 23256 14612
rect 24032 14560 24084 14612
rect 25136 14560 25188 14612
rect 33968 14560 34020 14612
rect 35348 14560 35400 14612
rect 24584 14492 24636 14544
rect 25504 14492 25556 14544
rect 17316 14356 17368 14408
rect 20720 14424 20772 14476
rect 21364 14467 21416 14476
rect 21364 14433 21373 14467
rect 21373 14433 21407 14467
rect 21407 14433 21416 14467
rect 21364 14424 21416 14433
rect 21732 14424 21784 14476
rect 24860 14424 24912 14476
rect 27160 14424 27212 14476
rect 27528 14424 27580 14476
rect 28264 14467 28316 14476
rect 28264 14433 28273 14467
rect 28273 14433 28307 14467
rect 28307 14433 28316 14467
rect 28264 14424 28316 14433
rect 28632 14424 28684 14476
rect 13176 14288 13228 14340
rect 11244 14263 11296 14272
rect 11244 14229 11253 14263
rect 11253 14229 11287 14263
rect 11287 14229 11296 14263
rect 11244 14220 11296 14229
rect 12624 14220 12676 14272
rect 13452 14263 13504 14272
rect 13452 14229 13461 14263
rect 13461 14229 13495 14263
rect 13495 14229 13504 14263
rect 13452 14220 13504 14229
rect 13728 14220 13780 14272
rect 16488 14220 16540 14272
rect 16948 14220 17000 14272
rect 19892 14331 19944 14340
rect 19892 14297 19901 14331
rect 19901 14297 19935 14331
rect 19935 14297 19944 14331
rect 19892 14288 19944 14297
rect 25320 14356 25372 14408
rect 30748 14424 30800 14476
rect 31944 14492 31996 14544
rect 32128 14424 32180 14476
rect 32496 14424 32548 14476
rect 32864 14492 32916 14544
rect 36636 14603 36688 14612
rect 36636 14569 36645 14603
rect 36645 14569 36679 14603
rect 36679 14569 36688 14603
rect 36636 14560 36688 14569
rect 38108 14560 38160 14612
rect 38384 14560 38436 14612
rect 38936 14560 38988 14612
rect 39764 14560 39816 14612
rect 21272 14288 21324 14340
rect 22652 14288 22704 14340
rect 23204 14288 23256 14340
rect 18512 14263 18564 14272
rect 18512 14229 18521 14263
rect 18521 14229 18555 14263
rect 18555 14229 18564 14263
rect 18512 14220 18564 14229
rect 19524 14263 19576 14272
rect 19524 14229 19533 14263
rect 19533 14229 19567 14263
rect 19567 14229 19576 14263
rect 19524 14220 19576 14229
rect 19800 14220 19852 14272
rect 20536 14263 20588 14272
rect 20536 14229 20545 14263
rect 20545 14229 20579 14263
rect 20579 14229 20588 14263
rect 20536 14220 20588 14229
rect 20720 14263 20772 14272
rect 20720 14229 20729 14263
rect 20729 14229 20763 14263
rect 20763 14229 20772 14263
rect 20720 14220 20772 14229
rect 22376 14220 22428 14272
rect 25504 14288 25556 14340
rect 23664 14220 23716 14272
rect 24400 14263 24452 14272
rect 24400 14229 24409 14263
rect 24409 14229 24443 14263
rect 24443 14229 24452 14263
rect 24400 14220 24452 14229
rect 24584 14263 24636 14272
rect 24584 14229 24593 14263
rect 24593 14229 24627 14263
rect 24627 14229 24636 14263
rect 24584 14220 24636 14229
rect 24952 14263 25004 14272
rect 24952 14229 24961 14263
rect 24961 14229 24995 14263
rect 24995 14229 25004 14263
rect 24952 14220 25004 14229
rect 26884 14288 26936 14340
rect 28448 14288 28500 14340
rect 28540 14288 28592 14340
rect 29736 14288 29788 14340
rect 31760 14356 31812 14408
rect 33416 14356 33468 14408
rect 34888 14467 34940 14476
rect 34888 14433 34897 14467
rect 34897 14433 34931 14467
rect 34931 14433 34940 14467
rect 34888 14424 34940 14433
rect 37464 14424 37516 14476
rect 37740 14424 37792 14476
rect 39580 14356 39632 14408
rect 49148 14399 49200 14408
rect 49148 14365 49157 14399
rect 49157 14365 49191 14399
rect 49191 14365 49200 14399
rect 49148 14356 49200 14365
rect 30380 14288 30432 14340
rect 25964 14220 26016 14272
rect 29000 14263 29052 14272
rect 29000 14229 29009 14263
rect 29009 14229 29043 14263
rect 29043 14229 29052 14263
rect 29000 14220 29052 14229
rect 29552 14220 29604 14272
rect 31116 14220 31168 14272
rect 32128 14263 32180 14272
rect 32128 14229 32137 14263
rect 32137 14229 32171 14263
rect 32171 14229 32180 14263
rect 32128 14220 32180 14229
rect 33600 14288 33652 14340
rect 33232 14220 33284 14272
rect 34612 14220 34664 14272
rect 35164 14331 35216 14340
rect 35164 14297 35173 14331
rect 35173 14297 35207 14331
rect 35207 14297 35216 14331
rect 35164 14288 35216 14297
rect 36452 14288 36504 14340
rect 37464 14288 37516 14340
rect 37832 14288 37884 14340
rect 37556 14220 37608 14272
rect 39304 14263 39356 14272
rect 39304 14229 39313 14263
rect 39313 14229 39347 14263
rect 39347 14229 39356 14263
rect 39304 14220 39356 14229
rect 48320 14220 48372 14272
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 27950 14118 28002 14170
rect 28014 14118 28066 14170
rect 28078 14118 28130 14170
rect 28142 14118 28194 14170
rect 28206 14118 28258 14170
rect 37950 14118 38002 14170
rect 38014 14118 38066 14170
rect 38078 14118 38130 14170
rect 38142 14118 38194 14170
rect 38206 14118 38258 14170
rect 47950 14118 48002 14170
rect 48014 14118 48066 14170
rect 48078 14118 48130 14170
rect 48142 14118 48194 14170
rect 48206 14118 48258 14170
rect 10232 14016 10284 14068
rect 10324 14016 10376 14068
rect 10692 14059 10744 14068
rect 10692 14025 10701 14059
rect 10701 14025 10735 14059
rect 10735 14025 10744 14059
rect 10692 14016 10744 14025
rect 12164 14016 12216 14068
rect 14648 14016 14700 14068
rect 15200 14016 15252 14068
rect 16580 14016 16632 14068
rect 17500 14059 17552 14068
rect 17500 14025 17509 14059
rect 17509 14025 17543 14059
rect 17543 14025 17552 14059
rect 17500 14016 17552 14025
rect 18420 14016 18472 14068
rect 18972 14016 19024 14068
rect 19800 14016 19852 14068
rect 22376 14016 22428 14068
rect 22652 14016 22704 14068
rect 23848 14016 23900 14068
rect 25504 14016 25556 14068
rect 11244 13948 11296 14000
rect 14004 13948 14056 14000
rect 3516 13923 3568 13932
rect 3516 13889 3525 13923
rect 3525 13889 3559 13923
rect 3559 13889 3568 13923
rect 3516 13880 3568 13889
rect 1308 13812 1360 13864
rect 9588 13812 9640 13864
rect 11520 13812 11572 13864
rect 12348 13880 12400 13932
rect 15844 13880 15896 13932
rect 19524 13948 19576 14000
rect 10048 13744 10100 13796
rect 12808 13812 12860 13864
rect 13360 13812 13412 13864
rect 14004 13812 14056 13864
rect 14924 13812 14976 13864
rect 16672 13880 16724 13932
rect 19432 13880 19484 13932
rect 16212 13855 16264 13864
rect 16212 13821 16221 13855
rect 16221 13821 16255 13855
rect 16255 13821 16264 13855
rect 16212 13812 16264 13821
rect 16488 13812 16540 13864
rect 17684 13855 17736 13864
rect 17684 13821 17693 13855
rect 17693 13821 17727 13855
rect 17727 13821 17736 13855
rect 17684 13812 17736 13821
rect 12532 13744 12584 13796
rect 10876 13676 10928 13728
rect 15752 13744 15804 13796
rect 15384 13676 15436 13728
rect 18788 13744 18840 13796
rect 18972 13812 19024 13864
rect 20720 13812 20772 13864
rect 24032 13948 24084 14000
rect 25136 13991 25188 14000
rect 25136 13957 25145 13991
rect 25145 13957 25179 13991
rect 25179 13957 25188 13991
rect 25136 13948 25188 13957
rect 26516 14016 26568 14068
rect 24860 13923 24912 13932
rect 24860 13889 24869 13923
rect 24869 13889 24903 13923
rect 24903 13889 24912 13923
rect 24860 13880 24912 13889
rect 26792 13880 26844 13932
rect 28080 13880 28132 13932
rect 28908 13991 28960 14000
rect 28908 13957 28917 13991
rect 28917 13957 28951 13991
rect 28951 13957 28960 13991
rect 28908 13948 28960 13957
rect 29276 13880 29328 13932
rect 30012 14016 30064 14068
rect 30472 14016 30524 14068
rect 31116 14059 31168 14068
rect 31116 14025 31125 14059
rect 31125 14025 31159 14059
rect 31159 14025 31168 14059
rect 31116 14016 31168 14025
rect 36452 14016 36504 14068
rect 41512 14016 41564 14068
rect 47032 14016 47084 14068
rect 48412 14059 48464 14068
rect 48412 14025 48421 14059
rect 48421 14025 48455 14059
rect 48455 14025 48464 14059
rect 48412 14016 48464 14025
rect 49240 14059 49292 14068
rect 49240 14025 49249 14059
rect 49249 14025 49283 14059
rect 49283 14025 49292 14059
rect 49240 14016 49292 14025
rect 31392 13948 31444 14000
rect 21364 13812 21416 13864
rect 22008 13855 22060 13864
rect 22008 13821 22017 13855
rect 22017 13821 22051 13855
rect 22051 13821 22060 13855
rect 22008 13812 22060 13821
rect 22284 13855 22336 13864
rect 22284 13821 22293 13855
rect 22293 13821 22327 13855
rect 22327 13821 22336 13855
rect 22284 13812 22336 13821
rect 24216 13855 24268 13864
rect 24216 13821 24225 13855
rect 24225 13821 24259 13855
rect 24259 13821 24268 13855
rect 24216 13812 24268 13821
rect 28632 13812 28684 13864
rect 32864 13948 32916 14000
rect 34336 13948 34388 14000
rect 32312 13855 32364 13864
rect 32312 13821 32321 13855
rect 32321 13821 32355 13855
rect 32355 13821 32364 13855
rect 32312 13812 32364 13821
rect 31300 13744 31352 13796
rect 32220 13744 32272 13796
rect 32680 13812 32732 13864
rect 34980 13923 35032 13932
rect 34980 13889 34989 13923
rect 34989 13889 35023 13923
rect 35023 13889 35032 13923
rect 34980 13880 35032 13889
rect 37556 13948 37608 14000
rect 37648 13948 37700 14000
rect 39304 13948 39356 14000
rect 49148 13991 49200 14000
rect 49148 13957 49157 13991
rect 49157 13957 49191 13991
rect 49191 13957 49200 13991
rect 49148 13948 49200 13957
rect 33876 13744 33928 13796
rect 35348 13744 35400 13796
rect 39396 13880 39448 13932
rect 39764 13880 39816 13932
rect 45836 13923 45888 13932
rect 45836 13889 45845 13923
rect 45845 13889 45879 13923
rect 45879 13889 45888 13923
rect 45836 13880 45888 13889
rect 48228 13880 48280 13932
rect 36176 13855 36228 13864
rect 36176 13821 36185 13855
rect 36185 13821 36219 13855
rect 36219 13821 36228 13855
rect 36176 13812 36228 13821
rect 36636 13812 36688 13864
rect 37740 13744 37792 13796
rect 46480 13812 46532 13864
rect 19800 13676 19852 13728
rect 20444 13676 20496 13728
rect 23848 13676 23900 13728
rect 30840 13676 30892 13728
rect 31208 13676 31260 13728
rect 33324 13676 33376 13728
rect 33692 13676 33744 13728
rect 38384 13676 38436 13728
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 32950 13574 33002 13626
rect 33014 13574 33066 13626
rect 33078 13574 33130 13626
rect 33142 13574 33194 13626
rect 33206 13574 33258 13626
rect 42950 13574 43002 13626
rect 43014 13574 43066 13626
rect 43078 13574 43130 13626
rect 43142 13574 43194 13626
rect 43206 13574 43258 13626
rect 14924 13515 14976 13524
rect 14924 13481 14933 13515
rect 14933 13481 14967 13515
rect 14967 13481 14976 13515
rect 14924 13472 14976 13481
rect 15108 13472 15160 13524
rect 12532 13447 12584 13456
rect 12532 13413 12541 13447
rect 12541 13413 12575 13447
rect 12575 13413 12584 13447
rect 12532 13404 12584 13413
rect 14832 13404 14884 13456
rect 15476 13404 15528 13456
rect 17408 13472 17460 13524
rect 17684 13472 17736 13524
rect 20260 13472 20312 13524
rect 20352 13472 20404 13524
rect 23388 13472 23440 13524
rect 23480 13472 23532 13524
rect 24124 13472 24176 13524
rect 25228 13472 25280 13524
rect 28080 13515 28132 13524
rect 28080 13481 28089 13515
rect 28089 13481 28123 13515
rect 28123 13481 28132 13515
rect 28080 13472 28132 13481
rect 28356 13472 28408 13524
rect 11060 13336 11112 13388
rect 14740 13336 14792 13388
rect 17776 13404 17828 13456
rect 2780 13311 2832 13320
rect 2780 13277 2789 13311
rect 2789 13277 2823 13311
rect 2823 13277 2832 13311
rect 2780 13268 2832 13277
rect 12808 13268 12860 13320
rect 13084 13268 13136 13320
rect 18972 13336 19024 13388
rect 19432 13447 19484 13456
rect 19432 13413 19441 13447
rect 19441 13413 19475 13447
rect 19475 13413 19484 13447
rect 19432 13404 19484 13413
rect 19892 13404 19944 13456
rect 20168 13379 20220 13388
rect 20168 13345 20177 13379
rect 20177 13345 20211 13379
rect 20211 13345 20220 13379
rect 20168 13336 20220 13345
rect 11704 13200 11756 13252
rect 11980 13132 12032 13184
rect 12716 13132 12768 13184
rect 14096 13132 14148 13184
rect 14188 13132 14240 13184
rect 15384 13132 15436 13184
rect 15568 13243 15620 13252
rect 15568 13209 15577 13243
rect 15577 13209 15611 13243
rect 15611 13209 15620 13243
rect 15568 13200 15620 13209
rect 16396 13200 16448 13252
rect 17132 13200 17184 13252
rect 19984 13268 20036 13320
rect 19064 13132 19116 13184
rect 19708 13132 19760 13184
rect 21456 13379 21508 13388
rect 21456 13345 21465 13379
rect 21465 13345 21499 13379
rect 21499 13345 21508 13379
rect 21456 13336 21508 13345
rect 27436 13404 27488 13456
rect 30840 13404 30892 13456
rect 32772 13515 32824 13524
rect 32772 13481 32781 13515
rect 32781 13481 32815 13515
rect 32815 13481 32824 13515
rect 32772 13472 32824 13481
rect 33324 13515 33376 13524
rect 33324 13481 33333 13515
rect 33333 13481 33367 13515
rect 33367 13481 33376 13515
rect 33324 13472 33376 13481
rect 35992 13472 36044 13524
rect 33692 13404 33744 13456
rect 37372 13472 37424 13524
rect 37832 13472 37884 13524
rect 38752 13472 38804 13524
rect 23756 13336 23808 13388
rect 22836 13268 22888 13320
rect 23664 13311 23716 13320
rect 23664 13277 23673 13311
rect 23673 13277 23707 13311
rect 23707 13277 23716 13311
rect 23664 13268 23716 13277
rect 24952 13268 25004 13320
rect 25964 13336 26016 13388
rect 29644 13336 29696 13388
rect 30288 13379 30340 13388
rect 30288 13345 30297 13379
rect 30297 13345 30331 13379
rect 30331 13345 30340 13379
rect 30288 13336 30340 13345
rect 32312 13336 32364 13388
rect 32496 13336 32548 13388
rect 32772 13336 32824 13388
rect 32864 13336 32916 13388
rect 35072 13336 35124 13388
rect 35348 13336 35400 13388
rect 25780 13268 25832 13320
rect 28816 13268 28868 13320
rect 29828 13268 29880 13320
rect 33324 13268 33376 13320
rect 33600 13268 33652 13320
rect 37096 13336 37148 13388
rect 24032 13200 24084 13252
rect 24400 13200 24452 13252
rect 20444 13132 20496 13184
rect 20904 13175 20956 13184
rect 20904 13141 20913 13175
rect 20913 13141 20947 13175
rect 20947 13141 20956 13175
rect 20904 13132 20956 13141
rect 21088 13132 21140 13184
rect 21364 13175 21416 13184
rect 21364 13141 21373 13175
rect 21373 13141 21407 13175
rect 21407 13141 21416 13175
rect 21364 13132 21416 13141
rect 21824 13132 21876 13184
rect 23664 13132 23716 13184
rect 24492 13175 24544 13184
rect 24492 13141 24501 13175
rect 24501 13141 24535 13175
rect 24535 13141 24544 13175
rect 26332 13200 26384 13252
rect 24492 13132 24544 13141
rect 26056 13175 26108 13184
rect 26056 13141 26065 13175
rect 26065 13141 26099 13175
rect 26099 13141 26108 13175
rect 26056 13132 26108 13141
rect 26792 13175 26844 13184
rect 26792 13141 26801 13175
rect 26801 13141 26835 13175
rect 26835 13141 26844 13175
rect 26792 13132 26844 13141
rect 28540 13132 28592 13184
rect 29000 13132 29052 13184
rect 29920 13132 29972 13184
rect 33876 13200 33928 13252
rect 34336 13243 34388 13252
rect 34336 13209 34345 13243
rect 34345 13209 34379 13243
rect 34379 13209 34388 13243
rect 34336 13200 34388 13209
rect 35348 13243 35400 13252
rect 35348 13209 35357 13243
rect 35357 13209 35391 13243
rect 35391 13209 35400 13243
rect 35348 13200 35400 13209
rect 36360 13200 36412 13252
rect 37832 13268 37884 13320
rect 41512 13311 41564 13320
rect 41512 13277 41521 13311
rect 41521 13277 41555 13311
rect 41555 13277 41564 13311
rect 41512 13268 41564 13277
rect 46480 13268 46532 13320
rect 36636 13200 36688 13252
rect 49148 13243 49200 13252
rect 49148 13209 49157 13243
rect 49157 13209 49191 13243
rect 49191 13209 49200 13243
rect 49148 13200 49200 13209
rect 34796 13132 34848 13184
rect 35992 13175 36044 13184
rect 35992 13141 36001 13175
rect 36001 13141 36035 13175
rect 36035 13141 36044 13175
rect 35992 13132 36044 13141
rect 36452 13132 36504 13184
rect 37372 13132 37424 13184
rect 37740 13132 37792 13184
rect 46112 13132 46164 13184
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 27950 13030 28002 13082
rect 28014 13030 28066 13082
rect 28078 13030 28130 13082
rect 28142 13030 28194 13082
rect 28206 13030 28258 13082
rect 37950 13030 38002 13082
rect 38014 13030 38066 13082
rect 38078 13030 38130 13082
rect 38142 13030 38194 13082
rect 38206 13030 38258 13082
rect 47950 13030 48002 13082
rect 48014 13030 48066 13082
rect 48078 13030 48130 13082
rect 48142 13030 48194 13082
rect 48206 13030 48258 13082
rect 5448 12928 5500 12980
rect 10968 12928 11020 12980
rect 13360 12928 13412 12980
rect 16028 12928 16080 12980
rect 16396 12928 16448 12980
rect 17132 12928 17184 12980
rect 1308 12860 1360 12912
rect 11704 12860 11756 12912
rect 12072 12903 12124 12912
rect 12072 12869 12081 12903
rect 12081 12869 12115 12903
rect 12115 12869 12124 12903
rect 12072 12860 12124 12869
rect 1216 12792 1268 12844
rect 12532 12792 12584 12844
rect 15108 12860 15160 12912
rect 20536 12928 20588 12980
rect 17960 12860 18012 12912
rect 18328 12860 18380 12912
rect 18788 12860 18840 12912
rect 20904 12928 20956 12980
rect 21824 12928 21876 12980
rect 22744 12928 22796 12980
rect 23112 12971 23164 12980
rect 23112 12937 23121 12971
rect 23121 12937 23155 12971
rect 23155 12937 23164 12971
rect 23112 12928 23164 12937
rect 23480 12928 23532 12980
rect 23848 12928 23900 12980
rect 20996 12860 21048 12912
rect 24768 12928 24820 12980
rect 25044 12928 25096 12980
rect 26332 12928 26384 12980
rect 27344 12928 27396 12980
rect 26792 12860 26844 12912
rect 28448 12928 28500 12980
rect 28724 12860 28776 12912
rect 29552 12903 29604 12912
rect 29552 12869 29561 12903
rect 29561 12869 29595 12903
rect 29595 12869 29604 12903
rect 29552 12860 29604 12869
rect 12716 12792 12768 12844
rect 13084 12835 13136 12844
rect 13084 12801 13093 12835
rect 13093 12801 13127 12835
rect 13127 12801 13136 12835
rect 13084 12792 13136 12801
rect 9864 12724 9916 12776
rect 12256 12767 12308 12776
rect 12256 12733 12265 12767
rect 12265 12733 12299 12767
rect 12299 12733 12308 12767
rect 12256 12724 12308 12733
rect 13360 12767 13412 12776
rect 13360 12733 13369 12767
rect 13369 12733 13403 12767
rect 13403 12733 13412 12767
rect 13360 12724 13412 12733
rect 14096 12724 14148 12776
rect 16212 12792 16264 12844
rect 16488 12792 16540 12844
rect 18972 12792 19024 12844
rect 19616 12835 19668 12844
rect 19616 12801 19625 12835
rect 19625 12801 19659 12835
rect 19659 12801 19668 12835
rect 19616 12792 19668 12801
rect 21916 12792 21968 12844
rect 23020 12835 23072 12844
rect 23020 12801 23029 12835
rect 23029 12801 23063 12835
rect 23063 12801 23072 12835
rect 23020 12792 23072 12801
rect 26240 12792 26292 12844
rect 26976 12792 27028 12844
rect 27160 12835 27212 12844
rect 27160 12801 27169 12835
rect 27169 12801 27203 12835
rect 27203 12801 27212 12835
rect 27160 12792 27212 12801
rect 29368 12792 29420 12844
rect 30012 12835 30064 12844
rect 30012 12801 30021 12835
rect 30021 12801 30055 12835
rect 30055 12801 30064 12835
rect 30012 12792 30064 12801
rect 31392 12792 31444 12844
rect 19524 12724 19576 12776
rect 19708 12767 19760 12776
rect 19708 12733 19717 12767
rect 19717 12733 19751 12767
rect 19751 12733 19760 12767
rect 19708 12724 19760 12733
rect 20904 12724 20956 12776
rect 21180 12724 21232 12776
rect 21364 12724 21416 12776
rect 22100 12724 22152 12776
rect 23388 12724 23440 12776
rect 23848 12767 23900 12776
rect 23848 12733 23857 12767
rect 23857 12733 23891 12767
rect 23891 12733 23900 12767
rect 23848 12724 23900 12733
rect 24124 12767 24176 12776
rect 24124 12733 24133 12767
rect 24133 12733 24167 12767
rect 24167 12733 24176 12767
rect 24124 12724 24176 12733
rect 26516 12724 26568 12776
rect 15660 12656 15712 12708
rect 16488 12656 16540 12708
rect 17684 12656 17736 12708
rect 12624 12588 12676 12640
rect 17408 12588 17460 12640
rect 18696 12588 18748 12640
rect 21456 12588 21508 12640
rect 23480 12588 23532 12640
rect 25872 12699 25924 12708
rect 25872 12665 25881 12699
rect 25881 12665 25915 12699
rect 25915 12665 25924 12699
rect 25872 12656 25924 12665
rect 29552 12724 29604 12776
rect 31760 12971 31812 12980
rect 31760 12937 31769 12971
rect 31769 12937 31803 12971
rect 31803 12937 31812 12971
rect 31760 12928 31812 12937
rect 32404 12928 32456 12980
rect 31760 12792 31812 12844
rect 32772 12971 32824 12980
rect 32772 12937 32781 12971
rect 32781 12937 32815 12971
rect 32815 12937 32824 12971
rect 32772 12928 32824 12937
rect 33784 12971 33836 12980
rect 33784 12937 33793 12971
rect 33793 12937 33827 12971
rect 33827 12937 33836 12971
rect 33784 12928 33836 12937
rect 34060 12928 34112 12980
rect 34428 12928 34480 12980
rect 35532 12928 35584 12980
rect 35808 12971 35860 12980
rect 35808 12937 35817 12971
rect 35817 12937 35851 12971
rect 35851 12937 35860 12971
rect 35808 12928 35860 12937
rect 36084 12928 36136 12980
rect 36820 12928 36872 12980
rect 34888 12903 34940 12912
rect 32312 12724 32364 12776
rect 34888 12869 34897 12903
rect 34897 12869 34931 12903
rect 34931 12869 34940 12903
rect 34888 12860 34940 12869
rect 36452 12860 36504 12912
rect 36728 12860 36780 12912
rect 37832 12928 37884 12980
rect 37740 12903 37792 12912
rect 37740 12869 37749 12903
rect 37749 12869 37783 12903
rect 37783 12869 37792 12903
rect 37740 12860 37792 12869
rect 38752 12860 38804 12912
rect 39948 12860 40000 12912
rect 34060 12835 34112 12844
rect 34060 12801 34069 12835
rect 34069 12801 34103 12835
rect 34103 12801 34112 12835
rect 34060 12792 34112 12801
rect 35164 12792 35216 12844
rect 33508 12724 33560 12776
rect 35624 12724 35676 12776
rect 37372 12792 37424 12844
rect 46112 12835 46164 12844
rect 46112 12801 46121 12835
rect 46121 12801 46155 12835
rect 46155 12801 46164 12835
rect 46112 12792 46164 12801
rect 47032 12792 47084 12844
rect 49148 12835 49200 12844
rect 49148 12801 49157 12835
rect 49157 12801 49191 12835
rect 49191 12801 49200 12835
rect 49148 12792 49200 12801
rect 27160 12588 27212 12640
rect 29368 12588 29420 12640
rect 34520 12656 34572 12708
rect 37372 12656 37424 12708
rect 47032 12656 47084 12708
rect 33324 12588 33376 12640
rect 34336 12588 34388 12640
rect 36084 12588 36136 12640
rect 39488 12588 39540 12640
rect 47952 12588 48004 12640
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 32950 12486 33002 12538
rect 33014 12486 33066 12538
rect 33078 12486 33130 12538
rect 33142 12486 33194 12538
rect 33206 12486 33258 12538
rect 42950 12486 43002 12538
rect 43014 12486 43066 12538
rect 43078 12486 43130 12538
rect 43142 12486 43194 12538
rect 43206 12486 43258 12538
rect 12440 12384 12492 12436
rect 13268 12384 13320 12436
rect 16120 12384 16172 12436
rect 19340 12384 19392 12436
rect 15936 12316 15988 12368
rect 22928 12384 22980 12436
rect 5448 12248 5500 12300
rect 11060 12248 11112 12300
rect 12716 12248 12768 12300
rect 14924 12248 14976 12300
rect 17224 12248 17276 12300
rect 1308 12180 1360 12232
rect 15844 12180 15896 12232
rect 17132 12223 17184 12232
rect 17132 12189 17141 12223
rect 17141 12189 17175 12223
rect 17175 12189 17184 12223
rect 17132 12180 17184 12189
rect 17960 12223 18012 12232
rect 17960 12189 17969 12223
rect 17969 12189 18003 12223
rect 18003 12189 18012 12223
rect 17960 12180 18012 12189
rect 10048 12112 10100 12164
rect 11704 12112 11756 12164
rect 11244 12087 11296 12096
rect 11244 12053 11253 12087
rect 11253 12053 11287 12087
rect 11287 12053 11296 12087
rect 11244 12044 11296 12053
rect 12532 12112 12584 12164
rect 13728 12155 13780 12164
rect 13728 12121 13737 12155
rect 13737 12121 13771 12155
rect 13771 12121 13780 12155
rect 13728 12112 13780 12121
rect 12716 12044 12768 12096
rect 14740 12044 14792 12096
rect 15016 12112 15068 12164
rect 16856 12112 16908 12164
rect 19340 12248 19392 12300
rect 19524 12180 19576 12232
rect 19984 12291 20036 12300
rect 19984 12257 19993 12291
rect 19993 12257 20027 12291
rect 20027 12257 20036 12291
rect 19984 12248 20036 12257
rect 20628 12291 20680 12300
rect 20628 12257 20637 12291
rect 20637 12257 20671 12291
rect 20671 12257 20680 12291
rect 20628 12248 20680 12257
rect 21456 12248 21508 12300
rect 22100 12248 22152 12300
rect 20996 12180 21048 12232
rect 22652 12291 22704 12300
rect 22652 12257 22661 12291
rect 22661 12257 22695 12291
rect 22695 12257 22704 12291
rect 22652 12248 22704 12257
rect 23572 12316 23624 12368
rect 26056 12384 26108 12436
rect 31760 12384 31812 12436
rect 24492 12248 24544 12300
rect 24952 12248 25004 12300
rect 25320 12248 25372 12300
rect 27436 12248 27488 12300
rect 29184 12316 29236 12368
rect 31024 12316 31076 12368
rect 34704 12384 34756 12436
rect 33876 12359 33928 12368
rect 33876 12325 33885 12359
rect 33885 12325 33919 12359
rect 33919 12325 33928 12359
rect 37648 12384 37700 12436
rect 33876 12316 33928 12325
rect 29368 12248 29420 12300
rect 34060 12248 34112 12300
rect 34796 12248 34848 12300
rect 35808 12248 35860 12300
rect 23572 12180 23624 12232
rect 24308 12180 24360 12232
rect 24584 12223 24636 12232
rect 24584 12189 24593 12223
rect 24593 12189 24627 12223
rect 24627 12189 24636 12223
rect 24584 12180 24636 12189
rect 26792 12180 26844 12232
rect 21732 12112 21784 12164
rect 15292 12044 15344 12096
rect 16396 12044 16448 12096
rect 16488 12044 16540 12096
rect 17316 12044 17368 12096
rect 20536 12044 20588 12096
rect 21272 12044 21324 12096
rect 21640 12044 21692 12096
rect 22468 12087 22520 12096
rect 22468 12053 22477 12087
rect 22477 12053 22511 12087
rect 22511 12053 22520 12087
rect 22468 12044 22520 12053
rect 22560 12087 22612 12096
rect 22560 12053 22569 12087
rect 22569 12053 22603 12087
rect 22603 12053 22612 12087
rect 22560 12044 22612 12053
rect 26700 12112 26752 12164
rect 27160 12112 27212 12164
rect 27528 12112 27580 12164
rect 28908 12180 28960 12232
rect 31392 12180 31444 12232
rect 34888 12223 34940 12232
rect 34888 12189 34897 12223
rect 34897 12189 34931 12223
rect 34931 12189 34940 12223
rect 34888 12180 34940 12189
rect 28724 12112 28776 12164
rect 29644 12112 29696 12164
rect 26332 12087 26384 12096
rect 26332 12053 26341 12087
rect 26341 12053 26375 12087
rect 26375 12053 26384 12087
rect 26332 12044 26384 12053
rect 27344 12087 27396 12096
rect 27344 12053 27353 12087
rect 27353 12053 27387 12087
rect 27387 12053 27396 12087
rect 27344 12044 27396 12053
rect 30932 12044 30984 12096
rect 32404 12155 32456 12164
rect 32404 12121 32413 12155
rect 32413 12121 32447 12155
rect 32447 12121 32456 12155
rect 32404 12112 32456 12121
rect 31392 12044 31444 12096
rect 31760 12044 31812 12096
rect 33324 12044 33376 12096
rect 35072 12112 35124 12164
rect 34336 12044 34388 12096
rect 36728 12112 36780 12164
rect 37464 12248 37516 12300
rect 37648 12291 37700 12300
rect 37648 12257 37657 12291
rect 37657 12257 37691 12291
rect 37691 12257 37700 12291
rect 37648 12248 37700 12257
rect 37740 12248 37792 12300
rect 37280 12180 37332 12232
rect 49148 12291 49200 12300
rect 49148 12257 49157 12291
rect 49157 12257 49191 12291
rect 49191 12257 49200 12291
rect 49148 12248 49200 12257
rect 39304 12112 39356 12164
rect 43352 12112 43404 12164
rect 36544 12044 36596 12096
rect 36820 12044 36872 12096
rect 37464 12087 37516 12096
rect 37464 12053 37473 12087
rect 37473 12053 37507 12087
rect 37507 12053 37516 12087
rect 37464 12044 37516 12053
rect 38660 12087 38712 12096
rect 38660 12053 38669 12087
rect 38669 12053 38703 12087
rect 38703 12053 38712 12087
rect 38660 12044 38712 12053
rect 40776 12087 40828 12096
rect 40776 12053 40785 12087
rect 40785 12053 40819 12087
rect 40819 12053 40828 12087
rect 40776 12044 40828 12053
rect 47952 12223 48004 12232
rect 47952 12189 47961 12223
rect 47961 12189 47995 12223
rect 47995 12189 48004 12223
rect 47952 12180 48004 12189
rect 45928 12087 45980 12096
rect 45928 12053 45937 12087
rect 45937 12053 45971 12087
rect 45971 12053 45980 12087
rect 45928 12044 45980 12053
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 27950 11942 28002 11994
rect 28014 11942 28066 11994
rect 28078 11942 28130 11994
rect 28142 11942 28194 11994
rect 28206 11942 28258 11994
rect 37950 11942 38002 11994
rect 38014 11942 38066 11994
rect 38078 11942 38130 11994
rect 38142 11942 38194 11994
rect 38206 11942 38258 11994
rect 47950 11942 48002 11994
rect 48014 11942 48066 11994
rect 48078 11942 48130 11994
rect 48142 11942 48194 11994
rect 48206 11942 48258 11994
rect 4160 11840 4212 11892
rect 11704 11840 11756 11892
rect 12164 11840 12216 11892
rect 13268 11840 13320 11892
rect 13636 11840 13688 11892
rect 15568 11883 15620 11892
rect 14188 11772 14240 11824
rect 15200 11772 15252 11824
rect 1216 11704 1268 11756
rect 1308 11636 1360 11688
rect 11888 11704 11940 11756
rect 15568 11849 15577 11883
rect 15577 11849 15611 11883
rect 15611 11849 15620 11883
rect 15568 11840 15620 11849
rect 16396 11883 16448 11892
rect 16396 11849 16405 11883
rect 16405 11849 16439 11883
rect 16439 11849 16448 11883
rect 16396 11840 16448 11849
rect 18788 11840 18840 11892
rect 19248 11840 19300 11892
rect 19340 11772 19392 11824
rect 19892 11815 19944 11824
rect 19892 11781 19901 11815
rect 19901 11781 19935 11815
rect 19935 11781 19944 11815
rect 19892 11772 19944 11781
rect 11244 11636 11296 11688
rect 12256 11636 12308 11688
rect 15936 11704 15988 11756
rect 20076 11772 20128 11824
rect 11796 11568 11848 11620
rect 14464 11568 14516 11620
rect 14740 11636 14792 11688
rect 16764 11636 16816 11688
rect 12532 11500 12584 11552
rect 14832 11500 14884 11552
rect 16212 11568 16264 11620
rect 15660 11500 15712 11552
rect 18144 11500 18196 11552
rect 18236 11500 18288 11552
rect 22192 11772 22244 11824
rect 21364 11704 21416 11756
rect 21640 11704 21692 11756
rect 22100 11747 22152 11756
rect 22100 11713 22109 11747
rect 22109 11713 22143 11747
rect 22143 11713 22152 11747
rect 22100 11704 22152 11713
rect 24492 11840 24544 11892
rect 27344 11840 27396 11892
rect 27528 11840 27580 11892
rect 31576 11840 31628 11892
rect 31760 11883 31812 11892
rect 31760 11849 31769 11883
rect 31769 11849 31803 11883
rect 31803 11849 31812 11883
rect 31760 11840 31812 11849
rect 32128 11840 32180 11892
rect 33692 11840 33744 11892
rect 34796 11840 34848 11892
rect 35348 11840 35400 11892
rect 36084 11840 36136 11892
rect 37740 11840 37792 11892
rect 37832 11840 37884 11892
rect 38660 11883 38712 11892
rect 38660 11849 38669 11883
rect 38669 11849 38703 11883
rect 38703 11849 38712 11883
rect 38660 11840 38712 11849
rect 22652 11772 22704 11824
rect 24308 11772 24360 11824
rect 25964 11772 26016 11824
rect 22560 11747 22612 11756
rect 22560 11713 22569 11747
rect 22569 11713 22603 11747
rect 22603 11713 22612 11747
rect 22560 11704 22612 11713
rect 26148 11747 26200 11756
rect 26148 11713 26157 11747
rect 26157 11713 26191 11747
rect 26191 11713 26200 11747
rect 26148 11704 26200 11713
rect 27344 11704 27396 11756
rect 20628 11636 20680 11688
rect 20076 11568 20128 11620
rect 20812 11568 20864 11620
rect 21456 11636 21508 11688
rect 22008 11636 22060 11688
rect 23480 11636 23532 11688
rect 23848 11636 23900 11688
rect 24308 11636 24360 11688
rect 26332 11636 26384 11688
rect 28816 11772 28868 11824
rect 30012 11772 30064 11824
rect 30932 11772 30984 11824
rect 21548 11568 21600 11620
rect 21732 11568 21784 11620
rect 21180 11500 21232 11552
rect 21640 11500 21692 11552
rect 23572 11568 23624 11620
rect 31392 11772 31444 11824
rect 31116 11747 31168 11756
rect 31116 11713 31125 11747
rect 31125 11713 31159 11747
rect 31159 11713 31168 11747
rect 31116 11704 31168 11713
rect 27252 11568 27304 11620
rect 31208 11679 31260 11688
rect 31208 11645 31217 11679
rect 31217 11645 31251 11679
rect 31251 11645 31260 11679
rect 31208 11636 31260 11645
rect 31300 11679 31352 11688
rect 31300 11645 31309 11679
rect 31309 11645 31343 11679
rect 31343 11645 31352 11679
rect 31300 11636 31352 11645
rect 31484 11636 31536 11688
rect 32864 11679 32916 11688
rect 32864 11645 32873 11679
rect 32873 11645 32907 11679
rect 32907 11645 32916 11679
rect 32864 11636 32916 11645
rect 36728 11772 36780 11824
rect 37372 11772 37424 11824
rect 40776 11772 40828 11824
rect 49148 11815 49200 11824
rect 49148 11781 49157 11815
rect 49157 11781 49191 11815
rect 49191 11781 49200 11815
rect 49148 11772 49200 11781
rect 36912 11704 36964 11756
rect 39028 11747 39080 11756
rect 39028 11713 39037 11747
rect 39037 11713 39071 11747
rect 39071 11713 39080 11747
rect 39028 11704 39080 11713
rect 39948 11747 40000 11756
rect 39948 11713 39957 11747
rect 39957 11713 39991 11747
rect 39991 11713 40000 11747
rect 39948 11704 40000 11713
rect 45928 11704 45980 11756
rect 30564 11568 30616 11620
rect 35072 11636 35124 11688
rect 36636 11636 36688 11688
rect 36820 11568 36872 11620
rect 43720 11568 43772 11620
rect 46296 11568 46348 11620
rect 29460 11500 29512 11552
rect 30104 11500 30156 11552
rect 33416 11500 33468 11552
rect 37372 11500 37424 11552
rect 40224 11500 40276 11552
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 32950 11398 33002 11450
rect 33014 11398 33066 11450
rect 33078 11398 33130 11450
rect 33142 11398 33194 11450
rect 33206 11398 33258 11450
rect 42950 11398 43002 11450
rect 43014 11398 43066 11450
rect 43078 11398 43130 11450
rect 43142 11398 43194 11450
rect 43206 11398 43258 11450
rect 1216 11296 1268 11348
rect 12440 11296 12492 11348
rect 13452 11296 13504 11348
rect 16672 11296 16724 11348
rect 19248 11339 19300 11348
rect 19248 11305 19257 11339
rect 19257 11305 19291 11339
rect 19291 11305 19300 11339
rect 19248 11296 19300 11305
rect 19892 11296 19944 11348
rect 21732 11296 21784 11348
rect 22008 11296 22060 11348
rect 22468 11296 22520 11348
rect 22560 11296 22612 11348
rect 24400 11296 24452 11348
rect 28908 11339 28960 11348
rect 28908 11305 28917 11339
rect 28917 11305 28951 11339
rect 28951 11305 28960 11339
rect 28908 11296 28960 11305
rect 1768 11271 1820 11280
rect 1768 11237 1777 11271
rect 1777 11237 1811 11271
rect 1811 11237 1820 11271
rect 1768 11228 1820 11237
rect 12716 11271 12768 11280
rect 12716 11237 12725 11271
rect 12725 11237 12759 11271
rect 12759 11237 12768 11271
rect 12716 11228 12768 11237
rect 14648 11228 14700 11280
rect 13820 11160 13872 11212
rect 14832 11203 14884 11212
rect 14832 11169 14841 11203
rect 14841 11169 14875 11203
rect 14875 11169 14884 11203
rect 14832 11160 14884 11169
rect 18788 11228 18840 11280
rect 23388 11228 23440 11280
rect 26608 11228 26660 11280
rect 28448 11228 28500 11280
rect 15476 11160 15528 11212
rect 17040 11160 17092 11212
rect 1584 11135 1636 11144
rect 1584 11101 1593 11135
rect 1593 11101 1627 11135
rect 1627 11101 1636 11135
rect 1584 11092 1636 11101
rect 12348 11092 12400 11144
rect 12900 11092 12952 11144
rect 14740 11135 14792 11144
rect 14740 11101 14749 11135
rect 14749 11101 14783 11135
rect 14783 11101 14792 11135
rect 14740 11092 14792 11101
rect 18328 11092 18380 11144
rect 18420 11135 18472 11144
rect 18420 11101 18429 11135
rect 18429 11101 18463 11135
rect 18463 11101 18472 11135
rect 18420 11092 18472 11101
rect 18604 11203 18656 11212
rect 18604 11169 18613 11203
rect 18613 11169 18647 11203
rect 18647 11169 18656 11203
rect 18604 11160 18656 11169
rect 18880 11160 18932 11212
rect 21456 11160 21508 11212
rect 21732 11160 21784 11212
rect 23848 11160 23900 11212
rect 24124 11160 24176 11212
rect 24492 11160 24544 11212
rect 29184 11160 29236 11212
rect 19524 11092 19576 11144
rect 23480 11092 23532 11144
rect 24584 11135 24636 11144
rect 24584 11101 24593 11135
rect 24593 11101 24627 11135
rect 24627 11101 24636 11135
rect 24584 11092 24636 11101
rect 25964 11092 26016 11144
rect 11244 11067 11296 11076
rect 11244 11033 11253 11067
rect 11253 11033 11287 11067
rect 11287 11033 11296 11067
rect 11244 11024 11296 11033
rect 1768 10956 1820 11008
rect 15844 11024 15896 11076
rect 16580 11024 16632 11076
rect 17776 11024 17828 11076
rect 18144 11024 18196 11076
rect 14004 10956 14056 11008
rect 15384 10956 15436 11008
rect 16396 10956 16448 11008
rect 17868 10956 17920 11008
rect 19064 11024 19116 11076
rect 20812 11024 20864 11076
rect 21180 11024 21232 11076
rect 18604 10956 18656 11008
rect 19892 10956 19944 11008
rect 22652 10999 22704 11008
rect 22652 10965 22661 10999
rect 22661 10965 22695 10999
rect 22695 10965 22704 10999
rect 22652 10956 22704 10965
rect 24216 11024 24268 11076
rect 28816 11024 28868 11076
rect 30012 11228 30064 11280
rect 33416 11296 33468 11348
rect 34980 11296 35032 11348
rect 36176 11296 36228 11348
rect 39304 11296 39356 11348
rect 39488 11296 39540 11348
rect 31024 11160 31076 11212
rect 31944 11160 31996 11212
rect 32128 11160 32180 11212
rect 32772 11160 32824 11212
rect 34060 11203 34112 11212
rect 34060 11169 34069 11203
rect 34069 11169 34103 11203
rect 34103 11169 34112 11203
rect 34060 11160 34112 11169
rect 34152 11160 34204 11212
rect 35716 11203 35768 11212
rect 35716 11169 35725 11203
rect 35725 11169 35759 11203
rect 35759 11169 35768 11203
rect 35716 11160 35768 11169
rect 41604 11296 41656 11348
rect 29552 11092 29604 11144
rect 33784 11092 33836 11144
rect 29368 11024 29420 11076
rect 30196 11067 30248 11076
rect 30196 11033 30205 11067
rect 30205 11033 30239 11067
rect 30239 11033 30248 11067
rect 30196 11024 30248 11033
rect 30748 11067 30800 11076
rect 26148 10956 26200 11008
rect 26976 10956 27028 11008
rect 27804 10956 27856 11008
rect 29736 10956 29788 11008
rect 30012 10956 30064 11008
rect 30748 11033 30757 11067
rect 30757 11033 30791 11067
rect 30791 11033 30800 11067
rect 30748 11024 30800 11033
rect 33232 11024 33284 11076
rect 36084 11024 36136 11076
rect 36728 11024 36780 11076
rect 37372 11024 37424 11076
rect 39488 11092 39540 11144
rect 40224 11092 40276 11144
rect 49148 11203 49200 11212
rect 49148 11169 49157 11203
rect 49157 11169 49191 11203
rect 49191 11169 49200 11203
rect 49148 11160 49200 11169
rect 47032 11092 47084 11144
rect 45744 11024 45796 11076
rect 46940 11024 46992 11076
rect 30380 10956 30432 11008
rect 32312 10956 32364 11008
rect 32956 10956 33008 11008
rect 37464 10956 37516 11008
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 27950 10854 28002 10906
rect 28014 10854 28066 10906
rect 28078 10854 28130 10906
rect 28142 10854 28194 10906
rect 28206 10854 28258 10906
rect 37950 10854 38002 10906
rect 38014 10854 38066 10906
rect 38078 10854 38130 10906
rect 38142 10854 38194 10906
rect 38206 10854 38258 10906
rect 47950 10854 48002 10906
rect 48014 10854 48066 10906
rect 48078 10854 48130 10906
rect 48142 10854 48194 10906
rect 48206 10854 48258 10906
rect 1768 10795 1820 10804
rect 1768 10761 1777 10795
rect 1777 10761 1811 10795
rect 1811 10761 1820 10795
rect 1768 10752 1820 10761
rect 1860 10752 1912 10804
rect 1216 10684 1268 10736
rect 12348 10752 12400 10804
rect 12808 10752 12860 10804
rect 14188 10752 14240 10804
rect 18052 10752 18104 10804
rect 1308 10616 1360 10668
rect 14556 10684 14608 10736
rect 13544 10659 13596 10668
rect 13544 10625 13553 10659
rect 13553 10625 13587 10659
rect 13587 10625 13596 10659
rect 13544 10616 13596 10625
rect 13636 10659 13688 10668
rect 13636 10625 13645 10659
rect 13645 10625 13679 10659
rect 13679 10625 13688 10659
rect 13636 10616 13688 10625
rect 13912 10616 13964 10668
rect 15752 10684 15804 10736
rect 15844 10684 15896 10736
rect 17592 10684 17644 10736
rect 16488 10616 16540 10668
rect 18236 10616 18288 10668
rect 14372 10548 14424 10600
rect 14924 10591 14976 10600
rect 14924 10557 14933 10591
rect 14933 10557 14967 10591
rect 14967 10557 14976 10591
rect 14924 10548 14976 10557
rect 16028 10591 16080 10600
rect 16028 10557 16037 10591
rect 16037 10557 16071 10591
rect 16071 10557 16080 10591
rect 16028 10548 16080 10557
rect 16120 10591 16172 10600
rect 16120 10557 16129 10591
rect 16129 10557 16163 10591
rect 16163 10557 16172 10591
rect 16120 10548 16172 10557
rect 16580 10548 16632 10600
rect 18696 10659 18748 10668
rect 18696 10625 18705 10659
rect 18705 10625 18739 10659
rect 18739 10625 18748 10659
rect 18696 10616 18748 10625
rect 19708 10752 19760 10804
rect 19892 10795 19944 10804
rect 19892 10761 19901 10795
rect 19901 10761 19935 10795
rect 19935 10761 19944 10795
rect 19892 10752 19944 10761
rect 22652 10752 22704 10804
rect 23664 10752 23716 10804
rect 26148 10752 26200 10804
rect 22284 10684 22336 10736
rect 28908 10752 28960 10804
rect 29736 10752 29788 10804
rect 15016 10480 15068 10532
rect 14280 10412 14332 10464
rect 15568 10455 15620 10464
rect 15568 10421 15577 10455
rect 15577 10421 15611 10455
rect 15611 10421 15620 10455
rect 15568 10412 15620 10421
rect 16396 10412 16448 10464
rect 18420 10412 18472 10464
rect 21456 10616 21508 10668
rect 23388 10616 23440 10668
rect 20812 10548 20864 10600
rect 21548 10548 21600 10600
rect 22008 10591 22060 10600
rect 22008 10557 22017 10591
rect 22017 10557 22051 10591
rect 22051 10557 22060 10591
rect 22008 10548 22060 10557
rect 21824 10480 21876 10532
rect 22836 10548 22888 10600
rect 27436 10616 27488 10668
rect 23940 10548 23992 10600
rect 24860 10591 24912 10600
rect 24860 10557 24869 10591
rect 24869 10557 24903 10591
rect 24903 10557 24912 10591
rect 24860 10548 24912 10557
rect 26608 10548 26660 10600
rect 27804 10591 27856 10600
rect 27804 10557 27813 10591
rect 27813 10557 27847 10591
rect 27847 10557 27856 10591
rect 27804 10548 27856 10557
rect 29552 10727 29604 10736
rect 29552 10693 29561 10727
rect 29561 10693 29595 10727
rect 29595 10693 29604 10727
rect 29552 10684 29604 10693
rect 30288 10684 30340 10736
rect 31116 10752 31168 10804
rect 32956 10752 33008 10804
rect 33324 10795 33376 10804
rect 33324 10761 33333 10795
rect 33333 10761 33367 10795
rect 33367 10761 33376 10795
rect 33324 10752 33376 10761
rect 29736 10616 29788 10668
rect 29092 10548 29144 10600
rect 30380 10548 30432 10600
rect 30472 10548 30524 10600
rect 31760 10684 31812 10736
rect 32220 10684 32272 10736
rect 32404 10684 32456 10736
rect 32680 10659 32732 10668
rect 32680 10625 32689 10659
rect 32689 10625 32723 10659
rect 32723 10625 32732 10659
rect 32680 10616 32732 10625
rect 35072 10752 35124 10804
rect 35716 10752 35768 10804
rect 36912 10752 36964 10804
rect 35348 10684 35400 10736
rect 35532 10616 35584 10668
rect 35716 10616 35768 10668
rect 22100 10412 22152 10464
rect 23664 10412 23716 10464
rect 25964 10455 26016 10464
rect 25964 10421 25973 10455
rect 25973 10421 26007 10455
rect 26007 10421 26016 10455
rect 25964 10412 26016 10421
rect 26148 10455 26200 10464
rect 26148 10421 26157 10455
rect 26157 10421 26191 10455
rect 26191 10421 26200 10455
rect 26148 10412 26200 10421
rect 26516 10455 26568 10464
rect 26516 10421 26525 10455
rect 26525 10421 26559 10455
rect 26559 10421 26568 10455
rect 26516 10412 26568 10421
rect 26792 10455 26844 10464
rect 26792 10421 26801 10455
rect 26801 10421 26835 10455
rect 26835 10421 26844 10455
rect 26792 10412 26844 10421
rect 32312 10480 32364 10532
rect 30012 10412 30064 10464
rect 31300 10412 31352 10464
rect 31944 10455 31996 10464
rect 31944 10421 31953 10455
rect 31953 10421 31987 10455
rect 31987 10421 31996 10455
rect 31944 10412 31996 10421
rect 32220 10412 32272 10464
rect 32864 10412 32916 10464
rect 35164 10480 35216 10532
rect 35900 10548 35952 10600
rect 36728 10684 36780 10736
rect 49240 10684 49292 10736
rect 39764 10659 39816 10668
rect 39764 10625 39773 10659
rect 39773 10625 39807 10659
rect 39807 10625 39816 10659
rect 39764 10616 39816 10625
rect 46940 10616 46992 10668
rect 46940 10480 46992 10532
rect 35348 10412 35400 10464
rect 36636 10412 36688 10464
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 32950 10310 33002 10362
rect 33014 10310 33066 10362
rect 33078 10310 33130 10362
rect 33142 10310 33194 10362
rect 33206 10310 33258 10362
rect 42950 10310 43002 10362
rect 43014 10310 43066 10362
rect 43078 10310 43130 10362
rect 43142 10310 43194 10362
rect 43206 10310 43258 10362
rect 16028 10208 16080 10260
rect 16212 10208 16264 10260
rect 18052 10208 18104 10260
rect 18328 10208 18380 10260
rect 13912 10183 13964 10192
rect 13912 10149 13921 10183
rect 13921 10149 13955 10183
rect 13955 10149 13964 10183
rect 13912 10140 13964 10149
rect 1860 10115 1912 10124
rect 1860 10081 1869 10115
rect 1869 10081 1903 10115
rect 1903 10081 1912 10115
rect 1860 10072 1912 10081
rect 1308 10004 1360 10056
rect 17960 10140 18012 10192
rect 16856 10072 16908 10124
rect 17408 10115 17460 10124
rect 17408 10081 17417 10115
rect 17417 10081 17451 10115
rect 17451 10081 17460 10115
rect 17408 10072 17460 10081
rect 17500 10115 17552 10124
rect 17500 10081 17509 10115
rect 17509 10081 17543 10115
rect 17543 10081 17552 10115
rect 17500 10072 17552 10081
rect 18236 10072 18288 10124
rect 13820 10004 13872 10056
rect 16672 10004 16724 10056
rect 21640 10208 21692 10260
rect 22836 10208 22888 10260
rect 23756 10208 23808 10260
rect 32128 10251 32180 10260
rect 32128 10217 32137 10251
rect 32137 10217 32171 10251
rect 32171 10217 32180 10251
rect 32128 10208 32180 10217
rect 34428 10208 34480 10260
rect 18512 10072 18564 10124
rect 19616 10072 19668 10124
rect 19708 10072 19760 10124
rect 21548 10072 21600 10124
rect 19800 10004 19852 10056
rect 23388 10140 23440 10192
rect 23848 10183 23900 10192
rect 23848 10149 23857 10183
rect 23857 10149 23891 10183
rect 23891 10149 23900 10183
rect 23848 10140 23900 10149
rect 26516 10140 26568 10192
rect 22008 10072 22060 10124
rect 24124 10072 24176 10124
rect 29092 10140 29144 10192
rect 30288 10140 30340 10192
rect 33048 10140 33100 10192
rect 35164 10208 35216 10260
rect 35348 10208 35400 10260
rect 14832 9936 14884 9988
rect 15292 9936 15344 9988
rect 15844 9936 15896 9988
rect 16212 9936 16264 9988
rect 12440 9911 12492 9920
rect 12440 9877 12449 9911
rect 12449 9877 12483 9911
rect 12483 9877 12492 9911
rect 13084 9911 13136 9920
rect 12440 9868 12492 9877
rect 13084 9877 13093 9911
rect 13093 9877 13127 9911
rect 13127 9877 13136 9911
rect 13084 9868 13136 9877
rect 13912 9868 13964 9920
rect 14464 9868 14516 9920
rect 16120 9868 16172 9920
rect 16948 9911 17000 9920
rect 16948 9877 16957 9911
rect 16957 9877 16991 9911
rect 16991 9877 17000 9911
rect 16948 9868 17000 9877
rect 17316 9911 17368 9920
rect 17316 9877 17325 9911
rect 17325 9877 17359 9911
rect 17359 9877 17368 9911
rect 17316 9868 17368 9877
rect 20812 9936 20864 9988
rect 21180 9936 21232 9988
rect 22560 10004 22612 10056
rect 25964 10004 26016 10056
rect 26516 10004 26568 10056
rect 26976 10047 27028 10056
rect 26976 10013 26985 10047
rect 26985 10013 27019 10047
rect 27019 10013 27028 10047
rect 26976 10004 27028 10013
rect 28816 10072 28868 10124
rect 29368 10115 29420 10124
rect 29368 10081 29377 10115
rect 29377 10081 29411 10115
rect 29411 10081 29420 10115
rect 29368 10072 29420 10081
rect 32680 10072 32732 10124
rect 33232 10115 33284 10124
rect 33232 10081 33241 10115
rect 33241 10081 33275 10115
rect 33275 10081 33284 10115
rect 33232 10072 33284 10081
rect 34060 10072 34112 10124
rect 35256 10072 35308 10124
rect 30380 10047 30432 10056
rect 30380 10013 30389 10047
rect 30389 10013 30423 10047
rect 30423 10013 30432 10047
rect 30380 10004 30432 10013
rect 31760 10004 31812 10056
rect 36636 10251 36688 10260
rect 36636 10217 36645 10251
rect 36645 10217 36679 10251
rect 36679 10217 36688 10251
rect 36636 10208 36688 10217
rect 36728 10208 36780 10260
rect 49148 10115 49200 10124
rect 49148 10081 49157 10115
rect 49157 10081 49191 10115
rect 49191 10081 49200 10115
rect 49148 10072 49200 10081
rect 21548 9868 21600 9920
rect 21824 9868 21876 9920
rect 23940 9868 23992 9920
rect 24860 9979 24912 9988
rect 24860 9945 24869 9979
rect 24869 9945 24903 9979
rect 24903 9945 24912 9979
rect 24860 9936 24912 9945
rect 26332 9936 26384 9988
rect 26148 9868 26200 9920
rect 30104 9936 30156 9988
rect 30656 9979 30708 9988
rect 30656 9945 30665 9979
rect 30665 9945 30699 9979
rect 30699 9945 30708 9979
rect 30656 9936 30708 9945
rect 29000 9868 29052 9920
rect 33140 9936 33192 9988
rect 32680 9868 32732 9920
rect 35808 9868 35860 9920
rect 36728 9936 36780 9988
rect 38568 9936 38620 9988
rect 41604 10004 41656 10056
rect 45744 10004 45796 10056
rect 46296 10004 46348 10056
rect 38384 9911 38436 9920
rect 38384 9877 38393 9911
rect 38393 9877 38427 9911
rect 38427 9877 38436 9911
rect 38384 9868 38436 9877
rect 46020 9936 46072 9988
rect 47308 9979 47360 9988
rect 47308 9945 47317 9979
rect 47317 9945 47351 9979
rect 47351 9945 47360 9979
rect 47308 9936 47360 9945
rect 45836 9868 45888 9920
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 27950 9766 28002 9818
rect 28014 9766 28066 9818
rect 28078 9766 28130 9818
rect 28142 9766 28194 9818
rect 28206 9766 28258 9818
rect 37950 9766 38002 9818
rect 38014 9766 38066 9818
rect 38078 9766 38130 9818
rect 38142 9766 38194 9818
rect 38206 9766 38258 9818
rect 47950 9766 48002 9818
rect 48014 9766 48066 9818
rect 48078 9766 48130 9818
rect 48142 9766 48194 9818
rect 48206 9766 48258 9818
rect 1308 9664 1360 9716
rect 16580 9664 16632 9716
rect 17316 9664 17368 9716
rect 20904 9664 20956 9716
rect 21180 9664 21232 9716
rect 21732 9664 21784 9716
rect 22284 9707 22336 9716
rect 22284 9673 22293 9707
rect 22293 9673 22327 9707
rect 22327 9673 22336 9707
rect 22284 9664 22336 9673
rect 31484 9707 31536 9716
rect 12532 9639 12584 9648
rect 12532 9605 12541 9639
rect 12541 9605 12575 9639
rect 12575 9605 12584 9639
rect 12532 9596 12584 9605
rect 12624 9639 12676 9648
rect 12624 9605 12633 9639
rect 12633 9605 12667 9639
rect 12667 9605 12676 9639
rect 12624 9596 12676 9605
rect 12716 9596 12768 9648
rect 15292 9596 15344 9648
rect 17224 9596 17276 9648
rect 17408 9596 17460 9648
rect 18880 9639 18932 9648
rect 18880 9605 18889 9639
rect 18889 9605 18923 9639
rect 18923 9605 18932 9639
rect 18880 9596 18932 9605
rect 19524 9596 19576 9648
rect 21456 9596 21508 9648
rect 23756 9639 23808 9648
rect 23756 9605 23765 9639
rect 23765 9605 23799 9639
rect 23799 9605 23808 9639
rect 23756 9596 23808 9605
rect 25596 9596 25648 9648
rect 1308 9528 1360 9580
rect 16212 9528 16264 9580
rect 16488 9571 16540 9580
rect 16488 9537 16497 9571
rect 16497 9537 16531 9571
rect 16531 9537 16540 9571
rect 16488 9528 16540 9537
rect 21088 9528 21140 9580
rect 22652 9571 22704 9580
rect 22652 9537 22661 9571
rect 22661 9537 22695 9571
rect 22695 9537 22704 9571
rect 22652 9528 22704 9537
rect 23480 9571 23532 9580
rect 23480 9537 23489 9571
rect 23489 9537 23523 9571
rect 23523 9537 23532 9571
rect 23480 9528 23532 9537
rect 1768 9435 1820 9444
rect 1768 9401 1777 9435
rect 1777 9401 1811 9435
rect 1811 9401 1820 9435
rect 1768 9392 1820 9401
rect 12808 9324 12860 9376
rect 13636 9503 13688 9512
rect 13636 9469 13645 9503
rect 13645 9469 13679 9503
rect 13679 9469 13688 9503
rect 13636 9460 13688 9469
rect 14188 9460 14240 9512
rect 16672 9460 16724 9512
rect 16764 9460 16816 9512
rect 14924 9392 14976 9444
rect 16580 9392 16632 9444
rect 13820 9324 13872 9376
rect 15292 9324 15344 9376
rect 18604 9460 18656 9512
rect 22560 9392 22612 9444
rect 21088 9324 21140 9376
rect 21732 9324 21784 9376
rect 23388 9324 23440 9376
rect 23848 9460 23900 9512
rect 25320 9528 25372 9580
rect 25964 9596 26016 9648
rect 28816 9596 28868 9648
rect 31484 9673 31493 9707
rect 31493 9673 31527 9707
rect 31527 9673 31536 9707
rect 31484 9664 31536 9673
rect 31760 9664 31812 9716
rect 32680 9664 32732 9716
rect 33324 9664 33376 9716
rect 35808 9664 35860 9716
rect 30564 9596 30616 9648
rect 31300 9596 31352 9648
rect 25780 9528 25832 9580
rect 26148 9571 26200 9580
rect 26148 9537 26157 9571
rect 26157 9537 26191 9571
rect 26191 9537 26200 9571
rect 26148 9528 26200 9537
rect 34060 9596 34112 9648
rect 34152 9639 34204 9648
rect 34152 9605 34161 9639
rect 34161 9605 34195 9639
rect 34195 9605 34204 9639
rect 34152 9596 34204 9605
rect 35532 9596 35584 9648
rect 38384 9664 38436 9716
rect 47032 9664 47084 9716
rect 49332 9596 49384 9648
rect 26332 9503 26384 9512
rect 26332 9469 26341 9503
rect 26341 9469 26375 9503
rect 26375 9469 26384 9503
rect 26332 9460 26384 9469
rect 26976 9460 27028 9512
rect 28816 9460 28868 9512
rect 29552 9460 29604 9512
rect 29184 9392 29236 9444
rect 29644 9392 29696 9444
rect 30656 9460 30708 9512
rect 31300 9460 31352 9512
rect 25688 9367 25740 9376
rect 25688 9333 25697 9367
rect 25697 9333 25731 9367
rect 25731 9333 25740 9367
rect 25688 9324 25740 9333
rect 30380 9324 30432 9376
rect 31668 9392 31720 9444
rect 43352 9528 43404 9580
rect 35256 9392 35308 9444
rect 35532 9324 35584 9376
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 32950 9222 33002 9274
rect 33014 9222 33066 9274
rect 33078 9222 33130 9274
rect 33142 9222 33194 9274
rect 33206 9222 33258 9274
rect 42950 9222 43002 9274
rect 43014 9222 43066 9274
rect 43078 9222 43130 9274
rect 43142 9222 43194 9274
rect 43206 9222 43258 9274
rect 14188 9120 14240 9172
rect 17868 9120 17920 9172
rect 19524 9120 19576 9172
rect 24400 9163 24452 9172
rect 24400 9129 24409 9163
rect 24409 9129 24443 9163
rect 24443 9129 24452 9163
rect 24400 9120 24452 9129
rect 25320 9163 25372 9172
rect 25320 9129 25329 9163
rect 25329 9129 25363 9163
rect 25363 9129 25372 9163
rect 25320 9120 25372 9129
rect 25596 9163 25648 9172
rect 25596 9129 25605 9163
rect 25605 9129 25639 9163
rect 25639 9129 25648 9163
rect 25596 9120 25648 9129
rect 26148 9120 26200 9172
rect 29000 9120 29052 9172
rect 29644 9120 29696 9172
rect 32680 9120 32732 9172
rect 35900 9120 35952 9172
rect 43628 9120 43680 9172
rect 2320 9052 2372 9104
rect 11152 9052 11204 9104
rect 13820 9052 13872 9104
rect 1216 8916 1268 8968
rect 13636 8984 13688 9036
rect 15384 8984 15436 9036
rect 25688 9052 25740 9104
rect 30472 9052 30524 9104
rect 32312 9052 32364 9104
rect 35716 9052 35768 9104
rect 16764 8984 16816 9036
rect 17040 8984 17092 9036
rect 18696 9027 18748 9036
rect 18696 8993 18705 9027
rect 18705 8993 18739 9027
rect 18739 8993 18748 9027
rect 18696 8984 18748 8993
rect 19708 8984 19760 9036
rect 22008 8984 22060 9036
rect 22560 9027 22612 9036
rect 22560 8993 22569 9027
rect 22569 8993 22603 9027
rect 22603 8993 22612 9027
rect 22560 8984 22612 8993
rect 22652 8984 22704 9036
rect 24860 8984 24912 9036
rect 29644 8984 29696 9036
rect 30380 8984 30432 9036
rect 32588 8984 32640 9036
rect 1308 8848 1360 8900
rect 11336 8916 11388 8968
rect 15292 8916 15344 8968
rect 15568 8959 15620 8968
rect 15568 8925 15577 8959
rect 15577 8925 15611 8959
rect 15611 8925 15620 8959
rect 15568 8916 15620 8925
rect 15660 8959 15712 8968
rect 15660 8925 15669 8959
rect 15669 8925 15703 8959
rect 15703 8925 15712 8959
rect 15660 8916 15712 8925
rect 32680 8916 32732 8968
rect 33876 8916 33928 8968
rect 34060 8984 34112 9036
rect 35532 8984 35584 9036
rect 15108 8848 15160 8900
rect 16580 8848 16632 8900
rect 17224 8848 17276 8900
rect 19800 8848 19852 8900
rect 21088 8848 21140 8900
rect 22100 8848 22152 8900
rect 17592 8780 17644 8832
rect 22376 8780 22428 8832
rect 23848 8848 23900 8900
rect 31024 8891 31076 8900
rect 31024 8857 31033 8891
rect 31033 8857 31067 8891
rect 31067 8857 31076 8891
rect 31024 8848 31076 8857
rect 32588 8848 32640 8900
rect 34152 8916 34204 8968
rect 34520 8916 34572 8968
rect 49240 8984 49292 9036
rect 34980 8848 35032 8900
rect 35808 8848 35860 8900
rect 43720 8916 43772 8968
rect 47492 8848 47544 8900
rect 24860 8823 24912 8832
rect 24860 8789 24869 8823
rect 24869 8789 24903 8823
rect 24903 8789 24912 8823
rect 24860 8780 24912 8789
rect 25688 8823 25740 8832
rect 25688 8789 25697 8823
rect 25697 8789 25731 8823
rect 25731 8789 25740 8823
rect 25688 8780 25740 8789
rect 27804 8823 27856 8832
rect 27804 8789 27813 8823
rect 27813 8789 27847 8823
rect 27847 8789 27856 8823
rect 28632 8823 28684 8832
rect 27804 8780 27856 8789
rect 28632 8789 28641 8823
rect 28641 8789 28675 8823
rect 28675 8789 28684 8823
rect 28632 8780 28684 8789
rect 30380 8780 30432 8832
rect 30564 8780 30616 8832
rect 31392 8780 31444 8832
rect 33784 8823 33836 8832
rect 33784 8789 33793 8823
rect 33793 8789 33827 8823
rect 33827 8789 33836 8823
rect 33784 8780 33836 8789
rect 34888 8823 34940 8832
rect 34888 8789 34897 8823
rect 34897 8789 34931 8823
rect 34931 8789 34940 8823
rect 34888 8780 34940 8789
rect 35256 8823 35308 8832
rect 35256 8789 35265 8823
rect 35265 8789 35299 8823
rect 35299 8789 35308 8823
rect 35256 8780 35308 8789
rect 39580 8780 39632 8832
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 27950 8678 28002 8730
rect 28014 8678 28066 8730
rect 28078 8678 28130 8730
rect 28142 8678 28194 8730
rect 28206 8678 28258 8730
rect 37950 8678 38002 8730
rect 38014 8678 38066 8730
rect 38078 8678 38130 8730
rect 38142 8678 38194 8730
rect 38206 8678 38258 8730
rect 47950 8678 48002 8730
rect 48014 8678 48066 8730
rect 48078 8678 48130 8730
rect 48142 8678 48194 8730
rect 48206 8678 48258 8730
rect 15384 8619 15436 8628
rect 15384 8585 15393 8619
rect 15393 8585 15427 8619
rect 15427 8585 15436 8619
rect 15384 8576 15436 8585
rect 16672 8576 16724 8628
rect 17224 8576 17276 8628
rect 13820 8508 13872 8560
rect 13912 8551 13964 8560
rect 13912 8517 13921 8551
rect 13921 8517 13955 8551
rect 13955 8517 13964 8551
rect 13912 8508 13964 8517
rect 15292 8508 15344 8560
rect 15752 8508 15804 8560
rect 17040 8508 17092 8560
rect 17408 8508 17460 8560
rect 18604 8619 18656 8628
rect 18604 8585 18613 8619
rect 18613 8585 18647 8619
rect 18647 8585 18656 8619
rect 18604 8576 18656 8585
rect 19984 8576 20036 8628
rect 22100 8576 22152 8628
rect 23848 8576 23900 8628
rect 30656 8576 30708 8628
rect 31024 8576 31076 8628
rect 34060 8619 34112 8628
rect 34060 8585 34069 8619
rect 34069 8585 34103 8619
rect 34103 8585 34112 8619
rect 34060 8576 34112 8585
rect 35624 8576 35676 8628
rect 40224 8576 40276 8628
rect 47676 8576 47728 8628
rect 29092 8551 29144 8560
rect 29092 8517 29101 8551
rect 29101 8517 29135 8551
rect 29135 8517 29144 8551
rect 29092 8508 29144 8517
rect 1400 8372 1452 8424
rect 16764 8440 16816 8492
rect 19708 8483 19760 8492
rect 19708 8449 19717 8483
rect 19717 8449 19751 8483
rect 19751 8449 19760 8483
rect 19708 8440 19760 8449
rect 21088 8440 21140 8492
rect 22008 8483 22060 8492
rect 22008 8449 22017 8483
rect 22017 8449 22051 8483
rect 22051 8449 22060 8483
rect 22008 8440 22060 8449
rect 30380 8440 30432 8492
rect 30656 8440 30708 8492
rect 30932 8440 30984 8492
rect 17776 8372 17828 8424
rect 15752 8347 15804 8356
rect 15752 8313 15761 8347
rect 15761 8313 15795 8347
rect 15795 8313 15804 8347
rect 15752 8304 15804 8313
rect 16672 8304 16724 8356
rect 16856 8304 16908 8356
rect 6920 8236 6972 8288
rect 15200 8236 15252 8288
rect 28816 8415 28868 8424
rect 28816 8381 28825 8415
rect 28825 8381 28859 8415
rect 28859 8381 28868 8415
rect 28816 8372 28868 8381
rect 31484 8415 31536 8424
rect 31484 8381 31493 8415
rect 31493 8381 31527 8415
rect 31527 8381 31536 8415
rect 31484 8372 31536 8381
rect 32588 8508 32640 8560
rect 32680 8508 32732 8560
rect 34888 8508 34940 8560
rect 31668 8440 31720 8492
rect 34428 8440 34480 8492
rect 39580 8508 39632 8560
rect 49148 8551 49200 8560
rect 49148 8517 49157 8551
rect 49157 8517 49191 8551
rect 49191 8517 49200 8551
rect 49148 8508 49200 8517
rect 32220 8372 32272 8424
rect 32680 8372 32732 8424
rect 33048 8372 33100 8424
rect 38752 8372 38804 8424
rect 45836 8483 45888 8492
rect 45836 8449 45845 8483
rect 45845 8449 45879 8483
rect 45879 8449 45888 8483
rect 45836 8440 45888 8449
rect 46020 8440 46072 8492
rect 22652 8236 22704 8288
rect 32312 8304 32364 8356
rect 33600 8304 33652 8356
rect 36268 8304 36320 8356
rect 46848 8415 46900 8424
rect 46848 8381 46857 8415
rect 46857 8381 46891 8415
rect 46891 8381 46900 8415
rect 46848 8372 46900 8381
rect 40132 8304 40184 8356
rect 47860 8304 47912 8356
rect 27160 8236 27212 8288
rect 33968 8236 34020 8288
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 32950 8134 33002 8186
rect 33014 8134 33066 8186
rect 33078 8134 33130 8186
rect 33142 8134 33194 8186
rect 33206 8134 33258 8186
rect 42950 8134 43002 8186
rect 43014 8134 43066 8186
rect 43078 8134 43130 8186
rect 43142 8134 43194 8186
rect 43206 8134 43258 8186
rect 1400 8032 1452 8084
rect 18880 8032 18932 8084
rect 19800 8032 19852 8084
rect 21916 8032 21968 8084
rect 17040 7964 17092 8016
rect 1308 7828 1360 7880
rect 2412 7828 2464 7880
rect 14004 7896 14056 7948
rect 16948 7896 17000 7948
rect 19248 7964 19300 8016
rect 24860 7964 24912 8016
rect 32772 7964 32824 8016
rect 18604 7896 18656 7948
rect 19708 7896 19760 7948
rect 23664 7896 23716 7948
rect 29736 7939 29788 7948
rect 29736 7905 29745 7939
rect 29745 7905 29779 7939
rect 29779 7905 29788 7939
rect 29736 7896 29788 7905
rect 30564 7939 30616 7948
rect 30564 7905 30573 7939
rect 30573 7905 30607 7939
rect 30607 7905 30616 7939
rect 30564 7896 30616 7905
rect 31484 7896 31536 7948
rect 32220 7896 32272 7948
rect 33416 7964 33468 8016
rect 33968 8032 34020 8084
rect 35256 7964 35308 8016
rect 12808 7828 12860 7880
rect 18420 7828 18472 7880
rect 22376 7871 22428 7880
rect 22376 7837 22385 7871
rect 22385 7837 22419 7871
rect 22419 7837 22428 7871
rect 22376 7828 22428 7837
rect 34796 7896 34848 7948
rect 49240 7896 49292 7948
rect 14188 7760 14240 7812
rect 18512 7760 18564 7812
rect 19984 7760 20036 7812
rect 21088 7760 21140 7812
rect 18788 7692 18840 7744
rect 21456 7735 21508 7744
rect 21456 7701 21465 7735
rect 21465 7701 21499 7735
rect 21499 7701 21508 7735
rect 21456 7692 21508 7701
rect 22284 7692 22336 7744
rect 25688 7692 25740 7744
rect 30656 7735 30708 7744
rect 30656 7701 30665 7735
rect 30665 7701 30699 7735
rect 30699 7701 30708 7735
rect 30656 7692 30708 7701
rect 31392 7735 31444 7744
rect 31392 7701 31401 7735
rect 31401 7701 31435 7735
rect 31435 7701 31444 7735
rect 31392 7692 31444 7701
rect 32864 7760 32916 7812
rect 39028 7828 39080 7880
rect 46940 7828 46992 7880
rect 38752 7803 38804 7812
rect 38752 7769 38761 7803
rect 38761 7769 38795 7803
rect 38795 7769 38804 7803
rect 38752 7760 38804 7769
rect 40040 7760 40092 7812
rect 32772 7735 32824 7744
rect 32772 7701 32781 7735
rect 32781 7701 32815 7735
rect 32815 7701 32824 7735
rect 32772 7692 32824 7701
rect 38660 7692 38712 7744
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 27950 7590 28002 7642
rect 28014 7590 28066 7642
rect 28078 7590 28130 7642
rect 28142 7590 28194 7642
rect 28206 7590 28258 7642
rect 37950 7590 38002 7642
rect 38014 7590 38066 7642
rect 38078 7590 38130 7642
rect 38142 7590 38194 7642
rect 38206 7590 38258 7642
rect 47950 7590 48002 7642
rect 48014 7590 48066 7642
rect 48078 7590 48130 7642
rect 48142 7590 48194 7642
rect 48206 7590 48258 7642
rect 17408 7488 17460 7540
rect 20536 7488 20588 7540
rect 22468 7531 22520 7540
rect 22468 7497 22477 7531
rect 22477 7497 22511 7531
rect 22511 7497 22520 7531
rect 22468 7488 22520 7497
rect 28540 7488 28592 7540
rect 17316 7420 17368 7472
rect 30564 7420 30616 7472
rect 30932 7531 30984 7540
rect 30932 7497 30941 7531
rect 30941 7497 30975 7531
rect 30975 7497 30984 7531
rect 30932 7488 30984 7497
rect 31392 7488 31444 7540
rect 38660 7488 38712 7540
rect 46940 7488 46992 7540
rect 40132 7420 40184 7472
rect 49332 7420 49384 7472
rect 1308 7352 1360 7404
rect 34336 7352 34388 7404
rect 47032 7352 47084 7404
rect 22652 7327 22704 7336
rect 22652 7293 22661 7327
rect 22661 7293 22695 7327
rect 22695 7293 22704 7327
rect 22652 7284 22704 7293
rect 19156 7216 19208 7268
rect 21456 7148 21508 7200
rect 22468 7148 22520 7200
rect 32772 7148 32824 7200
rect 37372 7148 37424 7200
rect 37924 7191 37976 7200
rect 37924 7157 37933 7191
rect 37933 7157 37967 7191
rect 37967 7157 37976 7191
rect 37924 7148 37976 7157
rect 47768 7216 47820 7268
rect 45836 7148 45888 7200
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 32950 7046 33002 7098
rect 33014 7046 33066 7098
rect 33078 7046 33130 7098
rect 33142 7046 33194 7098
rect 33206 7046 33258 7098
rect 42950 7046 43002 7098
rect 43014 7046 43066 7098
rect 43078 7046 43130 7098
rect 43142 7046 43194 7098
rect 43206 7046 43258 7098
rect 37924 6876 37976 6928
rect 47032 6876 47084 6928
rect 33784 6808 33836 6860
rect 40132 6808 40184 6860
rect 49148 6851 49200 6860
rect 49148 6817 49157 6851
rect 49157 6817 49191 6851
rect 49191 6817 49200 6851
rect 49148 6808 49200 6817
rect 1308 6740 1360 6792
rect 16580 6740 16632 6792
rect 19248 6740 19300 6792
rect 40040 6740 40092 6792
rect 47860 6740 47912 6792
rect 1216 6672 1268 6724
rect 27804 6672 27856 6724
rect 48872 6672 48924 6724
rect 2320 6647 2372 6656
rect 2320 6613 2329 6647
rect 2329 6613 2363 6647
rect 2363 6613 2372 6647
rect 2320 6604 2372 6613
rect 19156 6604 19208 6656
rect 21916 6604 21968 6656
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 27950 6502 28002 6554
rect 28014 6502 28066 6554
rect 28078 6502 28130 6554
rect 28142 6502 28194 6554
rect 28206 6502 28258 6554
rect 37950 6502 38002 6554
rect 38014 6502 38066 6554
rect 38078 6502 38130 6554
rect 38142 6502 38194 6554
rect 38206 6502 38258 6554
rect 47950 6502 48002 6554
rect 48014 6502 48066 6554
rect 48078 6502 48130 6554
rect 48142 6502 48194 6554
rect 48206 6502 48258 6554
rect 1216 6400 1268 6452
rect 40224 6332 40276 6384
rect 49240 6332 49292 6384
rect 1308 6264 1360 6316
rect 17868 6264 17920 6316
rect 18328 6196 18380 6248
rect 25688 6196 25740 6248
rect 36452 6196 36504 6248
rect 14096 6128 14148 6180
rect 7840 6060 7892 6112
rect 22560 6128 22612 6180
rect 28356 6128 28408 6180
rect 37280 6128 37332 6180
rect 47492 6264 47544 6316
rect 19616 6060 19668 6112
rect 30748 6060 30800 6112
rect 47124 6128 47176 6180
rect 37648 6103 37700 6112
rect 37648 6069 37657 6103
rect 37657 6069 37691 6103
rect 37691 6069 37700 6103
rect 37648 6060 37700 6069
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 32950 5958 33002 6010
rect 33014 5958 33066 6010
rect 33078 5958 33130 6010
rect 33142 5958 33194 6010
rect 33206 5958 33258 6010
rect 42950 5958 43002 6010
rect 43014 5958 43066 6010
rect 43078 5958 43130 6010
rect 43142 5958 43194 6010
rect 43206 5958 43258 6010
rect 6920 5856 6972 5908
rect 37648 5856 37700 5908
rect 47308 5856 47360 5908
rect 27436 5788 27488 5840
rect 35808 5788 35860 5840
rect 1308 5652 1360 5704
rect 49424 5720 49476 5772
rect 2780 5652 2832 5704
rect 19340 5652 19392 5704
rect 23940 5652 23992 5704
rect 27344 5652 27396 5704
rect 32772 5652 32824 5704
rect 43720 5695 43772 5704
rect 43720 5661 43729 5695
rect 43729 5661 43763 5695
rect 43763 5661 43772 5695
rect 43720 5652 43772 5661
rect 47676 5652 47728 5704
rect 45744 5584 45796 5636
rect 17684 5516 17736 5568
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 27950 5414 28002 5466
rect 28014 5414 28066 5466
rect 28078 5414 28130 5466
rect 28142 5414 28194 5466
rect 28206 5414 28258 5466
rect 37950 5414 38002 5466
rect 38014 5414 38066 5466
rect 38078 5414 38130 5466
rect 38142 5414 38194 5466
rect 38206 5414 38258 5466
rect 47950 5414 48002 5466
rect 48014 5414 48066 5466
rect 48078 5414 48130 5466
rect 48142 5414 48194 5466
rect 48206 5414 48258 5466
rect 31484 5244 31536 5296
rect 49148 5287 49200 5296
rect 49148 5253 49157 5287
rect 49157 5253 49191 5287
rect 49191 5253 49200 5287
rect 49148 5244 49200 5253
rect 18880 5219 18932 5228
rect 18880 5185 18889 5219
rect 18889 5185 18923 5219
rect 18923 5185 18932 5219
rect 18880 5176 18932 5185
rect 37372 5219 37424 5228
rect 37372 5185 37381 5219
rect 37381 5185 37415 5219
rect 37415 5185 37424 5219
rect 37372 5176 37424 5185
rect 45836 5219 45888 5228
rect 45836 5185 45845 5219
rect 45845 5185 45879 5219
rect 45879 5185 45888 5219
rect 45836 5176 45888 5185
rect 47768 5176 47820 5228
rect 1308 5108 1360 5160
rect 11796 5108 11848 5160
rect 19064 5151 19116 5160
rect 19064 5117 19073 5151
rect 19073 5117 19107 5151
rect 19107 5117 19116 5151
rect 19064 5108 19116 5117
rect 48320 5108 48372 5160
rect 40408 5040 40460 5092
rect 1860 4972 1912 5024
rect 12440 4972 12492 5024
rect 20812 4972 20864 5024
rect 37832 5015 37884 5024
rect 37832 4981 37841 5015
rect 37841 4981 37875 5015
rect 37875 4981 37884 5015
rect 37832 4972 37884 4981
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 32950 4870 33002 4922
rect 33014 4870 33066 4922
rect 33078 4870 33130 4922
rect 33142 4870 33194 4922
rect 33206 4870 33258 4922
rect 42950 4870 43002 4922
rect 43014 4870 43066 4922
rect 43078 4870 43130 4922
rect 43142 4870 43194 4922
rect 43206 4870 43258 4922
rect 1308 4768 1360 4820
rect 35808 4768 35860 4820
rect 11704 4700 11756 4752
rect 20996 4700 21048 4752
rect 19156 4632 19208 4684
rect 21916 4675 21968 4684
rect 21916 4641 21925 4675
rect 21925 4641 21959 4675
rect 21959 4641 21968 4675
rect 21916 4632 21968 4641
rect 1308 4564 1360 4616
rect 19524 4564 19576 4616
rect 22928 4632 22980 4684
rect 23204 4632 23256 4684
rect 22100 4607 22152 4616
rect 22100 4573 22109 4607
rect 22109 4573 22143 4607
rect 22143 4573 22152 4607
rect 22100 4564 22152 4573
rect 19064 4496 19116 4548
rect 24032 4564 24084 4616
rect 40132 4768 40184 4820
rect 37832 4700 37884 4752
rect 47216 4700 47268 4752
rect 37004 4632 37056 4684
rect 49424 4632 49476 4684
rect 24584 4496 24636 4548
rect 19340 4428 19392 4480
rect 21456 4428 21508 4480
rect 24400 4428 24452 4480
rect 32772 4496 32824 4548
rect 46940 4564 46992 4616
rect 39764 4496 39816 4548
rect 32864 4428 32916 4480
rect 37372 4471 37424 4480
rect 37372 4437 37381 4471
rect 37381 4437 37415 4471
rect 37415 4437 37424 4471
rect 37372 4428 37424 4437
rect 47676 4496 47728 4548
rect 49792 4428 49844 4480
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 27950 4326 28002 4378
rect 28014 4326 28066 4378
rect 28078 4326 28130 4378
rect 28142 4326 28194 4378
rect 28206 4326 28258 4378
rect 37950 4326 38002 4378
rect 38014 4326 38066 4378
rect 38078 4326 38130 4378
rect 38142 4326 38194 4378
rect 38206 4326 38258 4378
rect 47950 4326 48002 4378
rect 48014 4326 48066 4378
rect 48078 4326 48130 4378
rect 48142 4326 48194 4378
rect 48206 4326 48258 4378
rect 37372 4224 37424 4276
rect 45652 4224 45704 4276
rect 1400 4156 1452 4208
rect 1308 4088 1360 4140
rect 2504 4088 2556 4140
rect 22100 4156 22152 4208
rect 14924 4020 14976 4072
rect 2688 3884 2740 3936
rect 17960 3952 18012 4004
rect 18328 3952 18380 4004
rect 22928 4131 22980 4140
rect 22928 4097 22972 4131
rect 22972 4097 22980 4131
rect 22928 4088 22980 4097
rect 23204 4088 23256 4140
rect 23480 4020 23532 4072
rect 24216 4063 24268 4072
rect 24216 4029 24225 4063
rect 24225 4029 24259 4063
rect 24259 4029 24268 4063
rect 24216 4020 24268 4029
rect 24400 4063 24452 4072
rect 24400 4029 24409 4063
rect 24409 4029 24443 4063
rect 24443 4029 24452 4063
rect 24400 4020 24452 4029
rect 25412 4063 25464 4072
rect 25412 4029 25421 4063
rect 25421 4029 25455 4063
rect 25455 4029 25464 4063
rect 25412 4020 25464 4029
rect 7840 3884 7892 3936
rect 22836 3884 22888 3936
rect 37280 4088 37332 4140
rect 39212 4088 39264 4140
rect 45836 4131 45888 4140
rect 45836 4097 45845 4131
rect 45845 4097 45879 4131
rect 45879 4097 45888 4131
rect 45836 4088 45888 4097
rect 47032 4088 47084 4140
rect 49332 4088 49384 4140
rect 27620 4063 27672 4072
rect 27620 4029 27629 4063
rect 27629 4029 27663 4063
rect 27663 4029 27672 4063
rect 27620 4020 27672 4029
rect 46664 4063 46716 4072
rect 46664 4029 46673 4063
rect 46673 4029 46707 4063
rect 46707 4029 46716 4063
rect 46664 4020 46716 4029
rect 34428 3952 34480 4004
rect 27804 3884 27856 3936
rect 47676 3927 47728 3936
rect 47676 3893 47685 3927
rect 47685 3893 47719 3927
rect 47719 3893 47728 3927
rect 47676 3884 47728 3893
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 32950 3782 33002 3834
rect 33014 3782 33066 3834
rect 33078 3782 33130 3834
rect 33142 3782 33194 3834
rect 33206 3782 33258 3834
rect 42950 3782 43002 3834
rect 43014 3782 43066 3834
rect 43078 3782 43130 3834
rect 43142 3782 43194 3834
rect 43206 3782 43258 3834
rect 25964 3680 26016 3732
rect 26056 3680 26108 3732
rect 27620 3680 27672 3732
rect 22560 3612 22612 3664
rect 24032 3655 24084 3664
rect 24032 3621 24041 3655
rect 24041 3621 24075 3655
rect 24075 3621 24084 3655
rect 24032 3612 24084 3621
rect 24124 3612 24176 3664
rect 1860 3587 1912 3596
rect 1860 3553 1869 3587
rect 1869 3553 1903 3587
rect 1903 3553 1912 3587
rect 1860 3544 1912 3553
rect 7472 3544 7524 3596
rect 1308 3476 1360 3528
rect 3332 3476 3384 3528
rect 11704 3476 11756 3528
rect 17960 3476 18012 3528
rect 20996 3519 21048 3528
rect 20996 3485 21005 3519
rect 21005 3485 21039 3519
rect 21039 3485 21048 3519
rect 20996 3476 21048 3485
rect 21180 3408 21232 3460
rect 22560 3408 22612 3460
rect 22836 3544 22888 3596
rect 40408 3612 40460 3664
rect 45836 3544 45888 3596
rect 23572 3519 23624 3528
rect 23572 3485 23581 3519
rect 23581 3485 23615 3519
rect 23615 3485 23624 3519
rect 23572 3476 23624 3485
rect 24124 3408 24176 3460
rect 12808 3340 12860 3392
rect 23388 3340 23440 3392
rect 36452 3519 36504 3528
rect 36452 3485 36461 3519
rect 36461 3485 36495 3519
rect 36495 3485 36504 3519
rect 36452 3476 36504 3485
rect 45560 3476 45612 3528
rect 49148 3587 49200 3596
rect 49148 3553 49157 3587
rect 49157 3553 49191 3587
rect 49191 3553 49200 3587
rect 49148 3544 49200 3553
rect 47124 3476 47176 3528
rect 48688 3408 48740 3460
rect 27528 3340 27580 3392
rect 35440 3340 35492 3392
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 27950 3238 28002 3290
rect 28014 3238 28066 3290
rect 28078 3238 28130 3290
rect 28142 3238 28194 3290
rect 28206 3238 28258 3290
rect 37950 3238 38002 3290
rect 38014 3238 38066 3290
rect 38078 3238 38130 3290
rect 38142 3238 38194 3290
rect 38206 3238 38258 3290
rect 47950 3238 48002 3290
rect 48014 3238 48066 3290
rect 48078 3238 48130 3290
rect 48142 3238 48194 3290
rect 48206 3238 48258 3290
rect 1308 3136 1360 3188
rect 21180 3136 21232 3188
rect 23204 3136 23256 3188
rect 16672 3111 16724 3120
rect 16672 3077 16681 3111
rect 16681 3077 16715 3111
rect 16715 3077 16724 3111
rect 16672 3068 16724 3077
rect 1308 3000 1360 3052
rect 13820 3000 13872 3052
rect 19064 3068 19116 3120
rect 22100 3068 22152 3120
rect 22652 3068 22704 3120
rect 11060 2932 11112 2984
rect 2412 2864 2464 2916
rect 15844 2864 15896 2916
rect 20812 3043 20864 3052
rect 20812 3009 20821 3043
rect 20821 3009 20855 3043
rect 20855 3009 20864 3043
rect 20812 3000 20864 3009
rect 21456 3043 21508 3052
rect 21456 3009 21465 3043
rect 21465 3009 21499 3043
rect 21499 3009 21508 3043
rect 21456 3000 21508 3009
rect 23572 3136 23624 3188
rect 23388 3068 23440 3120
rect 26884 3068 26936 3120
rect 18420 2932 18472 2984
rect 20996 2932 21048 2984
rect 22008 2932 22060 2984
rect 24584 2932 24636 2984
rect 37740 3136 37792 3188
rect 27712 3068 27764 3120
rect 29644 3068 29696 3120
rect 49240 3068 49292 3120
rect 28816 3000 28868 3052
rect 39764 3000 39816 3052
rect 45744 3000 45796 3052
rect 47308 3000 47360 3052
rect 25964 2975 26016 2984
rect 25964 2941 25973 2975
rect 25973 2941 26007 2975
rect 26007 2941 26016 2975
rect 25964 2932 26016 2941
rect 29644 2932 29696 2984
rect 30656 2932 30708 2984
rect 46756 2932 46808 2984
rect 46848 2975 46900 2984
rect 46848 2941 46857 2975
rect 46857 2941 46891 2975
rect 46891 2941 46900 2975
rect 46848 2932 46900 2941
rect 22376 2864 22428 2916
rect 22652 2907 22704 2916
rect 22652 2873 22661 2907
rect 22661 2873 22695 2907
rect 22695 2873 22704 2907
rect 22652 2864 22704 2873
rect 23204 2864 23256 2916
rect 2320 2839 2372 2848
rect 2320 2805 2329 2839
rect 2329 2805 2363 2839
rect 2363 2805 2372 2839
rect 2320 2796 2372 2805
rect 2780 2839 2832 2848
rect 2780 2805 2789 2839
rect 2789 2805 2823 2839
rect 2823 2805 2832 2839
rect 2780 2796 2832 2805
rect 21180 2796 21232 2848
rect 23388 2839 23440 2848
rect 23388 2805 23397 2839
rect 23397 2805 23431 2839
rect 23431 2805 23440 2839
rect 23388 2796 23440 2805
rect 23480 2796 23532 2848
rect 26884 2864 26936 2916
rect 27712 2864 27764 2916
rect 24584 2796 24636 2848
rect 27160 2796 27212 2848
rect 27896 2796 27948 2848
rect 38292 2864 38344 2916
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 32950 2694 33002 2746
rect 33014 2694 33066 2746
rect 33078 2694 33130 2746
rect 33142 2694 33194 2746
rect 33206 2694 33258 2746
rect 42950 2694 43002 2746
rect 43014 2694 43066 2746
rect 43078 2694 43130 2746
rect 43142 2694 43194 2746
rect 43206 2694 43258 2746
rect 4344 2524 4396 2576
rect 11060 2592 11112 2644
rect 13544 2592 13596 2644
rect 22284 2592 22336 2644
rect 26884 2592 26936 2644
rect 27528 2592 27580 2644
rect 32864 2592 32916 2644
rect 34428 2592 34480 2644
rect 11704 2456 11756 2508
rect 13820 2456 13872 2508
rect 1308 2388 1360 2440
rect 2780 2388 2832 2440
rect 1216 2320 1268 2372
rect 2320 2320 2372 2372
rect 1308 2252 1360 2304
rect 9680 2388 9732 2440
rect 12808 2388 12860 2440
rect 15844 2388 15896 2440
rect 4344 2320 4396 2372
rect 15936 2320 15988 2372
rect 19524 2388 19576 2440
rect 19616 2431 19668 2440
rect 19616 2397 19625 2431
rect 19625 2397 19659 2431
rect 19659 2397 19668 2431
rect 19616 2388 19668 2397
rect 24216 2524 24268 2576
rect 35900 2524 35952 2576
rect 20168 2456 20220 2508
rect 22284 2456 22336 2508
rect 24400 2456 24452 2508
rect 26516 2456 26568 2508
rect 37740 2499 37792 2508
rect 37740 2465 37749 2499
rect 37749 2465 37783 2499
rect 37783 2465 37792 2499
rect 37740 2456 37792 2465
rect 41328 2456 41380 2508
rect 49148 2499 49200 2508
rect 49148 2465 49157 2499
rect 49157 2465 49191 2499
rect 49191 2465 49200 2499
rect 49148 2456 49200 2465
rect 22376 2431 22428 2440
rect 22376 2397 22385 2431
rect 22385 2397 22419 2431
rect 22419 2397 22428 2431
rect 22376 2388 22428 2397
rect 24584 2431 24636 2440
rect 24584 2397 24593 2431
rect 24593 2397 24627 2431
rect 24627 2397 24636 2431
rect 24584 2388 24636 2397
rect 27160 2431 27212 2440
rect 27160 2397 27169 2431
rect 27169 2397 27203 2431
rect 27203 2397 27212 2431
rect 27160 2388 27212 2397
rect 29000 2388 29052 2440
rect 30748 2388 30800 2440
rect 33140 2431 33192 2440
rect 33140 2397 33149 2431
rect 33149 2397 33183 2431
rect 33183 2397 33192 2431
rect 33140 2388 33192 2397
rect 34980 2388 35032 2440
rect 38292 2388 38344 2440
rect 45652 2388 45704 2440
rect 47216 2388 47268 2440
rect 48504 2320 48556 2372
rect 12716 2252 12768 2304
rect 37096 2295 37148 2304
rect 37096 2261 37105 2295
rect 37105 2261 37139 2295
rect 37139 2261 37148 2295
rect 37096 2252 37148 2261
rect 43444 2252 43496 2304
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 27950 2150 28002 2202
rect 28014 2150 28066 2202
rect 28078 2150 28130 2202
rect 28142 2150 28194 2202
rect 28206 2150 28258 2202
rect 37950 2150 38002 2202
rect 38014 2150 38066 2202
rect 38078 2150 38130 2202
rect 38142 2150 38194 2202
rect 38206 2150 38258 2202
rect 47950 2150 48002 2202
rect 48014 2150 48066 2202
rect 48078 2150 48130 2202
rect 48142 2150 48194 2202
rect 48206 2150 48258 2202
<< metal2 >>
rect 1582 26200 1638 27000
rect 2226 26200 2282 27000
rect 2870 26200 2926 27000
rect 3514 26200 3570 27000
rect 4158 26200 4214 27000
rect 4802 26330 4858 27000
rect 4802 26302 5028 26330
rect 4802 26200 4858 26302
rect 1596 23186 1624 26200
rect 2136 24132 2188 24138
rect 2136 24074 2188 24080
rect 2148 23866 2176 24074
rect 2136 23860 2188 23866
rect 2136 23802 2188 23808
rect 1584 23180 1636 23186
rect 1584 23122 1636 23128
rect 2240 22234 2268 26200
rect 2778 24440 2834 24449
rect 2778 24375 2780 24384
rect 2832 24375 2834 24384
rect 2780 24346 2832 24352
rect 2320 24200 2372 24206
rect 2320 24142 2372 24148
rect 2228 22228 2280 22234
rect 2228 22170 2280 22176
rect 1308 22092 1360 22098
rect 1308 22034 1360 22040
rect 1320 20777 1348 22034
rect 1306 20768 1362 20777
rect 1306 20703 1362 20712
rect 1952 20460 2004 20466
rect 1952 20402 2004 20408
rect 1768 20256 1820 20262
rect 1768 20198 1820 20204
rect 1780 19854 1808 20198
rect 1768 19848 1820 19854
rect 1768 19790 1820 19796
rect 1964 18737 1992 20402
rect 2332 19174 2360 24142
rect 2884 23322 2912 26200
rect 3422 25664 3478 25673
rect 3422 25599 3478 25608
rect 3436 25090 3464 25599
rect 3424 25084 3476 25090
rect 3424 25026 3476 25032
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2950 24443 3258 24452
rect 3528 24274 3556 26200
rect 4066 25256 4122 25265
rect 4066 25191 4122 25200
rect 4080 24954 4108 25191
rect 4068 24948 4120 24954
rect 4068 24890 4120 24896
rect 3882 24848 3938 24857
rect 3882 24783 3938 24792
rect 3896 24614 3924 24783
rect 3884 24608 3936 24614
rect 3884 24550 3936 24556
rect 3516 24268 3568 24274
rect 3516 24210 3568 24216
rect 3790 24032 3846 24041
rect 3790 23967 3846 23976
rect 3700 23724 3752 23730
rect 3700 23666 3752 23672
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 2872 23316 2924 23322
rect 2872 23258 2924 23264
rect 2780 23044 2832 23050
rect 2780 22986 2832 22992
rect 2792 22250 2820 22986
rect 3608 22976 3660 22982
rect 3608 22918 3660 22924
rect 2872 22568 2924 22574
rect 2872 22510 2924 22516
rect 2700 22222 2820 22250
rect 2700 21593 2728 22222
rect 2686 21584 2742 21593
rect 2686 21519 2742 21528
rect 2778 21176 2834 21185
rect 2884 21162 2912 22510
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 3620 21554 3648 22918
rect 3608 21548 3660 21554
rect 3608 21490 3660 21496
rect 3332 21480 3384 21486
rect 3332 21422 3384 21428
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2950 21179 3258 21188
rect 2834 21134 2912 21162
rect 2778 21111 2834 21120
rect 2780 20868 2832 20874
rect 2780 20810 2832 20816
rect 2792 19904 2820 20810
rect 2872 20392 2924 20398
rect 2872 20334 2924 20340
rect 2700 19876 2820 19904
rect 2700 19553 2728 19876
rect 2780 19780 2832 19786
rect 2780 19722 2832 19728
rect 2686 19544 2742 19553
rect 2686 19479 2742 19488
rect 2320 19168 2372 19174
rect 2320 19110 2372 19116
rect 2792 18873 2820 19722
rect 2884 19530 2912 20334
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 3344 19961 3372 21422
rect 3330 19952 3386 19961
rect 3330 19887 3386 19896
rect 2884 19502 3004 19530
rect 2872 19440 2924 19446
rect 2872 19382 2924 19388
rect 2778 18864 2834 18873
rect 2778 18799 2834 18808
rect 1950 18728 2006 18737
rect 1950 18663 2006 18672
rect 2780 18692 2832 18698
rect 2780 18634 2832 18640
rect 2792 18306 2820 18634
rect 2884 18329 2912 19382
rect 2976 19281 3004 19502
rect 2962 19272 3018 19281
rect 2962 19207 3018 19216
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 2700 18278 2820 18306
rect 2870 18320 2926 18329
rect 2700 17921 2728 18278
rect 3712 18290 3740 23666
rect 3804 18834 3832 23967
rect 4172 23798 4200 26200
rect 4160 23792 4212 23798
rect 4160 23734 4212 23740
rect 4712 23724 4764 23730
rect 4712 23666 4764 23672
rect 4066 23624 4122 23633
rect 4066 23559 4068 23568
rect 4120 23559 4122 23568
rect 4068 23530 4120 23536
rect 4724 23322 4752 23666
rect 4804 23520 4856 23526
rect 4804 23462 4856 23468
rect 4344 23316 4396 23322
rect 4344 23258 4396 23264
rect 4712 23316 4764 23322
rect 4712 23258 4764 23264
rect 4066 23216 4122 23225
rect 4066 23151 4122 23160
rect 3974 22808 4030 22817
rect 4080 22778 4108 23151
rect 3974 22743 4030 22752
rect 4068 22772 4120 22778
rect 3988 22166 4016 22743
rect 4068 22714 4120 22720
rect 4080 22596 4292 22624
rect 4080 22545 4108 22596
rect 4066 22536 4122 22545
rect 4066 22471 4122 22480
rect 4160 22500 4212 22506
rect 4160 22442 4212 22448
rect 3976 22160 4028 22166
rect 3976 22102 4028 22108
rect 3884 22092 3936 22098
rect 3884 22034 3936 22040
rect 3896 22001 3924 22034
rect 4068 22024 4120 22030
rect 3882 21992 3938 22001
rect 4068 21966 4120 21972
rect 3882 21927 3938 21936
rect 4080 21690 4108 21966
rect 4068 21684 4120 21690
rect 4068 21626 4120 21632
rect 4172 20398 4200 22442
rect 4264 21010 4292 22596
rect 4356 21622 4384 23258
rect 4436 23180 4488 23186
rect 4436 23122 4488 23128
rect 4344 21616 4396 21622
rect 4344 21558 4396 21564
rect 4344 21344 4396 21350
rect 4344 21286 4396 21292
rect 4252 21004 4304 21010
rect 4252 20946 4304 20952
rect 4356 20942 4384 21286
rect 4344 20936 4396 20942
rect 4344 20878 4396 20884
rect 3884 20392 3936 20398
rect 3882 20360 3884 20369
rect 4160 20392 4212 20398
rect 3936 20360 3938 20369
rect 4160 20334 4212 20340
rect 3882 20295 3938 20304
rect 4448 19446 4476 23122
rect 4528 23112 4580 23118
rect 4528 23054 4580 23060
rect 4436 19440 4488 19446
rect 4436 19382 4488 19388
rect 3792 18828 3844 18834
rect 3792 18770 3844 18776
rect 2870 18255 2926 18264
rect 3700 18284 3752 18290
rect 3700 18226 3752 18232
rect 2780 18216 2832 18222
rect 2780 18158 2832 18164
rect 4160 18216 4212 18222
rect 4160 18158 4212 18164
rect 2686 17912 2742 17921
rect 2686 17847 2742 17856
rect 1216 17740 1268 17746
rect 1216 17682 1268 17688
rect 1228 17105 1256 17682
rect 2792 17513 2820 18158
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 2778 17504 2834 17513
rect 2778 17439 2834 17448
rect 1308 17128 1360 17134
rect 1214 17096 1270 17105
rect 1308 17070 1360 17076
rect 1214 17031 1270 17040
rect 1320 16697 1348 17070
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 1306 16688 1362 16697
rect 1306 16623 1362 16632
rect 1308 16516 1360 16522
rect 1308 16458 1360 16464
rect 1320 16289 1348 16458
rect 1306 16280 1362 16289
rect 1306 16215 1362 16224
rect 4172 16046 4200 18158
rect 4540 16658 4568 23054
rect 4816 22642 4844 23462
rect 4804 22636 4856 22642
rect 4804 22578 4856 22584
rect 5000 22574 5028 26302
rect 5446 26200 5502 27000
rect 6090 26200 6146 27000
rect 6734 26200 6790 27000
rect 7378 26330 7434 27000
rect 8022 26330 8078 27000
rect 7378 26302 7696 26330
rect 7378 26200 7434 26302
rect 5460 23662 5488 26200
rect 5540 24064 5592 24070
rect 5540 24006 5592 24012
rect 5448 23656 5500 23662
rect 5448 23598 5500 23604
rect 5552 23118 5580 24006
rect 6104 23186 6132 26200
rect 6644 24608 6696 24614
rect 6644 24550 6696 24556
rect 6184 24404 6236 24410
rect 6184 24346 6236 24352
rect 6092 23180 6144 23186
rect 6092 23122 6144 23128
rect 5080 23112 5132 23118
rect 5080 23054 5132 23060
rect 5540 23112 5592 23118
rect 5540 23054 5592 23060
rect 4988 22568 5040 22574
rect 4988 22510 5040 22516
rect 4896 22228 4948 22234
rect 4896 22170 4948 22176
rect 4804 20256 4856 20262
rect 4804 20198 4856 20204
rect 4816 19990 4844 20198
rect 4804 19984 4856 19990
rect 4804 19926 4856 19932
rect 4908 19922 4936 22170
rect 4988 20256 5040 20262
rect 4988 20198 5040 20204
rect 4896 19916 4948 19922
rect 4896 19858 4948 19864
rect 5000 18358 5028 20198
rect 5092 18426 5120 23054
rect 5540 22772 5592 22778
rect 5540 22714 5592 22720
rect 5264 21480 5316 21486
rect 5264 21422 5316 21428
rect 5276 20602 5304 21422
rect 5552 21010 5580 22714
rect 5908 21548 5960 21554
rect 5908 21490 5960 21496
rect 5920 21457 5948 21490
rect 5906 21448 5962 21457
rect 5632 21412 5684 21418
rect 5906 21383 5962 21392
rect 5632 21354 5684 21360
rect 5540 21004 5592 21010
rect 5540 20946 5592 20952
rect 5264 20596 5316 20602
rect 5264 20538 5316 20544
rect 5356 19372 5408 19378
rect 5356 19314 5408 19320
rect 5080 18420 5132 18426
rect 5080 18362 5132 18368
rect 4988 18352 5040 18358
rect 4988 18294 5040 18300
rect 5368 16794 5396 19314
rect 5644 18426 5672 21354
rect 6196 19922 6224 24346
rect 6460 22024 6512 22030
rect 6460 21966 6512 21972
rect 6472 21078 6500 21966
rect 6460 21072 6512 21078
rect 6460 21014 6512 21020
rect 6656 20398 6684 24550
rect 6748 24342 6776 26200
rect 6736 24336 6788 24342
rect 6736 24278 6788 24284
rect 7378 24304 7434 24313
rect 7378 24239 7434 24248
rect 7392 24206 7420 24239
rect 7380 24200 7432 24206
rect 7380 24142 7432 24148
rect 7472 24064 7524 24070
rect 7472 24006 7524 24012
rect 6736 23588 6788 23594
rect 6736 23530 6788 23536
rect 6748 21486 6776 23530
rect 6920 22976 6972 22982
rect 6920 22918 6972 22924
rect 7012 22976 7064 22982
rect 7012 22918 7064 22924
rect 6932 22234 6960 22918
rect 6920 22228 6972 22234
rect 6920 22170 6972 22176
rect 6736 21480 6788 21486
rect 6736 21422 6788 21428
rect 6644 20392 6696 20398
rect 6644 20334 6696 20340
rect 7024 20058 7052 22918
rect 7484 22642 7512 24006
rect 7472 22636 7524 22642
rect 7472 22578 7524 22584
rect 7668 22574 7696 26302
rect 7852 26302 8078 26330
rect 7748 24404 7800 24410
rect 7748 24346 7800 24352
rect 7760 23730 7788 24346
rect 7748 23724 7800 23730
rect 7748 23666 7800 23672
rect 7852 23186 7880 26302
rect 8022 26200 8078 26302
rect 8666 26200 8722 27000
rect 9310 26200 9366 27000
rect 9954 26330 10010 27000
rect 10598 26330 10654 27000
rect 9954 26302 10272 26330
rect 9954 26200 10010 26302
rect 8680 24274 8708 26200
rect 8852 24948 8904 24954
rect 8852 24890 8904 24896
rect 8668 24268 8720 24274
rect 8668 24210 8720 24216
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 8392 23656 8444 23662
rect 8392 23598 8444 23604
rect 7840 23180 7892 23186
rect 7840 23122 7892 23128
rect 7748 23044 7800 23050
rect 7748 22986 7800 22992
rect 7656 22568 7708 22574
rect 7656 22510 7708 22516
rect 7104 22432 7156 22438
rect 7104 22374 7156 22380
rect 7012 20052 7064 20058
rect 7012 19994 7064 20000
rect 6184 19916 6236 19922
rect 6184 19858 6236 19864
rect 7116 19786 7144 22374
rect 7760 21146 7788 22986
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 8404 22234 8432 23598
rect 8668 22432 8720 22438
rect 8668 22374 8720 22380
rect 8392 22228 8444 22234
rect 8392 22170 8444 22176
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 8576 21548 8628 21554
rect 8576 21490 8628 21496
rect 8588 21418 8616 21490
rect 8576 21412 8628 21418
rect 8576 21354 8628 21360
rect 7748 21140 7800 21146
rect 7748 21082 7800 21088
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 8392 20528 8444 20534
rect 8392 20470 8444 20476
rect 7104 19780 7156 19786
rect 7104 19722 7156 19728
rect 7840 19780 7892 19786
rect 7840 19722 7892 19728
rect 5632 18420 5684 18426
rect 5632 18362 5684 18368
rect 5356 16788 5408 16794
rect 5356 16730 5408 16736
rect 4528 16652 4580 16658
rect 4528 16594 4580 16600
rect 1308 16040 1360 16046
rect 1308 15982 1360 15988
rect 4160 16040 4212 16046
rect 4160 15982 4212 15988
rect 1320 15881 1348 15982
rect 1306 15872 1362 15881
rect 1306 15807 1362 15816
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 1308 15564 1360 15570
rect 1308 15506 1360 15512
rect 1320 15473 1348 15506
rect 1306 15464 1362 15473
rect 1306 15399 1362 15408
rect 1306 15056 1362 15065
rect 1306 14991 1362 15000
rect 1320 14958 1348 14991
rect 1308 14952 1360 14958
rect 1308 14894 1360 14900
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 1306 14648 1362 14657
rect 2950 14651 3258 14660
rect 1306 14583 1362 14592
rect 1320 14482 1348 14583
rect 1308 14476 1360 14482
rect 1308 14418 1360 14424
rect 1306 14240 1362 14249
rect 1306 14175 1362 14184
rect 1320 13870 1348 14175
rect 3516 13932 3568 13938
rect 3516 13874 3568 13880
rect 1308 13864 1360 13870
rect 1308 13806 1360 13812
rect 2778 13832 2834 13841
rect 2778 13767 2834 13776
rect 2792 13326 2820 13767
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 3528 13433 3556 13874
rect 3514 13424 3570 13433
rect 3514 13359 3570 13368
rect 2780 13320 2832 13326
rect 2780 13262 2832 13268
rect 1306 13016 1362 13025
rect 1306 12951 1362 12960
rect 1320 12918 1348 12951
rect 1308 12912 1360 12918
rect 1308 12854 1360 12860
rect 1216 12844 1268 12850
rect 1216 12786 1268 12792
rect 1228 12617 1256 12786
rect 1214 12608 1270 12617
rect 1214 12543 1270 12552
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 1308 12232 1360 12238
rect 1214 12200 1270 12209
rect 1308 12174 1360 12180
rect 1214 12135 1270 12144
rect 1228 11762 1256 12135
rect 1320 11801 1348 12174
rect 4172 11898 4200 15982
rect 5368 12434 5396 16730
rect 5448 16652 5500 16658
rect 5448 16594 5500 16600
rect 5460 12986 5488 16594
rect 7852 16454 7880 19722
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 8404 19174 8432 20470
rect 8392 19168 8444 19174
rect 8392 19110 8444 19116
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 8312 17202 8340 18566
rect 8300 17196 8352 17202
rect 8300 17138 8352 17144
rect 7840 16448 7892 16454
rect 7840 16390 7892 16396
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 8404 16250 8432 19110
rect 8680 18834 8708 22374
rect 8864 21486 8892 24890
rect 9128 24064 9180 24070
rect 9128 24006 9180 24012
rect 9140 23118 9168 24006
rect 9324 23798 9352 26200
rect 10048 25084 10100 25090
rect 10048 25026 10100 25032
rect 9772 24064 9824 24070
rect 9772 24006 9824 24012
rect 9312 23792 9364 23798
rect 9312 23734 9364 23740
rect 9128 23112 9180 23118
rect 9128 23054 9180 23060
rect 9128 22500 9180 22506
rect 9128 22442 9180 22448
rect 9140 22030 9168 22442
rect 9128 22024 9180 22030
rect 9128 21966 9180 21972
rect 9680 21888 9732 21894
rect 9680 21830 9732 21836
rect 8852 21480 8904 21486
rect 8758 21448 8814 21457
rect 8852 21422 8904 21428
rect 8758 21383 8814 21392
rect 8772 21350 8800 21383
rect 8760 21344 8812 21350
rect 8760 21286 8812 21292
rect 9692 20602 9720 21830
rect 9784 21690 9812 24006
rect 10060 22098 10088 25026
rect 10140 24336 10192 24342
rect 10140 24278 10192 24284
rect 10048 22092 10100 22098
rect 10152 22094 10180 24278
rect 10244 22574 10272 26302
rect 10598 26302 10732 26330
rect 10598 26200 10654 26302
rect 10704 23798 10732 26302
rect 11242 26200 11298 27000
rect 11886 26200 11942 27000
rect 12530 26200 12586 27000
rect 13174 26330 13230 27000
rect 13174 26302 13400 26330
rect 13174 26200 13230 26302
rect 10876 24132 10928 24138
rect 10876 24074 10928 24080
rect 10888 23798 10916 24074
rect 10692 23792 10744 23798
rect 10692 23734 10744 23740
rect 10876 23792 10928 23798
rect 10876 23734 10928 23740
rect 10324 23588 10376 23594
rect 10324 23530 10376 23536
rect 10232 22568 10284 22574
rect 10232 22510 10284 22516
rect 10152 22066 10272 22094
rect 10048 22034 10100 22040
rect 9864 21888 9916 21894
rect 9864 21830 9916 21836
rect 9772 21684 9824 21690
rect 9772 21626 9824 21632
rect 9876 20942 9904 21830
rect 10048 21616 10100 21622
rect 10048 21558 10100 21564
rect 9956 21344 10008 21350
rect 9956 21286 10008 21292
rect 9864 20936 9916 20942
rect 9864 20878 9916 20884
rect 9680 20596 9732 20602
rect 9680 20538 9732 20544
rect 9968 20058 9996 21286
rect 10060 20262 10088 21558
rect 10048 20256 10100 20262
rect 10048 20198 10100 20204
rect 9956 20052 10008 20058
rect 9956 19994 10008 20000
rect 9772 19848 9824 19854
rect 9772 19790 9824 19796
rect 9312 19508 9364 19514
rect 9312 19450 9364 19456
rect 8668 18828 8720 18834
rect 8668 18770 8720 18776
rect 8576 17672 8628 17678
rect 8576 17614 8628 17620
rect 8588 16658 8616 17614
rect 8484 16652 8536 16658
rect 8484 16594 8536 16600
rect 8576 16652 8628 16658
rect 8576 16594 8628 16600
rect 8392 16244 8444 16250
rect 8392 16186 8444 16192
rect 8496 16046 8524 16594
rect 9324 16250 9352 19450
rect 9680 19304 9732 19310
rect 9680 19246 9732 19252
rect 9404 19236 9456 19242
rect 9404 19178 9456 19184
rect 9416 18698 9444 19178
rect 9404 18692 9456 18698
rect 9404 18634 9456 18640
rect 9692 18426 9720 19246
rect 9680 18420 9732 18426
rect 9680 18362 9732 18368
rect 9784 16561 9812 19790
rect 9968 17202 9996 19994
rect 10048 19780 10100 19786
rect 10048 19722 10100 19728
rect 10060 19514 10088 19722
rect 10048 19508 10100 19514
rect 10048 19450 10100 19456
rect 10244 18154 10272 22066
rect 10336 20602 10364 23530
rect 11256 23186 11284 26200
rect 11900 24342 11928 26200
rect 11888 24336 11940 24342
rect 11888 24278 11940 24284
rect 11704 24064 11756 24070
rect 11704 24006 11756 24012
rect 11796 24064 11848 24070
rect 11796 24006 11848 24012
rect 11244 23180 11296 23186
rect 11244 23122 11296 23128
rect 11060 22772 11112 22778
rect 11060 22714 11112 22720
rect 11072 22098 11100 22714
rect 11716 22642 11744 24006
rect 11808 23866 11836 24006
rect 11796 23860 11848 23866
rect 11796 23802 11848 23808
rect 12348 23792 12400 23798
rect 12348 23734 12400 23740
rect 12360 23526 12388 23734
rect 12440 23724 12492 23730
rect 12440 23666 12492 23672
rect 12348 23520 12400 23526
rect 12348 23462 12400 23468
rect 12348 23112 12400 23118
rect 12348 23054 12400 23060
rect 12256 22772 12308 22778
rect 12256 22714 12308 22720
rect 11704 22636 11756 22642
rect 11704 22578 11756 22584
rect 12268 22574 12296 22714
rect 12256 22568 12308 22574
rect 12256 22510 12308 22516
rect 12360 22234 12388 23054
rect 12348 22228 12400 22234
rect 12348 22170 12400 22176
rect 11152 22160 11204 22166
rect 11152 22102 11204 22108
rect 11060 22092 11112 22098
rect 11060 22034 11112 22040
rect 11164 21962 11192 22102
rect 11336 22024 11388 22030
rect 11336 21966 11388 21972
rect 11152 21956 11204 21962
rect 11152 21898 11204 21904
rect 11348 21457 11376 21966
rect 11980 21548 12032 21554
rect 11980 21490 12032 21496
rect 11334 21448 11390 21457
rect 11334 21383 11390 21392
rect 11888 21344 11940 21350
rect 11888 21286 11940 21292
rect 10508 21072 10560 21078
rect 10508 21014 10560 21020
rect 11334 21040 11390 21049
rect 10324 20596 10376 20602
rect 10324 20538 10376 20544
rect 10416 20392 10468 20398
rect 10416 20334 10468 20340
rect 10428 18154 10456 20334
rect 10520 19718 10548 21014
rect 11334 20975 11390 20984
rect 11796 21004 11848 21010
rect 11348 20942 11376 20975
rect 11796 20946 11848 20952
rect 11244 20936 11296 20942
rect 11244 20878 11296 20884
rect 11336 20936 11388 20942
rect 11336 20878 11388 20884
rect 11060 20800 11112 20806
rect 11256 20788 11284 20878
rect 11256 20760 11376 20788
rect 11060 20742 11112 20748
rect 10600 20528 10652 20534
rect 10600 20470 10652 20476
rect 10612 19854 10640 20470
rect 10968 20392 11020 20398
rect 10968 20334 11020 20340
rect 10876 20324 10928 20330
rect 10876 20266 10928 20272
rect 10888 19990 10916 20266
rect 10876 19984 10928 19990
rect 10876 19926 10928 19932
rect 10600 19848 10652 19854
rect 10980 19825 11008 20334
rect 10600 19790 10652 19796
rect 10966 19816 11022 19825
rect 10966 19751 11022 19760
rect 10508 19712 10560 19718
rect 10508 19654 10560 19660
rect 10232 18148 10284 18154
rect 10232 18090 10284 18096
rect 10416 18148 10468 18154
rect 10416 18090 10468 18096
rect 10324 18080 10376 18086
rect 10324 18022 10376 18028
rect 9956 17196 10008 17202
rect 9956 17138 10008 17144
rect 9864 16992 9916 16998
rect 9864 16934 9916 16940
rect 9770 16552 9826 16561
rect 9588 16516 9640 16522
rect 9770 16487 9826 16496
rect 9588 16458 9640 16464
rect 9312 16244 9364 16250
rect 9312 16186 9364 16192
rect 8484 16040 8536 16046
rect 8484 15982 8536 15988
rect 9220 15904 9272 15910
rect 9220 15846 9272 15852
rect 6552 15360 6604 15366
rect 6552 15302 6604 15308
rect 6564 15026 6592 15302
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 9232 15162 9260 15846
rect 9220 15156 9272 15162
rect 9220 15098 9272 15104
rect 9600 15094 9628 16458
rect 9588 15088 9640 15094
rect 9588 15030 9640 15036
rect 6552 15020 6604 15026
rect 6552 14962 6604 14968
rect 9588 14340 9640 14346
rect 9588 14282 9640 14288
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 9600 13870 9628 14282
rect 9588 13864 9640 13870
rect 9588 13806 9640 13812
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 5448 12980 5500 12986
rect 5448 12922 5500 12928
rect 9876 12782 9904 16934
rect 10336 16250 10364 18022
rect 10520 16697 10548 19654
rect 10876 19372 10928 19378
rect 10876 19314 10928 19320
rect 10888 18902 10916 19314
rect 11072 18970 11100 20742
rect 11152 19372 11204 19378
rect 11152 19314 11204 19320
rect 11060 18964 11112 18970
rect 11060 18906 11112 18912
rect 10876 18896 10928 18902
rect 10876 18838 10928 18844
rect 10600 18828 10652 18834
rect 10600 18770 10652 18776
rect 10612 18154 10640 18770
rect 10600 18148 10652 18154
rect 10600 18090 10652 18096
rect 10612 17746 10640 18090
rect 10600 17740 10652 17746
rect 10600 17682 10652 17688
rect 10506 16688 10562 16697
rect 10506 16623 10562 16632
rect 10508 16516 10560 16522
rect 10508 16458 10560 16464
rect 10324 16244 10376 16250
rect 10324 16186 10376 16192
rect 10232 15904 10284 15910
rect 10232 15846 10284 15852
rect 10048 14952 10100 14958
rect 10048 14894 10100 14900
rect 10060 13802 10088 14894
rect 10244 14074 10272 15846
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 10428 14618 10456 15438
rect 10520 15337 10548 16458
rect 10612 15570 10640 17682
rect 10690 17232 10746 17241
rect 10690 17167 10746 17176
rect 10704 17134 10732 17167
rect 10692 17128 10744 17134
rect 10692 17070 10744 17076
rect 10888 16658 10916 18838
rect 11060 18216 11112 18222
rect 11164 18193 11192 19314
rect 11348 19310 11376 20760
rect 11808 20482 11836 20946
rect 11900 20602 11928 21286
rect 11888 20596 11940 20602
rect 11888 20538 11940 20544
rect 11808 20466 11928 20482
rect 11428 20460 11480 20466
rect 11808 20460 11940 20466
rect 11808 20454 11888 20460
rect 11428 20402 11480 20408
rect 11888 20402 11940 20408
rect 11336 19304 11388 19310
rect 11336 19246 11388 19252
rect 11244 19236 11296 19242
rect 11244 19178 11296 19184
rect 11060 18158 11112 18164
rect 11150 18184 11206 18193
rect 11072 17882 11100 18158
rect 11150 18119 11206 18128
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 11060 17060 11112 17066
rect 11060 17002 11112 17008
rect 10876 16652 10928 16658
rect 10876 16594 10928 16600
rect 11072 16590 11100 17002
rect 11060 16584 11112 16590
rect 11060 16526 11112 16532
rect 11256 16182 11284 19178
rect 11440 18970 11468 20402
rect 11888 19168 11940 19174
rect 11888 19110 11940 19116
rect 11428 18964 11480 18970
rect 11428 18906 11480 18912
rect 11900 18902 11928 19110
rect 11888 18896 11940 18902
rect 11888 18838 11940 18844
rect 11520 18760 11572 18766
rect 11520 18702 11572 18708
rect 11888 18760 11940 18766
rect 11888 18702 11940 18708
rect 11428 18284 11480 18290
rect 11428 18226 11480 18232
rect 11336 16448 11388 16454
rect 11336 16390 11388 16396
rect 11152 16176 11204 16182
rect 11152 16118 11204 16124
rect 11244 16176 11296 16182
rect 11244 16118 11296 16124
rect 10784 16108 10836 16114
rect 10784 16050 10836 16056
rect 10876 16108 10928 16114
rect 10876 16050 10928 16056
rect 10796 15706 10824 16050
rect 10784 15700 10836 15706
rect 10784 15642 10836 15648
rect 10600 15564 10652 15570
rect 10600 15506 10652 15512
rect 10506 15328 10562 15337
rect 10506 15263 10562 15272
rect 10416 14612 10468 14618
rect 10416 14554 10468 14560
rect 10322 14512 10378 14521
rect 10322 14447 10378 14456
rect 10336 14414 10364 14447
rect 10324 14408 10376 14414
rect 10324 14350 10376 14356
rect 10692 14408 10744 14414
rect 10692 14350 10744 14356
rect 10336 14074 10364 14350
rect 10704 14074 10732 14350
rect 10232 14068 10284 14074
rect 10232 14010 10284 14016
rect 10324 14068 10376 14074
rect 10324 14010 10376 14016
rect 10692 14068 10744 14074
rect 10692 14010 10744 14016
rect 10048 13796 10100 13802
rect 10048 13738 10100 13744
rect 9864 12776 9916 12782
rect 9864 12718 9916 12724
rect 5368 12406 5488 12434
rect 5460 12306 5488 12406
rect 5448 12300 5500 12306
rect 5448 12242 5500 12248
rect 10060 12170 10088 13738
rect 10888 13734 10916 16050
rect 11060 16040 11112 16046
rect 11060 15982 11112 15988
rect 11072 15910 11100 15982
rect 11060 15904 11112 15910
rect 11060 15846 11112 15852
rect 11164 15094 11192 16118
rect 11152 15088 11204 15094
rect 11152 15030 11204 15036
rect 11152 14952 11204 14958
rect 11152 14894 11204 14900
rect 10968 14816 11020 14822
rect 10968 14758 11020 14764
rect 10876 13728 10928 13734
rect 10876 13670 10928 13676
rect 10980 12986 11008 14758
rect 11060 13388 11112 13394
rect 11060 13330 11112 13336
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 11072 12306 11100 13330
rect 11060 12300 11112 12306
rect 11060 12242 11112 12248
rect 10048 12164 10100 12170
rect 10048 12106 10100 12112
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 4160 11892 4212 11898
rect 4160 11834 4212 11840
rect 1306 11792 1362 11801
rect 1216 11756 1268 11762
rect 1306 11727 1362 11736
rect 1216 11698 1268 11704
rect 1228 11354 1256 11698
rect 1308 11688 1360 11694
rect 1308 11630 1360 11636
rect 1320 11393 1348 11630
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 1306 11384 1362 11393
rect 2950 11387 3258 11396
rect 1216 11348 1268 11354
rect 1306 11319 1362 11328
rect 1216 11290 1268 11296
rect 1768 11280 1820 11286
rect 1768 11222 1820 11228
rect 1584 11144 1636 11150
rect 1780 11121 1808 11222
rect 1584 11086 1636 11092
rect 1766 11112 1822 11121
rect 1596 10985 1624 11086
rect 1766 11047 1822 11056
rect 1768 11008 1820 11014
rect 1582 10976 1638 10985
rect 1768 10950 1820 10956
rect 1582 10911 1638 10920
rect 1780 10810 1808 10950
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 1768 10804 1820 10810
rect 1768 10746 1820 10752
rect 1860 10804 1912 10810
rect 1860 10746 1912 10752
rect 1216 10736 1268 10742
rect 1216 10678 1268 10684
rect 1228 10169 1256 10678
rect 1308 10668 1360 10674
rect 1308 10610 1360 10616
rect 1320 10577 1348 10610
rect 1306 10568 1362 10577
rect 1306 10503 1362 10512
rect 1214 10160 1270 10169
rect 1872 10130 1900 10746
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 1214 10095 1270 10104
rect 1860 10124 1912 10130
rect 1860 10066 1912 10072
rect 1308 10056 1360 10062
rect 1308 9998 1360 10004
rect 1320 9761 1348 9998
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 1306 9752 1362 9761
rect 7950 9755 8258 9764
rect 1306 9687 1308 9696
rect 1360 9687 1362 9696
rect 1308 9658 1360 9664
rect 1308 9580 1360 9586
rect 1308 9522 1360 9528
rect 1320 9353 1348 9522
rect 1766 9480 1822 9489
rect 1766 9415 1768 9424
rect 1820 9415 1822 9424
rect 1768 9386 1820 9392
rect 1306 9344 1362 9353
rect 1306 9279 1362 9288
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 11164 9110 11192 14894
rect 11244 14272 11296 14278
rect 11244 14214 11296 14220
rect 11256 14006 11284 14214
rect 11244 14000 11296 14006
rect 11244 13942 11296 13948
rect 11244 12096 11296 12102
rect 11244 12038 11296 12044
rect 11256 11694 11284 12038
rect 11244 11688 11296 11694
rect 11244 11630 11296 11636
rect 11256 11082 11284 11630
rect 11244 11076 11296 11082
rect 11244 11018 11296 11024
rect 2320 9104 2372 9110
rect 2320 9046 2372 9052
rect 11152 9104 11204 9110
rect 11152 9046 11204 9052
rect 1216 8968 1268 8974
rect 1216 8910 1268 8916
rect 1306 8936 1362 8945
rect 1228 8537 1256 8910
rect 1306 8871 1308 8880
rect 1360 8871 1362 8880
rect 1308 8842 1360 8848
rect 1214 8528 1270 8537
rect 1214 8463 1270 8472
rect 1400 8424 1452 8430
rect 1400 8366 1452 8372
rect 1412 8129 1440 8366
rect 1398 8120 1454 8129
rect 1398 8055 1400 8064
rect 1452 8055 1454 8064
rect 1400 8026 1452 8032
rect 1308 7880 1360 7886
rect 1308 7822 1360 7828
rect 1320 7721 1348 7822
rect 1306 7712 1362 7721
rect 1306 7647 1362 7656
rect 1308 7404 1360 7410
rect 1308 7346 1360 7352
rect 1320 7313 1348 7346
rect 1306 7304 1362 7313
rect 1306 7239 1362 7248
rect 1214 6896 1270 6905
rect 1214 6831 1270 6840
rect 1228 6730 1256 6831
rect 1308 6792 1360 6798
rect 1308 6734 1360 6740
rect 1216 6724 1268 6730
rect 1216 6666 1268 6672
rect 1228 6458 1256 6666
rect 1320 6497 1348 6734
rect 2332 6662 2360 9046
rect 11348 8974 11376 16390
rect 11440 14890 11468 18226
rect 11532 17610 11560 18702
rect 11704 18692 11756 18698
rect 11704 18634 11756 18640
rect 11612 18352 11664 18358
rect 11612 18294 11664 18300
rect 11520 17604 11572 17610
rect 11520 17546 11572 17552
rect 11532 16590 11560 17546
rect 11520 16584 11572 16590
rect 11520 16526 11572 16532
rect 11520 16448 11572 16454
rect 11520 16390 11572 16396
rect 11532 16250 11560 16390
rect 11520 16244 11572 16250
rect 11520 16186 11572 16192
rect 11428 14884 11480 14890
rect 11428 14826 11480 14832
rect 11624 14618 11652 18294
rect 11716 16998 11744 18634
rect 11900 18358 11928 18702
rect 11888 18352 11940 18358
rect 11888 18294 11940 18300
rect 11992 17814 12020 21490
rect 12452 21146 12480 23666
rect 12544 22574 12572 26200
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 12624 24132 12676 24138
rect 12624 24074 12676 24080
rect 12532 22568 12584 22574
rect 12532 22510 12584 22516
rect 12532 22024 12584 22030
rect 12532 21966 12584 21972
rect 12440 21140 12492 21146
rect 12440 21082 12492 21088
rect 12072 20868 12124 20874
rect 12072 20810 12124 20816
rect 12084 19530 12112 20810
rect 12440 20800 12492 20806
rect 12440 20742 12492 20748
rect 12452 20482 12480 20742
rect 12176 20454 12480 20482
rect 12176 19786 12204 20454
rect 12164 19780 12216 19786
rect 12164 19722 12216 19728
rect 12256 19780 12308 19786
rect 12256 19722 12308 19728
rect 12084 19502 12204 19530
rect 12072 19372 12124 19378
rect 12072 19314 12124 19320
rect 12084 18873 12112 19314
rect 12070 18864 12126 18873
rect 12070 18799 12126 18808
rect 12176 18170 12204 19502
rect 12084 18142 12204 18170
rect 11980 17808 12032 17814
rect 11980 17750 12032 17756
rect 11796 17264 11848 17270
rect 11796 17206 11848 17212
rect 11808 17105 11836 17206
rect 11980 17128 12032 17134
rect 11794 17096 11850 17105
rect 11980 17070 12032 17076
rect 11794 17031 11850 17040
rect 11704 16992 11756 16998
rect 11704 16934 11756 16940
rect 11992 16794 12020 17070
rect 11980 16788 12032 16794
rect 11980 16730 12032 16736
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 11716 15434 11744 16526
rect 12084 16096 12112 18142
rect 12164 18080 12216 18086
rect 12164 18022 12216 18028
rect 12176 17762 12204 18022
rect 12268 17882 12296 19722
rect 12348 18080 12400 18086
rect 12348 18022 12400 18028
rect 12256 17876 12308 17882
rect 12256 17818 12308 17824
rect 12176 17746 12296 17762
rect 12176 17740 12308 17746
rect 12176 17734 12256 17740
rect 12256 17682 12308 17688
rect 12256 17536 12308 17542
rect 12360 17524 12388 18022
rect 12544 17882 12572 21966
rect 12636 21690 12664 24074
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 13372 23186 13400 26302
rect 13818 26200 13874 27000
rect 14462 26200 14518 27000
rect 15106 26200 15162 27000
rect 15750 26200 15806 27000
rect 16394 26330 16450 27000
rect 16132 26302 16450 26330
rect 13832 24274 13860 26200
rect 13820 24268 13872 24274
rect 13820 24210 13872 24216
rect 13728 24200 13780 24206
rect 13728 24142 13780 24148
rect 14372 24200 14424 24206
rect 14372 24142 14424 24148
rect 13360 23180 13412 23186
rect 13360 23122 13412 23128
rect 12716 22772 12768 22778
rect 12716 22714 12768 22720
rect 13544 22772 13596 22778
rect 13544 22714 13596 22720
rect 12728 22642 12756 22714
rect 12716 22636 12768 22642
rect 12716 22578 12768 22584
rect 13556 22574 13584 22714
rect 13544 22568 13596 22574
rect 13544 22510 13596 22516
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 12716 21956 12768 21962
rect 12716 21898 12768 21904
rect 12624 21684 12676 21690
rect 12624 21626 12676 21632
rect 12728 20534 12756 21898
rect 12808 21548 12860 21554
rect 12808 21490 12860 21496
rect 12820 21078 12848 21490
rect 13452 21480 13504 21486
rect 13452 21422 13504 21428
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 12992 21140 13044 21146
rect 12992 21082 13044 21088
rect 12808 21072 12860 21078
rect 12808 21014 12860 21020
rect 12808 20868 12860 20874
rect 12808 20810 12860 20816
rect 12716 20528 12768 20534
rect 12716 20470 12768 20476
rect 12624 19440 12676 19446
rect 12624 19382 12676 19388
rect 12636 18766 12664 19382
rect 12716 19372 12768 19378
rect 12716 19314 12768 19320
rect 12624 18760 12676 18766
rect 12624 18702 12676 18708
rect 12728 18426 12756 19314
rect 12716 18420 12768 18426
rect 12716 18362 12768 18368
rect 12532 17876 12584 17882
rect 12532 17818 12584 17824
rect 12820 17660 12848 20810
rect 13004 20806 13032 21082
rect 12992 20800 13044 20806
rect 12992 20742 13044 20748
rect 13360 20596 13412 20602
rect 13360 20538 13412 20544
rect 13268 20528 13320 20534
rect 13268 20470 13320 20476
rect 13280 20262 13308 20470
rect 13268 20256 13320 20262
rect 13268 20198 13320 20204
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 13372 19961 13400 20538
rect 13358 19952 13414 19961
rect 13358 19887 13414 19896
rect 13360 19508 13412 19514
rect 13360 19450 13412 19456
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 13372 18834 13400 19450
rect 13360 18828 13412 18834
rect 13360 18770 13412 18776
rect 13268 18760 13320 18766
rect 13268 18702 13320 18708
rect 13280 18154 13308 18702
rect 13372 18222 13400 18770
rect 13464 18766 13492 21422
rect 13556 20448 13584 22510
rect 13740 22098 13768 24142
rect 14188 23792 14240 23798
rect 14188 23734 14240 23740
rect 14200 23322 14228 23734
rect 14188 23316 14240 23322
rect 14188 23258 14240 23264
rect 13912 23112 13964 23118
rect 13912 23054 13964 23060
rect 13728 22092 13780 22098
rect 13728 22034 13780 22040
rect 13924 21690 13952 23054
rect 14188 22432 14240 22438
rect 14188 22374 14240 22380
rect 13912 21684 13964 21690
rect 13912 21626 13964 21632
rect 14004 21548 14056 21554
rect 14004 21490 14056 21496
rect 13728 21072 13780 21078
rect 13728 21014 13780 21020
rect 13636 21004 13688 21010
rect 13636 20946 13688 20952
rect 13648 20602 13676 20946
rect 13636 20596 13688 20602
rect 13740 20584 13768 21014
rect 13740 20556 13860 20584
rect 13636 20538 13688 20544
rect 13556 20420 13768 20448
rect 13544 20256 13596 20262
rect 13544 20198 13596 20204
rect 13556 19786 13584 20198
rect 13634 19816 13690 19825
rect 13544 19780 13596 19786
rect 13634 19751 13690 19760
rect 13544 19722 13596 19728
rect 13556 19446 13584 19722
rect 13544 19440 13596 19446
rect 13544 19382 13596 19388
rect 13452 18760 13504 18766
rect 13452 18702 13504 18708
rect 13452 18624 13504 18630
rect 13452 18566 13504 18572
rect 13464 18358 13492 18566
rect 13648 18426 13676 19751
rect 13544 18420 13596 18426
rect 13544 18362 13596 18368
rect 13636 18420 13688 18426
rect 13636 18362 13688 18368
rect 13452 18352 13504 18358
rect 13452 18294 13504 18300
rect 13360 18216 13412 18222
rect 13360 18158 13412 18164
rect 13268 18148 13320 18154
rect 13268 18090 13320 18096
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 13556 17746 13584 18362
rect 12900 17740 12952 17746
rect 12900 17682 12952 17688
rect 13544 17740 13596 17746
rect 13544 17682 13596 17688
rect 12308 17496 12388 17524
rect 12256 17478 12308 17484
rect 11808 16068 12112 16096
rect 11704 15428 11756 15434
rect 11704 15370 11756 15376
rect 11716 14822 11744 15370
rect 11808 15366 11836 16068
rect 12084 16028 12112 16068
rect 11886 16008 11942 16017
rect 12084 16000 12296 16028
rect 11886 15943 11942 15952
rect 11980 15972 12032 15978
rect 11900 15910 11928 15943
rect 11980 15914 12032 15920
rect 11888 15904 11940 15910
rect 11888 15846 11940 15852
rect 11796 15360 11848 15366
rect 11796 15302 11848 15308
rect 11704 14816 11756 14822
rect 11704 14758 11756 14764
rect 11612 14612 11664 14618
rect 11612 14554 11664 14560
rect 11520 13864 11572 13870
rect 11518 13832 11520 13841
rect 11572 13832 11574 13841
rect 11518 13767 11574 13776
rect 11716 13258 11744 14758
rect 11704 13252 11756 13258
rect 11704 13194 11756 13200
rect 11716 12918 11744 13194
rect 11704 12912 11756 12918
rect 11704 12854 11756 12860
rect 11716 12170 11744 12854
rect 11704 12164 11756 12170
rect 11704 12106 11756 12112
rect 11716 11898 11744 12106
rect 11704 11892 11756 11898
rect 11704 11834 11756 11840
rect 11900 11762 11928 15846
rect 11992 14890 12020 15914
rect 12072 15632 12124 15638
rect 12072 15574 12124 15580
rect 11980 14884 12032 14890
rect 11980 14826 12032 14832
rect 11992 13190 12020 14826
rect 11980 13184 12032 13190
rect 11980 13126 12032 13132
rect 12084 12918 12112 15574
rect 12268 14090 12296 16000
rect 12360 15094 12388 17496
rect 12544 17632 12848 17660
rect 12544 16454 12572 17632
rect 12912 17542 12940 17682
rect 13084 17672 13136 17678
rect 13084 17614 13136 17620
rect 12900 17536 12952 17542
rect 12900 17478 12952 17484
rect 13096 16998 13124 17614
rect 13452 17332 13504 17338
rect 13452 17274 13504 17280
rect 12716 16992 12768 16998
rect 12716 16934 12768 16940
rect 13084 16992 13136 16998
rect 13084 16934 13136 16940
rect 12624 16516 12676 16522
rect 12624 16458 12676 16464
rect 12532 16448 12584 16454
rect 12532 16390 12584 16396
rect 12440 16108 12492 16114
rect 12440 16050 12492 16056
rect 12452 15473 12480 16050
rect 12532 16040 12584 16046
rect 12532 15982 12584 15988
rect 12438 15464 12494 15473
rect 12438 15399 12494 15408
rect 12544 15366 12572 15982
rect 12532 15360 12584 15366
rect 12438 15328 12494 15337
rect 12532 15302 12584 15308
rect 12438 15263 12494 15272
rect 12348 15088 12400 15094
rect 12348 15030 12400 15036
rect 12348 14952 12400 14958
rect 12346 14920 12348 14929
rect 12400 14920 12402 14929
rect 12346 14855 12402 14864
rect 12164 14068 12216 14074
rect 12268 14062 12388 14090
rect 12164 14010 12216 14016
rect 12072 12912 12124 12918
rect 12072 12854 12124 12860
rect 12176 11898 12204 14010
rect 12360 13938 12388 14062
rect 12348 13932 12400 13938
rect 12348 13874 12400 13880
rect 12256 12776 12308 12782
rect 12256 12718 12308 12724
rect 12164 11892 12216 11898
rect 12164 11834 12216 11840
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 12268 11694 12296 12718
rect 12452 12442 12480 15263
rect 12544 14482 12572 15302
rect 12636 14618 12664 16458
rect 12728 15502 12756 16934
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 13360 16584 13412 16590
rect 13360 16526 13412 16532
rect 12992 16448 13044 16454
rect 12992 16390 13044 16396
rect 13004 16182 13032 16390
rect 12992 16176 13044 16182
rect 12992 16118 13044 16124
rect 12900 16040 12952 16046
rect 12900 15982 12952 15988
rect 12912 15892 12940 15982
rect 12820 15864 12940 15892
rect 12820 15570 12848 15864
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 12808 15564 12860 15570
rect 12808 15506 12860 15512
rect 12716 15496 12768 15502
rect 12716 15438 12768 15444
rect 12992 15156 13044 15162
rect 12992 15098 13044 15104
rect 12808 14884 12860 14890
rect 12808 14826 12860 14832
rect 12624 14612 12676 14618
rect 12624 14554 12676 14560
rect 12532 14476 12584 14482
rect 12532 14418 12584 14424
rect 12820 14414 12848 14826
rect 13004 14822 13032 15098
rect 12992 14816 13044 14822
rect 12992 14758 13044 14764
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 13176 14612 13228 14618
rect 13176 14554 13228 14560
rect 12808 14408 12860 14414
rect 12544 14346 12756 14362
rect 12808 14350 12860 14356
rect 13188 14346 13216 14554
rect 13268 14544 13320 14550
rect 13268 14486 13320 14492
rect 13372 14498 13400 16526
rect 13464 15570 13492 17274
rect 13452 15564 13504 15570
rect 13452 15506 13504 15512
rect 13556 15094 13584 17682
rect 13636 17536 13688 17542
rect 13636 17478 13688 17484
rect 13648 17116 13676 17478
rect 13740 17270 13768 20420
rect 13832 20262 13860 20556
rect 13820 20256 13872 20262
rect 13820 20198 13872 20204
rect 13912 19984 13964 19990
rect 13912 19926 13964 19932
rect 13924 19786 13952 19926
rect 13912 19780 13964 19786
rect 13912 19722 13964 19728
rect 14016 17338 14044 21490
rect 14096 19848 14148 19854
rect 14096 19790 14148 19796
rect 14108 19417 14136 19790
rect 14094 19408 14150 19417
rect 14094 19343 14150 19352
rect 14108 18902 14136 19343
rect 14096 18896 14148 18902
rect 14096 18838 14148 18844
rect 14200 18290 14228 22374
rect 14280 21548 14332 21554
rect 14280 21490 14332 21496
rect 14292 20942 14320 21490
rect 14280 20936 14332 20942
rect 14280 20878 14332 20884
rect 14292 19922 14320 20878
rect 14384 20058 14412 24142
rect 14476 23798 14504 26200
rect 14924 24336 14976 24342
rect 14924 24278 14976 24284
rect 14464 23792 14516 23798
rect 14464 23734 14516 23740
rect 14648 22976 14700 22982
rect 14648 22918 14700 22924
rect 14660 22642 14688 22918
rect 14648 22636 14700 22642
rect 14648 22578 14700 22584
rect 14464 22568 14516 22574
rect 14462 22536 14464 22545
rect 14516 22536 14518 22545
rect 14462 22471 14518 22480
rect 14740 21956 14792 21962
rect 14740 21898 14792 21904
rect 14556 20868 14608 20874
rect 14556 20810 14608 20816
rect 14372 20052 14424 20058
rect 14372 19994 14424 20000
rect 14280 19916 14332 19922
rect 14280 19858 14332 19864
rect 14292 18834 14320 19858
rect 14568 19786 14596 20810
rect 14556 19780 14608 19786
rect 14556 19722 14608 19728
rect 14280 18828 14332 18834
rect 14280 18770 14332 18776
rect 14188 18284 14240 18290
rect 14188 18226 14240 18232
rect 14004 17332 14056 17338
rect 14004 17274 14056 17280
rect 13728 17264 13780 17270
rect 13728 17206 13780 17212
rect 13648 17088 13768 17116
rect 13636 16448 13688 16454
rect 13636 16390 13688 16396
rect 13648 15978 13676 16390
rect 13636 15972 13688 15978
rect 13636 15914 13688 15920
rect 13636 15428 13688 15434
rect 13636 15370 13688 15376
rect 13544 15088 13596 15094
rect 13544 15030 13596 15036
rect 12532 14340 12756 14346
rect 12584 14334 12756 14340
rect 12532 14282 12584 14288
rect 12624 14272 12676 14278
rect 12624 14214 12676 14220
rect 12532 13796 12584 13802
rect 12532 13738 12584 13744
rect 12544 13462 12572 13738
rect 12532 13456 12584 13462
rect 12532 13398 12584 13404
rect 12636 13002 12664 14214
rect 12728 13190 12756 14334
rect 13176 14340 13228 14346
rect 13176 14282 13228 14288
rect 12808 13864 12860 13870
rect 13280 13852 13308 14486
rect 13372 14470 13584 14498
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 13360 13864 13412 13870
rect 13280 13824 13360 13852
rect 12808 13806 12860 13812
rect 13360 13806 13412 13812
rect 12820 13326 12848 13806
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 12808 13320 12860 13326
rect 12808 13262 12860 13268
rect 13084 13320 13136 13326
rect 13084 13262 13136 13268
rect 12716 13184 12768 13190
rect 12716 13126 12768 13132
rect 12636 12974 12848 13002
rect 12532 12844 12584 12850
rect 12532 12786 12584 12792
rect 12716 12844 12768 12850
rect 12716 12786 12768 12792
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 12544 12170 12572 12786
rect 12624 12640 12676 12646
rect 12624 12582 12676 12588
rect 12532 12164 12584 12170
rect 12452 12124 12532 12152
rect 12256 11688 12308 11694
rect 12256 11630 12308 11636
rect 11796 11620 11848 11626
rect 11796 11562 11848 11568
rect 11336 8968 11388 8974
rect 11336 8910 11388 8916
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 6920 8288 6972 8294
rect 6920 8230 6972 8236
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 2412 7880 2464 7886
rect 2412 7822 2464 7828
rect 2320 6656 2372 6662
rect 2320 6598 2372 6604
rect 1306 6488 1362 6497
rect 1216 6452 1268 6458
rect 1306 6423 1362 6432
rect 1216 6394 1268 6400
rect 1308 6316 1360 6322
rect 1308 6258 1360 6264
rect 1320 6089 1348 6258
rect 1306 6080 1362 6089
rect 1306 6015 1362 6024
rect 1308 5704 1360 5710
rect 1306 5672 1308 5681
rect 1360 5672 1362 5681
rect 1306 5607 1362 5616
rect 1308 5160 1360 5166
rect 1308 5102 1360 5108
rect 1320 4865 1348 5102
rect 1860 5024 1912 5030
rect 1860 4966 1912 4972
rect 1306 4856 1362 4865
rect 1306 4791 1308 4800
rect 1360 4791 1362 4800
rect 1308 4762 1360 4768
rect 1308 4616 1360 4622
rect 1308 4558 1360 4564
rect 1320 4457 1348 4558
rect 1306 4448 1362 4457
rect 1306 4383 1362 4392
rect 1400 4208 1452 4214
rect 1400 4150 1452 4156
rect 1308 4140 1360 4146
rect 1308 4082 1360 4088
rect 1320 3641 1348 4082
rect 1412 4049 1440 4150
rect 1398 4040 1454 4049
rect 1398 3975 1454 3984
rect 1306 3632 1362 3641
rect 1872 3602 1900 4966
rect 1306 3567 1362 3576
rect 1860 3596 1912 3602
rect 1860 3538 1912 3544
rect 1308 3528 1360 3534
rect 1122 3496 1178 3505
rect 1308 3470 1360 3476
rect 1122 3431 1178 3440
rect 1136 800 1164 3431
rect 1320 3233 1348 3470
rect 1306 3224 1362 3233
rect 1306 3159 1308 3168
rect 1360 3159 1362 3168
rect 1308 3130 1360 3136
rect 1308 3052 1360 3058
rect 1308 2994 1360 3000
rect 1320 2825 1348 2994
rect 2424 2922 2452 7822
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 6932 5914 6960 8230
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 2780 5704 2832 5710
rect 2780 5646 2832 5652
rect 2792 5273 2820 5646
rect 2778 5264 2834 5273
rect 2778 5199 2834 5208
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 2950 4859 3258 4868
rect 2504 4140 2556 4146
rect 2504 4082 2556 4088
rect 2516 3924 2544 4082
rect 5354 4040 5410 4049
rect 5354 3975 5410 3984
rect 2688 3936 2740 3942
rect 2516 3896 2688 3924
rect 2688 3878 2740 3884
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 3332 3528 3384 3534
rect 3332 3470 3384 3476
rect 2412 2916 2464 2922
rect 2412 2858 2464 2864
rect 2320 2848 2372 2854
rect 1306 2816 1362 2825
rect 2320 2790 2372 2796
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 1306 2751 1362 2760
rect 1308 2440 1360 2446
rect 1306 2408 1308 2417
rect 1360 2408 1362 2417
rect 1216 2372 1268 2378
rect 2332 2378 2360 2790
rect 2792 2446 2820 2790
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 1306 2343 1362 2352
rect 2320 2372 2372 2378
rect 1216 2314 1268 2320
rect 2320 2314 2372 2320
rect 1228 2009 1256 2314
rect 1308 2304 1360 2310
rect 1308 2246 1360 2252
rect 1214 2000 1270 2009
rect 1214 1935 1270 1944
rect 1320 1601 1348 2246
rect 3344 1850 3372 3470
rect 4344 2576 4396 2582
rect 4344 2518 4396 2524
rect 4356 2378 4384 2518
rect 4344 2372 4396 2378
rect 4344 2314 4396 2320
rect 3252 1822 3372 1850
rect 1306 1592 1362 1601
rect 1306 1527 1362 1536
rect 3252 800 3280 1822
rect 5368 800 5396 3975
rect 7852 3942 7880 6054
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 11808 5166 11836 11562
rect 12452 11354 12480 12124
rect 12532 12106 12584 12112
rect 12532 11552 12584 11558
rect 12532 11494 12584 11500
rect 12440 11348 12492 11354
rect 12360 11308 12440 11336
rect 12360 11150 12388 11308
rect 12440 11290 12492 11296
rect 12348 11144 12400 11150
rect 12348 11086 12400 11092
rect 12360 10810 12388 11086
rect 12348 10804 12400 10810
rect 12348 10746 12400 10752
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 11796 5160 11848 5166
rect 11796 5102 11848 5108
rect 12452 5030 12480 9862
rect 12544 9654 12572 11494
rect 12636 9654 12664 12582
rect 12728 12306 12756 12786
rect 12716 12300 12768 12306
rect 12716 12242 12768 12248
rect 12716 12096 12768 12102
rect 12716 12038 12768 12044
rect 12728 11286 12756 12038
rect 12716 11280 12768 11286
rect 12716 11222 12768 11228
rect 12728 9654 12756 11222
rect 12820 10810 12848 12974
rect 13096 12850 13124 13262
rect 13372 12986 13400 13806
rect 13360 12980 13412 12986
rect 13360 12922 13412 12928
rect 13084 12844 13136 12850
rect 13084 12786 13136 12792
rect 13360 12776 13412 12782
rect 13360 12718 13412 12724
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 13268 12436 13320 12442
rect 13268 12378 13320 12384
rect 13280 11898 13308 12378
rect 13268 11892 13320 11898
rect 13268 11834 13320 11840
rect 13372 11529 13400 12718
rect 13358 11520 13414 11529
rect 12950 11452 13258 11461
rect 13358 11455 13414 11464
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 13464 11354 13492 14214
rect 13556 11393 13584 14470
rect 13648 11898 13676 15370
rect 13740 14278 13768 17088
rect 13912 16652 13964 16658
rect 13912 16594 13964 16600
rect 13924 14958 13952 16594
rect 14200 16590 14228 18226
rect 14648 17604 14700 17610
rect 14648 17546 14700 17552
rect 14278 17368 14334 17377
rect 14278 17303 14334 17312
rect 14292 17270 14320 17303
rect 14280 17264 14332 17270
rect 14280 17206 14332 17212
rect 14372 17196 14424 17202
rect 14372 17138 14424 17144
rect 14280 16788 14332 16794
rect 14280 16730 14332 16736
rect 14188 16584 14240 16590
rect 14188 16526 14240 16532
rect 14292 16153 14320 16730
rect 14278 16144 14334 16153
rect 14278 16079 14334 16088
rect 14004 15088 14056 15094
rect 14384 15065 14412 17138
rect 14554 16552 14610 16561
rect 14554 16487 14610 16496
rect 14568 16250 14596 16487
rect 14556 16244 14608 16250
rect 14556 16186 14608 16192
rect 14556 16040 14608 16046
rect 14556 15982 14608 15988
rect 14464 15360 14516 15366
rect 14464 15302 14516 15308
rect 14004 15030 14056 15036
rect 14370 15056 14426 15065
rect 13912 14952 13964 14958
rect 13912 14894 13964 14900
rect 13728 14272 13780 14278
rect 13728 14214 13780 14220
rect 13924 14090 13952 14894
rect 13740 14062 13952 14090
rect 13740 12170 13768 14062
rect 14016 14006 14044 15030
rect 14370 14991 14426 15000
rect 14476 14550 14504 15302
rect 14568 15162 14596 15982
rect 14660 15609 14688 17546
rect 14752 16794 14780 21898
rect 14832 21616 14884 21622
rect 14832 21558 14884 21564
rect 14844 20806 14872 21558
rect 14832 20800 14884 20806
rect 14832 20742 14884 20748
rect 14844 20398 14872 20742
rect 14936 20602 14964 24278
rect 15120 22574 15148 26200
rect 15384 23520 15436 23526
rect 15384 23462 15436 23468
rect 15292 22704 15344 22710
rect 15292 22646 15344 22652
rect 15108 22568 15160 22574
rect 15108 22510 15160 22516
rect 15200 22024 15252 22030
rect 15200 21966 15252 21972
rect 14924 20596 14976 20602
rect 14924 20538 14976 20544
rect 15108 20596 15160 20602
rect 15108 20538 15160 20544
rect 14924 20460 14976 20466
rect 14924 20402 14976 20408
rect 14832 20392 14884 20398
rect 14832 20334 14884 20340
rect 14936 20058 14964 20402
rect 14924 20052 14976 20058
rect 14924 19994 14976 20000
rect 15016 19780 15068 19786
rect 15120 19768 15148 20538
rect 15068 19740 15148 19768
rect 15016 19722 15068 19728
rect 15028 19514 15056 19722
rect 15016 19508 15068 19514
rect 15016 19450 15068 19456
rect 15106 19408 15162 19417
rect 15106 19343 15162 19352
rect 15120 18970 15148 19343
rect 15108 18964 15160 18970
rect 15108 18906 15160 18912
rect 15016 18420 15068 18426
rect 15016 18362 15068 18368
rect 15028 18329 15056 18362
rect 15014 18320 15070 18329
rect 14844 18278 15014 18306
rect 14740 16788 14792 16794
rect 14740 16730 14792 16736
rect 14844 16454 14872 18278
rect 15014 18255 15070 18264
rect 14922 18184 14978 18193
rect 14922 18119 14978 18128
rect 14740 16448 14792 16454
rect 14740 16390 14792 16396
rect 14832 16448 14884 16454
rect 14832 16390 14884 16396
rect 14646 15600 14702 15609
rect 14646 15535 14702 15544
rect 14556 15156 14608 15162
rect 14556 15098 14608 15104
rect 14464 14544 14516 14550
rect 14464 14486 14516 14492
rect 14188 14408 14240 14414
rect 14186 14376 14188 14385
rect 14240 14376 14242 14385
rect 14186 14311 14242 14320
rect 14004 14000 14056 14006
rect 14004 13942 14056 13948
rect 14568 13954 14596 15098
rect 14660 14074 14688 15535
rect 14648 14068 14700 14074
rect 14648 14010 14700 14016
rect 14016 13870 14044 13942
rect 14568 13926 14688 13954
rect 14004 13864 14056 13870
rect 14004 13806 14056 13812
rect 14554 13696 14610 13705
rect 14554 13631 14610 13640
rect 14278 13560 14334 13569
rect 14278 13495 14334 13504
rect 14016 13246 14228 13274
rect 13728 12164 13780 12170
rect 13728 12106 13780 12112
rect 13636 11892 13688 11898
rect 13636 11834 13688 11840
rect 13542 11384 13598 11393
rect 13452 11348 13504 11354
rect 13542 11319 13598 11328
rect 13452 11290 13504 11296
rect 13820 11212 13872 11218
rect 13820 11154 13872 11160
rect 12900 11144 12952 11150
rect 12900 11086 12952 11092
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 12912 10690 12940 11086
rect 12820 10662 12940 10690
rect 13634 10704 13690 10713
rect 13544 10668 13596 10674
rect 12532 9648 12584 9654
rect 12532 9590 12584 9596
rect 12624 9648 12676 9654
rect 12624 9590 12676 9596
rect 12716 9648 12768 9654
rect 12716 9590 12768 9596
rect 12820 9466 12848 10662
rect 13634 10639 13636 10648
rect 13544 10610 13596 10616
rect 13688 10639 13690 10648
rect 13636 10610 13688 10616
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 13082 10160 13138 10169
rect 13082 10095 13138 10104
rect 13096 9926 13124 10095
rect 13084 9920 13136 9926
rect 13084 9862 13136 9868
rect 12728 9438 12848 9466
rect 12440 5024 12492 5030
rect 12440 4966 12492 4972
rect 11704 4752 11756 4758
rect 11704 4694 11756 4700
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 7840 3936 7892 3942
rect 7840 3878 7892 3884
rect 7472 3596 7524 3602
rect 7472 3538 7524 3544
rect 7484 800 7512 3538
rect 11716 3534 11744 4694
rect 11704 3528 11756 3534
rect 11704 3470 11756 3476
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 11060 2984 11112 2990
rect 11060 2926 11112 2932
rect 11072 2650 11100 2926
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 11704 2508 11756 2514
rect 11704 2450 11756 2456
rect 9680 2440 9732 2446
rect 9600 2388 9680 2394
rect 9600 2382 9732 2388
rect 9600 2366 9720 2382
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 9600 800 9628 2366
rect 11716 800 11744 2450
rect 12728 2310 12756 9438
rect 12808 9376 12860 9382
rect 12808 9318 12860 9324
rect 12820 7886 12848 9318
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 12808 7880 12860 7886
rect 12808 7822 12860 7828
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 12808 3392 12860 3398
rect 12808 3334 12860 3340
rect 12820 2446 12848 3334
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 13556 2650 13584 10610
rect 13832 10062 13860 11154
rect 14016 11014 14044 13246
rect 14200 13190 14228 13246
rect 14096 13184 14148 13190
rect 14096 13126 14148 13132
rect 14188 13184 14240 13190
rect 14188 13126 14240 13132
rect 14108 12782 14136 13126
rect 14096 12776 14148 12782
rect 14096 12718 14148 12724
rect 14004 11008 14056 11014
rect 14004 10950 14056 10956
rect 13912 10668 13964 10674
rect 13912 10610 13964 10616
rect 13924 10198 13952 10610
rect 13912 10192 13964 10198
rect 13912 10134 13964 10140
rect 13820 10056 13872 10062
rect 13820 9998 13872 10004
rect 13924 10010 13952 10134
rect 13636 9512 13688 9518
rect 13636 9454 13688 9460
rect 13648 9042 13676 9454
rect 13832 9382 13860 9998
rect 13924 9982 14044 10010
rect 13912 9920 13964 9926
rect 13912 9862 13964 9868
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 13832 9110 13860 9318
rect 13820 9104 13872 9110
rect 13820 9046 13872 9052
rect 13636 9036 13688 9042
rect 13636 8978 13688 8984
rect 13832 8566 13860 9046
rect 13924 8566 13952 9862
rect 13820 8560 13872 8566
rect 13820 8502 13872 8508
rect 13912 8560 13964 8566
rect 13912 8502 13964 8508
rect 13832 3058 13860 8502
rect 14016 7954 14044 9982
rect 14004 7948 14056 7954
rect 14004 7890 14056 7896
rect 14108 6186 14136 12718
rect 14188 11824 14240 11830
rect 14188 11766 14240 11772
rect 14200 10810 14228 11766
rect 14188 10804 14240 10810
rect 14188 10746 14240 10752
rect 14292 10470 14320 13495
rect 14464 11620 14516 11626
rect 14464 11562 14516 11568
rect 14370 11520 14426 11529
rect 14370 11455 14426 11464
rect 14384 10606 14412 11455
rect 14372 10600 14424 10606
rect 14372 10542 14424 10548
rect 14280 10464 14332 10470
rect 14280 10406 14332 10412
rect 14476 9926 14504 11562
rect 14568 10742 14596 13631
rect 14660 11286 14688 13926
rect 14752 13394 14780 16390
rect 14936 16250 14964 18119
rect 15016 17876 15068 17882
rect 15016 17818 15068 17824
rect 15028 17270 15056 17818
rect 15120 17610 15148 18906
rect 15212 17746 15240 21966
rect 15304 19310 15332 22646
rect 15396 20602 15424 23462
rect 15764 23186 15792 26200
rect 16028 24744 16080 24750
rect 16028 24686 16080 24692
rect 15844 23248 15896 23254
rect 15844 23190 15896 23196
rect 15752 23180 15804 23186
rect 15752 23122 15804 23128
rect 15856 20602 15884 23190
rect 16040 20602 16068 24686
rect 16132 23798 16160 26302
rect 16394 26200 16450 26302
rect 17038 26330 17094 27000
rect 17038 26302 17264 26330
rect 17038 26200 17094 26302
rect 17040 24608 17092 24614
rect 17040 24550 17092 24556
rect 17052 23866 17080 24550
rect 17040 23860 17092 23866
rect 17040 23802 17092 23808
rect 16120 23792 16172 23798
rect 16120 23734 16172 23740
rect 17040 23112 17092 23118
rect 17040 23054 17092 23060
rect 17052 22710 17080 23054
rect 17040 22704 17092 22710
rect 17040 22646 17092 22652
rect 16672 22636 16724 22642
rect 16672 22578 16724 22584
rect 16120 22094 16172 22098
rect 16120 22092 16344 22094
rect 16172 22066 16344 22092
rect 16488 22092 16540 22098
rect 16120 22034 16172 22040
rect 16210 21992 16266 22001
rect 16210 21927 16266 21936
rect 16120 21480 16172 21486
rect 16120 21422 16172 21428
rect 15384 20596 15436 20602
rect 15384 20538 15436 20544
rect 15844 20596 15896 20602
rect 15844 20538 15896 20544
rect 16028 20596 16080 20602
rect 16028 20538 16080 20544
rect 15936 20460 15988 20466
rect 15936 20402 15988 20408
rect 15476 20392 15528 20398
rect 15476 20334 15528 20340
rect 15382 19408 15438 19417
rect 15382 19343 15384 19352
rect 15436 19343 15438 19352
rect 15384 19314 15436 19320
rect 15292 19304 15344 19310
rect 15292 19246 15344 19252
rect 15292 18828 15344 18834
rect 15292 18770 15344 18776
rect 15304 18222 15332 18770
rect 15292 18216 15344 18222
rect 15292 18158 15344 18164
rect 15382 18184 15438 18193
rect 15304 17882 15332 18158
rect 15382 18119 15384 18128
rect 15436 18119 15438 18128
rect 15384 18090 15436 18096
rect 15292 17876 15344 17882
rect 15292 17818 15344 17824
rect 15200 17740 15252 17746
rect 15200 17682 15252 17688
rect 15108 17604 15160 17610
rect 15108 17546 15160 17552
rect 15396 17377 15424 18090
rect 15382 17368 15438 17377
rect 15382 17303 15438 17312
rect 15016 17264 15068 17270
rect 15016 17206 15068 17212
rect 15108 17196 15160 17202
rect 15108 17138 15160 17144
rect 15016 16516 15068 16522
rect 15016 16458 15068 16464
rect 14924 16244 14976 16250
rect 14924 16186 14976 16192
rect 15028 16046 15056 16458
rect 14832 16040 14884 16046
rect 14830 16008 14832 16017
rect 15016 16040 15068 16046
rect 14884 16008 14886 16017
rect 15016 15982 15068 15988
rect 14830 15943 14886 15952
rect 14844 15706 14872 15943
rect 14832 15700 14884 15706
rect 14832 15642 14884 15648
rect 14832 15564 14884 15570
rect 14832 15506 14884 15512
rect 14844 13462 14872 15506
rect 15028 15178 15056 15982
rect 14936 15150 15056 15178
rect 14936 14550 14964 15150
rect 15014 15056 15070 15065
rect 15014 14991 15070 15000
rect 14924 14544 14976 14550
rect 14924 14486 14976 14492
rect 14924 13864 14976 13870
rect 14924 13806 14976 13812
rect 14936 13530 14964 13806
rect 14924 13524 14976 13530
rect 14924 13466 14976 13472
rect 14832 13456 14884 13462
rect 15028 13410 15056 14991
rect 15120 14804 15148 17138
rect 15200 16720 15252 16726
rect 15200 16662 15252 16668
rect 15212 16046 15240 16662
rect 15488 16522 15516 20334
rect 15752 20256 15804 20262
rect 15752 20198 15804 20204
rect 15568 19916 15620 19922
rect 15620 19876 15700 19904
rect 15568 19858 15620 19864
rect 15568 18624 15620 18630
rect 15568 18566 15620 18572
rect 15580 17338 15608 18566
rect 15568 17332 15620 17338
rect 15568 17274 15620 17280
rect 15672 16561 15700 19876
rect 15764 19310 15792 20198
rect 15752 19304 15804 19310
rect 15752 19246 15804 19252
rect 15948 18902 15976 20402
rect 16028 19236 16080 19242
rect 16028 19178 16080 19184
rect 16040 18970 16068 19178
rect 16028 18964 16080 18970
rect 16028 18906 16080 18912
rect 15936 18896 15988 18902
rect 15936 18838 15988 18844
rect 15752 17196 15804 17202
rect 15752 17138 15804 17144
rect 15658 16552 15714 16561
rect 15476 16516 15528 16522
rect 15658 16487 15714 16496
rect 15476 16458 15528 16464
rect 15660 16448 15712 16454
rect 15660 16390 15712 16396
rect 15200 16040 15252 16046
rect 15200 15982 15252 15988
rect 15476 15632 15528 15638
rect 15476 15574 15528 15580
rect 15384 15564 15436 15570
rect 15384 15506 15436 15512
rect 15120 14776 15332 14804
rect 15200 14068 15252 14074
rect 15200 14010 15252 14016
rect 15108 13524 15160 13530
rect 15108 13466 15160 13472
rect 14832 13398 14884 13404
rect 14740 13388 14792 13394
rect 14740 13330 14792 13336
rect 14740 12096 14792 12102
rect 14740 12038 14792 12044
rect 14752 11694 14780 12038
rect 14740 11688 14792 11694
rect 14740 11630 14792 11636
rect 14844 11642 14872 13398
rect 14936 13382 15056 13410
rect 14936 12306 14964 13382
rect 15120 13308 15148 13466
rect 15028 13280 15148 13308
rect 14924 12300 14976 12306
rect 14924 12242 14976 12248
rect 15028 12170 15056 13280
rect 15108 12912 15160 12918
rect 15108 12854 15160 12860
rect 15016 12164 15068 12170
rect 15016 12106 15068 12112
rect 15014 11792 15070 11801
rect 15014 11727 15070 11736
rect 14844 11614 14964 11642
rect 14832 11552 14884 11558
rect 14832 11494 14884 11500
rect 14648 11280 14700 11286
rect 14648 11222 14700 11228
rect 14844 11218 14872 11494
rect 14832 11212 14884 11218
rect 14832 11154 14884 11160
rect 14740 11144 14792 11150
rect 14738 11112 14740 11121
rect 14792 11112 14794 11121
rect 14738 11047 14794 11056
rect 14556 10736 14608 10742
rect 14556 10678 14608 10684
rect 14936 10606 14964 11614
rect 14924 10600 14976 10606
rect 14924 10542 14976 10548
rect 15028 10538 15056 11727
rect 15016 10532 15068 10538
rect 15016 10474 15068 10480
rect 14832 9988 14884 9994
rect 15028 9976 15056 10474
rect 14884 9948 15056 9976
rect 14832 9930 14884 9936
rect 14464 9920 14516 9926
rect 14464 9862 14516 9868
rect 14188 9512 14240 9518
rect 14188 9454 14240 9460
rect 14200 9178 14228 9454
rect 14924 9444 14976 9450
rect 14924 9386 14976 9392
rect 14188 9172 14240 9178
rect 14188 9114 14240 9120
rect 14186 9072 14242 9081
rect 14186 9007 14242 9016
rect 14200 7818 14228 9007
rect 14188 7812 14240 7818
rect 14188 7754 14240 7760
rect 14096 6180 14148 6186
rect 14096 6122 14148 6128
rect 14936 4078 14964 9386
rect 15120 8906 15148 12854
rect 15212 11830 15240 14010
rect 15304 12434 15332 14776
rect 15396 14260 15424 15506
rect 15488 15366 15516 15574
rect 15566 15464 15622 15473
rect 15566 15399 15622 15408
rect 15476 15360 15528 15366
rect 15476 15302 15528 15308
rect 15580 15162 15608 15399
rect 15568 15156 15620 15162
rect 15568 15098 15620 15104
rect 15672 15094 15700 16390
rect 15660 15088 15712 15094
rect 15660 15030 15712 15036
rect 15764 14940 15792 17138
rect 16040 17134 16068 18906
rect 16132 18154 16160 21422
rect 16224 20398 16252 21927
rect 16316 21350 16344 22066
rect 16408 22052 16488 22080
rect 16304 21344 16356 21350
rect 16304 21286 16356 21292
rect 16212 20392 16264 20398
rect 16212 20334 16264 20340
rect 16212 19168 16264 19174
rect 16212 19110 16264 19116
rect 16224 18737 16252 19110
rect 16316 18834 16344 21286
rect 16408 19718 16436 22052
rect 16488 22034 16540 22040
rect 16488 21888 16540 21894
rect 16488 21830 16540 21836
rect 16396 19712 16448 19718
rect 16396 19654 16448 19660
rect 16500 18970 16528 21830
rect 16684 21593 16712 22578
rect 16764 22568 16816 22574
rect 16764 22510 16816 22516
rect 16776 22234 16804 22510
rect 17052 22234 17080 22646
rect 16764 22228 16816 22234
rect 16764 22170 16816 22176
rect 17040 22228 17092 22234
rect 17040 22170 17092 22176
rect 16764 21956 16816 21962
rect 16764 21898 16816 21904
rect 16776 21622 16804 21898
rect 17052 21690 17080 22170
rect 17236 22166 17264 26302
rect 17682 26200 17738 27000
rect 18326 26200 18382 27000
rect 18970 26200 19026 27000
rect 19614 26200 19670 27000
rect 20258 26330 20314 27000
rect 20258 26302 20576 26330
rect 20258 26200 20314 26302
rect 17696 24274 17724 26200
rect 17868 24676 17920 24682
rect 17868 24618 17920 24624
rect 17684 24268 17736 24274
rect 17684 24210 17736 24216
rect 17316 23044 17368 23050
rect 17316 22986 17368 22992
rect 17408 23044 17460 23050
rect 17408 22986 17460 22992
rect 17224 22160 17276 22166
rect 17224 22102 17276 22108
rect 17040 21684 17092 21690
rect 17040 21626 17092 21632
rect 16764 21616 16816 21622
rect 16670 21584 16726 21593
rect 16764 21558 16816 21564
rect 16670 21519 16726 21528
rect 16578 21176 16634 21185
rect 16578 21111 16580 21120
rect 16632 21111 16634 21120
rect 16580 21082 16632 21088
rect 16776 20874 16804 21558
rect 17052 20942 17080 21626
rect 17130 21176 17186 21185
rect 17130 21111 17186 21120
rect 17040 20936 17092 20942
rect 17040 20878 17092 20884
rect 16764 20868 16816 20874
rect 16684 20828 16764 20856
rect 16488 18964 16540 18970
rect 16488 18906 16540 18912
rect 16304 18828 16356 18834
rect 16304 18770 16356 18776
rect 16684 18766 16712 20828
rect 16764 20810 16816 20816
rect 17052 20398 17080 20878
rect 16764 20392 16816 20398
rect 16762 20360 16764 20369
rect 17040 20392 17092 20398
rect 16816 20360 16818 20369
rect 17040 20334 17092 20340
rect 16762 20295 16818 20304
rect 16856 20324 16908 20330
rect 16776 19446 16804 20295
rect 16856 20266 16908 20272
rect 16868 19514 16896 20266
rect 17040 19780 17092 19786
rect 17040 19722 17092 19728
rect 16856 19508 16908 19514
rect 16856 19450 16908 19456
rect 16764 19440 16816 19446
rect 16764 19382 16816 19388
rect 16764 19304 16816 19310
rect 16764 19246 16816 19252
rect 16672 18760 16724 18766
rect 16210 18728 16266 18737
rect 16672 18702 16724 18708
rect 16210 18663 16266 18672
rect 16684 18358 16712 18702
rect 16776 18630 16804 19246
rect 17052 18970 17080 19722
rect 17040 18964 17092 18970
rect 17040 18906 17092 18912
rect 16948 18692 17000 18698
rect 16948 18634 17000 18640
rect 16764 18624 16816 18630
rect 16764 18566 16816 18572
rect 16672 18352 16724 18358
rect 16672 18294 16724 18300
rect 16212 18216 16264 18222
rect 16212 18158 16264 18164
rect 16120 18148 16172 18154
rect 16120 18090 16172 18096
rect 16120 17808 16172 17814
rect 16120 17750 16172 17756
rect 16132 17338 16160 17750
rect 16224 17678 16252 18158
rect 16580 18080 16632 18086
rect 16580 18022 16632 18028
rect 16304 17740 16356 17746
rect 16304 17682 16356 17688
rect 16212 17672 16264 17678
rect 16212 17614 16264 17620
rect 16120 17332 16172 17338
rect 16120 17274 16172 17280
rect 16028 17128 16080 17134
rect 16028 17070 16080 17076
rect 15934 16688 15990 16697
rect 15934 16623 15990 16632
rect 16118 16688 16174 16697
rect 16316 16658 16344 17682
rect 16488 17332 16540 17338
rect 16488 17274 16540 17280
rect 16118 16623 16120 16632
rect 15948 16182 15976 16623
rect 16172 16623 16174 16632
rect 16304 16652 16356 16658
rect 16120 16594 16172 16600
rect 16304 16594 16356 16600
rect 16500 16590 16528 17274
rect 16488 16584 16540 16590
rect 16488 16526 16540 16532
rect 15936 16176 15988 16182
rect 15936 16118 15988 16124
rect 15844 16040 15896 16046
rect 15842 16008 15844 16017
rect 15936 16040 15988 16046
rect 15896 16008 15898 16017
rect 15936 15982 15988 15988
rect 15842 15943 15898 15952
rect 15856 15910 15884 15943
rect 15844 15904 15896 15910
rect 15844 15846 15896 15852
rect 15948 15638 15976 15982
rect 16488 15972 16540 15978
rect 16488 15914 16540 15920
rect 15936 15632 15988 15638
rect 15936 15574 15988 15580
rect 16500 15570 16528 15914
rect 16592 15706 16620 18022
rect 16672 15904 16724 15910
rect 16672 15846 16724 15852
rect 16776 15892 16804 18566
rect 16960 16726 16988 18634
rect 17040 17128 17092 17134
rect 17040 17070 17092 17076
rect 16948 16720 17000 16726
rect 16948 16662 17000 16668
rect 17052 16114 17080 17070
rect 17144 16266 17172 21111
rect 17224 19712 17276 19718
rect 17224 19654 17276 19660
rect 17236 17882 17264 19654
rect 17328 17882 17356 22986
rect 17420 22778 17448 22986
rect 17500 22976 17552 22982
rect 17500 22918 17552 22924
rect 17408 22772 17460 22778
rect 17408 22714 17460 22720
rect 17408 19848 17460 19854
rect 17408 19790 17460 19796
rect 17420 19310 17448 19790
rect 17512 19718 17540 22918
rect 17684 22024 17736 22030
rect 17684 21966 17736 21972
rect 17696 21690 17724 21966
rect 17880 21690 17908 24618
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 18340 23798 18368 26200
rect 18420 24132 18472 24138
rect 18420 24074 18472 24080
rect 18328 23792 18380 23798
rect 18328 23734 18380 23740
rect 17960 23656 18012 23662
rect 17960 23598 18012 23604
rect 17972 23322 18000 23598
rect 17960 23316 18012 23322
rect 17960 23258 18012 23264
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 18236 22636 18288 22642
rect 18236 22578 18288 22584
rect 18248 22030 18276 22578
rect 18432 22137 18460 24074
rect 18512 24064 18564 24070
rect 18512 24006 18564 24012
rect 18418 22128 18474 22137
rect 18418 22063 18474 22072
rect 18236 22024 18288 22030
rect 18236 21966 18288 21972
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 17684 21684 17736 21690
rect 17684 21626 17736 21632
rect 17868 21684 17920 21690
rect 17868 21626 17920 21632
rect 18328 21548 18380 21554
rect 18328 21490 18380 21496
rect 17776 20800 17828 20806
rect 17776 20742 17828 20748
rect 17684 20392 17736 20398
rect 17684 20334 17736 20340
rect 17500 19712 17552 19718
rect 17500 19654 17552 19660
rect 17408 19304 17460 19310
rect 17408 19246 17460 19252
rect 17696 18902 17724 20334
rect 17684 18896 17736 18902
rect 17684 18838 17736 18844
rect 17408 18760 17460 18766
rect 17406 18728 17408 18737
rect 17460 18728 17462 18737
rect 17406 18663 17462 18672
rect 17224 17876 17276 17882
rect 17224 17818 17276 17824
rect 17316 17876 17368 17882
rect 17316 17818 17368 17824
rect 17696 17746 17724 18838
rect 17788 18766 17816 20742
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 18052 20392 18104 20398
rect 18052 20334 18104 20340
rect 18064 20058 18092 20334
rect 18340 20058 18368 21490
rect 18052 20052 18104 20058
rect 18052 19994 18104 20000
rect 18328 20052 18380 20058
rect 18328 19994 18380 20000
rect 18524 19854 18552 24006
rect 18880 22976 18932 22982
rect 18880 22918 18932 22924
rect 18788 22704 18840 22710
rect 18788 22646 18840 22652
rect 18604 22568 18656 22574
rect 18604 22510 18656 22516
rect 18616 22234 18644 22510
rect 18696 22500 18748 22506
rect 18696 22442 18748 22448
rect 18708 22234 18736 22442
rect 18604 22228 18656 22234
rect 18604 22170 18656 22176
rect 18696 22228 18748 22234
rect 18696 22170 18748 22176
rect 18616 21486 18644 22170
rect 18694 22128 18750 22137
rect 18694 22063 18750 22072
rect 18604 21480 18656 21486
rect 18604 21422 18656 21428
rect 18512 19848 18564 19854
rect 18512 19790 18564 19796
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 18616 19446 18644 21422
rect 18708 21350 18736 22063
rect 18696 21344 18748 21350
rect 18696 21286 18748 21292
rect 18800 20806 18828 22646
rect 18892 22001 18920 22918
rect 18984 22166 19012 26200
rect 19628 24342 19656 26200
rect 19616 24336 19668 24342
rect 19616 24278 19668 24284
rect 20548 24206 20576 26302
rect 20902 26200 20958 27000
rect 21546 26200 21602 27000
rect 22190 26200 22246 27000
rect 22834 26200 22890 27000
rect 23478 26330 23534 27000
rect 23478 26302 23980 26330
rect 23478 26200 23534 26302
rect 20720 24404 20772 24410
rect 20720 24346 20772 24352
rect 19340 24200 19392 24206
rect 19340 24142 19392 24148
rect 20536 24200 20588 24206
rect 20536 24142 20588 24148
rect 19352 24041 19380 24142
rect 20444 24132 20496 24138
rect 20444 24074 20496 24080
rect 19432 24064 19484 24070
rect 19338 24032 19394 24041
rect 19432 24006 19484 24012
rect 19338 23967 19394 23976
rect 19064 23656 19116 23662
rect 19064 23598 19116 23604
rect 18972 22160 19024 22166
rect 18972 22102 19024 22108
rect 18878 21992 18934 22001
rect 18878 21927 18934 21936
rect 18880 21480 18932 21486
rect 18880 21422 18932 21428
rect 18788 20800 18840 20806
rect 18788 20742 18840 20748
rect 18800 20398 18828 20742
rect 18892 20602 18920 21422
rect 18972 21140 19024 21146
rect 18972 21082 19024 21088
rect 18880 20596 18932 20602
rect 18880 20538 18932 20544
rect 18788 20392 18840 20398
rect 18788 20334 18840 20340
rect 18788 20256 18840 20262
rect 18788 20198 18840 20204
rect 18604 19440 18656 19446
rect 18604 19382 18656 19388
rect 18696 18828 18748 18834
rect 18696 18770 18748 18776
rect 17776 18760 17828 18766
rect 17776 18702 17828 18708
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 17776 18216 17828 18222
rect 17776 18158 17828 18164
rect 17684 17740 17736 17746
rect 17684 17682 17736 17688
rect 17500 17536 17552 17542
rect 17500 17478 17552 17484
rect 17512 16998 17540 17478
rect 17408 16992 17460 16998
rect 17500 16992 17552 16998
rect 17408 16934 17460 16940
rect 17498 16960 17500 16969
rect 17552 16960 17554 16969
rect 17224 16788 17276 16794
rect 17224 16730 17276 16736
rect 17236 16454 17264 16730
rect 17224 16448 17276 16454
rect 17224 16390 17276 16396
rect 17144 16238 17264 16266
rect 17040 16108 17092 16114
rect 17040 16050 17092 16056
rect 16948 15972 17000 15978
rect 16948 15914 17000 15920
rect 16856 15904 16908 15910
rect 16776 15864 16856 15892
rect 16580 15700 16632 15706
rect 16580 15642 16632 15648
rect 16488 15564 16540 15570
rect 16488 15506 16540 15512
rect 15844 15496 15896 15502
rect 15896 15456 16252 15484
rect 15844 15438 15896 15444
rect 16028 15360 16080 15366
rect 16028 15302 16080 15308
rect 15672 14912 15792 14940
rect 15396 14232 15608 14260
rect 15384 13728 15436 13734
rect 15384 13670 15436 13676
rect 15396 13190 15424 13670
rect 15476 13456 15528 13462
rect 15476 13398 15528 13404
rect 15384 13184 15436 13190
rect 15384 13126 15436 13132
rect 15304 12406 15424 12434
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 15200 11824 15252 11830
rect 15200 11766 15252 11772
rect 15198 11656 15254 11665
rect 15198 11591 15254 11600
rect 15108 8900 15160 8906
rect 15108 8842 15160 8848
rect 15212 8294 15240 11591
rect 15304 9994 15332 12038
rect 15396 11014 15424 12406
rect 15488 11218 15516 13398
rect 15580 13258 15608 14232
rect 15568 13252 15620 13258
rect 15568 13194 15620 13200
rect 15672 13138 15700 14912
rect 15936 14884 15988 14890
rect 15936 14826 15988 14832
rect 15844 14816 15896 14822
rect 15844 14758 15896 14764
rect 15856 13938 15884 14758
rect 15844 13932 15896 13938
rect 15844 13874 15896 13880
rect 15752 13796 15804 13802
rect 15752 13738 15804 13744
rect 15580 13110 15700 13138
rect 15580 11898 15608 13110
rect 15660 12708 15712 12714
rect 15660 12650 15712 12656
rect 15568 11892 15620 11898
rect 15568 11834 15620 11840
rect 15672 11665 15700 12650
rect 15764 12434 15792 13738
rect 15948 12434 15976 14826
rect 16040 12986 16068 15302
rect 16120 14952 16172 14958
rect 16120 14894 16172 14900
rect 16132 14482 16160 14894
rect 16120 14476 16172 14482
rect 16120 14418 16172 14424
rect 16224 13870 16252 15456
rect 16500 15094 16528 15506
rect 16488 15088 16540 15094
rect 16316 15048 16488 15076
rect 16212 13864 16264 13870
rect 16132 13824 16212 13852
rect 16028 12980 16080 12986
rect 16028 12922 16080 12928
rect 16132 12442 16160 13824
rect 16212 13806 16264 13812
rect 16316 13546 16344 15048
rect 16488 15030 16540 15036
rect 16578 15056 16634 15065
rect 16578 14991 16634 15000
rect 16592 14890 16620 14991
rect 16580 14884 16632 14890
rect 16580 14826 16632 14832
rect 16488 14272 16540 14278
rect 16488 14214 16540 14220
rect 16500 13870 16528 14214
rect 16580 14068 16632 14074
rect 16580 14010 16632 14016
rect 16488 13864 16540 13870
rect 16486 13832 16488 13841
rect 16540 13832 16542 13841
rect 16486 13767 16542 13776
rect 16316 13518 16436 13546
rect 16408 13258 16436 13518
rect 16396 13252 16448 13258
rect 16448 13212 16528 13240
rect 16396 13194 16448 13200
rect 16396 12980 16448 12986
rect 16396 12922 16448 12928
rect 16210 12880 16266 12889
rect 16210 12815 16212 12824
rect 16264 12815 16266 12824
rect 16212 12786 16264 12792
rect 16210 12744 16266 12753
rect 16210 12679 16266 12688
rect 16120 12436 16172 12442
rect 15764 12406 15884 12434
rect 15948 12406 16068 12434
rect 15856 12238 15884 12406
rect 15936 12368 15988 12374
rect 15936 12310 15988 12316
rect 15844 12232 15896 12238
rect 15844 12174 15896 12180
rect 15948 11762 15976 12310
rect 15936 11756 15988 11762
rect 15936 11698 15988 11704
rect 15658 11656 15714 11665
rect 15658 11591 15714 11600
rect 15660 11552 15712 11558
rect 15660 11494 15712 11500
rect 15476 11212 15528 11218
rect 15476 11154 15528 11160
rect 15384 11008 15436 11014
rect 15384 10950 15436 10956
rect 15568 10464 15620 10470
rect 15568 10406 15620 10412
rect 15292 9988 15344 9994
rect 15292 9930 15344 9936
rect 15292 9648 15344 9654
rect 15292 9590 15344 9596
rect 15304 9382 15332 9590
rect 15292 9376 15344 9382
rect 15292 9318 15344 9324
rect 15304 8974 15332 9318
rect 15384 9036 15436 9042
rect 15384 8978 15436 8984
rect 15292 8968 15344 8974
rect 15292 8910 15344 8916
rect 15304 8566 15332 8910
rect 15396 8634 15424 8978
rect 15580 8974 15608 10406
rect 15672 8974 15700 11494
rect 15844 11076 15896 11082
rect 15844 11018 15896 11024
rect 15856 10742 15884 11018
rect 15752 10736 15804 10742
rect 15752 10678 15804 10684
rect 15844 10736 15896 10742
rect 15844 10678 15896 10684
rect 16040 10690 16068 12406
rect 16120 12378 16172 12384
rect 16132 11801 16160 12378
rect 16118 11792 16174 11801
rect 16118 11727 16174 11736
rect 16224 11626 16252 12679
rect 16408 12102 16436 12922
rect 16500 12850 16528 13212
rect 16488 12844 16540 12850
rect 16488 12786 16540 12792
rect 16488 12708 16540 12714
rect 16488 12650 16540 12656
rect 16500 12209 16528 12650
rect 16486 12200 16542 12209
rect 16486 12135 16542 12144
rect 16396 12096 16448 12102
rect 16396 12038 16448 12044
rect 16488 12096 16540 12102
rect 16488 12038 16540 12044
rect 16408 11898 16436 12038
rect 16396 11892 16448 11898
rect 16396 11834 16448 11840
rect 16212 11620 16264 11626
rect 16212 11562 16264 11568
rect 16396 11008 16448 11014
rect 16396 10950 16448 10956
rect 15764 10554 15792 10678
rect 16040 10662 16252 10690
rect 16028 10600 16080 10606
rect 15764 10526 15884 10554
rect 16028 10542 16080 10548
rect 16120 10600 16172 10606
rect 16120 10542 16172 10548
rect 15856 9994 15884 10526
rect 16040 10266 16068 10542
rect 16028 10260 16080 10266
rect 16028 10202 16080 10208
rect 15844 9988 15896 9994
rect 15844 9930 15896 9936
rect 16132 9926 16160 10542
rect 16224 10266 16252 10662
rect 16408 10470 16436 10950
rect 16500 10674 16528 12038
rect 16592 11082 16620 14010
rect 16684 13938 16712 15846
rect 16776 14958 16804 15864
rect 16960 15881 16988 15914
rect 17132 15904 17184 15910
rect 16856 15846 16908 15852
rect 16946 15872 17002 15881
rect 17132 15846 17184 15852
rect 16946 15807 17002 15816
rect 16960 15638 16988 15807
rect 17144 15706 17172 15846
rect 17132 15700 17184 15706
rect 17132 15642 17184 15648
rect 16948 15632 17000 15638
rect 16948 15574 17000 15580
rect 17236 15026 17264 16238
rect 17314 15600 17370 15609
rect 17314 15535 17316 15544
rect 17368 15535 17370 15544
rect 17316 15506 17368 15512
rect 17224 15020 17276 15026
rect 17224 14962 17276 14968
rect 16764 14952 16816 14958
rect 16764 14894 16816 14900
rect 16672 13932 16724 13938
rect 16672 13874 16724 13880
rect 16776 12434 16804 14894
rect 17236 14618 17264 14962
rect 17420 14822 17448 16934
rect 17498 16895 17554 16904
rect 17590 15056 17646 15065
rect 17590 14991 17646 15000
rect 17500 14884 17552 14890
rect 17500 14826 17552 14832
rect 17408 14816 17460 14822
rect 17408 14758 17460 14764
rect 17132 14612 17184 14618
rect 17132 14554 17184 14560
rect 17224 14612 17276 14618
rect 17224 14554 17276 14560
rect 17144 14482 17172 14554
rect 17132 14476 17184 14482
rect 17132 14418 17184 14424
rect 17316 14408 17368 14414
rect 17316 14350 17368 14356
rect 16948 14272 17000 14278
rect 16948 14214 17000 14220
rect 16960 13569 16988 14214
rect 16946 13560 17002 13569
rect 16946 13495 17002 13504
rect 17132 13252 17184 13258
rect 17132 13194 17184 13200
rect 17144 12986 17172 13194
rect 17132 12980 17184 12986
rect 17132 12922 17184 12928
rect 17328 12434 17356 14350
rect 17512 14074 17540 14826
rect 17604 14482 17632 14991
rect 17592 14476 17644 14482
rect 17592 14418 17644 14424
rect 17500 14068 17552 14074
rect 17500 14010 17552 14016
rect 17408 13524 17460 13530
rect 17460 13484 17540 13512
rect 17408 13466 17460 13472
rect 17408 12640 17460 12646
rect 17408 12582 17460 12588
rect 16776 12406 16988 12434
rect 16856 12164 16908 12170
rect 16776 12124 16856 12152
rect 16776 11694 16804 12124
rect 16856 12106 16908 12112
rect 16764 11688 16816 11694
rect 16764 11630 16816 11636
rect 16670 11384 16726 11393
rect 16670 11319 16672 11328
rect 16724 11319 16726 11328
rect 16672 11290 16724 11296
rect 16580 11076 16632 11082
rect 16580 11018 16632 11024
rect 16488 10668 16540 10674
rect 16488 10610 16540 10616
rect 16580 10600 16632 10606
rect 16580 10542 16632 10548
rect 16396 10464 16448 10470
rect 16396 10406 16448 10412
rect 16212 10260 16264 10266
rect 16212 10202 16264 10208
rect 16592 10033 16620 10542
rect 16672 10056 16724 10062
rect 16578 10024 16634 10033
rect 16212 9988 16264 9994
rect 16672 9998 16724 10004
rect 16578 9959 16634 9968
rect 16212 9930 16264 9936
rect 16120 9920 16172 9926
rect 16120 9862 16172 9868
rect 16224 9586 16252 9930
rect 16592 9874 16620 9959
rect 16500 9846 16620 9874
rect 16500 9586 16528 9846
rect 16580 9716 16632 9722
rect 16580 9658 16632 9664
rect 16212 9580 16264 9586
rect 16212 9522 16264 9528
rect 16488 9580 16540 9586
rect 16488 9522 16540 9528
rect 16592 9450 16620 9658
rect 16684 9518 16712 9998
rect 16776 9518 16804 11630
rect 16854 11112 16910 11121
rect 16854 11047 16910 11056
rect 16868 10130 16896 11047
rect 16856 10124 16908 10130
rect 16856 10066 16908 10072
rect 16960 10010 16988 12406
rect 17236 12406 17356 12434
rect 17130 12336 17186 12345
rect 17236 12306 17264 12406
rect 17130 12271 17186 12280
rect 17224 12300 17276 12306
rect 17144 12238 17172 12271
rect 17224 12242 17276 12248
rect 17132 12232 17184 12238
rect 17132 12174 17184 12180
rect 17040 11212 17092 11218
rect 17040 11154 17092 11160
rect 16868 9982 16988 10010
rect 16672 9512 16724 9518
rect 16672 9454 16724 9460
rect 16764 9512 16816 9518
rect 16764 9454 16816 9460
rect 16580 9444 16632 9450
rect 16580 9386 16632 9392
rect 16776 9042 16804 9454
rect 16764 9036 16816 9042
rect 16764 8978 16816 8984
rect 15568 8968 15620 8974
rect 15568 8910 15620 8916
rect 15660 8968 15712 8974
rect 15660 8910 15712 8916
rect 16580 8900 16632 8906
rect 16580 8842 16632 8848
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 15292 8560 15344 8566
rect 15292 8502 15344 8508
rect 15752 8560 15804 8566
rect 15752 8502 15804 8508
rect 15764 8362 15792 8502
rect 15752 8356 15804 8362
rect 15752 8298 15804 8304
rect 15200 8288 15252 8294
rect 15200 8230 15252 8236
rect 16592 6798 16620 8842
rect 16672 8628 16724 8634
rect 16672 8570 16724 8576
rect 16684 8362 16712 8570
rect 16776 8498 16804 8978
rect 16764 8492 16816 8498
rect 16764 8434 16816 8440
rect 16868 8362 16896 9982
rect 16948 9920 17000 9926
rect 16948 9862 17000 9868
rect 16672 8356 16724 8362
rect 16672 8298 16724 8304
rect 16856 8356 16908 8362
rect 16856 8298 16908 8304
rect 16580 6792 16632 6798
rect 16580 6734 16632 6740
rect 14924 4072 14976 4078
rect 14924 4014 14976 4020
rect 16684 3126 16712 8298
rect 16960 7954 16988 9862
rect 17052 9042 17080 11154
rect 17236 9654 17264 12242
rect 17314 12200 17370 12209
rect 17314 12135 17370 12144
rect 17328 12102 17356 12135
rect 17316 12096 17368 12102
rect 17316 12038 17368 12044
rect 17420 10130 17448 12582
rect 17512 10130 17540 13484
rect 17604 10742 17632 14418
rect 17684 13864 17736 13870
rect 17684 13806 17736 13812
rect 17696 13530 17724 13806
rect 17684 13524 17736 13530
rect 17684 13466 17736 13472
rect 17788 13462 17816 18158
rect 18328 17672 18380 17678
rect 18328 17614 18380 17620
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 18340 17270 18368 17614
rect 18512 17536 18564 17542
rect 18512 17478 18564 17484
rect 18420 17332 18472 17338
rect 18420 17274 18472 17280
rect 18328 17264 18380 17270
rect 18328 17206 18380 17212
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 18340 16250 18368 17206
rect 18432 16726 18460 17274
rect 18524 17202 18552 17478
rect 18512 17196 18564 17202
rect 18512 17138 18564 17144
rect 18420 16720 18472 16726
rect 18420 16662 18472 16668
rect 18328 16244 18380 16250
rect 18328 16186 18380 16192
rect 17868 15428 17920 15434
rect 17868 15370 17920 15376
rect 17880 14618 17908 15370
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 17868 14612 17920 14618
rect 17868 14554 17920 14560
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 17776 13456 17828 13462
rect 17776 13398 17828 13404
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 18340 12918 18368 16186
rect 18420 16108 18472 16114
rect 18420 16050 18472 16056
rect 18432 14074 18460 16050
rect 18524 15706 18552 17138
rect 18604 17128 18656 17134
rect 18604 17070 18656 17076
rect 18616 16658 18644 17070
rect 18604 16652 18656 16658
rect 18604 16594 18656 16600
rect 18616 16114 18644 16594
rect 18604 16108 18656 16114
rect 18604 16050 18656 16056
rect 18512 15700 18564 15706
rect 18512 15642 18564 15648
rect 18524 14278 18552 15642
rect 18604 15020 18656 15026
rect 18604 14962 18656 14968
rect 18616 14618 18644 14962
rect 18604 14612 18656 14618
rect 18604 14554 18656 14560
rect 18512 14272 18564 14278
rect 18512 14214 18564 14220
rect 18420 14068 18472 14074
rect 18420 14010 18472 14016
rect 18510 13832 18566 13841
rect 18510 13767 18566 13776
rect 17960 12912 18012 12918
rect 17960 12854 18012 12860
rect 18328 12912 18380 12918
rect 18328 12854 18380 12860
rect 17684 12708 17736 12714
rect 17684 12650 17736 12656
rect 17696 11257 17724 12650
rect 17972 12238 18000 12854
rect 17960 12232 18012 12238
rect 17960 12174 18012 12180
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 18144 11552 18196 11558
rect 18236 11552 18288 11558
rect 18144 11494 18196 11500
rect 18234 11520 18236 11529
rect 18288 11520 18290 11529
rect 17682 11248 17738 11257
rect 17682 11183 17738 11192
rect 17592 10736 17644 10742
rect 17592 10678 17644 10684
rect 17408 10124 17460 10130
rect 17408 10066 17460 10072
rect 17500 10124 17552 10130
rect 17552 10084 17632 10112
rect 17500 10066 17552 10072
rect 17316 9920 17368 9926
rect 17316 9862 17368 9868
rect 17328 9722 17356 9862
rect 17316 9716 17368 9722
rect 17316 9658 17368 9664
rect 17224 9648 17276 9654
rect 17224 9590 17276 9596
rect 17040 9036 17092 9042
rect 17040 8978 17092 8984
rect 17052 8566 17080 8978
rect 17224 8900 17276 8906
rect 17224 8842 17276 8848
rect 17236 8634 17264 8842
rect 17224 8628 17276 8634
rect 17224 8570 17276 8576
rect 17040 8560 17092 8566
rect 17040 8502 17092 8508
rect 17052 8022 17080 8502
rect 17040 8016 17092 8022
rect 17040 7958 17092 7964
rect 16948 7948 17000 7954
rect 16948 7890 17000 7896
rect 17328 7478 17356 9658
rect 17408 9648 17460 9654
rect 17408 9590 17460 9596
rect 17420 8566 17448 9590
rect 17604 8838 17632 10084
rect 17592 8832 17644 8838
rect 17592 8774 17644 8780
rect 17408 8560 17460 8566
rect 17408 8502 17460 8508
rect 17420 7546 17448 8502
rect 17408 7540 17460 7546
rect 17408 7482 17460 7488
rect 17316 7472 17368 7478
rect 17316 7414 17368 7420
rect 17696 5574 17724 11183
rect 18156 11082 18184 11494
rect 18234 11455 18290 11464
rect 18418 11248 18474 11257
rect 18418 11183 18474 11192
rect 18432 11150 18460 11183
rect 18328 11144 18380 11150
rect 18328 11086 18380 11092
rect 18420 11144 18472 11150
rect 18420 11086 18472 11092
rect 17776 11076 17828 11082
rect 17776 11018 17828 11024
rect 18144 11076 18196 11082
rect 18144 11018 18196 11024
rect 17788 8430 17816 11018
rect 17868 11008 17920 11014
rect 17868 10950 17920 10956
rect 17880 10724 17908 10950
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 18052 10804 18104 10810
rect 18052 10746 18104 10752
rect 17880 10696 18000 10724
rect 17972 10198 18000 10696
rect 18064 10266 18092 10746
rect 18236 10668 18288 10674
rect 18236 10610 18288 10616
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 17960 10192 18012 10198
rect 17960 10134 18012 10140
rect 18248 10130 18276 10610
rect 18340 10266 18368 11086
rect 18420 10464 18472 10470
rect 18420 10406 18472 10412
rect 18328 10260 18380 10266
rect 18328 10202 18380 10208
rect 18236 10124 18288 10130
rect 18236 10066 18288 10072
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 17868 9172 17920 9178
rect 17868 9114 17920 9120
rect 17776 8424 17828 8430
rect 17776 8366 17828 8372
rect 17880 6322 17908 9114
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 18432 7886 18460 10406
rect 18524 10130 18552 13767
rect 18616 11218 18644 14554
rect 18708 12646 18736 18770
rect 18800 17746 18828 20198
rect 18892 19990 18920 20538
rect 18984 20398 19012 21082
rect 18972 20392 19024 20398
rect 18972 20334 19024 20340
rect 18880 19984 18932 19990
rect 18880 19926 18932 19932
rect 18984 18834 19012 20334
rect 19076 19922 19104 23598
rect 19340 23180 19392 23186
rect 19340 23122 19392 23128
rect 19248 23112 19300 23118
rect 19248 23054 19300 23060
rect 19156 21140 19208 21146
rect 19156 21082 19208 21088
rect 19168 20874 19196 21082
rect 19260 21049 19288 23054
rect 19352 22642 19380 23122
rect 19340 22636 19392 22642
rect 19340 22578 19392 22584
rect 19444 22030 19472 24006
rect 20168 23724 20220 23730
rect 20168 23666 20220 23672
rect 20180 23594 20208 23666
rect 20168 23588 20220 23594
rect 20168 23530 20220 23536
rect 20180 23186 20208 23530
rect 20352 23520 20404 23526
rect 20352 23462 20404 23468
rect 20364 23186 20392 23462
rect 20168 23180 20220 23186
rect 20168 23122 20220 23128
rect 20352 23180 20404 23186
rect 20352 23122 20404 23128
rect 19708 23044 19760 23050
rect 19708 22986 19760 22992
rect 19432 22024 19484 22030
rect 19432 21966 19484 21972
rect 19338 21720 19394 21729
rect 19338 21655 19394 21664
rect 19246 21040 19302 21049
rect 19246 20975 19302 20984
rect 19156 20868 19208 20874
rect 19156 20810 19208 20816
rect 19168 20602 19196 20810
rect 19156 20596 19208 20602
rect 19156 20538 19208 20544
rect 19168 20466 19196 20538
rect 19352 20534 19380 21655
rect 19720 20913 19748 22986
rect 20364 22438 20392 23122
rect 20456 22778 20484 24074
rect 20732 23594 20760 24346
rect 20916 24274 20944 26200
rect 20996 24336 21048 24342
rect 20996 24278 21048 24284
rect 20904 24268 20956 24274
rect 20904 24210 20956 24216
rect 21008 23866 21036 24278
rect 21272 24200 21324 24206
rect 21272 24142 21324 24148
rect 21284 23866 21312 24142
rect 20996 23860 21048 23866
rect 20996 23802 21048 23808
rect 21272 23860 21324 23866
rect 21272 23802 21324 23808
rect 20720 23588 20772 23594
rect 20720 23530 20772 23536
rect 20536 23520 20588 23526
rect 20536 23462 20588 23468
rect 21088 23520 21140 23526
rect 21088 23462 21140 23468
rect 20548 22982 20576 23462
rect 21100 23050 21128 23462
rect 20720 23044 20772 23050
rect 20720 22986 20772 22992
rect 21088 23044 21140 23050
rect 21088 22986 21140 22992
rect 20536 22976 20588 22982
rect 20536 22918 20588 22924
rect 20444 22772 20496 22778
rect 20444 22714 20496 22720
rect 20352 22432 20404 22438
rect 20352 22374 20404 22380
rect 20548 21690 20576 22918
rect 20732 22506 20760 22986
rect 21100 22710 21128 22986
rect 21088 22704 21140 22710
rect 21088 22646 21140 22652
rect 20720 22500 20772 22506
rect 20720 22442 20772 22448
rect 21100 22098 21128 22646
rect 21560 22574 21588 26200
rect 22100 23656 22152 23662
rect 22100 23598 22152 23604
rect 22008 23588 22060 23594
rect 22008 23530 22060 23536
rect 22020 23254 22048 23530
rect 22112 23254 22140 23598
rect 22008 23248 22060 23254
rect 22008 23190 22060 23196
rect 22100 23248 22152 23254
rect 22100 23190 22152 23196
rect 22008 23112 22060 23118
rect 21928 23072 22008 23100
rect 21548 22568 21600 22574
rect 21548 22510 21600 22516
rect 21180 22500 21232 22506
rect 21180 22442 21232 22448
rect 21192 22137 21220 22442
rect 21456 22160 21508 22166
rect 21178 22128 21234 22137
rect 20720 22092 20772 22098
rect 20720 22034 20772 22040
rect 21088 22092 21140 22098
rect 21456 22102 21508 22108
rect 21638 22128 21694 22137
rect 21178 22063 21234 22072
rect 21088 22034 21140 22040
rect 20536 21684 20588 21690
rect 20536 21626 20588 21632
rect 20732 21622 20760 22034
rect 21270 21856 21326 21865
rect 21270 21791 21326 21800
rect 20720 21616 20772 21622
rect 20720 21558 20772 21564
rect 20732 21350 20760 21558
rect 20352 21344 20404 21350
rect 20352 21286 20404 21292
rect 20720 21344 20772 21350
rect 20720 21286 20772 21292
rect 19706 20904 19762 20913
rect 19706 20839 19762 20848
rect 19982 20632 20038 20641
rect 19982 20567 20038 20576
rect 20260 20596 20312 20602
rect 19996 20534 20024 20567
rect 20260 20538 20312 20544
rect 19340 20528 19392 20534
rect 19340 20470 19392 20476
rect 19984 20528 20036 20534
rect 19984 20470 20036 20476
rect 19156 20460 19208 20466
rect 19156 20402 19208 20408
rect 19064 19916 19116 19922
rect 19064 19858 19116 19864
rect 19340 19916 19392 19922
rect 19340 19858 19392 19864
rect 19352 19689 19380 19858
rect 19616 19780 19668 19786
rect 19616 19722 19668 19728
rect 20168 19780 20220 19786
rect 20168 19722 20220 19728
rect 19338 19680 19394 19689
rect 19338 19615 19394 19624
rect 19352 19514 19380 19615
rect 19340 19508 19392 19514
rect 19340 19450 19392 19456
rect 19628 18970 19656 19722
rect 19708 19508 19760 19514
rect 19708 19450 19760 19456
rect 19616 18964 19668 18970
rect 19616 18906 19668 18912
rect 19430 18864 19486 18873
rect 18972 18828 19024 18834
rect 19430 18799 19486 18808
rect 18972 18770 19024 18776
rect 19064 18760 19116 18766
rect 18878 18728 18934 18737
rect 19064 18702 19116 18708
rect 18878 18663 18880 18672
rect 18932 18663 18934 18672
rect 18880 18634 18932 18640
rect 19076 18329 19104 18702
rect 19156 18624 19208 18630
rect 19156 18566 19208 18572
rect 19340 18624 19392 18630
rect 19340 18566 19392 18572
rect 19062 18320 19118 18329
rect 19062 18255 19118 18264
rect 18972 18080 19024 18086
rect 18972 18022 19024 18028
rect 18788 17740 18840 17746
rect 18788 17682 18840 17688
rect 18984 17678 19012 18022
rect 18972 17672 19024 17678
rect 18972 17614 19024 17620
rect 18788 16788 18840 16794
rect 18788 16730 18840 16736
rect 18800 13802 18828 16730
rect 18880 16448 18932 16454
rect 18880 16390 18932 16396
rect 18972 16448 19024 16454
rect 18972 16390 19024 16396
rect 18892 16182 18920 16390
rect 18880 16176 18932 16182
rect 18880 16118 18932 16124
rect 18880 14952 18932 14958
rect 18880 14894 18932 14900
rect 18892 14550 18920 14894
rect 18880 14544 18932 14550
rect 18880 14486 18932 14492
rect 18984 14074 19012 16390
rect 19064 16244 19116 16250
rect 19064 16186 19116 16192
rect 19076 15978 19104 16186
rect 19064 15972 19116 15978
rect 19064 15914 19116 15920
rect 19168 15638 19196 18566
rect 19352 18465 19380 18566
rect 19338 18456 19394 18465
rect 19338 18391 19394 18400
rect 19444 15706 19472 18799
rect 19524 18284 19576 18290
rect 19524 18226 19576 18232
rect 19432 15700 19484 15706
rect 19432 15642 19484 15648
rect 19156 15632 19208 15638
rect 19156 15574 19208 15580
rect 19444 15162 19472 15642
rect 19536 15162 19564 18226
rect 19616 18148 19668 18154
rect 19616 18090 19668 18096
rect 19628 17882 19656 18090
rect 19616 17876 19668 17882
rect 19616 17818 19668 17824
rect 19720 17610 19748 19450
rect 20076 19372 20128 19378
rect 20076 19314 20128 19320
rect 19800 19168 19852 19174
rect 19800 19110 19852 19116
rect 19812 18737 19840 19110
rect 19798 18728 19854 18737
rect 19798 18663 19854 18672
rect 19708 17604 19760 17610
rect 19708 17546 19760 17552
rect 19812 17490 19840 18663
rect 19892 18352 19944 18358
rect 19892 18294 19944 18300
rect 19904 17746 19932 18294
rect 19892 17740 19944 17746
rect 19892 17682 19944 17688
rect 19904 17610 19932 17682
rect 19892 17604 19944 17610
rect 19892 17546 19944 17552
rect 19628 17462 19840 17490
rect 19432 15156 19484 15162
rect 19432 15098 19484 15104
rect 19524 15156 19576 15162
rect 19524 15098 19576 15104
rect 19248 15020 19300 15026
rect 19248 14962 19300 14968
rect 19064 14612 19116 14618
rect 19064 14554 19116 14560
rect 18972 14068 19024 14074
rect 18972 14010 19024 14016
rect 18972 13864 19024 13870
rect 19076 13841 19104 14554
rect 18972 13806 19024 13812
rect 19062 13832 19118 13841
rect 18788 13796 18840 13802
rect 18788 13738 18840 13744
rect 18984 13394 19012 13806
rect 19062 13767 19118 13776
rect 18972 13388 19024 13394
rect 18972 13330 19024 13336
rect 18788 12912 18840 12918
rect 18788 12854 18840 12860
rect 18696 12640 18748 12646
rect 18696 12582 18748 12588
rect 18800 11898 18828 12854
rect 18984 12850 19012 13330
rect 19260 13297 19288 14962
rect 19628 14822 19656 17462
rect 20088 17218 20116 19314
rect 20180 19310 20208 19722
rect 20168 19304 20220 19310
rect 20168 19246 20220 19252
rect 20272 17746 20300 20538
rect 20364 19553 20392 21286
rect 20732 21146 20760 21286
rect 21284 21146 21312 21791
rect 20720 21140 20772 21146
rect 20720 21082 20772 21088
rect 21272 21140 21324 21146
rect 21272 21082 21324 21088
rect 21086 21040 21142 21049
rect 20444 21004 20496 21010
rect 21086 20975 21142 20984
rect 20444 20946 20496 20952
rect 20350 19544 20406 19553
rect 20350 19479 20406 19488
rect 20260 17740 20312 17746
rect 20260 17682 20312 17688
rect 20168 17672 20220 17678
rect 20168 17614 20220 17620
rect 19996 17190 20116 17218
rect 19892 16992 19944 16998
rect 19892 16934 19944 16940
rect 19706 16688 19762 16697
rect 19706 16623 19762 16632
rect 19340 14816 19392 14822
rect 19340 14758 19392 14764
rect 19616 14816 19668 14822
rect 19616 14758 19668 14764
rect 19246 13288 19302 13297
rect 19246 13223 19302 13232
rect 19064 13184 19116 13190
rect 19064 13126 19116 13132
rect 18972 12844 19024 12850
rect 18972 12786 19024 12792
rect 18788 11892 18840 11898
rect 18788 11834 18840 11840
rect 18788 11280 18840 11286
rect 18788 11222 18840 11228
rect 18604 11212 18656 11218
rect 18604 11154 18656 11160
rect 18602 11112 18658 11121
rect 18602 11047 18658 11056
rect 18616 11014 18644 11047
rect 18604 11008 18656 11014
rect 18604 10950 18656 10956
rect 18696 10668 18748 10674
rect 18696 10610 18748 10616
rect 18512 10124 18564 10130
rect 18512 10066 18564 10072
rect 18420 7880 18472 7886
rect 18420 7822 18472 7828
rect 18524 7818 18552 10066
rect 18604 9512 18656 9518
rect 18604 9454 18656 9460
rect 18616 8634 18644 9454
rect 18708 9042 18736 10610
rect 18696 9036 18748 9042
rect 18696 8978 18748 8984
rect 18604 8628 18656 8634
rect 18604 8570 18656 8576
rect 18616 7954 18644 8570
rect 18604 7948 18656 7954
rect 18604 7890 18656 7896
rect 18512 7812 18564 7818
rect 18512 7754 18564 7760
rect 18800 7750 18828 11222
rect 18880 11212 18932 11218
rect 18880 11154 18932 11160
rect 18892 9654 18920 11154
rect 19076 11082 19104 13126
rect 19260 12434 19288 13223
rect 19352 12442 19380 14758
rect 19524 14272 19576 14278
rect 19524 14214 19576 14220
rect 19536 14006 19564 14214
rect 19524 14000 19576 14006
rect 19524 13942 19576 13948
rect 19432 13932 19484 13938
rect 19432 13874 19484 13880
rect 19444 13462 19472 13874
rect 19432 13456 19484 13462
rect 19432 13398 19484 13404
rect 19720 13190 19748 16623
rect 19798 16144 19854 16153
rect 19798 16079 19854 16088
rect 19812 15502 19840 16079
rect 19904 15706 19932 16934
rect 19892 15700 19944 15706
rect 19892 15642 19944 15648
rect 19800 15496 19852 15502
rect 19800 15438 19852 15444
rect 19996 15162 20024 17190
rect 20076 17128 20128 17134
rect 20076 17070 20128 17076
rect 19984 15156 20036 15162
rect 19984 15098 20036 15104
rect 20088 14958 20116 17070
rect 20180 15450 20208 17614
rect 20272 17338 20300 17682
rect 20364 17626 20392 19479
rect 20456 19242 20484 20946
rect 21100 20942 21128 20975
rect 21088 20936 21140 20942
rect 21088 20878 21140 20884
rect 21180 20936 21232 20942
rect 21180 20878 21232 20884
rect 21192 20482 21220 20878
rect 21272 20528 21324 20534
rect 21192 20476 21272 20482
rect 21192 20470 21324 20476
rect 21192 20454 21312 20470
rect 20536 20052 20588 20058
rect 20536 19994 20588 20000
rect 20548 19446 20576 19994
rect 21192 19922 21220 20454
rect 21468 20398 21496 22102
rect 21638 22063 21694 22072
rect 21548 21140 21600 21146
rect 21548 21082 21600 21088
rect 21560 21049 21588 21082
rect 21546 21040 21602 21049
rect 21546 20975 21602 20984
rect 21548 20868 21600 20874
rect 21548 20810 21600 20816
rect 21560 20466 21588 20810
rect 21548 20460 21600 20466
rect 21548 20402 21600 20408
rect 21456 20392 21508 20398
rect 21456 20334 21508 20340
rect 21180 19916 21232 19922
rect 21180 19858 21232 19864
rect 21364 19916 21416 19922
rect 21364 19858 21416 19864
rect 21088 19712 21140 19718
rect 21088 19654 21140 19660
rect 21180 19712 21232 19718
rect 21180 19654 21232 19660
rect 20536 19440 20588 19446
rect 20536 19382 20588 19388
rect 20444 19236 20496 19242
rect 20444 19178 20496 19184
rect 20548 19174 20576 19382
rect 20536 19168 20588 19174
rect 20536 19110 20588 19116
rect 21100 18970 21128 19654
rect 21088 18964 21140 18970
rect 21088 18906 21140 18912
rect 21192 18630 21220 19654
rect 21376 18834 21404 19858
rect 21560 19786 21588 20402
rect 21548 19780 21600 19786
rect 21548 19722 21600 19728
rect 21560 19174 21588 19722
rect 21548 19168 21600 19174
rect 21548 19110 21600 19116
rect 21364 18828 21416 18834
rect 21364 18770 21416 18776
rect 21180 18624 21232 18630
rect 21456 18624 21508 18630
rect 21180 18566 21232 18572
rect 21270 18592 21326 18601
rect 21456 18566 21508 18572
rect 21270 18527 21326 18536
rect 20904 18216 20956 18222
rect 20904 18158 20956 18164
rect 20364 17610 20576 17626
rect 20364 17604 20588 17610
rect 20364 17598 20536 17604
rect 20536 17546 20588 17552
rect 20352 17536 20404 17542
rect 20352 17478 20404 17484
rect 20720 17536 20772 17542
rect 20720 17478 20772 17484
rect 20364 17338 20392 17478
rect 20260 17332 20312 17338
rect 20260 17274 20312 17280
rect 20352 17332 20404 17338
rect 20352 17274 20404 17280
rect 20272 16640 20300 17274
rect 20536 17196 20588 17202
rect 20536 17138 20588 17144
rect 20352 16652 20404 16658
rect 20272 16612 20352 16640
rect 20352 16594 20404 16600
rect 20548 16454 20576 17138
rect 20536 16448 20588 16454
rect 20536 16390 20588 16396
rect 20536 15904 20588 15910
rect 20536 15846 20588 15852
rect 20180 15422 20392 15450
rect 20260 15360 20312 15366
rect 20260 15302 20312 15308
rect 20076 14952 20128 14958
rect 20076 14894 20128 14900
rect 19892 14816 19944 14822
rect 19892 14758 19944 14764
rect 19904 14346 19932 14758
rect 19892 14340 19944 14346
rect 19892 14282 19944 14288
rect 19800 14272 19852 14278
rect 19800 14214 19852 14220
rect 19982 14240 20038 14249
rect 19812 14074 19840 14214
rect 19982 14175 20038 14184
rect 19800 14068 19852 14074
rect 19800 14010 19852 14016
rect 19812 13734 19840 14010
rect 19800 13728 19852 13734
rect 19800 13670 19852 13676
rect 19892 13456 19944 13462
rect 19892 13398 19944 13404
rect 19708 13184 19760 13190
rect 19708 13126 19760 13132
rect 19616 12844 19668 12850
rect 19616 12786 19668 12792
rect 19524 12776 19576 12782
rect 19524 12718 19576 12724
rect 19168 12406 19288 12434
rect 19340 12436 19392 12442
rect 19064 11076 19116 11082
rect 19064 11018 19116 11024
rect 18880 9648 18932 9654
rect 18880 9590 18932 9596
rect 18880 8084 18932 8090
rect 18880 8026 18932 8032
rect 18788 7744 18840 7750
rect 18788 7686 18840 7692
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 17868 6316 17920 6322
rect 17868 6258 17920 6264
rect 18328 6248 18380 6254
rect 18328 6190 18380 6196
rect 17684 5568 17736 5574
rect 17684 5510 17736 5516
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 18340 4010 18368 6190
rect 18892 5234 18920 8026
rect 19168 7274 19196 12406
rect 19340 12378 19392 12384
rect 19340 12300 19392 12306
rect 19340 12242 19392 12248
rect 19248 11892 19300 11898
rect 19248 11834 19300 11840
rect 19260 11354 19288 11834
rect 19352 11830 19380 12242
rect 19536 12238 19564 12718
rect 19524 12232 19576 12238
rect 19524 12174 19576 12180
rect 19340 11824 19392 11830
rect 19340 11766 19392 11772
rect 19248 11348 19300 11354
rect 19248 11290 19300 11296
rect 19524 11144 19576 11150
rect 19524 11086 19576 11092
rect 19536 9654 19564 11086
rect 19628 10130 19656 12786
rect 19708 12776 19760 12782
rect 19708 12718 19760 12724
rect 19720 10810 19748 12718
rect 19904 11830 19932 13398
rect 19996 13326 20024 14175
rect 20272 13530 20300 15302
rect 20364 13530 20392 15422
rect 20548 15201 20576 15846
rect 20534 15192 20590 15201
rect 20534 15127 20590 15136
rect 20536 14952 20588 14958
rect 20536 14894 20588 14900
rect 20548 14278 20576 14894
rect 20732 14482 20760 17478
rect 20916 17338 20944 18158
rect 21180 17536 21232 17542
rect 21180 17478 21232 17484
rect 20904 17332 20956 17338
rect 20904 17274 20956 17280
rect 20996 17332 21048 17338
rect 20996 17274 21048 17280
rect 21008 16794 21036 17274
rect 21192 16969 21220 17478
rect 21178 16960 21234 16969
rect 21178 16895 21234 16904
rect 20996 16788 21048 16794
rect 20996 16730 21048 16736
rect 20994 16552 21050 16561
rect 20994 16487 21050 16496
rect 20812 16448 20864 16454
rect 20812 16390 20864 16396
rect 20824 16182 20852 16390
rect 20812 16176 20864 16182
rect 20812 16118 20864 16124
rect 20812 15088 20864 15094
rect 20812 15030 20864 15036
rect 20720 14476 20772 14482
rect 20720 14418 20772 14424
rect 20536 14272 20588 14278
rect 20536 14214 20588 14220
rect 20720 14272 20772 14278
rect 20720 14214 20772 14220
rect 20444 13728 20496 13734
rect 20444 13670 20496 13676
rect 20260 13524 20312 13530
rect 20260 13466 20312 13472
rect 20352 13524 20404 13530
rect 20352 13466 20404 13472
rect 20168 13388 20220 13394
rect 20168 13330 20220 13336
rect 19984 13320 20036 13326
rect 19984 13262 20036 13268
rect 20074 12744 20130 12753
rect 20074 12679 20130 12688
rect 19984 12300 20036 12306
rect 19984 12242 20036 12248
rect 19892 11824 19944 11830
rect 19890 11792 19892 11801
rect 19944 11792 19946 11801
rect 19890 11727 19946 11736
rect 19904 11354 19932 11727
rect 19892 11348 19944 11354
rect 19892 11290 19944 11296
rect 19892 11008 19944 11014
rect 19892 10950 19944 10956
rect 19904 10810 19932 10950
rect 19708 10804 19760 10810
rect 19708 10746 19760 10752
rect 19892 10804 19944 10810
rect 19892 10746 19944 10752
rect 19616 10124 19668 10130
rect 19616 10066 19668 10072
rect 19708 10124 19760 10130
rect 19708 10066 19760 10072
rect 19524 9648 19576 9654
rect 19524 9590 19576 9596
rect 19536 9178 19564 9590
rect 19524 9172 19576 9178
rect 19524 9114 19576 9120
rect 19720 9042 19748 10066
rect 19800 10056 19852 10062
rect 19800 9998 19852 10004
rect 19708 9036 19760 9042
rect 19708 8978 19760 8984
rect 19720 8498 19748 8978
rect 19812 8906 19840 9998
rect 19800 8900 19852 8906
rect 19800 8842 19852 8848
rect 19708 8492 19760 8498
rect 19708 8434 19760 8440
rect 19248 8016 19300 8022
rect 19248 7958 19300 7964
rect 19156 7268 19208 7274
rect 19156 7210 19208 7216
rect 19260 6798 19288 7958
rect 19720 7954 19748 8434
rect 19812 8090 19840 8842
rect 19996 8634 20024 12242
rect 20088 11830 20116 12679
rect 20076 11824 20128 11830
rect 20076 11766 20128 11772
rect 20076 11620 20128 11626
rect 20180 11608 20208 13330
rect 20456 13190 20484 13670
rect 20444 13184 20496 13190
rect 20444 13126 20496 13132
rect 20548 12986 20576 14214
rect 20732 13870 20760 14214
rect 20720 13864 20772 13870
rect 20720 13806 20772 13812
rect 20536 12980 20588 12986
rect 20536 12922 20588 12928
rect 20628 12300 20680 12306
rect 20628 12242 20680 12248
rect 20536 12096 20588 12102
rect 20536 12038 20588 12044
rect 20128 11580 20208 11608
rect 20076 11562 20128 11568
rect 19984 8628 20036 8634
rect 19984 8570 20036 8576
rect 19800 8084 19852 8090
rect 19800 8026 19852 8032
rect 19708 7948 19760 7954
rect 19708 7890 19760 7896
rect 19996 7818 20024 8570
rect 19984 7812 20036 7818
rect 19984 7754 20036 7760
rect 20548 7546 20576 12038
rect 20640 11694 20668 12242
rect 20628 11688 20680 11694
rect 20628 11630 20680 11636
rect 20824 11626 20852 15030
rect 20904 15020 20956 15026
rect 20904 14962 20956 14968
rect 20916 13190 20944 14962
rect 20904 13184 20956 13190
rect 20904 13126 20956 13132
rect 20904 12980 20956 12986
rect 20904 12922 20956 12928
rect 20916 12782 20944 12922
rect 21008 12918 21036 16487
rect 21088 15496 21140 15502
rect 21088 15438 21140 15444
rect 21100 14618 21128 15438
rect 21088 14612 21140 14618
rect 21088 14554 21140 14560
rect 21192 14498 21220 16895
rect 21284 16658 21312 18527
rect 21468 17542 21496 18566
rect 21560 18358 21588 19110
rect 21652 18834 21680 22063
rect 21928 22030 21956 23072
rect 22008 23054 22060 23060
rect 22204 22234 22232 26200
rect 22560 24064 22612 24070
rect 22560 24006 22612 24012
rect 22284 22976 22336 22982
rect 22284 22918 22336 22924
rect 22296 22710 22324 22918
rect 22284 22704 22336 22710
rect 22284 22646 22336 22652
rect 22468 22432 22520 22438
rect 22468 22374 22520 22380
rect 22192 22228 22244 22234
rect 22192 22170 22244 22176
rect 21916 22024 21968 22030
rect 21916 21966 21968 21972
rect 21916 21888 21968 21894
rect 21916 21830 21968 21836
rect 21928 21690 21956 21830
rect 21916 21684 21968 21690
rect 21916 21626 21968 21632
rect 22284 21684 22336 21690
rect 22284 21626 22336 21632
rect 22296 21418 22324 21626
rect 22480 21486 22508 22374
rect 22468 21480 22520 21486
rect 22468 21422 22520 21428
rect 22284 21412 22336 21418
rect 22284 21354 22336 21360
rect 21916 21344 21968 21350
rect 21916 21286 21968 21292
rect 21928 20874 21956 21286
rect 21916 20868 21968 20874
rect 21916 20810 21968 20816
rect 21914 20632 21970 20641
rect 22480 20602 22508 21422
rect 22572 20754 22600 24006
rect 22848 23322 22876 26200
rect 23296 24676 23348 24682
rect 23296 24618 23348 24624
rect 23388 24676 23440 24682
rect 23388 24618 23440 24624
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 23308 23866 23336 24618
rect 23296 23860 23348 23866
rect 23296 23802 23348 23808
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 22836 23316 22888 23322
rect 22836 23258 22888 23264
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 23204 22092 23256 22098
rect 23204 22034 23256 22040
rect 22742 21992 22798 22001
rect 22742 21927 22798 21936
rect 22652 21888 22704 21894
rect 22652 21830 22704 21836
rect 22664 21146 22692 21830
rect 22756 21622 22784 21927
rect 23216 21865 23244 22034
rect 23202 21856 23258 21865
rect 23202 21791 23258 21800
rect 22744 21616 22796 21622
rect 23204 21616 23256 21622
rect 22744 21558 22796 21564
rect 22834 21584 22890 21593
rect 23204 21558 23256 21564
rect 22834 21519 22890 21528
rect 22848 21146 22876 21519
rect 23216 21350 23244 21558
rect 23204 21344 23256 21350
rect 23204 21286 23256 21292
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 22652 21140 22704 21146
rect 22652 21082 22704 21088
rect 22836 21140 22888 21146
rect 22836 21082 22888 21088
rect 22572 20726 22876 20754
rect 22848 20602 22876 20726
rect 21914 20567 21970 20576
rect 22468 20596 22520 20602
rect 21822 19952 21878 19961
rect 21822 19887 21878 19896
rect 21732 19440 21784 19446
rect 21732 19382 21784 19388
rect 21640 18828 21692 18834
rect 21640 18770 21692 18776
rect 21640 18624 21692 18630
rect 21640 18566 21692 18572
rect 21548 18352 21600 18358
rect 21548 18294 21600 18300
rect 21560 17610 21588 18294
rect 21652 17785 21680 18566
rect 21744 17882 21772 19382
rect 21732 17876 21784 17882
rect 21732 17818 21784 17824
rect 21638 17776 21694 17785
rect 21638 17711 21694 17720
rect 21548 17604 21600 17610
rect 21548 17546 21600 17552
rect 21456 17536 21508 17542
rect 21456 17478 21508 17484
rect 21560 16998 21588 17546
rect 21548 16992 21600 16998
rect 21548 16934 21600 16940
rect 21272 16652 21324 16658
rect 21324 16612 21496 16640
rect 21272 16594 21324 16600
rect 21364 15564 21416 15570
rect 21364 15506 21416 15512
rect 21272 15088 21324 15094
rect 21272 15030 21324 15036
rect 21100 14470 21220 14498
rect 21100 13190 21128 14470
rect 21284 14346 21312 15030
rect 21376 14482 21404 15506
rect 21468 14618 21496 16612
rect 21560 16182 21588 16934
rect 21548 16176 21600 16182
rect 21548 16118 21600 16124
rect 21548 15496 21600 15502
rect 21548 15438 21600 15444
rect 21456 14612 21508 14618
rect 21456 14554 21508 14560
rect 21364 14476 21416 14482
rect 21364 14418 21416 14424
rect 21272 14340 21324 14346
rect 21272 14282 21324 14288
rect 21376 13870 21404 14418
rect 21364 13864 21416 13870
rect 21364 13806 21416 13812
rect 21468 13394 21496 14554
rect 21560 13852 21588 15438
rect 21652 15065 21680 17711
rect 21732 15700 21784 15706
rect 21732 15642 21784 15648
rect 21744 15570 21772 15642
rect 21732 15564 21784 15570
rect 21732 15506 21784 15512
rect 21836 15162 21864 19887
rect 21928 18086 21956 20567
rect 22468 20538 22520 20544
rect 22744 20596 22796 20602
rect 22744 20538 22796 20544
rect 22836 20596 22888 20602
rect 22836 20538 22888 20544
rect 22468 20392 22520 20398
rect 22468 20334 22520 20340
rect 22192 20324 22244 20330
rect 22192 20266 22244 20272
rect 22008 20256 22060 20262
rect 22008 20198 22060 20204
rect 21916 18080 21968 18086
rect 21916 18022 21968 18028
rect 21928 15570 21956 18022
rect 22020 16250 22048 20198
rect 22204 17746 22232 20266
rect 22480 20058 22508 20334
rect 22468 20052 22520 20058
rect 22468 19994 22520 20000
rect 22376 19848 22428 19854
rect 22376 19790 22428 19796
rect 22284 18692 22336 18698
rect 22284 18634 22336 18640
rect 22296 18086 22324 18634
rect 22388 18630 22416 19790
rect 22756 19446 22784 20538
rect 23400 20466 23428 24618
rect 23952 23882 23980 26302
rect 24122 26200 24178 27000
rect 24766 26200 24822 27000
rect 25410 26330 25466 27000
rect 25240 26302 25466 26330
rect 24032 24336 24084 24342
rect 24032 24278 24084 24284
rect 23768 23854 23980 23882
rect 23768 23662 23796 23854
rect 23952 23798 23980 23854
rect 23848 23792 23900 23798
rect 23848 23734 23900 23740
rect 23940 23792 23992 23798
rect 23940 23734 23992 23740
rect 23756 23656 23808 23662
rect 23756 23598 23808 23604
rect 23756 23316 23808 23322
rect 23756 23258 23808 23264
rect 23480 22568 23532 22574
rect 23480 22510 23532 22516
rect 23492 21185 23520 22510
rect 23768 22234 23796 23258
rect 23756 22228 23808 22234
rect 23756 22170 23808 22176
rect 23572 22092 23624 22098
rect 23572 22034 23624 22040
rect 23584 21894 23612 22034
rect 23756 22024 23808 22030
rect 23756 21966 23808 21972
rect 23572 21888 23624 21894
rect 23572 21830 23624 21836
rect 23478 21176 23534 21185
rect 23478 21111 23534 21120
rect 23388 20460 23440 20466
rect 23388 20402 23440 20408
rect 23480 20460 23532 20466
rect 23480 20402 23532 20408
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 23386 20088 23442 20097
rect 23386 20023 23442 20032
rect 23400 19990 23428 20023
rect 23388 19984 23440 19990
rect 23388 19926 23440 19932
rect 22928 19712 22980 19718
rect 22928 19654 22980 19660
rect 22744 19440 22796 19446
rect 22744 19382 22796 19388
rect 22940 19378 22968 19654
rect 23492 19378 23520 20402
rect 22928 19372 22980 19378
rect 22928 19314 22980 19320
rect 23480 19372 23532 19378
rect 23480 19314 23532 19320
rect 22940 19258 22968 19314
rect 22848 19230 22968 19258
rect 22652 18828 22704 18834
rect 22652 18770 22704 18776
rect 22376 18624 22428 18630
rect 22376 18566 22428 18572
rect 22284 18080 22336 18086
rect 22284 18022 22336 18028
rect 22192 17740 22244 17746
rect 22192 17682 22244 17688
rect 22204 17338 22232 17682
rect 22192 17332 22244 17338
rect 22192 17274 22244 17280
rect 22664 17202 22692 18770
rect 22848 18358 22876 19230
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 23296 18828 23348 18834
rect 23492 18816 23520 19314
rect 23348 18788 23520 18816
rect 23296 18770 23348 18776
rect 23492 18358 23520 18788
rect 22836 18352 22888 18358
rect 22836 18294 22888 18300
rect 23480 18352 23532 18358
rect 23480 18294 23532 18300
rect 22744 18216 22796 18222
rect 22744 18158 22796 18164
rect 22652 17196 22704 17202
rect 22652 17138 22704 17144
rect 22652 17060 22704 17066
rect 22756 17048 22784 18158
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 22704 17020 22784 17048
rect 22652 17002 22704 17008
rect 22560 16992 22612 16998
rect 22560 16934 22612 16940
rect 22466 16552 22522 16561
rect 22572 16522 22600 16934
rect 22756 16726 22784 17020
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 22744 16720 22796 16726
rect 23584 16697 23612 21830
rect 23768 21162 23796 21966
rect 23860 21894 23888 23734
rect 24044 23322 24072 24278
rect 24032 23316 24084 23322
rect 24032 23258 24084 23264
rect 24030 22536 24086 22545
rect 24030 22471 24086 22480
rect 23848 21888 23900 21894
rect 23848 21830 23900 21836
rect 23768 21134 23980 21162
rect 23848 21072 23900 21078
rect 23848 21014 23900 21020
rect 23756 20392 23808 20398
rect 23756 20334 23808 20340
rect 23664 19916 23716 19922
rect 23664 19858 23716 19864
rect 23676 18902 23704 19858
rect 23664 18896 23716 18902
rect 23664 18838 23716 18844
rect 23768 18154 23796 20334
rect 23860 19514 23888 21014
rect 23952 19922 23980 21134
rect 24044 20806 24072 22471
rect 24136 20942 24164 26200
rect 24584 24744 24636 24750
rect 24584 24686 24636 24692
rect 24308 24608 24360 24614
rect 24308 24550 24360 24556
rect 24320 22778 24348 24550
rect 24596 24410 24624 24686
rect 24780 24614 24808 26200
rect 24768 24608 24820 24614
rect 24768 24550 24820 24556
rect 24584 24404 24636 24410
rect 24584 24346 24636 24352
rect 25044 24200 25096 24206
rect 25240 24188 25268 26302
rect 25410 26200 25466 26302
rect 26054 26200 26110 27000
rect 26698 26330 26754 27000
rect 26698 26302 27016 26330
rect 26698 26200 26754 26302
rect 25596 24880 25648 24886
rect 25596 24822 25648 24828
rect 25096 24160 25268 24188
rect 25044 24142 25096 24148
rect 24676 24064 24728 24070
rect 24676 24006 24728 24012
rect 24952 24064 25004 24070
rect 24952 24006 25004 24012
rect 24492 23588 24544 23594
rect 24492 23530 24544 23536
rect 24400 23112 24452 23118
rect 24400 23054 24452 23060
rect 24504 23066 24532 23530
rect 24584 23520 24636 23526
rect 24688 23497 24716 24006
rect 24964 23866 24992 24006
rect 24952 23860 25004 23866
rect 24952 23802 25004 23808
rect 24860 23656 24912 23662
rect 24860 23598 24912 23604
rect 24584 23462 24636 23468
rect 24674 23488 24730 23497
rect 24596 23254 24624 23462
rect 24674 23423 24730 23432
rect 24584 23248 24636 23254
rect 24584 23190 24636 23196
rect 24674 23080 24730 23089
rect 24216 22772 24268 22778
rect 24216 22714 24268 22720
rect 24308 22772 24360 22778
rect 24308 22714 24360 22720
rect 24228 22012 24256 22714
rect 24412 22234 24440 23054
rect 24504 23038 24624 23066
rect 24492 22976 24544 22982
rect 24492 22918 24544 22924
rect 24504 22574 24532 22918
rect 24596 22624 24624 23038
rect 24674 23015 24676 23024
rect 24728 23015 24730 23024
rect 24676 22986 24728 22992
rect 24872 22778 24900 23598
rect 25240 23322 25268 24160
rect 25412 23792 25464 23798
rect 25412 23734 25464 23740
rect 25424 23322 25452 23734
rect 25228 23316 25280 23322
rect 25228 23258 25280 23264
rect 25412 23316 25464 23322
rect 25412 23258 25464 23264
rect 25504 23248 25556 23254
rect 25504 23190 25556 23196
rect 25320 23112 25372 23118
rect 25320 23054 25372 23060
rect 25136 22976 25188 22982
rect 25136 22918 25188 22924
rect 24860 22772 24912 22778
rect 24860 22714 24912 22720
rect 24872 22642 24900 22714
rect 25148 22710 25176 22918
rect 25044 22704 25096 22710
rect 25044 22646 25096 22652
rect 25136 22704 25188 22710
rect 25136 22646 25188 22652
rect 24860 22636 24912 22642
rect 24596 22596 24716 22624
rect 24492 22568 24544 22574
rect 24492 22510 24544 22516
rect 24584 22500 24636 22506
rect 24584 22442 24636 22448
rect 24400 22228 24452 22234
rect 24400 22170 24452 22176
rect 24596 22098 24624 22442
rect 24584 22092 24636 22098
rect 24584 22034 24636 22040
rect 24228 21984 24532 22012
rect 24124 20936 24176 20942
rect 24124 20878 24176 20884
rect 24032 20800 24084 20806
rect 24032 20742 24084 20748
rect 23940 19916 23992 19922
rect 23940 19858 23992 19864
rect 24044 19786 24072 20742
rect 24504 20398 24532 21984
rect 24688 21146 24716 22596
rect 24860 22578 24912 22584
rect 24952 22024 25004 22030
rect 24952 21966 25004 21972
rect 24768 21956 24820 21962
rect 24768 21898 24820 21904
rect 24780 21418 24808 21898
rect 24860 21888 24912 21894
rect 24860 21830 24912 21836
rect 24768 21412 24820 21418
rect 24768 21354 24820 21360
rect 24676 21140 24728 21146
rect 24676 21082 24728 21088
rect 24688 20534 24716 21082
rect 24872 21049 24900 21830
rect 24858 21040 24914 21049
rect 24858 20975 24914 20984
rect 24676 20528 24728 20534
rect 24676 20470 24728 20476
rect 24492 20392 24544 20398
rect 24492 20334 24544 20340
rect 24122 20224 24178 20233
rect 24122 20159 24178 20168
rect 24136 19990 24164 20159
rect 24124 19984 24176 19990
rect 24124 19926 24176 19932
rect 24032 19780 24084 19786
rect 24032 19722 24084 19728
rect 23848 19508 23900 19514
rect 23848 19450 23900 19456
rect 24032 19440 24084 19446
rect 24032 19382 24084 19388
rect 23940 18624 23992 18630
rect 23940 18566 23992 18572
rect 23756 18148 23808 18154
rect 23756 18090 23808 18096
rect 23756 17740 23808 17746
rect 23756 17682 23808 17688
rect 23664 17128 23716 17134
rect 23664 17070 23716 17076
rect 22744 16662 22796 16668
rect 23570 16688 23626 16697
rect 23570 16623 23626 16632
rect 22466 16487 22522 16496
rect 22560 16516 22612 16522
rect 22008 16244 22060 16250
rect 22008 16186 22060 16192
rect 22284 15904 22336 15910
rect 22284 15846 22336 15852
rect 21916 15564 21968 15570
rect 21916 15506 21968 15512
rect 21824 15156 21876 15162
rect 21824 15098 21876 15104
rect 21638 15056 21694 15065
rect 21638 14991 21694 15000
rect 21732 14884 21784 14890
rect 21732 14826 21784 14832
rect 21744 14482 21772 14826
rect 21822 14512 21878 14521
rect 21732 14476 21784 14482
rect 21822 14447 21878 14456
rect 21732 14418 21784 14424
rect 21730 14376 21786 14385
rect 21730 14311 21786 14320
rect 21560 13824 21680 13852
rect 21456 13388 21508 13394
rect 21508 13348 21588 13376
rect 21456 13330 21508 13336
rect 21088 13184 21140 13190
rect 21364 13184 21416 13190
rect 21088 13126 21140 13132
rect 21284 13132 21364 13138
rect 21284 13126 21416 13132
rect 20996 12912 21048 12918
rect 20996 12854 21048 12860
rect 20904 12776 20956 12782
rect 20904 12718 20956 12724
rect 21100 12594 21128 13126
rect 21284 13110 21404 13126
rect 21180 12776 21232 12782
rect 21180 12718 21232 12724
rect 20916 12566 21128 12594
rect 20916 12434 20944 12566
rect 20916 12406 21036 12434
rect 21008 12238 21036 12406
rect 20996 12232 21048 12238
rect 20996 12174 21048 12180
rect 20812 11620 20864 11626
rect 20812 11562 20864 11568
rect 20810 11112 20866 11121
rect 20810 11047 20812 11056
rect 20864 11047 20866 11056
rect 20812 11018 20864 11024
rect 20812 10600 20864 10606
rect 20812 10542 20864 10548
rect 20824 9994 20852 10542
rect 20812 9988 20864 9994
rect 20812 9930 20864 9936
rect 20824 9704 20852 9930
rect 20904 9716 20956 9722
rect 20824 9676 20904 9704
rect 20904 9658 20956 9664
rect 20536 7540 20588 7546
rect 20536 7482 20588 7488
rect 19248 6792 19300 6798
rect 19248 6734 19300 6740
rect 19156 6656 19208 6662
rect 19156 6598 19208 6604
rect 18880 5228 18932 5234
rect 18880 5170 18932 5176
rect 19064 5160 19116 5166
rect 19064 5102 19116 5108
rect 19076 4554 19104 5102
rect 19168 4690 19196 6598
rect 19616 6112 19668 6118
rect 19616 6054 19668 6060
rect 19340 5704 19392 5710
rect 19340 5646 19392 5652
rect 19156 4684 19208 4690
rect 19156 4626 19208 4632
rect 19064 4548 19116 4554
rect 19064 4490 19116 4496
rect 17960 4004 18012 4010
rect 17960 3946 18012 3952
rect 18328 4004 18380 4010
rect 18328 3946 18380 3952
rect 17972 3534 18000 3946
rect 17960 3528 18012 3534
rect 17960 3470 18012 3476
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 19076 3126 19104 4490
rect 19352 4486 19380 5646
rect 19524 4616 19576 4622
rect 19524 4558 19576 4564
rect 19340 4480 19392 4486
rect 19340 4422 19392 4428
rect 16672 3120 16724 3126
rect 16672 3062 16724 3068
rect 19064 3120 19116 3126
rect 19064 3062 19116 3068
rect 13820 3052 13872 3058
rect 13820 2994 13872 3000
rect 18420 2984 18472 2990
rect 18420 2926 18472 2932
rect 15844 2916 15896 2922
rect 15844 2858 15896 2864
rect 13544 2644 13596 2650
rect 13544 2586 13596 2592
rect 13820 2508 13872 2514
rect 13820 2450 13872 2456
rect 12808 2440 12860 2446
rect 12808 2382 12860 2388
rect 12716 2304 12768 2310
rect 12716 2246 12768 2252
rect 13832 800 13860 2450
rect 15856 2446 15884 2858
rect 15844 2440 15896 2446
rect 15844 2382 15896 2388
rect 15936 2372 15988 2378
rect 15936 2314 15988 2320
rect 15948 800 15976 2314
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 18064 870 18184 898
rect 18064 800 18092 870
rect 1122 0 1178 800
rect 3238 0 3294 800
rect 5354 0 5410 800
rect 7470 0 7526 800
rect 9586 0 9642 800
rect 11702 0 11758 800
rect 13818 0 13874 800
rect 15934 0 15990 800
rect 18050 0 18106 800
rect 18156 762 18184 870
rect 18432 762 18460 2926
rect 19536 2446 19564 4558
rect 19628 2446 19656 6054
rect 20812 5024 20864 5030
rect 20812 4966 20864 4972
rect 20824 3058 20852 4966
rect 21008 4758 21036 12174
rect 21192 11558 21220 12718
rect 21284 12102 21312 13110
rect 21364 12776 21416 12782
rect 21364 12718 21416 12724
rect 21272 12096 21324 12102
rect 21272 12038 21324 12044
rect 21180 11552 21232 11558
rect 21180 11494 21232 11500
rect 21180 11076 21232 11082
rect 21180 11018 21232 11024
rect 21192 9994 21220 11018
rect 21284 10033 21312 12038
rect 21376 11762 21404 12718
rect 21456 12640 21508 12646
rect 21456 12582 21508 12588
rect 21468 12306 21496 12582
rect 21456 12300 21508 12306
rect 21456 12242 21508 12248
rect 21364 11756 21416 11762
rect 21364 11698 21416 11704
rect 21456 11688 21508 11694
rect 21456 11630 21508 11636
rect 21468 11218 21496 11630
rect 21560 11626 21588 13348
rect 21652 12753 21680 13824
rect 21638 12744 21694 12753
rect 21638 12679 21694 12688
rect 21744 12170 21772 14311
rect 21836 13190 21864 14447
rect 22296 13870 22324 15846
rect 22480 15706 22508 16487
rect 22560 16458 22612 16464
rect 22836 16516 22888 16522
rect 22836 16458 22888 16464
rect 22652 16448 22704 16454
rect 22652 16390 22704 16396
rect 22468 15700 22520 15706
rect 22468 15642 22520 15648
rect 22664 15162 22692 16390
rect 22744 16040 22796 16046
rect 22744 15982 22796 15988
rect 22652 15156 22704 15162
rect 22652 15098 22704 15104
rect 22652 14340 22704 14346
rect 22652 14282 22704 14288
rect 22376 14272 22428 14278
rect 22376 14214 22428 14220
rect 22388 14074 22416 14214
rect 22664 14074 22692 14282
rect 22376 14068 22428 14074
rect 22376 14010 22428 14016
rect 22652 14068 22704 14074
rect 22652 14010 22704 14016
rect 22008 13864 22060 13870
rect 22008 13806 22060 13812
rect 22284 13864 22336 13870
rect 22284 13806 22336 13812
rect 21824 13184 21876 13190
rect 21824 13126 21876 13132
rect 21824 12980 21876 12986
rect 21824 12922 21876 12928
rect 21732 12164 21784 12170
rect 21732 12106 21784 12112
rect 21640 12096 21692 12102
rect 21640 12038 21692 12044
rect 21652 11762 21680 12038
rect 21640 11756 21692 11762
rect 21640 11698 21692 11704
rect 21548 11620 21600 11626
rect 21548 11562 21600 11568
rect 21732 11620 21784 11626
rect 21732 11562 21784 11568
rect 21640 11552 21692 11558
rect 21640 11494 21692 11500
rect 21652 11234 21680 11494
rect 21744 11354 21772 11562
rect 21732 11348 21784 11354
rect 21732 11290 21784 11296
rect 21652 11218 21772 11234
rect 21456 11212 21508 11218
rect 21652 11212 21784 11218
rect 21652 11206 21732 11212
rect 21456 11154 21508 11160
rect 21732 11154 21784 11160
rect 21456 10668 21508 10674
rect 21456 10610 21508 10616
rect 21270 10024 21326 10033
rect 21180 9988 21232 9994
rect 21270 9959 21326 9968
rect 21180 9930 21232 9936
rect 21192 9722 21220 9930
rect 21180 9716 21232 9722
rect 21180 9658 21232 9664
rect 21468 9654 21496 10610
rect 21548 10600 21600 10606
rect 21548 10542 21600 10548
rect 21560 10130 21588 10542
rect 21836 10538 21864 12922
rect 21916 12844 21968 12850
rect 21916 12786 21968 12792
rect 21824 10532 21876 10538
rect 21824 10474 21876 10480
rect 21640 10260 21692 10266
rect 21640 10202 21692 10208
rect 21548 10124 21600 10130
rect 21548 10066 21600 10072
rect 21652 10010 21680 10202
rect 21560 9982 21680 10010
rect 21560 9926 21588 9982
rect 21836 9926 21864 10474
rect 21548 9920 21600 9926
rect 21548 9862 21600 9868
rect 21824 9920 21876 9926
rect 21824 9862 21876 9868
rect 21732 9716 21784 9722
rect 21732 9658 21784 9664
rect 21456 9648 21508 9654
rect 21456 9590 21508 9596
rect 21088 9580 21140 9586
rect 21088 9522 21140 9528
rect 21100 9382 21128 9522
rect 21744 9382 21772 9658
rect 21088 9376 21140 9382
rect 21088 9318 21140 9324
rect 21732 9376 21784 9382
rect 21732 9318 21784 9324
rect 21100 8906 21128 9318
rect 21088 8900 21140 8906
rect 21088 8842 21140 8848
rect 21100 8498 21128 8842
rect 21088 8492 21140 8498
rect 21088 8434 21140 8440
rect 21100 7818 21128 8434
rect 21928 8090 21956 12786
rect 22020 11694 22048 13806
rect 22100 12776 22152 12782
rect 22100 12718 22152 12724
rect 22112 12306 22140 12718
rect 22296 12458 22324 13806
rect 22650 13016 22706 13025
rect 22756 12986 22784 15982
rect 22848 15978 22876 16458
rect 23296 16448 23348 16454
rect 23296 16390 23348 16396
rect 23388 16448 23440 16454
rect 23388 16390 23440 16396
rect 23308 16153 23336 16390
rect 23294 16144 23350 16153
rect 23294 16079 23350 16088
rect 22836 15972 22888 15978
rect 22836 15914 22888 15920
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 23296 15020 23348 15026
rect 23296 14962 23348 14968
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 23204 14612 23256 14618
rect 23204 14554 23256 14560
rect 23216 14346 23244 14554
rect 23204 14340 23256 14346
rect 23204 14282 23256 14288
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 22836 13320 22888 13326
rect 22836 13262 22888 13268
rect 22650 12951 22706 12960
rect 22744 12980 22796 12986
rect 22664 12481 22692 12951
rect 22744 12922 22796 12928
rect 22204 12430 22324 12458
rect 22650 12472 22706 12481
rect 22100 12300 22152 12306
rect 22100 12242 22152 12248
rect 22098 12200 22154 12209
rect 22098 12135 22154 12144
rect 22112 11762 22140 12135
rect 22204 11830 22232 12430
rect 22650 12407 22706 12416
rect 22848 12424 22876 13262
rect 23110 13016 23166 13025
rect 23110 12951 23112 12960
rect 23164 12951 23166 12960
rect 23112 12922 23164 12928
rect 23020 12844 23072 12850
rect 23020 12786 23072 12792
rect 23032 12753 23060 12786
rect 23018 12744 23074 12753
rect 23018 12679 23074 12688
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 22928 12436 22980 12442
rect 22848 12396 22928 12424
rect 22928 12378 22980 12384
rect 22652 12300 22704 12306
rect 22652 12242 22704 12248
rect 22558 12200 22614 12209
rect 22558 12135 22614 12144
rect 22572 12102 22600 12135
rect 22468 12096 22520 12102
rect 22468 12038 22520 12044
rect 22560 12096 22612 12102
rect 22560 12038 22612 12044
rect 22192 11824 22244 11830
rect 22192 11766 22244 11772
rect 22100 11756 22152 11762
rect 22100 11698 22152 11704
rect 22008 11688 22060 11694
rect 22008 11630 22060 11636
rect 22480 11354 22508 12038
rect 22664 11830 22692 12242
rect 23308 11880 23336 14962
rect 23400 14090 23428 16390
rect 23676 16182 23704 17070
rect 23572 16176 23624 16182
rect 23572 16118 23624 16124
rect 23664 16176 23716 16182
rect 23664 16118 23716 16124
rect 23480 15700 23532 15706
rect 23480 15642 23532 15648
rect 23492 15162 23520 15642
rect 23480 15156 23532 15162
rect 23480 15098 23532 15104
rect 23400 14062 23520 14090
rect 23492 13818 23520 14062
rect 23400 13790 23520 13818
rect 23400 13530 23428 13790
rect 23388 13524 23440 13530
rect 23388 13466 23440 13472
rect 23480 13524 23532 13530
rect 23480 13466 23532 13472
rect 23492 13410 23520 13466
rect 23400 13382 23520 13410
rect 23400 12782 23428 13382
rect 23480 12980 23532 12986
rect 23480 12922 23532 12928
rect 23388 12776 23440 12782
rect 23388 12718 23440 12724
rect 23492 12646 23520 12922
rect 23480 12640 23532 12646
rect 23480 12582 23532 12588
rect 23584 12374 23612 16118
rect 23768 15162 23796 17682
rect 23952 17678 23980 18566
rect 24044 17746 24072 19382
rect 24124 18692 24176 18698
rect 24124 18634 24176 18640
rect 24032 17740 24084 17746
rect 24032 17682 24084 17688
rect 23940 17672 23992 17678
rect 23940 17614 23992 17620
rect 23952 17338 23980 17614
rect 23940 17332 23992 17338
rect 23940 17274 23992 17280
rect 24032 17196 24084 17202
rect 24136 17184 24164 18634
rect 24400 18624 24452 18630
rect 24400 18566 24452 18572
rect 24412 17610 24440 18566
rect 24400 17604 24452 17610
rect 24400 17546 24452 17552
rect 24084 17156 24164 17184
rect 24032 17138 24084 17144
rect 23940 16788 23992 16794
rect 23940 16730 23992 16736
rect 23952 15570 23980 16730
rect 24044 16454 24072 17138
rect 24032 16448 24084 16454
rect 24032 16390 24084 16396
rect 24044 15978 24072 16390
rect 24124 16040 24176 16046
rect 24124 15982 24176 15988
rect 24032 15972 24084 15978
rect 24032 15914 24084 15920
rect 23848 15564 23900 15570
rect 23848 15506 23900 15512
rect 23940 15564 23992 15570
rect 23940 15506 23992 15512
rect 23756 15156 23808 15162
rect 23756 15098 23808 15104
rect 23664 14272 23716 14278
rect 23664 14214 23716 14220
rect 23676 13326 23704 14214
rect 23860 14074 23888 15506
rect 24044 14618 24072 15914
rect 24032 14612 24084 14618
rect 24032 14554 24084 14560
rect 23848 14068 23900 14074
rect 23848 14010 23900 14016
rect 23860 13734 23888 14010
rect 24044 14006 24072 14554
rect 24032 14000 24084 14006
rect 24032 13942 24084 13948
rect 23848 13728 23900 13734
rect 23848 13670 23900 13676
rect 24136 13530 24164 15982
rect 24308 14884 24360 14890
rect 24308 14826 24360 14832
rect 24216 13864 24268 13870
rect 24216 13806 24268 13812
rect 24124 13524 24176 13530
rect 24124 13466 24176 13472
rect 23756 13388 23808 13394
rect 23756 13330 23808 13336
rect 23664 13320 23716 13326
rect 23664 13262 23716 13268
rect 23664 13184 23716 13190
rect 23664 13126 23716 13132
rect 23572 12368 23624 12374
rect 23572 12310 23624 12316
rect 23572 12232 23624 12238
rect 23572 12174 23624 12180
rect 23308 11852 23428 11880
rect 22652 11824 22704 11830
rect 22652 11766 22704 11772
rect 22560 11756 22612 11762
rect 22560 11698 22612 11704
rect 22572 11354 22600 11698
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 22008 11348 22060 11354
rect 22008 11290 22060 11296
rect 22468 11348 22520 11354
rect 22468 11290 22520 11296
rect 22560 11348 22612 11354
rect 22560 11290 22612 11296
rect 22020 11121 22048 11290
rect 22006 11112 22062 11121
rect 22006 11047 22062 11056
rect 22284 10736 22336 10742
rect 22284 10678 22336 10684
rect 22008 10600 22060 10606
rect 22008 10542 22060 10548
rect 22020 10130 22048 10542
rect 22100 10464 22152 10470
rect 22100 10406 22152 10412
rect 22008 10124 22060 10130
rect 22008 10066 22060 10072
rect 22020 9042 22048 10066
rect 22008 9036 22060 9042
rect 22008 8978 22060 8984
rect 22020 8498 22048 8978
rect 22112 8906 22140 10406
rect 22296 9722 22324 10678
rect 22572 10062 22600 11290
rect 23400 11286 23428 11852
rect 23480 11688 23532 11694
rect 23480 11630 23532 11636
rect 23388 11280 23440 11286
rect 23388 11222 23440 11228
rect 23492 11150 23520 11630
rect 23584 11626 23612 12174
rect 23572 11620 23624 11626
rect 23572 11562 23624 11568
rect 23480 11144 23532 11150
rect 23480 11086 23532 11092
rect 22652 11008 22704 11014
rect 22652 10950 22704 10956
rect 22664 10810 22692 10950
rect 22652 10804 22704 10810
rect 22652 10746 22704 10752
rect 23388 10668 23440 10674
rect 23388 10610 23440 10616
rect 22836 10600 22888 10606
rect 22836 10542 22888 10548
rect 22848 10266 22876 10542
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 22836 10260 22888 10266
rect 22836 10202 22888 10208
rect 23400 10198 23428 10610
rect 23388 10192 23440 10198
rect 23388 10134 23440 10140
rect 22560 10056 22612 10062
rect 22466 10024 22522 10033
rect 22560 9998 22612 10004
rect 22466 9959 22522 9968
rect 22284 9716 22336 9722
rect 22284 9658 22336 9664
rect 22100 8900 22152 8906
rect 22100 8842 22152 8848
rect 22112 8634 22140 8842
rect 22376 8832 22428 8838
rect 22376 8774 22428 8780
rect 22100 8628 22152 8634
rect 22100 8570 22152 8576
rect 22008 8492 22060 8498
rect 22008 8434 22060 8440
rect 21916 8084 21968 8090
rect 21916 8026 21968 8032
rect 21088 7812 21140 7818
rect 21088 7754 21140 7760
rect 21456 7744 21508 7750
rect 21456 7686 21508 7692
rect 21468 7206 21496 7686
rect 21456 7200 21508 7206
rect 21456 7142 21508 7148
rect 21916 6656 21968 6662
rect 21916 6598 21968 6604
rect 20996 4752 21048 4758
rect 20996 4694 21048 4700
rect 21928 4690 21956 6598
rect 21916 4684 21968 4690
rect 21916 4626 21968 4632
rect 21456 4480 21508 4486
rect 21456 4422 21508 4428
rect 20996 3528 21048 3534
rect 20996 3470 21048 3476
rect 20812 3052 20864 3058
rect 20812 2994 20864 3000
rect 21008 2990 21036 3470
rect 21180 3460 21232 3466
rect 21180 3402 21232 3408
rect 21192 3194 21220 3402
rect 21180 3188 21232 3194
rect 21180 3130 21232 3136
rect 20996 2984 21048 2990
rect 20996 2926 21048 2932
rect 21192 2854 21220 3130
rect 21468 3058 21496 4422
rect 21456 3052 21508 3058
rect 21456 2994 21508 3000
rect 22020 2990 22048 8434
rect 22388 7886 22416 8774
rect 22376 7880 22428 7886
rect 22376 7822 22428 7828
rect 22284 7744 22336 7750
rect 22284 7686 22336 7692
rect 22100 4616 22152 4622
rect 22100 4558 22152 4564
rect 22112 4214 22140 4558
rect 22100 4208 22152 4214
rect 22100 4150 22152 4156
rect 22112 3126 22140 4150
rect 22100 3120 22152 3126
rect 22100 3062 22152 3068
rect 22008 2984 22060 2990
rect 22008 2926 22060 2932
rect 21180 2848 21232 2854
rect 21180 2790 21232 2796
rect 22296 2650 22324 7686
rect 22480 7546 22508 9959
rect 22652 9580 22704 9586
rect 22652 9522 22704 9528
rect 22560 9444 22612 9450
rect 22560 9386 22612 9392
rect 22572 9042 22600 9386
rect 22664 9042 22692 9522
rect 23400 9382 23428 10134
rect 23492 9586 23520 11086
rect 23584 10452 23612 11562
rect 23676 10810 23704 13126
rect 23664 10804 23716 10810
rect 23664 10746 23716 10752
rect 23664 10464 23716 10470
rect 23584 10424 23664 10452
rect 23664 10406 23716 10412
rect 23480 9580 23532 9586
rect 23480 9522 23532 9528
rect 23388 9376 23440 9382
rect 23388 9318 23440 9324
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 22560 9036 22612 9042
rect 22560 8978 22612 8984
rect 22652 9036 22704 9042
rect 22652 8978 22704 8984
rect 22664 8378 22692 8978
rect 22572 8350 22692 8378
rect 22468 7540 22520 7546
rect 22468 7482 22520 7488
rect 22468 7200 22520 7206
rect 22468 7142 22520 7148
rect 22480 3652 22508 7142
rect 22572 6186 22600 8350
rect 22652 8288 22704 8294
rect 22652 8230 22704 8236
rect 22664 7342 22692 8230
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 23676 7954 23704 10406
rect 23768 10266 23796 13330
rect 24032 13252 24084 13258
rect 24032 13194 24084 13200
rect 23848 12980 23900 12986
rect 24044 12968 24072 13194
rect 23900 12940 24072 12968
rect 23848 12922 23900 12928
rect 23848 12776 23900 12782
rect 23848 12718 23900 12724
rect 23860 11694 23888 12718
rect 23848 11688 23900 11694
rect 23848 11630 23900 11636
rect 23848 11212 23900 11218
rect 23848 11154 23900 11160
rect 23860 11121 23888 11154
rect 23846 11112 23902 11121
rect 23846 11047 23902 11056
rect 23940 10600 23992 10606
rect 23940 10542 23992 10548
rect 23756 10260 23808 10266
rect 23756 10202 23808 10208
rect 23768 9654 23796 10202
rect 23848 10192 23900 10198
rect 23848 10134 23900 10140
rect 23756 9648 23808 9654
rect 23756 9590 23808 9596
rect 23860 9518 23888 10134
rect 23952 9926 23980 10542
rect 23940 9920 23992 9926
rect 23940 9862 23992 9868
rect 23848 9512 23900 9518
rect 23848 9454 23900 9460
rect 23860 8906 23888 9454
rect 23848 8900 23900 8906
rect 23848 8842 23900 8848
rect 23860 8634 23888 8842
rect 23848 8628 23900 8634
rect 23848 8570 23900 8576
rect 23664 7948 23716 7954
rect 23664 7890 23716 7896
rect 22652 7336 22704 7342
rect 22652 7278 22704 7284
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 22560 6180 22612 6186
rect 22560 6122 22612 6128
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 23952 5710 23980 9862
rect 23940 5704 23992 5710
rect 23940 5646 23992 5652
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 24044 4706 24072 12940
rect 24124 12776 24176 12782
rect 24124 12718 24176 12724
rect 24136 11218 24164 12718
rect 24124 11212 24176 11218
rect 24124 11154 24176 11160
rect 24122 11112 24178 11121
rect 24228 11082 24256 13806
rect 24320 12238 24348 14826
rect 24412 14385 24440 17546
rect 24504 15994 24532 20334
rect 24688 19990 24716 20470
rect 24676 19984 24728 19990
rect 24728 19944 24808 19972
rect 24676 19926 24728 19932
rect 24780 19446 24808 19944
rect 24768 19440 24820 19446
rect 24768 19382 24820 19388
rect 24780 18698 24808 19382
rect 24768 18692 24820 18698
rect 24768 18634 24820 18640
rect 24676 18284 24728 18290
rect 24676 18226 24728 18232
rect 24688 17882 24716 18226
rect 24676 17876 24728 17882
rect 24676 17818 24728 17824
rect 24584 16652 24636 16658
rect 24584 16594 24636 16600
rect 24596 16114 24624 16594
rect 24688 16522 24716 17818
rect 24768 17536 24820 17542
rect 24768 17478 24820 17484
rect 24860 17536 24912 17542
rect 24860 17478 24912 17484
rect 24780 17270 24808 17478
rect 24768 17264 24820 17270
rect 24768 17206 24820 17212
rect 24676 16516 24728 16522
rect 24676 16458 24728 16464
rect 24872 16250 24900 17478
rect 24964 17338 24992 21966
rect 25056 21894 25084 22646
rect 25134 22128 25190 22137
rect 25134 22063 25136 22072
rect 25188 22063 25190 22072
rect 25136 22034 25188 22040
rect 25332 22030 25360 23054
rect 25320 22024 25372 22030
rect 25320 21966 25372 21972
rect 25044 21888 25096 21894
rect 25044 21830 25096 21836
rect 25056 21622 25084 21830
rect 25044 21616 25096 21622
rect 25044 21558 25096 21564
rect 25228 21480 25280 21486
rect 25226 21448 25228 21457
rect 25320 21480 25372 21486
rect 25280 21448 25282 21457
rect 25320 21422 25372 21428
rect 25226 21383 25282 21392
rect 25332 20641 25360 21422
rect 25412 21344 25464 21350
rect 25412 21286 25464 21292
rect 25318 20632 25374 20641
rect 25318 20567 25374 20576
rect 25424 20330 25452 21286
rect 25516 20534 25544 23190
rect 25608 22545 25636 24822
rect 25872 24812 25924 24818
rect 25872 24754 25924 24760
rect 25884 24206 25912 24754
rect 25964 24404 26016 24410
rect 25964 24346 26016 24352
rect 25976 24313 26004 24346
rect 25962 24304 26018 24313
rect 25962 24239 26018 24248
rect 26068 24206 26096 26200
rect 26700 24676 26752 24682
rect 26700 24618 26752 24624
rect 25872 24200 25924 24206
rect 25872 24142 25924 24148
rect 26056 24200 26108 24206
rect 26056 24142 26108 24148
rect 26146 24168 26202 24177
rect 26146 24103 26202 24112
rect 26160 24070 26188 24103
rect 26148 24064 26200 24070
rect 26148 24006 26200 24012
rect 26240 24064 26292 24070
rect 26240 24006 26292 24012
rect 26424 24064 26476 24070
rect 26424 24006 26476 24012
rect 26252 23882 26280 24006
rect 26160 23866 26280 23882
rect 26148 23860 26280 23866
rect 26200 23854 26280 23860
rect 26148 23802 26200 23808
rect 25688 23112 25740 23118
rect 25688 23054 25740 23060
rect 25594 22536 25650 22545
rect 25594 22471 25650 22480
rect 25596 21004 25648 21010
rect 25596 20946 25648 20952
rect 25504 20528 25556 20534
rect 25504 20470 25556 20476
rect 25412 20324 25464 20330
rect 25412 20266 25464 20272
rect 25504 20256 25556 20262
rect 25504 20198 25556 20204
rect 25412 19916 25464 19922
rect 25412 19858 25464 19864
rect 25228 19780 25280 19786
rect 25228 19722 25280 19728
rect 25240 19446 25268 19722
rect 25318 19544 25374 19553
rect 25318 19479 25374 19488
rect 25228 19440 25280 19446
rect 25228 19382 25280 19388
rect 25136 19304 25188 19310
rect 25136 19246 25188 19252
rect 25148 18970 25176 19246
rect 25228 19168 25280 19174
rect 25228 19110 25280 19116
rect 25136 18964 25188 18970
rect 25136 18906 25188 18912
rect 25042 18728 25098 18737
rect 25240 18698 25268 19110
rect 25042 18663 25044 18672
rect 25096 18663 25098 18672
rect 25228 18692 25280 18698
rect 25044 18634 25096 18640
rect 25228 18634 25280 18640
rect 25134 18320 25190 18329
rect 25044 18284 25096 18290
rect 25134 18255 25136 18264
rect 25044 18226 25096 18232
rect 25188 18255 25190 18264
rect 25136 18226 25188 18232
rect 25056 18193 25084 18226
rect 25332 18222 25360 19479
rect 25320 18216 25372 18222
rect 25042 18184 25098 18193
rect 25320 18158 25372 18164
rect 25042 18119 25098 18128
rect 25044 18080 25096 18086
rect 25044 18022 25096 18028
rect 25056 17746 25084 18022
rect 25044 17740 25096 17746
rect 25044 17682 25096 17688
rect 24952 17332 25004 17338
rect 24952 17274 25004 17280
rect 25424 17241 25452 19858
rect 25516 19378 25544 20198
rect 25504 19372 25556 19378
rect 25504 19314 25556 19320
rect 25504 18148 25556 18154
rect 25504 18090 25556 18096
rect 25410 17232 25466 17241
rect 25228 17196 25280 17202
rect 25410 17167 25466 17176
rect 25228 17138 25280 17144
rect 25136 17128 25188 17134
rect 25136 17070 25188 17076
rect 25044 16448 25096 16454
rect 25044 16390 25096 16396
rect 24860 16244 24912 16250
rect 24860 16186 24912 16192
rect 24584 16108 24636 16114
rect 24584 16050 24636 16056
rect 24504 15966 24716 15994
rect 24688 14958 24716 15966
rect 25056 15570 25084 16390
rect 25044 15564 25096 15570
rect 25044 15506 25096 15512
rect 25056 15094 25084 15506
rect 25044 15088 25096 15094
rect 25044 15030 25096 15036
rect 24584 14952 24636 14958
rect 24584 14894 24636 14900
rect 24676 14952 24728 14958
rect 24676 14894 24728 14900
rect 24768 14952 24820 14958
rect 24768 14894 24820 14900
rect 24596 14550 24624 14894
rect 24584 14544 24636 14550
rect 24584 14486 24636 14492
rect 24398 14376 24454 14385
rect 24398 14311 24454 14320
rect 24596 14278 24624 14486
rect 24400 14272 24452 14278
rect 24584 14272 24636 14278
rect 24400 14214 24452 14220
rect 24582 14240 24584 14249
rect 24636 14240 24638 14249
rect 24412 13258 24440 14214
rect 24582 14175 24638 14184
rect 24400 13252 24452 13258
rect 24400 13194 24452 13200
rect 24492 13184 24544 13190
rect 24492 13126 24544 13132
rect 24504 12889 24532 13126
rect 24780 12986 24808 14894
rect 25044 14816 25096 14822
rect 25044 14758 25096 14764
rect 24860 14476 24912 14482
rect 24860 14418 24912 14424
rect 24872 13938 24900 14418
rect 24952 14272 25004 14278
rect 24952 14214 25004 14220
rect 24860 13932 24912 13938
rect 24860 13874 24912 13880
rect 24964 13326 24992 14214
rect 24952 13320 25004 13326
rect 24952 13262 25004 13268
rect 25056 12986 25084 14758
rect 25148 14618 25176 17070
rect 25136 14612 25188 14618
rect 25136 14554 25188 14560
rect 25148 14006 25176 14554
rect 25136 14000 25188 14006
rect 25136 13942 25188 13948
rect 25240 13530 25268 17138
rect 25516 16726 25544 18090
rect 25608 17814 25636 20946
rect 25700 20602 25728 23054
rect 26160 22094 26188 23802
rect 26436 23798 26464 24006
rect 26516 23860 26568 23866
rect 26516 23802 26568 23808
rect 26424 23792 26476 23798
rect 26424 23734 26476 23740
rect 26330 23488 26386 23497
rect 26330 23423 26386 23432
rect 26344 22094 26372 23423
rect 26436 23050 26464 23734
rect 26528 23526 26556 23802
rect 26712 23526 26740 24618
rect 26988 23798 27016 26302
rect 27342 26200 27398 27000
rect 27986 26200 28042 27000
rect 28630 26200 28686 27000
rect 29274 26200 29330 27000
rect 29918 26200 29974 27000
rect 30562 26200 30618 27000
rect 30656 26376 30708 26382
rect 30656 26318 30708 26324
rect 27252 24336 27304 24342
rect 27252 24278 27304 24284
rect 27160 24132 27212 24138
rect 27160 24074 27212 24080
rect 26976 23792 27028 23798
rect 26976 23734 27028 23740
rect 26516 23520 26568 23526
rect 26516 23462 26568 23468
rect 26608 23520 26660 23526
rect 26608 23462 26660 23468
rect 26700 23520 26752 23526
rect 26700 23462 26752 23468
rect 26620 23186 26648 23462
rect 26608 23180 26660 23186
rect 26608 23122 26660 23128
rect 26700 23180 26752 23186
rect 26700 23122 26752 23128
rect 26424 23044 26476 23050
rect 26424 22986 26476 22992
rect 26436 22710 26464 22986
rect 26424 22704 26476 22710
rect 26424 22646 26476 22652
rect 26712 22522 26740 23122
rect 26436 22494 26740 22522
rect 27172 22506 27200 24074
rect 27160 22500 27212 22506
rect 26436 22098 26464 22494
rect 27160 22442 27212 22448
rect 26608 22432 26660 22438
rect 26608 22374 26660 22380
rect 26620 22166 26648 22374
rect 27264 22216 27292 24278
rect 27356 24274 27384 26200
rect 28000 24750 28028 26200
rect 27988 24744 28040 24750
rect 27988 24686 28040 24692
rect 28644 24342 28672 26200
rect 29184 24744 29236 24750
rect 29184 24686 29236 24692
rect 29092 24676 29144 24682
rect 29092 24618 29144 24624
rect 28632 24336 28684 24342
rect 28632 24278 28684 24284
rect 27344 24268 27396 24274
rect 27344 24210 27396 24216
rect 27344 24064 27396 24070
rect 27342 24032 27344 24041
rect 28632 24064 28684 24070
rect 27396 24032 27398 24041
rect 28632 24006 28684 24012
rect 27342 23967 27398 23976
rect 27950 23964 28258 23973
rect 27950 23962 27956 23964
rect 28012 23962 28036 23964
rect 28092 23962 28116 23964
rect 28172 23962 28196 23964
rect 28252 23962 28258 23964
rect 28012 23910 28014 23962
rect 28194 23910 28196 23962
rect 27950 23908 27956 23910
rect 28012 23908 28036 23910
rect 28092 23908 28116 23910
rect 28172 23908 28196 23910
rect 28252 23908 28258 23910
rect 27950 23899 28258 23908
rect 27988 23724 28040 23730
rect 27988 23666 28040 23672
rect 27804 23656 27856 23662
rect 27804 23598 27856 23604
rect 27620 23520 27672 23526
rect 27620 23462 27672 23468
rect 27712 23520 27764 23526
rect 27712 23462 27764 23468
rect 27528 23248 27580 23254
rect 27528 23190 27580 23196
rect 27540 22710 27568 23190
rect 27632 23118 27660 23462
rect 27620 23112 27672 23118
rect 27620 23054 27672 23060
rect 27528 22704 27580 22710
rect 27528 22646 27580 22652
rect 27344 22636 27396 22642
rect 27344 22578 27396 22584
rect 27172 22188 27292 22216
rect 26608 22160 26660 22166
rect 26608 22102 26660 22108
rect 27068 22160 27120 22166
rect 27068 22102 27120 22108
rect 26068 22066 26188 22094
rect 26252 22066 26372 22094
rect 26424 22092 26476 22098
rect 25778 21992 25834 22001
rect 25778 21927 25780 21936
rect 25832 21927 25834 21936
rect 25780 21898 25832 21904
rect 25964 21888 26016 21894
rect 25964 21830 26016 21836
rect 25872 21548 25924 21554
rect 25872 21490 25924 21496
rect 25884 21350 25912 21490
rect 25872 21344 25924 21350
rect 25872 21286 25924 21292
rect 25780 20936 25832 20942
rect 25780 20878 25832 20884
rect 25688 20596 25740 20602
rect 25688 20538 25740 20544
rect 25700 18834 25728 20538
rect 25792 20398 25820 20878
rect 25780 20392 25832 20398
rect 25780 20334 25832 20340
rect 25792 19514 25820 20334
rect 25884 19961 25912 21286
rect 25976 20874 26004 21830
rect 25964 20868 26016 20874
rect 25964 20810 26016 20816
rect 25870 19952 25926 19961
rect 26068 19922 26096 22066
rect 26252 21978 26280 22066
rect 26424 22034 26476 22040
rect 26160 21962 26648 21978
rect 26148 21956 26648 21962
rect 26200 21950 26648 21956
rect 26148 21898 26200 21904
rect 26516 21888 26568 21894
rect 26252 21848 26516 21876
rect 26146 21448 26202 21457
rect 26146 21383 26202 21392
rect 26160 21350 26188 21383
rect 26148 21344 26200 21350
rect 26148 21286 26200 21292
rect 25870 19887 25926 19896
rect 26056 19916 26108 19922
rect 26056 19858 26108 19864
rect 26148 19916 26200 19922
rect 26148 19858 26200 19864
rect 26054 19816 26110 19825
rect 25872 19780 25924 19786
rect 26054 19751 26110 19760
rect 25872 19722 25924 19728
rect 25780 19508 25832 19514
rect 25780 19450 25832 19456
rect 25780 19168 25832 19174
rect 25780 19110 25832 19116
rect 25688 18828 25740 18834
rect 25688 18770 25740 18776
rect 25792 18426 25820 19110
rect 25884 18873 25912 19722
rect 26068 19718 26096 19751
rect 25964 19712 26016 19718
rect 25964 19654 26016 19660
rect 26056 19712 26108 19718
rect 26056 19654 26108 19660
rect 25976 19514 26004 19654
rect 26160 19553 26188 19858
rect 26146 19544 26202 19553
rect 25964 19508 26016 19514
rect 26146 19479 26202 19488
rect 25964 19450 26016 19456
rect 25976 19378 26188 19394
rect 25964 19372 26188 19378
rect 26016 19366 26188 19372
rect 25964 19314 26016 19320
rect 26054 19136 26110 19145
rect 26054 19071 26110 19080
rect 25870 18864 25926 18873
rect 25870 18799 25926 18808
rect 25780 18420 25832 18426
rect 25780 18362 25832 18368
rect 25962 18320 26018 18329
rect 25962 18255 26018 18264
rect 25596 17808 25648 17814
rect 25596 17750 25648 17756
rect 25596 17672 25648 17678
rect 25596 17614 25648 17620
rect 25504 16720 25556 16726
rect 25504 16662 25556 16668
rect 25608 16658 25636 17614
rect 25976 17270 26004 18255
rect 25964 17264 26016 17270
rect 25964 17206 26016 17212
rect 25872 17060 25924 17066
rect 25872 17002 25924 17008
rect 25884 16658 25912 17002
rect 25976 16998 26004 17206
rect 25964 16992 26016 16998
rect 25964 16934 26016 16940
rect 25596 16652 25648 16658
rect 25596 16594 25648 16600
rect 25872 16652 25924 16658
rect 25872 16594 25924 16600
rect 25884 16538 25912 16594
rect 25792 16510 25912 16538
rect 25964 16516 26016 16522
rect 25594 16144 25650 16153
rect 25594 16079 25650 16088
rect 25320 15904 25372 15910
rect 25320 15846 25372 15852
rect 25332 15570 25360 15846
rect 25320 15564 25372 15570
rect 25320 15506 25372 15512
rect 25608 15434 25636 16079
rect 25596 15428 25648 15434
rect 25596 15370 25648 15376
rect 25412 15020 25464 15026
rect 25412 14962 25464 14968
rect 25504 15020 25556 15026
rect 25504 14962 25556 14968
rect 25320 14408 25372 14414
rect 25320 14350 25372 14356
rect 25228 13524 25280 13530
rect 25228 13466 25280 13472
rect 24768 12980 24820 12986
rect 24768 12922 24820 12928
rect 25044 12980 25096 12986
rect 25044 12922 25096 12928
rect 24490 12880 24546 12889
rect 24490 12815 24546 12824
rect 25056 12434 25084 12922
rect 24964 12406 25084 12434
rect 24964 12306 24992 12406
rect 25332 12306 25360 14350
rect 24492 12300 24544 12306
rect 24492 12242 24544 12248
rect 24952 12300 25004 12306
rect 24952 12242 25004 12248
rect 25320 12300 25372 12306
rect 25320 12242 25372 12248
rect 24308 12232 24360 12238
rect 24308 12174 24360 12180
rect 24504 11898 24532 12242
rect 24584 12232 24636 12238
rect 24584 12174 24636 12180
rect 24492 11892 24544 11898
rect 24492 11834 24544 11840
rect 24308 11824 24360 11830
rect 24308 11766 24360 11772
rect 24320 11694 24348 11766
rect 24308 11688 24360 11694
rect 24308 11630 24360 11636
rect 24400 11348 24452 11354
rect 24400 11290 24452 11296
rect 24122 11047 24178 11056
rect 24216 11076 24268 11082
rect 24136 10130 24164 11047
rect 24216 11018 24268 11024
rect 24124 10124 24176 10130
rect 24124 10066 24176 10072
rect 24412 9178 24440 11290
rect 24504 11218 24532 11834
rect 24492 11212 24544 11218
rect 24492 11154 24544 11160
rect 24596 11150 24624 12174
rect 25424 11801 25452 14962
rect 25516 14550 25544 14962
rect 25608 14822 25636 15370
rect 25596 14816 25648 14822
rect 25596 14758 25648 14764
rect 25504 14544 25556 14550
rect 25504 14486 25556 14492
rect 25504 14340 25556 14346
rect 25504 14282 25556 14288
rect 25516 14074 25544 14282
rect 25504 14068 25556 14074
rect 25504 14010 25556 14016
rect 25410 11792 25466 11801
rect 25410 11727 25466 11736
rect 24584 11144 24636 11150
rect 24584 11086 24636 11092
rect 24860 10600 24912 10606
rect 24860 10542 24912 10548
rect 24872 9994 24900 10542
rect 24860 9988 24912 9994
rect 24860 9930 24912 9936
rect 25320 9580 25372 9586
rect 25320 9522 25372 9528
rect 25332 9178 25360 9522
rect 24400 9172 24452 9178
rect 24400 9114 24452 9120
rect 25320 9172 25372 9178
rect 25320 9114 25372 9120
rect 24860 9036 24912 9042
rect 24860 8978 24912 8984
rect 24872 8838 24900 8978
rect 24860 8832 24912 8838
rect 24860 8774 24912 8780
rect 24872 8022 24900 8774
rect 24860 8016 24912 8022
rect 24860 7958 24912 7964
rect 22928 4684 22980 4690
rect 22928 4626 22980 4632
rect 23204 4684 23256 4690
rect 24044 4678 24164 4706
rect 23204 4626 23256 4632
rect 22940 4146 22968 4626
rect 23216 4146 23244 4626
rect 24032 4616 24084 4622
rect 24032 4558 24084 4564
rect 22928 4140 22980 4146
rect 22928 4082 22980 4088
rect 23204 4140 23256 4146
rect 23204 4082 23256 4088
rect 23480 4072 23532 4078
rect 23480 4014 23532 4020
rect 22836 3936 22888 3942
rect 22836 3878 22888 3884
rect 22560 3664 22612 3670
rect 22480 3624 22560 3652
rect 22560 3606 22612 3612
rect 22572 3466 22600 3606
rect 22848 3602 22876 3878
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 22836 3596 22888 3602
rect 22836 3538 22888 3544
rect 22560 3460 22612 3466
rect 22560 3402 22612 3408
rect 23388 3392 23440 3398
rect 23388 3334 23440 3340
rect 23204 3188 23256 3194
rect 23204 3130 23256 3136
rect 22652 3120 22704 3126
rect 22652 3062 22704 3068
rect 22664 2922 22692 3062
rect 23216 2922 23244 3130
rect 23400 3126 23428 3334
rect 23388 3120 23440 3126
rect 23388 3062 23440 3068
rect 22376 2916 22428 2922
rect 22376 2858 22428 2864
rect 22652 2916 22704 2922
rect 22652 2858 22704 2864
rect 23204 2916 23256 2922
rect 23204 2858 23256 2864
rect 22284 2644 22336 2650
rect 22284 2586 22336 2592
rect 20168 2508 20220 2514
rect 20168 2450 20220 2456
rect 22284 2508 22336 2514
rect 22284 2450 22336 2456
rect 19524 2440 19576 2446
rect 19524 2382 19576 2388
rect 19616 2440 19668 2446
rect 19616 2382 19668 2388
rect 20180 800 20208 2450
rect 22296 800 22324 2450
rect 22388 2446 22416 2858
rect 23400 2854 23428 3062
rect 23492 2854 23520 4014
rect 24044 3670 24072 4558
rect 24136 3670 24164 4678
rect 24584 4548 24636 4554
rect 24584 4490 24636 4496
rect 24400 4480 24452 4486
rect 24400 4422 24452 4428
rect 24412 4078 24440 4422
rect 24216 4072 24268 4078
rect 24216 4014 24268 4020
rect 24400 4072 24452 4078
rect 24400 4014 24452 4020
rect 24032 3664 24084 3670
rect 24032 3606 24084 3612
rect 24124 3664 24176 3670
rect 24124 3606 24176 3612
rect 23572 3528 23624 3534
rect 23572 3470 23624 3476
rect 23584 3194 23612 3470
rect 24136 3466 24164 3606
rect 24124 3460 24176 3466
rect 24124 3402 24176 3408
rect 23572 3188 23624 3194
rect 23572 3130 23624 3136
rect 23388 2848 23440 2854
rect 23388 2790 23440 2796
rect 23480 2848 23532 2854
rect 23480 2790 23532 2796
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 24228 2582 24256 4014
rect 24596 2990 24624 4490
rect 25424 4078 25452 11727
rect 25608 9654 25636 14758
rect 25792 13326 25820 16510
rect 25964 16458 26016 16464
rect 25976 16114 26004 16458
rect 25964 16108 26016 16114
rect 25964 16050 26016 16056
rect 25976 15910 26004 16050
rect 26068 16046 26096 19071
rect 26056 16040 26108 16046
rect 26056 15982 26108 15988
rect 25964 15904 26016 15910
rect 26160 15881 26188 19366
rect 26252 18222 26280 21848
rect 26516 21830 26568 21836
rect 26332 21344 26384 21350
rect 26332 21286 26384 21292
rect 26344 18442 26372 21286
rect 26620 20346 26648 21950
rect 26976 21616 27028 21622
rect 26976 21558 27028 21564
rect 26884 21548 26936 21554
rect 26884 21490 26936 21496
rect 26698 21176 26754 21185
rect 26698 21111 26700 21120
rect 26752 21111 26754 21120
rect 26700 21082 26752 21088
rect 26712 20466 26740 21082
rect 26896 21049 26924 21490
rect 26882 21040 26938 21049
rect 26882 20975 26938 20984
rect 26792 20868 26844 20874
rect 26792 20810 26844 20816
rect 26700 20460 26752 20466
rect 26700 20402 26752 20408
rect 26620 20318 26740 20346
rect 26608 20256 26660 20262
rect 26608 20198 26660 20204
rect 26424 19984 26476 19990
rect 26424 19926 26476 19932
rect 26436 19352 26464 19926
rect 26620 19417 26648 20198
rect 26606 19408 26662 19417
rect 26424 19346 26476 19352
rect 26606 19343 26662 19352
rect 26620 19310 26648 19343
rect 26424 19288 26476 19294
rect 26608 19304 26660 19310
rect 26436 18601 26464 19288
rect 26608 19246 26660 19252
rect 26422 18592 26478 18601
rect 26422 18527 26478 18536
rect 26344 18414 26556 18442
rect 26240 18216 26292 18222
rect 26424 18216 26476 18222
rect 26240 18158 26292 18164
rect 26330 18184 26386 18193
rect 26424 18158 26476 18164
rect 26330 18119 26386 18128
rect 26344 17814 26372 18119
rect 26332 17808 26384 17814
rect 26332 17750 26384 17756
rect 26344 16998 26372 17750
rect 26332 16992 26384 16998
rect 26332 16934 26384 16940
rect 26436 16250 26464 18158
rect 26528 17649 26556 18414
rect 26514 17640 26570 17649
rect 26514 17575 26570 17584
rect 26608 17536 26660 17542
rect 26608 17478 26660 17484
rect 26620 16658 26648 17478
rect 26712 17105 26740 20318
rect 26804 20058 26832 20810
rect 26884 20528 26936 20534
rect 26884 20470 26936 20476
rect 26792 20052 26844 20058
rect 26792 19994 26844 20000
rect 26896 19718 26924 20470
rect 26884 19712 26936 19718
rect 26790 19680 26846 19689
rect 26884 19654 26936 19660
rect 26790 19615 26846 19624
rect 26698 17096 26754 17105
rect 26698 17031 26754 17040
rect 26608 16652 26660 16658
rect 26608 16594 26660 16600
rect 26424 16244 26476 16250
rect 26424 16186 26476 16192
rect 26620 16114 26648 16594
rect 26804 16182 26832 19615
rect 26896 16250 26924 19654
rect 26988 18737 27016 21558
rect 27080 18834 27108 22102
rect 27172 21146 27200 22188
rect 27250 22128 27306 22137
rect 27250 22063 27252 22072
rect 27304 22063 27306 22072
rect 27252 22034 27304 22040
rect 27356 21185 27384 22578
rect 27528 22568 27580 22574
rect 27528 22510 27580 22516
rect 27436 21888 27488 21894
rect 27540 21876 27568 22510
rect 27620 21888 27672 21894
rect 27540 21848 27620 21876
rect 27436 21830 27488 21836
rect 27620 21830 27672 21836
rect 27448 21706 27476 21830
rect 27724 21706 27752 23462
rect 27816 22778 27844 23598
rect 28000 23322 28028 23666
rect 27988 23316 28040 23322
rect 27988 23258 28040 23264
rect 28540 23112 28592 23118
rect 28540 23054 28592 23060
rect 28448 23044 28500 23050
rect 28448 22986 28500 22992
rect 28264 22976 28316 22982
rect 28316 22936 28396 22964
rect 28264 22918 28316 22924
rect 27950 22876 28258 22885
rect 27950 22874 27956 22876
rect 28012 22874 28036 22876
rect 28092 22874 28116 22876
rect 28172 22874 28196 22876
rect 28252 22874 28258 22876
rect 28012 22822 28014 22874
rect 28194 22822 28196 22874
rect 27950 22820 27956 22822
rect 28012 22820 28036 22822
rect 28092 22820 28116 22822
rect 28172 22820 28196 22822
rect 28252 22820 28258 22822
rect 27950 22811 28258 22820
rect 27804 22772 27856 22778
rect 27804 22714 27856 22720
rect 27816 22642 27844 22714
rect 28368 22710 28396 22936
rect 28356 22704 28408 22710
rect 28356 22646 28408 22652
rect 27804 22636 27856 22642
rect 27804 22578 27856 22584
rect 28460 22574 28488 22986
rect 28356 22568 28408 22574
rect 28356 22510 28408 22516
rect 28448 22568 28500 22574
rect 28448 22510 28500 22516
rect 28368 22234 28396 22510
rect 27804 22228 27856 22234
rect 27804 22170 27856 22176
rect 28356 22228 28408 22234
rect 28356 22170 28408 22176
rect 27448 21678 27752 21706
rect 27816 21690 27844 22170
rect 28552 22098 28580 23054
rect 28540 22092 28592 22098
rect 28540 22034 28592 22040
rect 27950 21788 28258 21797
rect 27950 21786 27956 21788
rect 28012 21786 28036 21788
rect 28092 21786 28116 21788
rect 28172 21786 28196 21788
rect 28252 21786 28258 21788
rect 28012 21734 28014 21786
rect 28194 21734 28196 21786
rect 27950 21732 27956 21734
rect 28012 21732 28036 21734
rect 28092 21732 28116 21734
rect 28172 21732 28196 21734
rect 28252 21732 28258 21734
rect 27950 21723 28258 21732
rect 27724 21622 27752 21678
rect 27804 21684 27856 21690
rect 27804 21626 27856 21632
rect 27436 21616 27488 21622
rect 27436 21558 27488 21564
rect 27712 21616 27764 21622
rect 27712 21558 27764 21564
rect 27448 21457 27476 21558
rect 27434 21448 27490 21457
rect 27434 21383 27490 21392
rect 27342 21176 27398 21185
rect 27160 21140 27212 21146
rect 27342 21111 27398 21120
rect 27804 21140 27856 21146
rect 27160 21082 27212 21088
rect 27804 21082 27856 21088
rect 27344 20936 27396 20942
rect 27344 20878 27396 20884
rect 27160 20868 27212 20874
rect 27160 20810 27212 20816
rect 27172 20398 27200 20810
rect 27160 20392 27212 20398
rect 27160 20334 27212 20340
rect 27172 19922 27200 20334
rect 27160 19916 27212 19922
rect 27160 19858 27212 19864
rect 27356 19514 27384 20878
rect 27528 20392 27580 20398
rect 27528 20334 27580 20340
rect 27620 20392 27672 20398
rect 27672 20352 27752 20380
rect 27620 20334 27672 20340
rect 27344 19508 27396 19514
rect 27344 19450 27396 19456
rect 27252 19168 27304 19174
rect 27252 19110 27304 19116
rect 27068 18828 27120 18834
rect 27068 18770 27120 18776
rect 26974 18728 27030 18737
rect 26974 18663 27030 18672
rect 27066 18456 27122 18465
rect 27264 18426 27292 19110
rect 27344 18828 27396 18834
rect 27344 18770 27396 18776
rect 27066 18391 27122 18400
rect 27252 18420 27304 18426
rect 27080 18057 27108 18391
rect 27252 18362 27304 18368
rect 27252 18216 27304 18222
rect 27250 18184 27252 18193
rect 27304 18184 27306 18193
rect 27250 18119 27306 18128
rect 27160 18080 27212 18086
rect 27066 18048 27122 18057
rect 27160 18022 27212 18028
rect 27066 17983 27122 17992
rect 27080 16969 27108 17983
rect 27066 16960 27122 16969
rect 27066 16895 27122 16904
rect 26976 16584 27028 16590
rect 26976 16526 27028 16532
rect 26884 16244 26936 16250
rect 26884 16186 26936 16192
rect 26792 16176 26844 16182
rect 26792 16118 26844 16124
rect 26608 16108 26660 16114
rect 26608 16050 26660 16056
rect 26240 16040 26292 16046
rect 26240 15982 26292 15988
rect 25964 15846 26016 15852
rect 26146 15872 26202 15881
rect 26146 15807 26202 15816
rect 26252 15570 26280 15982
rect 26424 15972 26476 15978
rect 26424 15914 26476 15920
rect 26240 15564 26292 15570
rect 26240 15506 26292 15512
rect 26332 15428 26384 15434
rect 26332 15370 26384 15376
rect 26344 14929 26372 15370
rect 26330 14920 26386 14929
rect 26330 14855 26386 14864
rect 25964 14272 26016 14278
rect 25964 14214 26016 14220
rect 25976 13394 26004 14214
rect 25964 13388 26016 13394
rect 25964 13330 26016 13336
rect 25780 13320 25832 13326
rect 25780 13262 25832 13268
rect 26332 13252 26384 13258
rect 26332 13194 26384 13200
rect 26056 13184 26108 13190
rect 26056 13126 26108 13132
rect 25870 12744 25926 12753
rect 25870 12679 25872 12688
rect 25924 12679 25926 12688
rect 25872 12650 25924 12656
rect 25596 9648 25648 9654
rect 25596 9590 25648 9596
rect 25780 9580 25832 9586
rect 25780 9522 25832 9528
rect 25688 9376 25740 9382
rect 25688 9318 25740 9324
rect 25596 9172 25648 9178
rect 25596 9114 25648 9120
rect 25608 9081 25636 9114
rect 25700 9110 25728 9318
rect 25688 9104 25740 9110
rect 25594 9072 25650 9081
rect 25688 9046 25740 9052
rect 25594 9007 25650 9016
rect 25792 8922 25820 9522
rect 25884 9466 25912 12650
rect 26068 12442 26096 13126
rect 26238 13016 26294 13025
rect 26344 12986 26372 13194
rect 26238 12951 26294 12960
rect 26332 12980 26384 12986
rect 26252 12850 26280 12951
rect 26332 12922 26384 12928
rect 26240 12844 26292 12850
rect 26240 12786 26292 12792
rect 26056 12436 26108 12442
rect 26436 12434 26464 15914
rect 26608 15904 26660 15910
rect 26608 15846 26660 15852
rect 26700 15904 26752 15910
rect 26700 15846 26752 15852
rect 26620 15706 26648 15846
rect 26608 15700 26660 15706
rect 26608 15642 26660 15648
rect 26516 15564 26568 15570
rect 26516 15506 26568 15512
rect 26608 15564 26660 15570
rect 26608 15506 26660 15512
rect 26528 14074 26556 15506
rect 26516 14068 26568 14074
rect 26516 14010 26568 14016
rect 26528 12782 26556 14010
rect 26516 12776 26568 12782
rect 26516 12718 26568 12724
rect 26056 12378 26108 12384
rect 26344 12406 26464 12434
rect 26344 12102 26372 12406
rect 26332 12096 26384 12102
rect 26332 12038 26384 12044
rect 25964 11824 26016 11830
rect 25964 11766 26016 11772
rect 25976 11150 26004 11766
rect 26148 11756 26200 11762
rect 26148 11698 26200 11704
rect 25964 11144 26016 11150
rect 25964 11086 26016 11092
rect 25976 10470 26004 11086
rect 26160 11014 26188 11698
rect 26344 11694 26372 12038
rect 26332 11688 26384 11694
rect 26332 11630 26384 11636
rect 26620 11286 26648 15506
rect 26712 12170 26740 15846
rect 26884 15700 26936 15706
rect 26988 15688 27016 16526
rect 26936 15660 27016 15688
rect 26884 15642 26936 15648
rect 26896 14822 26924 15642
rect 27172 15502 27200 18022
rect 27356 17610 27384 18770
rect 27436 18760 27488 18766
rect 27436 18702 27488 18708
rect 27448 18290 27476 18702
rect 27436 18284 27488 18290
rect 27436 18226 27488 18232
rect 27436 18080 27488 18086
rect 27436 18022 27488 18028
rect 27344 17604 27396 17610
rect 27344 17546 27396 17552
rect 27344 17196 27396 17202
rect 27344 17138 27396 17144
rect 27252 17128 27304 17134
rect 27252 17070 27304 17076
rect 27264 16697 27292 17070
rect 27356 16794 27384 17138
rect 27344 16788 27396 16794
rect 27344 16730 27396 16736
rect 27250 16688 27306 16697
rect 27250 16623 27306 16632
rect 27264 16522 27292 16623
rect 27252 16516 27304 16522
rect 27252 16458 27304 16464
rect 27448 16046 27476 18022
rect 27540 17202 27568 20334
rect 27620 19712 27672 19718
rect 27724 19689 27752 20352
rect 27620 19654 27672 19660
rect 27710 19680 27766 19689
rect 27632 18358 27660 19654
rect 27710 19615 27766 19624
rect 27712 19508 27764 19514
rect 27712 19450 27764 19456
rect 27620 18352 27672 18358
rect 27620 18294 27672 18300
rect 27618 17912 27674 17921
rect 27618 17847 27674 17856
rect 27632 17610 27660 17847
rect 27620 17604 27672 17610
rect 27620 17546 27672 17552
rect 27528 17196 27580 17202
rect 27528 17138 27580 17144
rect 27632 16810 27660 17546
rect 27724 17218 27752 19450
rect 27816 19242 27844 21082
rect 28644 20942 28672 24006
rect 28908 22432 28960 22438
rect 28908 22374 28960 22380
rect 28920 22098 28948 22374
rect 29000 22228 29052 22234
rect 29000 22170 29052 22176
rect 28908 22092 28960 22098
rect 28908 22034 28960 22040
rect 28814 21584 28870 21593
rect 28724 21548 28776 21554
rect 28814 21519 28816 21528
rect 28724 21490 28776 21496
rect 28868 21519 28870 21528
rect 28816 21490 28868 21496
rect 28736 21010 28764 21490
rect 28724 21004 28776 21010
rect 28724 20946 28776 20952
rect 28828 20942 28856 21490
rect 28920 21486 28948 22034
rect 28908 21480 28960 21486
rect 28908 21422 28960 21428
rect 28632 20936 28684 20942
rect 28632 20878 28684 20884
rect 28816 20936 28868 20942
rect 28816 20878 28868 20884
rect 28632 20800 28684 20806
rect 28446 20768 28502 20777
rect 28724 20800 28776 20806
rect 28632 20742 28684 20748
rect 28722 20768 28724 20777
rect 28816 20800 28868 20806
rect 28776 20768 28778 20777
rect 27950 20700 28258 20709
rect 28446 20703 28502 20712
rect 27950 20698 27956 20700
rect 28012 20698 28036 20700
rect 28092 20698 28116 20700
rect 28172 20698 28196 20700
rect 28252 20698 28258 20700
rect 28012 20646 28014 20698
rect 28194 20646 28196 20698
rect 27950 20644 27956 20646
rect 28012 20644 28036 20646
rect 28092 20644 28116 20646
rect 28172 20644 28196 20646
rect 28252 20644 28258 20646
rect 27950 20635 28258 20644
rect 28264 20528 28316 20534
rect 28316 20488 28396 20516
rect 28264 20470 28316 20476
rect 28368 20058 28396 20488
rect 28356 20052 28408 20058
rect 28356 19994 28408 20000
rect 27950 19612 28258 19621
rect 27950 19610 27956 19612
rect 28012 19610 28036 19612
rect 28092 19610 28116 19612
rect 28172 19610 28196 19612
rect 28252 19610 28258 19612
rect 28012 19558 28014 19610
rect 28194 19558 28196 19610
rect 27950 19556 27956 19558
rect 28012 19556 28036 19558
rect 28092 19556 28116 19558
rect 28172 19556 28196 19558
rect 28252 19556 28258 19558
rect 27950 19547 28258 19556
rect 28264 19440 28316 19446
rect 28264 19382 28316 19388
rect 27804 19236 27856 19242
rect 27804 19178 27856 19184
rect 27988 19168 28040 19174
rect 27988 19110 28040 19116
rect 27804 18692 27856 18698
rect 27804 18634 27856 18640
rect 27816 17921 27844 18634
rect 28000 18630 28028 19110
rect 27988 18624 28040 18630
rect 28276 18612 28304 19382
rect 28368 18902 28396 19994
rect 28460 19514 28488 20703
rect 28644 20074 28672 20742
rect 28816 20742 28868 20748
rect 28722 20703 28778 20712
rect 28828 20233 28856 20742
rect 29012 20398 29040 22170
rect 29104 21418 29132 24618
rect 29196 23730 29224 24686
rect 29184 23724 29236 23730
rect 29184 23666 29236 23672
rect 29184 23520 29236 23526
rect 29184 23462 29236 23468
rect 29092 21412 29144 21418
rect 29092 21354 29144 21360
rect 29196 20482 29224 23462
rect 29288 23254 29316 26200
rect 29368 25084 29420 25090
rect 29368 25026 29420 25032
rect 29276 23248 29328 23254
rect 29276 23190 29328 23196
rect 29380 23100 29408 25026
rect 29644 24948 29696 24954
rect 29644 24890 29696 24896
rect 29460 23792 29512 23798
rect 29460 23734 29512 23740
rect 29472 23186 29500 23734
rect 29460 23180 29512 23186
rect 29460 23122 29512 23128
rect 29288 23072 29408 23100
rect 29288 22094 29316 23072
rect 29472 22982 29500 23122
rect 29460 22976 29512 22982
rect 29460 22918 29512 22924
rect 29472 22642 29500 22918
rect 29460 22636 29512 22642
rect 29460 22578 29512 22584
rect 29368 22500 29420 22506
rect 29368 22442 29420 22448
rect 29380 22234 29408 22442
rect 29472 22234 29500 22578
rect 29368 22228 29420 22234
rect 29368 22170 29420 22176
rect 29460 22228 29512 22234
rect 29460 22170 29512 22176
rect 29288 22066 29408 22094
rect 29276 21480 29328 21486
rect 29276 21422 29328 21428
rect 29288 20874 29316 21422
rect 29276 20868 29328 20874
rect 29276 20810 29328 20816
rect 29380 20806 29408 22066
rect 29368 20800 29420 20806
rect 29368 20742 29420 20748
rect 29196 20454 29408 20482
rect 29000 20392 29052 20398
rect 29000 20334 29052 20340
rect 29276 20392 29328 20398
rect 29276 20334 29328 20340
rect 29000 20256 29052 20262
rect 28814 20224 28870 20233
rect 29000 20198 29052 20204
rect 28814 20159 28870 20168
rect 28644 20046 28764 20074
rect 28736 19836 28764 20046
rect 29012 19922 29040 20198
rect 29000 19916 29052 19922
rect 29000 19858 29052 19864
rect 28908 19848 28960 19854
rect 28736 19808 28908 19836
rect 29288 19836 29316 20334
rect 28908 19790 28960 19796
rect 29104 19808 29316 19836
rect 28724 19712 28776 19718
rect 28538 19680 28594 19689
rect 28908 19712 28960 19718
rect 28776 19672 28908 19700
rect 28724 19654 28776 19660
rect 28908 19654 28960 19660
rect 28538 19615 28594 19624
rect 28448 19508 28500 19514
rect 28448 19450 28500 19456
rect 28552 19446 28580 19615
rect 28814 19544 28870 19553
rect 28814 19479 28870 19488
rect 28540 19440 28592 19446
rect 28540 19382 28592 19388
rect 28632 19372 28684 19378
rect 28460 19320 28632 19334
rect 28460 19314 28684 19320
rect 28828 19334 28856 19479
rect 28460 19306 28672 19314
rect 28356 18896 28408 18902
rect 28356 18838 28408 18844
rect 28460 18766 28488 19306
rect 28724 19304 28776 19310
rect 28828 19306 28948 19334
rect 28724 19246 28776 19252
rect 28540 19236 28592 19242
rect 28540 19178 28592 19184
rect 28632 19236 28684 19242
rect 28632 19178 28684 19184
rect 28448 18760 28500 18766
rect 28448 18702 28500 18708
rect 28276 18584 28488 18612
rect 27988 18566 28040 18572
rect 27950 18524 28258 18533
rect 27950 18522 27956 18524
rect 28012 18522 28036 18524
rect 28092 18522 28116 18524
rect 28172 18522 28196 18524
rect 28252 18522 28258 18524
rect 28012 18470 28014 18522
rect 28194 18470 28196 18522
rect 27950 18468 27956 18470
rect 28012 18468 28036 18470
rect 28092 18468 28116 18470
rect 28172 18468 28196 18470
rect 28252 18468 28258 18470
rect 27950 18459 28258 18468
rect 27802 17912 27858 17921
rect 27802 17847 27858 17856
rect 28356 17740 28408 17746
rect 28356 17682 28408 17688
rect 27950 17436 28258 17445
rect 27950 17434 27956 17436
rect 28012 17434 28036 17436
rect 28092 17434 28116 17436
rect 28172 17434 28196 17436
rect 28252 17434 28258 17436
rect 28012 17382 28014 17434
rect 28194 17382 28196 17434
rect 27950 17380 27956 17382
rect 28012 17380 28036 17382
rect 28092 17380 28116 17382
rect 28172 17380 28196 17382
rect 28252 17380 28258 17382
rect 27950 17371 28258 17380
rect 27896 17264 27948 17270
rect 27724 17212 27896 17218
rect 27724 17206 27948 17212
rect 28262 17232 28318 17241
rect 27724 17190 27936 17206
rect 28080 17196 28132 17202
rect 28262 17167 28318 17176
rect 28080 17138 28132 17144
rect 27804 16992 27856 16998
rect 27710 16960 27766 16969
rect 27804 16934 27856 16940
rect 27710 16895 27766 16904
rect 27540 16782 27660 16810
rect 27540 16590 27568 16782
rect 27620 16720 27672 16726
rect 27620 16662 27672 16668
rect 27528 16584 27580 16590
rect 27528 16526 27580 16532
rect 27632 16182 27660 16662
rect 27620 16176 27672 16182
rect 27620 16118 27672 16124
rect 27436 16040 27488 16046
rect 27342 16008 27398 16017
rect 27436 15982 27488 15988
rect 27342 15943 27398 15952
rect 27356 15706 27384 15943
rect 27344 15700 27396 15706
rect 27344 15642 27396 15648
rect 27160 15496 27212 15502
rect 26974 15464 27030 15473
rect 27160 15438 27212 15444
rect 27356 15434 27384 15642
rect 27724 15434 27752 16895
rect 27816 15502 27844 16934
rect 28092 16454 28120 17138
rect 28276 16522 28304 17167
rect 28264 16516 28316 16522
rect 28264 16458 28316 16464
rect 28080 16448 28132 16454
rect 28080 16390 28132 16396
rect 27950 16348 28258 16357
rect 27950 16346 27956 16348
rect 28012 16346 28036 16348
rect 28092 16346 28116 16348
rect 28172 16346 28196 16348
rect 28252 16346 28258 16348
rect 28012 16294 28014 16346
rect 28194 16294 28196 16346
rect 27950 16292 27956 16294
rect 28012 16292 28036 16294
rect 28092 16292 28116 16294
rect 28172 16292 28196 16294
rect 28252 16292 28258 16294
rect 27950 16283 28258 16292
rect 28368 16114 28396 17682
rect 28356 16108 28408 16114
rect 28356 16050 28408 16056
rect 27804 15496 27856 15502
rect 27804 15438 27856 15444
rect 26974 15399 27030 15408
rect 27344 15428 27396 15434
rect 26988 15366 27016 15399
rect 27344 15370 27396 15376
rect 27712 15428 27764 15434
rect 27712 15370 27764 15376
rect 26976 15360 27028 15366
rect 26976 15302 27028 15308
rect 27436 15360 27488 15366
rect 27436 15302 27488 15308
rect 26884 14816 26936 14822
rect 26884 14758 26936 14764
rect 26896 14346 26924 14758
rect 26884 14340 26936 14346
rect 26804 14300 26884 14328
rect 26804 13938 26832 14300
rect 26884 14282 26936 14288
rect 26792 13932 26844 13938
rect 26792 13874 26844 13880
rect 26804 13190 26832 13874
rect 26792 13184 26844 13190
rect 26792 13126 26844 13132
rect 26804 12918 26832 13126
rect 26792 12912 26844 12918
rect 26792 12854 26844 12860
rect 26804 12238 26832 12854
rect 26988 12850 27016 15302
rect 27066 15056 27122 15065
rect 27066 14991 27068 15000
rect 27120 14991 27122 15000
rect 27068 14962 27120 14968
rect 27344 14952 27396 14958
rect 27264 14900 27344 14906
rect 27264 14894 27396 14900
rect 27264 14878 27384 14894
rect 27160 14476 27212 14482
rect 27160 14418 27212 14424
rect 27172 12850 27200 14418
rect 26976 12844 27028 12850
rect 26976 12786 27028 12792
rect 27160 12844 27212 12850
rect 27160 12786 27212 12792
rect 27172 12646 27200 12786
rect 27160 12640 27212 12646
rect 27160 12582 27212 12588
rect 26792 12232 26844 12238
rect 26792 12174 26844 12180
rect 26700 12164 26752 12170
rect 26700 12106 26752 12112
rect 27160 12164 27212 12170
rect 27160 12106 27212 12112
rect 26608 11280 26660 11286
rect 26608 11222 26660 11228
rect 26148 11008 26200 11014
rect 26148 10950 26200 10956
rect 26148 10804 26200 10810
rect 26148 10746 26200 10752
rect 26160 10470 26188 10746
rect 26620 10606 26648 11222
rect 26976 11008 27028 11014
rect 26976 10950 27028 10956
rect 26608 10600 26660 10606
rect 26608 10542 26660 10548
rect 25964 10464 26016 10470
rect 25964 10406 26016 10412
rect 26148 10464 26200 10470
rect 26148 10406 26200 10412
rect 26516 10464 26568 10470
rect 26516 10406 26568 10412
rect 26792 10464 26844 10470
rect 26792 10406 26844 10412
rect 25976 10062 26004 10406
rect 25964 10056 26016 10062
rect 25964 9998 26016 10004
rect 25976 9654 26004 9998
rect 26160 9926 26188 10406
rect 26528 10198 26556 10406
rect 26516 10192 26568 10198
rect 26804 10169 26832 10406
rect 26516 10134 26568 10140
rect 26790 10160 26846 10169
rect 26528 10062 26556 10134
rect 26790 10095 26846 10104
rect 26988 10062 27016 10950
rect 26516 10056 26568 10062
rect 26516 9998 26568 10004
rect 26976 10056 27028 10062
rect 26976 9998 27028 10004
rect 26332 9988 26384 9994
rect 26332 9930 26384 9936
rect 26148 9920 26200 9926
rect 26148 9862 26200 9868
rect 25964 9648 26016 9654
rect 25964 9590 26016 9596
rect 26146 9616 26202 9625
rect 26146 9551 26148 9560
rect 26200 9551 26202 9560
rect 26148 9522 26200 9528
rect 25884 9438 26096 9466
rect 25700 8894 25820 8922
rect 25700 8838 25728 8894
rect 25688 8832 25740 8838
rect 25688 8774 25740 8780
rect 25700 7750 25728 8774
rect 25688 7744 25740 7750
rect 25688 7686 25740 7692
rect 25700 6254 25728 7686
rect 25688 6248 25740 6254
rect 25688 6190 25740 6196
rect 25412 4072 25464 4078
rect 25410 4040 25412 4049
rect 25464 4040 25466 4049
rect 25410 3975 25466 3984
rect 26068 3738 26096 9438
rect 26160 9178 26188 9522
rect 26344 9518 26372 9930
rect 26988 9518 27016 9998
rect 26332 9512 26384 9518
rect 26332 9454 26384 9460
rect 26976 9512 27028 9518
rect 26976 9454 27028 9460
rect 26148 9172 26200 9178
rect 26148 9114 26200 9120
rect 27172 8294 27200 12106
rect 27264 11626 27292 14878
rect 27448 13462 27476 15302
rect 27950 15260 28258 15269
rect 27950 15258 27956 15260
rect 28012 15258 28036 15260
rect 28092 15258 28116 15260
rect 28172 15258 28196 15260
rect 28252 15258 28258 15260
rect 28012 15206 28014 15258
rect 28194 15206 28196 15258
rect 27950 15204 27956 15206
rect 28012 15204 28036 15206
rect 28092 15204 28116 15206
rect 28172 15204 28196 15206
rect 28252 15204 28258 15206
rect 27526 15192 27582 15201
rect 27950 15195 28258 15204
rect 27526 15127 27582 15136
rect 27540 15094 27568 15127
rect 28368 15094 28396 16050
rect 27528 15088 27580 15094
rect 27528 15030 27580 15036
rect 28356 15088 28408 15094
rect 28356 15030 28408 15036
rect 27540 14482 27568 15030
rect 28460 14822 28488 18584
rect 28552 18086 28580 19178
rect 28644 19145 28672 19178
rect 28630 19136 28686 19145
rect 28630 19071 28686 19080
rect 28736 18630 28764 19246
rect 28920 18902 28948 19306
rect 28998 19000 29054 19009
rect 28998 18935 29054 18944
rect 28908 18896 28960 18902
rect 28908 18838 28960 18844
rect 29012 18698 29040 18935
rect 29000 18692 29052 18698
rect 29000 18634 29052 18640
rect 28724 18624 28776 18630
rect 28724 18566 28776 18572
rect 28540 18080 28592 18086
rect 28540 18022 28592 18028
rect 28538 17912 28594 17921
rect 28538 17847 28594 17856
rect 28552 17814 28580 17847
rect 28540 17808 28592 17814
rect 28540 17750 28592 17756
rect 28540 17332 28592 17338
rect 28540 17274 28592 17280
rect 28552 17218 28580 17274
rect 28552 17190 28672 17218
rect 28540 17128 28592 17134
rect 28540 17070 28592 17076
rect 28448 14816 28500 14822
rect 28448 14758 28500 14764
rect 27528 14476 27580 14482
rect 27528 14418 27580 14424
rect 28264 14476 28316 14482
rect 28264 14418 28316 14424
rect 28276 14385 28304 14418
rect 28262 14376 28318 14385
rect 28552 14346 28580 17070
rect 28644 16833 28672 17190
rect 28630 16824 28686 16833
rect 28630 16759 28632 16768
rect 28684 16759 28686 16768
rect 28632 16730 28684 16736
rect 28632 16040 28684 16046
rect 28632 15982 28684 15988
rect 28644 14482 28672 15982
rect 28632 14476 28684 14482
rect 28632 14418 28684 14424
rect 28262 14311 28318 14320
rect 28448 14340 28500 14346
rect 28448 14282 28500 14288
rect 28540 14340 28592 14346
rect 28540 14282 28592 14288
rect 27950 14172 28258 14181
rect 27950 14170 27956 14172
rect 28012 14170 28036 14172
rect 28092 14170 28116 14172
rect 28172 14170 28196 14172
rect 28252 14170 28258 14172
rect 28012 14118 28014 14170
rect 28194 14118 28196 14170
rect 27950 14116 27956 14118
rect 28012 14116 28036 14118
rect 28092 14116 28116 14118
rect 28172 14116 28196 14118
rect 28252 14116 28258 14118
rect 27950 14107 28258 14116
rect 28080 13932 28132 13938
rect 28080 13874 28132 13880
rect 28092 13530 28120 13874
rect 28080 13524 28132 13530
rect 28080 13466 28132 13472
rect 28356 13524 28408 13530
rect 28356 13466 28408 13472
rect 27436 13456 27488 13462
rect 27436 13398 27488 13404
rect 27950 13084 28258 13093
rect 27950 13082 27956 13084
rect 28012 13082 28036 13084
rect 28092 13082 28116 13084
rect 28172 13082 28196 13084
rect 28252 13082 28258 13084
rect 28012 13030 28014 13082
rect 28194 13030 28196 13082
rect 27950 13028 27956 13030
rect 28012 13028 28036 13030
rect 28092 13028 28116 13030
rect 28172 13028 28196 13030
rect 28252 13028 28258 13030
rect 27950 13019 28258 13028
rect 27344 12980 27396 12986
rect 27396 12940 27568 12968
rect 27344 12922 27396 12928
rect 27436 12300 27488 12306
rect 27436 12242 27488 12248
rect 27344 12096 27396 12102
rect 27344 12038 27396 12044
rect 27356 11898 27384 12038
rect 27344 11892 27396 11898
rect 27448 11880 27476 12242
rect 27540 12170 27568 12940
rect 27528 12164 27580 12170
rect 27528 12106 27580 12112
rect 27950 11996 28258 12005
rect 27950 11994 27956 11996
rect 28012 11994 28036 11996
rect 28092 11994 28116 11996
rect 28172 11994 28196 11996
rect 28252 11994 28258 11996
rect 28012 11942 28014 11994
rect 28194 11942 28196 11994
rect 27950 11940 27956 11942
rect 28012 11940 28036 11942
rect 28092 11940 28116 11942
rect 28172 11940 28196 11942
rect 28252 11940 28258 11942
rect 27950 11931 28258 11940
rect 27528 11892 27580 11898
rect 27448 11852 27528 11880
rect 27344 11834 27396 11840
rect 27528 11834 27580 11840
rect 27344 11756 27396 11762
rect 27344 11698 27396 11704
rect 27252 11620 27304 11626
rect 27252 11562 27304 11568
rect 27160 8288 27212 8294
rect 27160 8230 27212 8236
rect 27356 5710 27384 11698
rect 27436 10668 27488 10674
rect 27436 10610 27488 10616
rect 27448 5846 27476 10610
rect 27540 10169 27568 11834
rect 27804 11008 27856 11014
rect 27804 10950 27856 10956
rect 27816 10606 27844 10950
rect 27950 10908 28258 10917
rect 27950 10906 27956 10908
rect 28012 10906 28036 10908
rect 28092 10906 28116 10908
rect 28172 10906 28196 10908
rect 28252 10906 28258 10908
rect 28012 10854 28014 10906
rect 28194 10854 28196 10906
rect 27950 10852 27956 10854
rect 28012 10852 28036 10854
rect 28092 10852 28116 10854
rect 28172 10852 28196 10854
rect 28252 10852 28258 10854
rect 27950 10843 28258 10852
rect 27804 10600 27856 10606
rect 27804 10542 27856 10548
rect 27526 10160 27582 10169
rect 27526 10095 27582 10104
rect 27950 9820 28258 9829
rect 27950 9818 27956 9820
rect 28012 9818 28036 9820
rect 28092 9818 28116 9820
rect 28172 9818 28196 9820
rect 28252 9818 28258 9820
rect 28012 9766 28014 9818
rect 28194 9766 28196 9818
rect 27950 9764 27956 9766
rect 28012 9764 28036 9766
rect 28092 9764 28116 9766
rect 28172 9764 28196 9766
rect 28252 9764 28258 9766
rect 27950 9755 28258 9764
rect 27804 8832 27856 8838
rect 27804 8774 27856 8780
rect 27816 6730 27844 8774
rect 27950 8732 28258 8741
rect 27950 8730 27956 8732
rect 28012 8730 28036 8732
rect 28092 8730 28116 8732
rect 28172 8730 28196 8732
rect 28252 8730 28258 8732
rect 28012 8678 28014 8730
rect 28194 8678 28196 8730
rect 27950 8676 27956 8678
rect 28012 8676 28036 8678
rect 28092 8676 28116 8678
rect 28172 8676 28196 8678
rect 28252 8676 28258 8678
rect 27950 8667 28258 8676
rect 27950 7644 28258 7653
rect 27950 7642 27956 7644
rect 28012 7642 28036 7644
rect 28092 7642 28116 7644
rect 28172 7642 28196 7644
rect 28252 7642 28258 7644
rect 28012 7590 28014 7642
rect 28194 7590 28196 7642
rect 27950 7588 27956 7590
rect 28012 7588 28036 7590
rect 28092 7588 28116 7590
rect 28172 7588 28196 7590
rect 28252 7588 28258 7590
rect 27950 7579 28258 7588
rect 27804 6724 27856 6730
rect 27804 6666 27856 6672
rect 27950 6556 28258 6565
rect 27950 6554 27956 6556
rect 28012 6554 28036 6556
rect 28092 6554 28116 6556
rect 28172 6554 28196 6556
rect 28252 6554 28258 6556
rect 28012 6502 28014 6554
rect 28194 6502 28196 6554
rect 27950 6500 27956 6502
rect 28012 6500 28036 6502
rect 28092 6500 28116 6502
rect 28172 6500 28196 6502
rect 28252 6500 28258 6502
rect 27950 6491 28258 6500
rect 28368 6186 28396 13466
rect 28460 13172 28488 14282
rect 28644 13870 28672 14418
rect 28736 14385 28764 18566
rect 28998 18456 29054 18465
rect 28998 18391 29000 18400
rect 29052 18391 29054 18400
rect 29000 18362 29052 18368
rect 28816 18216 28868 18222
rect 28816 18158 28868 18164
rect 28828 17542 28856 18158
rect 28908 17876 28960 17882
rect 28908 17818 28960 17824
rect 28920 17678 28948 17818
rect 28908 17672 28960 17678
rect 28908 17614 28960 17620
rect 28816 17536 28868 17542
rect 28816 17478 28868 17484
rect 28828 17066 28856 17478
rect 28816 17060 28868 17066
rect 28816 17002 28868 17008
rect 28816 16584 28868 16590
rect 28816 16526 28868 16532
rect 28828 15638 28856 16526
rect 28816 15632 28868 15638
rect 28816 15574 28868 15580
rect 28722 14376 28778 14385
rect 28722 14311 28778 14320
rect 28920 14006 28948 17614
rect 29012 16522 29040 18362
rect 29000 16516 29052 16522
rect 29000 16458 29052 16464
rect 29104 16046 29132 19808
rect 29274 19680 29330 19689
rect 29274 19615 29330 19624
rect 29184 19304 29236 19310
rect 29182 19272 29184 19281
rect 29236 19272 29238 19281
rect 29182 19207 29238 19216
rect 29184 18760 29236 18766
rect 29184 18702 29236 18708
rect 29196 18426 29224 18702
rect 29184 18420 29236 18426
rect 29184 18362 29236 18368
rect 29288 17270 29316 19615
rect 29380 18465 29408 20454
rect 29472 20058 29500 22170
rect 29656 21457 29684 24890
rect 29932 24410 29960 26200
rect 30576 26058 30604 26200
rect 30668 26058 30696 26318
rect 31206 26200 31262 27000
rect 31850 26200 31906 27000
rect 32494 26200 32550 27000
rect 33138 26200 33194 27000
rect 33782 26200 33838 27000
rect 34426 26200 34482 27000
rect 35070 26200 35126 27000
rect 35714 26200 35770 27000
rect 36358 26330 36414 27000
rect 36358 26302 36768 26330
rect 36358 26200 36414 26302
rect 30576 26030 30696 26058
rect 30564 24608 30616 24614
rect 30564 24550 30616 24556
rect 30102 24440 30158 24449
rect 29920 24404 29972 24410
rect 30102 24375 30158 24384
rect 29920 24346 29972 24352
rect 30010 24304 30066 24313
rect 30010 24239 30066 24248
rect 29736 23588 29788 23594
rect 29736 23530 29788 23536
rect 29748 23322 29776 23530
rect 29736 23316 29788 23322
rect 29736 23258 29788 23264
rect 29920 22432 29972 22438
rect 29920 22374 29972 22380
rect 29932 22094 29960 22374
rect 30024 22137 30052 24239
rect 30116 24206 30144 24375
rect 30576 24206 30604 24550
rect 30104 24200 30156 24206
rect 30104 24142 30156 24148
rect 30564 24200 30616 24206
rect 30564 24142 30616 24148
rect 31116 24200 31168 24206
rect 31116 24142 31168 24148
rect 30748 24132 30800 24138
rect 30748 24074 30800 24080
rect 30380 24064 30432 24070
rect 30380 24006 30432 24012
rect 30194 23216 30250 23225
rect 30194 23151 30196 23160
rect 30248 23151 30250 23160
rect 30196 23122 30248 23128
rect 30104 22976 30156 22982
rect 30104 22918 30156 22924
rect 29840 22066 29960 22094
rect 30010 22128 30066 22137
rect 29840 21962 29868 22066
rect 30010 22063 30066 22072
rect 29828 21956 29880 21962
rect 29828 21898 29880 21904
rect 29828 21616 29880 21622
rect 29828 21558 29880 21564
rect 29642 21448 29698 21457
rect 29642 21383 29698 21392
rect 29552 21344 29604 21350
rect 29552 21286 29604 21292
rect 29564 21078 29592 21286
rect 29552 21072 29604 21078
rect 29552 21014 29604 21020
rect 29552 20800 29604 20806
rect 29552 20742 29604 20748
rect 29460 20052 29512 20058
rect 29460 19994 29512 20000
rect 29460 19916 29512 19922
rect 29460 19858 29512 19864
rect 29472 18834 29500 19858
rect 29460 18828 29512 18834
rect 29460 18770 29512 18776
rect 29366 18456 29422 18465
rect 29366 18391 29422 18400
rect 29564 18193 29592 20742
rect 29656 18834 29684 21383
rect 29734 20904 29790 20913
rect 29734 20839 29790 20848
rect 29748 20806 29776 20839
rect 29736 20800 29788 20806
rect 29736 20742 29788 20748
rect 29840 20534 29868 21558
rect 29920 21412 29972 21418
rect 29920 21354 29972 21360
rect 29828 20528 29880 20534
rect 29828 20470 29880 20476
rect 29736 19712 29788 19718
rect 29736 19654 29788 19660
rect 29644 18828 29696 18834
rect 29644 18770 29696 18776
rect 29642 18728 29698 18737
rect 29642 18663 29698 18672
rect 29550 18184 29606 18193
rect 29368 18148 29420 18154
rect 29550 18119 29606 18128
rect 29368 18090 29420 18096
rect 29276 17264 29328 17270
rect 29276 17206 29328 17212
rect 29184 17128 29236 17134
rect 29184 17070 29236 17076
rect 29092 16040 29144 16046
rect 29092 15982 29144 15988
rect 29000 14272 29052 14278
rect 29000 14214 29052 14220
rect 28908 14000 28960 14006
rect 28908 13942 28960 13948
rect 28632 13864 28684 13870
rect 28632 13806 28684 13812
rect 28816 13320 28868 13326
rect 28816 13262 28868 13268
rect 28540 13184 28592 13190
rect 28460 13144 28540 13172
rect 28540 13126 28592 13132
rect 28448 12980 28500 12986
rect 28448 12922 28500 12928
rect 28460 11286 28488 12922
rect 28448 11280 28500 11286
rect 28448 11222 28500 11228
rect 28552 11121 28580 13126
rect 28724 12912 28776 12918
rect 28724 12854 28776 12860
rect 28736 12170 28764 12854
rect 28724 12164 28776 12170
rect 28724 12106 28776 12112
rect 28538 11112 28594 11121
rect 28538 11047 28594 11056
rect 28736 11064 28764 12106
rect 28828 11830 28856 13262
rect 28920 12238 28948 13942
rect 29012 13190 29040 14214
rect 29000 13184 29052 13190
rect 29000 13126 29052 13132
rect 29196 12374 29224 17070
rect 29274 16688 29330 16697
rect 29274 16623 29276 16632
rect 29328 16623 29330 16632
rect 29276 16594 29328 16600
rect 29276 16040 29328 16046
rect 29276 15982 29328 15988
rect 29288 15366 29316 15982
rect 29276 15360 29328 15366
rect 29276 15302 29328 15308
rect 29288 15094 29316 15302
rect 29276 15088 29328 15094
rect 29276 15030 29328 15036
rect 29380 14906 29408 18090
rect 29460 17876 29512 17882
rect 29460 17818 29512 17824
rect 29472 17202 29500 17818
rect 29656 17542 29684 18663
rect 29748 18290 29776 19654
rect 29932 18766 29960 21354
rect 30024 20534 30052 22063
rect 30116 21146 30144 22918
rect 30392 22098 30420 24006
rect 30760 23798 30788 24074
rect 31128 24070 31156 24142
rect 30932 24064 30984 24070
rect 30932 24006 30984 24012
rect 31116 24064 31168 24070
rect 31116 24006 31168 24012
rect 30748 23792 30800 23798
rect 30748 23734 30800 23740
rect 30656 23656 30708 23662
rect 30484 23616 30656 23644
rect 30380 22092 30432 22098
rect 30380 22034 30432 22040
rect 30392 21146 30420 22034
rect 30104 21140 30156 21146
rect 30104 21082 30156 21088
rect 30380 21140 30432 21146
rect 30380 21082 30432 21088
rect 30484 21078 30512 23616
rect 30656 23598 30708 23604
rect 30746 22808 30802 22817
rect 30746 22743 30748 22752
rect 30800 22743 30802 22752
rect 30748 22714 30800 22720
rect 30656 22636 30708 22642
rect 30656 22578 30708 22584
rect 30564 22024 30616 22030
rect 30564 21966 30616 21972
rect 30472 21072 30524 21078
rect 30472 21014 30524 21020
rect 30196 21004 30248 21010
rect 30196 20946 30248 20952
rect 30104 20868 30156 20874
rect 30104 20810 30156 20816
rect 30012 20528 30064 20534
rect 30012 20470 30064 20476
rect 30010 20360 30066 20369
rect 30010 20295 30066 20304
rect 30024 19786 30052 20295
rect 30012 19780 30064 19786
rect 30012 19722 30064 19728
rect 30024 19514 30052 19722
rect 30012 19508 30064 19514
rect 30012 19450 30064 19456
rect 30024 18873 30052 19450
rect 30010 18864 30066 18873
rect 30010 18799 30066 18808
rect 29920 18760 29972 18766
rect 29920 18702 29972 18708
rect 29920 18624 29972 18630
rect 29920 18566 29972 18572
rect 29736 18284 29788 18290
rect 29736 18226 29788 18232
rect 29644 17536 29696 17542
rect 29644 17478 29696 17484
rect 29656 17202 29684 17478
rect 29460 17196 29512 17202
rect 29460 17138 29512 17144
rect 29644 17196 29696 17202
rect 29644 17138 29696 17144
rect 29828 17128 29880 17134
rect 29828 17070 29880 17076
rect 29460 16652 29512 16658
rect 29460 16594 29512 16600
rect 29288 14878 29408 14906
rect 29288 13938 29316 14878
rect 29276 13932 29328 13938
rect 29276 13874 29328 13880
rect 29184 12368 29236 12374
rect 29184 12310 29236 12316
rect 28908 12232 28960 12238
rect 28908 12174 28960 12180
rect 28816 11824 28868 11830
rect 28816 11766 28868 11772
rect 28920 11354 28948 12174
rect 28908 11348 28960 11354
rect 28908 11290 28960 11296
rect 28816 11076 28868 11082
rect 28552 7546 28580 11047
rect 28736 11036 28816 11064
rect 28816 11018 28868 11024
rect 28828 10130 28856 11018
rect 28920 10810 28948 11290
rect 29196 11218 29224 12310
rect 29184 11212 29236 11218
rect 29184 11154 29236 11160
rect 29090 10976 29146 10985
rect 29090 10911 29146 10920
rect 28908 10804 28960 10810
rect 28908 10746 28960 10752
rect 29104 10606 29132 10911
rect 29092 10600 29144 10606
rect 29092 10542 29144 10548
rect 29092 10192 29144 10198
rect 29092 10134 29144 10140
rect 28816 10124 28868 10130
rect 28816 10066 28868 10072
rect 28828 9654 28856 10066
rect 29000 9920 29052 9926
rect 29000 9862 29052 9868
rect 28816 9648 28868 9654
rect 28816 9590 28868 9596
rect 28816 9512 28868 9518
rect 28816 9454 28868 9460
rect 28630 9072 28686 9081
rect 28630 9007 28686 9016
rect 28644 8838 28672 9007
rect 28632 8832 28684 8838
rect 28632 8774 28684 8780
rect 28828 8430 28856 9454
rect 29012 9178 29040 9862
rect 29000 9172 29052 9178
rect 29000 9114 29052 9120
rect 29104 8566 29132 10134
rect 29196 9450 29224 11154
rect 29288 11064 29316 13874
rect 29368 12844 29420 12850
rect 29368 12786 29420 12792
rect 29380 12646 29408 12786
rect 29368 12640 29420 12646
rect 29368 12582 29420 12588
rect 29380 12306 29408 12582
rect 29368 12300 29420 12306
rect 29368 12242 29420 12248
rect 29472 11642 29500 16594
rect 29736 15904 29788 15910
rect 29736 15846 29788 15852
rect 29550 15600 29606 15609
rect 29550 15535 29606 15544
rect 29564 14278 29592 15535
rect 29748 15162 29776 15846
rect 29736 15156 29788 15162
rect 29656 15116 29736 15144
rect 29552 14272 29604 14278
rect 29552 14214 29604 14220
rect 29564 12918 29592 14214
rect 29656 13394 29684 15116
rect 29736 15098 29788 15104
rect 29840 14958 29868 17070
rect 29828 14952 29880 14958
rect 29828 14894 29880 14900
rect 29828 14816 29880 14822
rect 29828 14758 29880 14764
rect 29736 14340 29788 14346
rect 29736 14282 29788 14288
rect 29748 14113 29776 14282
rect 29734 14104 29790 14113
rect 29734 14039 29790 14048
rect 29644 13388 29696 13394
rect 29644 13330 29696 13336
rect 29552 12912 29604 12918
rect 29550 12880 29552 12889
rect 29604 12880 29606 12889
rect 29550 12815 29606 12824
rect 29552 12776 29604 12782
rect 29552 12718 29604 12724
rect 29564 11744 29592 12718
rect 29656 12170 29684 13330
rect 29840 13326 29868 14758
rect 29828 13320 29880 13326
rect 29828 13262 29880 13268
rect 29932 13190 29960 18566
rect 30116 18154 30144 20810
rect 30208 20777 30236 20946
rect 30576 20942 30604 21966
rect 30668 21729 30696 22578
rect 30748 21956 30800 21962
rect 30748 21898 30800 21904
rect 30654 21720 30710 21729
rect 30654 21655 30710 21664
rect 30656 21344 30708 21350
rect 30656 21286 30708 21292
rect 30288 20936 30340 20942
rect 30288 20878 30340 20884
rect 30564 20936 30616 20942
rect 30564 20878 30616 20884
rect 30194 20768 30250 20777
rect 30194 20703 30250 20712
rect 30300 19530 30328 20878
rect 30564 20256 30616 20262
rect 30564 20198 30616 20204
rect 30380 20052 30432 20058
rect 30380 19994 30432 20000
rect 30392 19922 30420 19994
rect 30380 19916 30432 19922
rect 30380 19858 30432 19864
rect 30300 19502 30512 19530
rect 30380 19372 30432 19378
rect 30380 19314 30432 19320
rect 30392 19174 30420 19314
rect 30380 19168 30432 19174
rect 30380 19110 30432 19116
rect 30288 18828 30340 18834
rect 30288 18770 30340 18776
rect 30194 18184 30250 18193
rect 30104 18148 30156 18154
rect 30194 18119 30250 18128
rect 30104 18090 30156 18096
rect 30104 17604 30156 17610
rect 30104 17546 30156 17552
rect 30010 16688 30066 16697
rect 30010 16623 30066 16632
rect 30024 15094 30052 16623
rect 30116 15552 30144 17546
rect 30208 16522 30236 18119
rect 30196 16516 30248 16522
rect 30196 16458 30248 16464
rect 30116 15524 30236 15552
rect 30208 15094 30236 15524
rect 30300 15162 30328 18770
rect 30392 17814 30420 19110
rect 30484 18737 30512 19502
rect 30470 18728 30526 18737
rect 30470 18663 30526 18672
rect 30472 18624 30524 18630
rect 30472 18566 30524 18572
rect 30380 17808 30432 17814
rect 30380 17750 30432 17756
rect 30392 17678 30420 17750
rect 30380 17672 30432 17678
rect 30380 17614 30432 17620
rect 30380 17536 30432 17542
rect 30380 17478 30432 17484
rect 30392 17134 30420 17478
rect 30380 17128 30432 17134
rect 30380 17070 30432 17076
rect 30484 15609 30512 18566
rect 30576 17134 30604 20198
rect 30668 19009 30696 21286
rect 30760 19514 30788 21898
rect 30838 21176 30894 21185
rect 30838 21111 30894 21120
rect 30852 21078 30880 21111
rect 30840 21072 30892 21078
rect 30840 21014 30892 21020
rect 30838 20496 30894 20505
rect 30838 20431 30840 20440
rect 30892 20431 30894 20440
rect 30840 20402 30892 20408
rect 30840 19712 30892 19718
rect 30944 19700 30972 24006
rect 31022 23624 31078 23633
rect 31022 23559 31078 23568
rect 31036 22982 31064 23559
rect 31220 23236 31248 26200
rect 31300 25016 31352 25022
rect 31300 24958 31352 24964
rect 31128 23208 31248 23236
rect 31128 22982 31156 23208
rect 31024 22976 31076 22982
rect 31024 22918 31076 22924
rect 31116 22976 31168 22982
rect 31116 22918 31168 22924
rect 31036 22094 31064 22918
rect 31208 22772 31260 22778
rect 31208 22714 31260 22720
rect 31220 22098 31248 22714
rect 31036 22066 31156 22094
rect 31128 20534 31156 22066
rect 31208 22092 31260 22098
rect 31208 22034 31260 22040
rect 31208 21616 31260 21622
rect 31206 21584 31208 21593
rect 31260 21584 31262 21593
rect 31206 21519 31262 21528
rect 31116 20528 31168 20534
rect 31116 20470 31168 20476
rect 31208 20392 31260 20398
rect 31208 20334 31260 20340
rect 31024 20256 31076 20262
rect 31024 20198 31076 20204
rect 30892 19672 30972 19700
rect 30840 19654 30892 19660
rect 30748 19508 30800 19514
rect 30748 19450 30800 19456
rect 30654 19000 30710 19009
rect 30654 18935 30710 18944
rect 30852 17678 30880 19654
rect 30932 17740 30984 17746
rect 30932 17682 30984 17688
rect 30840 17672 30892 17678
rect 30654 17640 30710 17649
rect 30840 17614 30892 17620
rect 30654 17575 30710 17584
rect 30564 17128 30616 17134
rect 30564 17070 30616 17076
rect 30564 15904 30616 15910
rect 30564 15846 30616 15852
rect 30470 15600 30526 15609
rect 30470 15535 30526 15544
rect 30472 15496 30524 15502
rect 30472 15438 30524 15444
rect 30380 15428 30432 15434
rect 30380 15370 30432 15376
rect 30288 15156 30340 15162
rect 30288 15098 30340 15104
rect 30012 15088 30064 15094
rect 30012 15030 30064 15036
rect 30196 15088 30248 15094
rect 30196 15030 30248 15036
rect 30300 14090 30328 15098
rect 30392 14346 30420 15370
rect 30380 14340 30432 14346
rect 30380 14282 30432 14288
rect 30012 14068 30064 14074
rect 30012 14010 30064 14016
rect 30116 14062 30328 14090
rect 29920 13184 29972 13190
rect 29920 13126 29972 13132
rect 30024 12850 30052 14010
rect 30012 12844 30064 12850
rect 30012 12786 30064 12792
rect 29644 12164 29696 12170
rect 29644 12106 29696 12112
rect 30012 11824 30064 11830
rect 30012 11766 30064 11772
rect 29564 11716 29776 11744
rect 29472 11614 29684 11642
rect 29460 11552 29512 11558
rect 29512 11512 29592 11540
rect 29460 11494 29512 11500
rect 29564 11150 29592 11512
rect 29552 11144 29604 11150
rect 29552 11086 29604 11092
rect 29368 11076 29420 11082
rect 29288 11036 29368 11064
rect 29368 11018 29420 11024
rect 29380 10130 29408 11018
rect 29564 10742 29592 11086
rect 29552 10736 29604 10742
rect 29552 10678 29604 10684
rect 29368 10124 29420 10130
rect 29368 10066 29420 10072
rect 29564 9518 29592 10678
rect 29552 9512 29604 9518
rect 29552 9454 29604 9460
rect 29656 9450 29684 11614
rect 29748 11014 29776 11716
rect 30024 11286 30052 11766
rect 30116 11558 30144 14062
rect 30288 13388 30340 13394
rect 30288 13330 30340 13336
rect 30104 11552 30156 11558
rect 30104 11494 30156 11500
rect 30012 11280 30064 11286
rect 30012 11222 30064 11228
rect 29736 11008 29788 11014
rect 29736 10950 29788 10956
rect 30012 11008 30064 11014
rect 30012 10950 30064 10956
rect 29748 10810 29776 10950
rect 29736 10804 29788 10810
rect 29736 10746 29788 10752
rect 29736 10668 29788 10674
rect 29736 10610 29788 10616
rect 29184 9444 29236 9450
rect 29184 9386 29236 9392
rect 29644 9444 29696 9450
rect 29644 9386 29696 9392
rect 29656 9178 29684 9386
rect 29644 9172 29696 9178
rect 29644 9114 29696 9120
rect 29656 9042 29684 9114
rect 29644 9036 29696 9042
rect 29644 8978 29696 8984
rect 29092 8560 29144 8566
rect 29092 8502 29144 8508
rect 28816 8424 28868 8430
rect 28816 8366 28868 8372
rect 28540 7540 28592 7546
rect 28540 7482 28592 7488
rect 28356 6180 28408 6186
rect 28356 6122 28408 6128
rect 27436 5840 27488 5846
rect 27436 5782 27488 5788
rect 27344 5704 27396 5710
rect 27344 5646 27396 5652
rect 27950 5468 28258 5477
rect 27950 5466 27956 5468
rect 28012 5466 28036 5468
rect 28092 5466 28116 5468
rect 28172 5466 28196 5468
rect 28252 5466 28258 5468
rect 28012 5414 28014 5466
rect 28194 5414 28196 5466
rect 27950 5412 27956 5414
rect 28012 5412 28036 5414
rect 28092 5412 28116 5414
rect 28172 5412 28196 5414
rect 28252 5412 28258 5414
rect 27950 5403 28258 5412
rect 27950 4380 28258 4389
rect 27950 4378 27956 4380
rect 28012 4378 28036 4380
rect 28092 4378 28116 4380
rect 28172 4378 28196 4380
rect 28252 4378 28258 4380
rect 28012 4326 28014 4378
rect 28194 4326 28196 4378
rect 27950 4324 27956 4326
rect 28012 4324 28036 4326
rect 28092 4324 28116 4326
rect 28172 4324 28196 4326
rect 28252 4324 28258 4326
rect 27950 4315 28258 4324
rect 27620 4072 27672 4078
rect 27620 4014 27672 4020
rect 27632 3738 27660 4014
rect 27804 3936 27856 3942
rect 27804 3878 27856 3884
rect 25964 3732 26016 3738
rect 25964 3674 26016 3680
rect 26056 3732 26108 3738
rect 26056 3674 26108 3680
rect 27620 3732 27672 3738
rect 27620 3674 27672 3680
rect 25976 2990 26004 3674
rect 26068 3505 26096 3674
rect 26054 3496 26110 3505
rect 26054 3431 26110 3440
rect 27528 3392 27580 3398
rect 27528 3334 27580 3340
rect 26884 3120 26936 3126
rect 26884 3062 26936 3068
rect 24584 2984 24636 2990
rect 24584 2926 24636 2932
rect 25964 2984 26016 2990
rect 25964 2926 26016 2932
rect 26896 2922 26924 3062
rect 26884 2916 26936 2922
rect 26884 2858 26936 2864
rect 24584 2848 24636 2854
rect 24584 2790 24636 2796
rect 24216 2576 24268 2582
rect 24216 2518 24268 2524
rect 24400 2508 24452 2514
rect 24400 2450 24452 2456
rect 22376 2440 22428 2446
rect 22376 2382 22428 2388
rect 24412 800 24440 2450
rect 24596 2446 24624 2790
rect 26896 2650 26924 2858
rect 27160 2848 27212 2854
rect 27160 2790 27212 2796
rect 26884 2644 26936 2650
rect 26884 2586 26936 2592
rect 26516 2508 26568 2514
rect 26516 2450 26568 2456
rect 24584 2440 24636 2446
rect 24584 2382 24636 2388
rect 26528 800 26556 2450
rect 27172 2446 27200 2790
rect 27540 2650 27568 3334
rect 27712 3120 27764 3126
rect 27712 3062 27764 3068
rect 27724 2922 27752 3062
rect 27712 2916 27764 2922
rect 27712 2858 27764 2864
rect 27816 2836 27844 3878
rect 27950 3292 28258 3301
rect 27950 3290 27956 3292
rect 28012 3290 28036 3292
rect 28092 3290 28116 3292
rect 28172 3290 28196 3292
rect 28252 3290 28258 3292
rect 28012 3238 28014 3290
rect 28194 3238 28196 3290
rect 27950 3236 27956 3238
rect 28012 3236 28036 3238
rect 28092 3236 28116 3238
rect 28172 3236 28196 3238
rect 28252 3236 28258 3238
rect 27950 3227 28258 3236
rect 28828 3058 28856 8366
rect 29748 7954 29776 10610
rect 30024 10470 30052 10950
rect 30012 10464 30064 10470
rect 30012 10406 30064 10412
rect 30116 9994 30144 11494
rect 30194 11112 30250 11121
rect 30194 11047 30196 11056
rect 30248 11047 30250 11056
rect 30196 11018 30248 11024
rect 30300 10742 30328 13330
rect 30392 12209 30420 14282
rect 30484 14074 30512 15438
rect 30472 14068 30524 14074
rect 30472 14010 30524 14016
rect 30378 12200 30434 12209
rect 30378 12135 30434 12144
rect 30576 11626 30604 15846
rect 30668 15162 30696 17575
rect 30944 17202 30972 17682
rect 30932 17196 30984 17202
rect 30932 17138 30984 17144
rect 30748 17060 30800 17066
rect 30748 17002 30800 17008
rect 30760 16250 30788 17002
rect 30932 16992 30984 16998
rect 30932 16934 30984 16940
rect 30840 16448 30892 16454
rect 30840 16390 30892 16396
rect 30748 16244 30800 16250
rect 30748 16186 30800 16192
rect 30760 15570 30788 16186
rect 30852 15978 30880 16390
rect 30944 16250 30972 16934
rect 31036 16250 31064 20198
rect 31116 19848 31168 19854
rect 31116 19790 31168 19796
rect 31128 19242 31156 19790
rect 31116 19236 31168 19242
rect 31116 19178 31168 19184
rect 31220 17542 31248 20334
rect 31312 19922 31340 24958
rect 31864 24682 31892 26200
rect 31852 24676 31904 24682
rect 31852 24618 31904 24624
rect 32312 24608 32364 24614
rect 32312 24550 32364 24556
rect 32324 24410 32352 24550
rect 32402 24440 32458 24449
rect 32312 24404 32364 24410
rect 32402 24375 32404 24384
rect 32312 24346 32364 24352
rect 32456 24375 32458 24384
rect 32404 24346 32456 24352
rect 31484 24336 31536 24342
rect 31484 24278 31536 24284
rect 31496 24206 31524 24278
rect 31484 24200 31536 24206
rect 31484 24142 31536 24148
rect 32128 24200 32180 24206
rect 32128 24142 32180 24148
rect 31944 24132 31996 24138
rect 31944 24074 31996 24080
rect 31576 23860 31628 23866
rect 31576 23802 31628 23808
rect 31668 23860 31720 23866
rect 31668 23802 31720 23808
rect 31588 23594 31616 23802
rect 31576 23588 31628 23594
rect 31576 23530 31628 23536
rect 31392 23520 31444 23526
rect 31392 23462 31444 23468
rect 31404 23186 31432 23462
rect 31392 23180 31444 23186
rect 31392 23122 31444 23128
rect 31404 22778 31432 23122
rect 31482 23080 31538 23089
rect 31482 23015 31538 23024
rect 31496 22778 31524 23015
rect 31392 22772 31444 22778
rect 31392 22714 31444 22720
rect 31484 22772 31536 22778
rect 31484 22714 31536 22720
rect 31576 22704 31628 22710
rect 31482 22672 31538 22681
rect 31680 22692 31708 23802
rect 31760 23520 31812 23526
rect 31760 23462 31812 23468
rect 31772 23186 31800 23462
rect 31760 23180 31812 23186
rect 31760 23122 31812 23128
rect 31956 23050 31984 24074
rect 32140 23322 32168 24142
rect 32128 23316 32180 23322
rect 32128 23258 32180 23264
rect 31944 23044 31996 23050
rect 31944 22986 31996 22992
rect 31628 22664 31708 22692
rect 31576 22646 31628 22652
rect 31482 22607 31538 22616
rect 31390 22128 31446 22137
rect 31390 22063 31446 22072
rect 31404 21962 31432 22063
rect 31392 21956 31444 21962
rect 31392 21898 31444 21904
rect 31392 21140 31444 21146
rect 31392 21082 31444 21088
rect 31404 20874 31432 21082
rect 31392 20868 31444 20874
rect 31392 20810 31444 20816
rect 31392 20460 31444 20466
rect 31392 20402 31444 20408
rect 31300 19916 31352 19922
rect 31300 19858 31352 19864
rect 31312 17626 31340 19858
rect 31404 18222 31432 20402
rect 31496 19922 31524 22607
rect 31576 22228 31628 22234
rect 31576 22170 31628 22176
rect 31588 21962 31616 22170
rect 31576 21956 31628 21962
rect 31576 21898 31628 21904
rect 31588 21622 31616 21898
rect 31576 21616 31628 21622
rect 31576 21558 31628 21564
rect 31576 21480 31628 21486
rect 31576 21422 31628 21428
rect 31484 19916 31536 19922
rect 31484 19858 31536 19864
rect 31588 19334 31616 21422
rect 31680 20534 31708 22664
rect 31852 22432 31904 22438
rect 31852 22374 31904 22380
rect 31864 21894 31892 22374
rect 32312 22092 32364 22098
rect 32312 22034 32364 22040
rect 31852 21888 31904 21894
rect 31852 21830 31904 21836
rect 32324 20942 32352 22034
rect 32404 21684 32456 21690
rect 32404 21626 32456 21632
rect 32312 20936 32364 20942
rect 32416 20913 32444 21626
rect 32508 21049 32536 26200
rect 33152 24698 33180 26200
rect 33152 24670 33364 24698
rect 32950 24508 33258 24517
rect 32950 24506 32956 24508
rect 33012 24506 33036 24508
rect 33092 24506 33116 24508
rect 33172 24506 33196 24508
rect 33252 24506 33258 24508
rect 33012 24454 33014 24506
rect 33194 24454 33196 24506
rect 32950 24452 32956 24454
rect 33012 24452 33036 24454
rect 33092 24452 33116 24454
rect 33172 24452 33196 24454
rect 33252 24452 33258 24454
rect 32950 24443 33258 24452
rect 32956 24064 33008 24070
rect 32956 24006 33008 24012
rect 32968 23866 32996 24006
rect 32956 23860 33008 23866
rect 32956 23802 33008 23808
rect 32680 23724 32732 23730
rect 32680 23666 32732 23672
rect 32588 23656 32640 23662
rect 32588 23598 32640 23604
rect 32600 22953 32628 23598
rect 32586 22944 32642 22953
rect 32586 22879 32642 22888
rect 32600 22234 32628 22879
rect 32588 22228 32640 22234
rect 32588 22170 32640 22176
rect 32692 21894 32720 23666
rect 32950 23420 33258 23429
rect 32950 23418 32956 23420
rect 33012 23418 33036 23420
rect 33092 23418 33116 23420
rect 33172 23418 33196 23420
rect 33252 23418 33258 23420
rect 33012 23366 33014 23418
rect 33194 23366 33196 23418
rect 32950 23364 32956 23366
rect 33012 23364 33036 23366
rect 33092 23364 33116 23366
rect 33172 23364 33196 23366
rect 33252 23364 33258 23366
rect 32950 23355 33258 23364
rect 32864 22432 32916 22438
rect 32864 22374 32916 22380
rect 32680 21888 32732 21894
rect 32680 21830 32732 21836
rect 32876 21622 32904 22374
rect 32950 22332 33258 22341
rect 32950 22330 32956 22332
rect 33012 22330 33036 22332
rect 33092 22330 33116 22332
rect 33172 22330 33196 22332
rect 33252 22330 33258 22332
rect 33012 22278 33014 22330
rect 33194 22278 33196 22330
rect 32950 22276 32956 22278
rect 33012 22276 33036 22278
rect 33092 22276 33116 22278
rect 33172 22276 33196 22278
rect 33252 22276 33258 22278
rect 32950 22267 33258 22276
rect 33336 22234 33364 24670
rect 33796 24449 33824 26200
rect 34060 24608 34112 24614
rect 34060 24550 34112 24556
rect 33782 24440 33838 24449
rect 33782 24375 33838 24384
rect 34072 24274 34100 24550
rect 34440 24342 34468 26200
rect 34796 24744 34848 24750
rect 34796 24686 34848 24692
rect 34886 24712 34942 24721
rect 34428 24336 34480 24342
rect 34428 24278 34480 24284
rect 34060 24268 34112 24274
rect 34060 24210 34112 24216
rect 34152 24132 34204 24138
rect 34152 24074 34204 24080
rect 33600 23656 33652 23662
rect 33600 23598 33652 23604
rect 33612 23168 33640 23598
rect 33966 23488 34022 23497
rect 33966 23423 34022 23432
rect 33980 23322 34008 23423
rect 33968 23316 34020 23322
rect 33968 23258 34020 23264
rect 33692 23180 33744 23186
rect 33612 23140 33692 23168
rect 33692 23122 33744 23128
rect 33600 23044 33652 23050
rect 33600 22986 33652 22992
rect 33612 22438 33640 22986
rect 33704 22642 33732 23122
rect 33784 22976 33836 22982
rect 33784 22918 33836 22924
rect 33876 22976 33928 22982
rect 33876 22918 33928 22924
rect 33692 22636 33744 22642
rect 33692 22578 33744 22584
rect 33600 22432 33652 22438
rect 33600 22374 33652 22380
rect 33324 22228 33376 22234
rect 33324 22170 33376 22176
rect 33048 22024 33100 22030
rect 33046 21992 33048 22001
rect 33100 21992 33102 22001
rect 33046 21927 33102 21936
rect 33416 21888 33468 21894
rect 33416 21830 33468 21836
rect 33508 21888 33560 21894
rect 33508 21830 33560 21836
rect 33428 21690 33456 21830
rect 33416 21684 33468 21690
rect 33416 21626 33468 21632
rect 32864 21616 32916 21622
rect 32864 21558 32916 21564
rect 32680 21344 32732 21350
rect 32680 21286 32732 21292
rect 32494 21040 32550 21049
rect 32494 20975 32550 20984
rect 32312 20878 32364 20884
rect 32402 20904 32458 20913
rect 32324 20602 32352 20878
rect 32402 20839 32458 20848
rect 32312 20596 32364 20602
rect 32312 20538 32364 20544
rect 31668 20528 31720 20534
rect 31668 20470 31720 20476
rect 32324 20398 32352 20538
rect 32312 20392 32364 20398
rect 31850 20360 31906 20369
rect 32312 20334 32364 20340
rect 31850 20295 31852 20304
rect 31904 20295 31906 20304
rect 31852 20266 31904 20272
rect 31864 19854 31892 20266
rect 31944 19984 31996 19990
rect 31944 19926 31996 19932
rect 31852 19848 31904 19854
rect 31852 19790 31904 19796
rect 31668 19712 31720 19718
rect 31668 19654 31720 19660
rect 31496 19310 31616 19334
rect 31484 19306 31616 19310
rect 31484 19304 31536 19306
rect 31484 19246 31536 19252
rect 31680 18630 31708 19654
rect 31956 18834 31984 19926
rect 32220 19780 32272 19786
rect 32220 19722 32272 19728
rect 32128 19712 32180 19718
rect 32128 19654 32180 19660
rect 31944 18828 31996 18834
rect 31944 18770 31996 18776
rect 31668 18624 31720 18630
rect 31668 18566 31720 18572
rect 31852 18624 31904 18630
rect 31852 18566 31904 18572
rect 32036 18624 32088 18630
rect 32036 18566 32088 18572
rect 31392 18216 31444 18222
rect 31392 18158 31444 18164
rect 31312 17598 31524 17626
rect 31496 17542 31524 17598
rect 31208 17536 31260 17542
rect 31208 17478 31260 17484
rect 31392 17536 31444 17542
rect 31392 17478 31444 17484
rect 31484 17536 31536 17542
rect 31484 17478 31536 17484
rect 31208 17196 31260 17202
rect 31208 17138 31260 17144
rect 30932 16244 30984 16250
rect 30932 16186 30984 16192
rect 31024 16244 31076 16250
rect 31024 16186 31076 16192
rect 30840 15972 30892 15978
rect 30840 15914 30892 15920
rect 30748 15564 30800 15570
rect 30748 15506 30800 15512
rect 30656 15156 30708 15162
rect 30656 15098 30708 15104
rect 30760 14482 30788 15506
rect 31116 15360 31168 15366
rect 31116 15302 31168 15308
rect 30932 15156 30984 15162
rect 30932 15098 30984 15104
rect 30944 15026 30972 15098
rect 30932 15020 30984 15026
rect 30932 14962 30984 14968
rect 30840 14952 30892 14958
rect 30840 14894 30892 14900
rect 30748 14476 30800 14482
rect 30748 14418 30800 14424
rect 30852 13734 30880 14894
rect 31128 14278 31156 15302
rect 31116 14272 31168 14278
rect 31116 14214 31168 14220
rect 31114 14104 31170 14113
rect 31114 14039 31116 14048
rect 31168 14039 31170 14048
rect 31116 14010 31168 14016
rect 31220 13734 31248 17138
rect 31300 16448 31352 16454
rect 31300 16390 31352 16396
rect 31312 15162 31340 16390
rect 31300 15156 31352 15162
rect 31300 15098 31352 15104
rect 31404 14906 31432 17478
rect 31668 17128 31720 17134
rect 31668 17070 31720 17076
rect 31680 16658 31708 17070
rect 31668 16652 31720 16658
rect 31668 16594 31720 16600
rect 31864 16522 31892 18566
rect 31944 17740 31996 17746
rect 31944 17682 31996 17688
rect 31852 16516 31904 16522
rect 31852 16458 31904 16464
rect 31484 16108 31536 16114
rect 31484 16050 31536 16056
rect 31496 15910 31524 16050
rect 31852 16040 31904 16046
rect 31772 15988 31852 15994
rect 31772 15982 31904 15988
rect 31772 15966 31892 15982
rect 31484 15904 31536 15910
rect 31484 15846 31536 15852
rect 31668 15904 31720 15910
rect 31668 15846 31720 15852
rect 31496 15570 31524 15846
rect 31484 15564 31536 15570
rect 31484 15506 31536 15512
rect 31680 15366 31708 15846
rect 31484 15360 31536 15366
rect 31484 15302 31536 15308
rect 31668 15360 31720 15366
rect 31772 15348 31800 15966
rect 31772 15320 31892 15348
rect 31668 15302 31720 15308
rect 31496 15094 31524 15302
rect 31576 15156 31628 15162
rect 31576 15098 31628 15104
rect 31484 15088 31536 15094
rect 31484 15030 31536 15036
rect 31404 14878 31524 14906
rect 31392 14000 31444 14006
rect 31392 13942 31444 13948
rect 31300 13796 31352 13802
rect 31300 13738 31352 13744
rect 30840 13728 30892 13734
rect 30840 13670 30892 13676
rect 31208 13728 31260 13734
rect 31208 13670 31260 13676
rect 30840 13456 30892 13462
rect 30840 13398 30892 13404
rect 30564 11620 30616 11626
rect 30564 11562 30616 11568
rect 30748 11076 30800 11082
rect 30748 11018 30800 11024
rect 30380 11008 30432 11014
rect 30380 10950 30432 10956
rect 30288 10736 30340 10742
rect 30288 10678 30340 10684
rect 30300 10198 30328 10678
rect 30392 10606 30420 10950
rect 30380 10600 30432 10606
rect 30380 10542 30432 10548
rect 30472 10600 30524 10606
rect 30472 10542 30524 10548
rect 30288 10192 30340 10198
rect 30288 10134 30340 10140
rect 30380 10056 30432 10062
rect 30380 9998 30432 10004
rect 30104 9988 30156 9994
rect 30104 9930 30156 9936
rect 30392 9382 30420 9998
rect 30380 9376 30432 9382
rect 30380 9318 30432 9324
rect 30392 9042 30420 9318
rect 30484 9110 30512 10542
rect 30656 9988 30708 9994
rect 30656 9930 30708 9936
rect 30564 9648 30616 9654
rect 30564 9590 30616 9596
rect 30472 9104 30524 9110
rect 30472 9046 30524 9052
rect 30380 9036 30432 9042
rect 30380 8978 30432 8984
rect 30576 8838 30604 9590
rect 30668 9518 30696 9930
rect 30656 9512 30708 9518
rect 30656 9454 30708 9460
rect 30380 8832 30432 8838
rect 30380 8774 30432 8780
rect 30564 8832 30616 8838
rect 30564 8774 30616 8780
rect 30392 8498 30420 8774
rect 30668 8634 30696 9454
rect 30656 8628 30708 8634
rect 30656 8570 30708 8576
rect 30380 8492 30432 8498
rect 30380 8434 30432 8440
rect 30656 8492 30708 8498
rect 30656 8434 30708 8440
rect 29736 7948 29788 7954
rect 29736 7890 29788 7896
rect 30564 7948 30616 7954
rect 30564 7890 30616 7896
rect 30576 7478 30604 7890
rect 30668 7750 30696 8434
rect 30656 7744 30708 7750
rect 30656 7686 30708 7692
rect 30564 7472 30616 7478
rect 30564 7414 30616 7420
rect 29644 3120 29696 3126
rect 29644 3062 29696 3068
rect 28816 3052 28868 3058
rect 28816 2994 28868 3000
rect 29656 2990 29684 3062
rect 30668 2990 30696 7686
rect 30760 6118 30788 11018
rect 30852 9466 30880 13398
rect 31024 12368 31076 12374
rect 31024 12310 31076 12316
rect 30932 12096 30984 12102
rect 30932 12038 30984 12044
rect 30944 11830 30972 12038
rect 30932 11824 30984 11830
rect 30932 11766 30984 11772
rect 31036 11218 31064 12310
rect 31116 11756 31168 11762
rect 31116 11698 31168 11704
rect 31024 11212 31076 11218
rect 31024 11154 31076 11160
rect 31128 10810 31156 11698
rect 31312 11694 31340 13738
rect 31404 12850 31432 13942
rect 31392 12844 31444 12850
rect 31392 12786 31444 12792
rect 31404 12238 31432 12786
rect 31392 12232 31444 12238
rect 31392 12174 31444 12180
rect 31392 12096 31444 12102
rect 31392 12038 31444 12044
rect 31404 11830 31432 12038
rect 31392 11824 31444 11830
rect 31392 11766 31444 11772
rect 31496 11694 31524 14878
rect 31588 11898 31616 15098
rect 31760 14408 31812 14414
rect 31760 14350 31812 14356
rect 31772 12986 31800 14350
rect 31760 12980 31812 12986
rect 31760 12922 31812 12928
rect 31760 12844 31812 12850
rect 31760 12786 31812 12792
rect 31772 12442 31800 12786
rect 31760 12436 31812 12442
rect 31760 12378 31812 12384
rect 31760 12096 31812 12102
rect 31760 12038 31812 12044
rect 31772 11898 31800 12038
rect 31576 11892 31628 11898
rect 31576 11834 31628 11840
rect 31760 11892 31812 11898
rect 31760 11834 31812 11840
rect 31208 11688 31260 11694
rect 31206 11656 31208 11665
rect 31300 11688 31352 11694
rect 31260 11656 31262 11665
rect 31300 11630 31352 11636
rect 31484 11688 31536 11694
rect 31484 11630 31536 11636
rect 31206 11591 31262 11600
rect 31864 11234 31892 15320
rect 31956 14550 31984 17682
rect 32048 16697 32076 18566
rect 32140 18358 32168 19654
rect 32128 18352 32180 18358
rect 32128 18294 32180 18300
rect 32128 17536 32180 17542
rect 32128 17478 32180 17484
rect 32140 17202 32168 17478
rect 32128 17196 32180 17202
rect 32128 17138 32180 17144
rect 32034 16688 32090 16697
rect 32034 16623 32090 16632
rect 32128 16516 32180 16522
rect 32128 16458 32180 16464
rect 31944 14544 31996 14550
rect 31944 14486 31996 14492
rect 31772 11206 31892 11234
rect 31956 11218 31984 14486
rect 32140 14482 32168 16458
rect 32232 15570 32260 19722
rect 32324 19378 32352 20334
rect 32416 19718 32444 20839
rect 32404 19712 32456 19718
rect 32404 19654 32456 19660
rect 32692 19446 32720 21286
rect 32876 20874 32904 21558
rect 33416 21480 33468 21486
rect 33416 21422 33468 21428
rect 32950 21244 33258 21253
rect 32950 21242 32956 21244
rect 33012 21242 33036 21244
rect 33092 21242 33116 21244
rect 33172 21242 33196 21244
rect 33252 21242 33258 21244
rect 33012 21190 33014 21242
rect 33194 21190 33196 21242
rect 32950 21188 32956 21190
rect 33012 21188 33036 21190
rect 33092 21188 33116 21190
rect 33172 21188 33196 21190
rect 33252 21188 33258 21190
rect 32950 21179 33258 21188
rect 32772 20868 32824 20874
rect 32772 20810 32824 20816
rect 32864 20868 32916 20874
rect 32864 20810 32916 20816
rect 33232 20868 33284 20874
rect 33232 20810 33284 20816
rect 32784 20754 32812 20810
rect 32784 20726 33180 20754
rect 33152 20346 33180 20726
rect 33244 20534 33272 20810
rect 33232 20528 33284 20534
rect 33232 20470 33284 20476
rect 33152 20318 33364 20346
rect 32950 20156 33258 20165
rect 32950 20154 32956 20156
rect 33012 20154 33036 20156
rect 33092 20154 33116 20156
rect 33172 20154 33196 20156
rect 33252 20154 33258 20156
rect 33012 20102 33014 20154
rect 33194 20102 33196 20154
rect 32950 20100 32956 20102
rect 33012 20100 33036 20102
rect 33092 20100 33116 20102
rect 33172 20100 33196 20102
rect 33252 20100 33258 20102
rect 32950 20091 33258 20100
rect 32772 19712 32824 19718
rect 32772 19654 32824 19660
rect 32784 19446 32812 19654
rect 32864 19508 32916 19514
rect 32864 19450 32916 19456
rect 32680 19440 32732 19446
rect 32680 19382 32732 19388
rect 32772 19440 32824 19446
rect 32772 19382 32824 19388
rect 32312 19372 32364 19378
rect 32312 19314 32364 19320
rect 32588 19372 32640 19378
rect 32588 19314 32640 19320
rect 32600 18766 32628 19314
rect 32772 19168 32824 19174
rect 32772 19110 32824 19116
rect 32588 18760 32640 18766
rect 32588 18702 32640 18708
rect 32588 18352 32640 18358
rect 32588 18294 32640 18300
rect 32496 18148 32548 18154
rect 32496 18090 32548 18096
rect 32508 17610 32536 18090
rect 32600 17882 32628 18294
rect 32680 18284 32732 18290
rect 32680 18226 32732 18232
rect 32588 17876 32640 17882
rect 32588 17818 32640 17824
rect 32496 17604 32548 17610
rect 32496 17546 32548 17552
rect 32312 17332 32364 17338
rect 32312 17274 32364 17280
rect 32404 17332 32456 17338
rect 32404 17274 32456 17280
rect 32220 15564 32272 15570
rect 32220 15506 32272 15512
rect 32128 14476 32180 14482
rect 32128 14418 32180 14424
rect 32128 14272 32180 14278
rect 32128 14214 32180 14220
rect 32140 11898 32168 14214
rect 32324 13954 32352 17274
rect 32416 16522 32444 17274
rect 32508 17270 32536 17546
rect 32692 17542 32720 18226
rect 32680 17536 32732 17542
rect 32680 17478 32732 17484
rect 32496 17264 32548 17270
rect 32496 17206 32548 17212
rect 32588 17264 32640 17270
rect 32588 17206 32640 17212
rect 32508 16658 32536 17206
rect 32496 16652 32548 16658
rect 32496 16594 32548 16600
rect 32404 16516 32456 16522
rect 32404 16458 32456 16464
rect 32600 15978 32628 17206
rect 32404 15972 32456 15978
rect 32404 15914 32456 15920
rect 32588 15972 32640 15978
rect 32588 15914 32640 15920
rect 32416 14362 32444 15914
rect 32494 15872 32550 15881
rect 32494 15807 32550 15816
rect 32508 14482 32536 15807
rect 32600 15706 32628 15914
rect 32588 15700 32640 15706
rect 32588 15642 32640 15648
rect 32692 15502 32720 17478
rect 32784 16046 32812 19110
rect 32772 16040 32824 16046
rect 32772 15982 32824 15988
rect 32680 15496 32732 15502
rect 32680 15438 32732 15444
rect 32680 15360 32732 15366
rect 32680 15302 32732 15308
rect 32496 14476 32548 14482
rect 32496 14418 32548 14424
rect 32416 14334 32628 14362
rect 32324 13926 32536 13954
rect 32312 13864 32364 13870
rect 32218 13832 32274 13841
rect 32312 13806 32364 13812
rect 32218 13767 32220 13776
rect 32272 13767 32274 13776
rect 32220 13738 32272 13744
rect 32324 13394 32352 13806
rect 32508 13394 32536 13926
rect 32312 13388 32364 13394
rect 32312 13330 32364 13336
rect 32496 13388 32548 13394
rect 32496 13330 32548 13336
rect 32324 12782 32352 13330
rect 32404 12980 32456 12986
rect 32404 12922 32456 12928
rect 32312 12776 32364 12782
rect 32312 12718 32364 12724
rect 32416 12170 32444 12922
rect 32404 12164 32456 12170
rect 32404 12106 32456 12112
rect 32128 11892 32180 11898
rect 32128 11834 32180 11840
rect 32034 11656 32090 11665
rect 32034 11591 32090 11600
rect 31944 11212 31996 11218
rect 31116 10804 31168 10810
rect 31116 10746 31168 10752
rect 31772 10742 31800 11206
rect 31944 11154 31996 11160
rect 31760 10736 31812 10742
rect 31760 10678 31812 10684
rect 31300 10464 31352 10470
rect 31300 10406 31352 10412
rect 31944 10464 31996 10470
rect 32048 10452 32076 11591
rect 32128 11212 32180 11218
rect 32128 11154 32180 11160
rect 31996 10424 32076 10452
rect 31944 10406 31996 10412
rect 31312 9654 31340 10406
rect 31760 10056 31812 10062
rect 31760 9998 31812 10004
rect 31482 9752 31538 9761
rect 31772 9722 31800 9998
rect 31482 9687 31484 9696
rect 31536 9687 31538 9696
rect 31760 9716 31812 9722
rect 31484 9658 31536 9664
rect 31588 9664 31760 9674
rect 31588 9658 31812 9664
rect 31300 9648 31352 9654
rect 31588 9646 31800 9658
rect 31588 9602 31616 9646
rect 31300 9590 31352 9596
rect 31404 9574 31616 9602
rect 31300 9512 31352 9518
rect 30852 9460 31300 9466
rect 30852 9454 31352 9460
rect 30852 9438 31340 9454
rect 31024 8900 31076 8906
rect 31024 8842 31076 8848
rect 31036 8634 31064 8842
rect 31404 8838 31432 9574
rect 31668 9444 31720 9450
rect 31668 9386 31720 9392
rect 31392 8832 31444 8838
rect 31392 8774 31444 8780
rect 31024 8628 31076 8634
rect 31024 8570 31076 8576
rect 31680 8498 31708 9386
rect 31956 9081 31984 10406
rect 32140 10266 32168 11154
rect 32312 11008 32364 11014
rect 32312 10950 32364 10956
rect 32220 10736 32272 10742
rect 32220 10678 32272 10684
rect 32232 10470 32260 10678
rect 32324 10538 32352 10950
rect 32416 10742 32444 12106
rect 32404 10736 32456 10742
rect 32404 10678 32456 10684
rect 32312 10532 32364 10538
rect 32312 10474 32364 10480
rect 32220 10464 32272 10470
rect 32220 10406 32272 10412
rect 32128 10260 32180 10266
rect 32128 10202 32180 10208
rect 32600 9908 32628 14334
rect 32692 13870 32720 15302
rect 32772 14816 32824 14822
rect 32772 14758 32824 14764
rect 32680 13864 32732 13870
rect 32680 13806 32732 13812
rect 32784 13530 32812 14758
rect 32876 14550 32904 19450
rect 32950 19068 33258 19077
rect 32950 19066 32956 19068
rect 33012 19066 33036 19068
rect 33092 19066 33116 19068
rect 33172 19066 33196 19068
rect 33252 19066 33258 19068
rect 33012 19014 33014 19066
rect 33194 19014 33196 19066
rect 32950 19012 32956 19014
rect 33012 19012 33036 19014
rect 33092 19012 33116 19014
rect 33172 19012 33196 19014
rect 33252 19012 33258 19014
rect 32950 19003 33258 19012
rect 33048 18964 33100 18970
rect 33048 18906 33100 18912
rect 32956 18624 33008 18630
rect 32954 18592 32956 18601
rect 33008 18592 33010 18601
rect 32954 18527 33010 18536
rect 33060 18290 33088 18906
rect 33140 18624 33192 18630
rect 33140 18566 33192 18572
rect 33152 18358 33180 18566
rect 33140 18352 33192 18358
rect 33140 18294 33192 18300
rect 33048 18284 33100 18290
rect 33048 18226 33100 18232
rect 32950 17980 33258 17989
rect 32950 17978 32956 17980
rect 33012 17978 33036 17980
rect 33092 17978 33116 17980
rect 33172 17978 33196 17980
rect 33252 17978 33258 17980
rect 33012 17926 33014 17978
rect 33194 17926 33196 17978
rect 32950 17924 32956 17926
rect 33012 17924 33036 17926
rect 33092 17924 33116 17926
rect 33172 17924 33196 17926
rect 33252 17924 33258 17926
rect 32950 17915 33258 17924
rect 33232 17740 33284 17746
rect 33336 17728 33364 20318
rect 33428 18222 33456 21422
rect 33520 20058 33548 21830
rect 33690 21584 33746 21593
rect 33600 21548 33652 21554
rect 33690 21519 33692 21528
rect 33600 21490 33652 21496
rect 33744 21519 33746 21528
rect 33692 21490 33744 21496
rect 33612 21321 33640 21490
rect 33598 21312 33654 21321
rect 33598 21247 33654 21256
rect 33508 20052 33560 20058
rect 33508 19994 33560 20000
rect 33508 19916 33560 19922
rect 33508 19858 33560 19864
rect 33416 18216 33468 18222
rect 33416 18158 33468 18164
rect 33284 17700 33364 17728
rect 33232 17682 33284 17688
rect 33428 17660 33456 18158
rect 33336 17632 33456 17660
rect 33336 17338 33364 17632
rect 33416 17536 33468 17542
rect 33416 17478 33468 17484
rect 33324 17332 33376 17338
rect 33324 17274 33376 17280
rect 32950 16892 33258 16901
rect 32950 16890 32956 16892
rect 33012 16890 33036 16892
rect 33092 16890 33116 16892
rect 33172 16890 33196 16892
rect 33252 16890 33258 16892
rect 33012 16838 33014 16890
rect 33194 16838 33196 16890
rect 32950 16836 32956 16838
rect 33012 16836 33036 16838
rect 33092 16836 33116 16838
rect 33172 16836 33196 16838
rect 33252 16836 33258 16838
rect 32950 16827 33258 16836
rect 33428 16182 33456 17478
rect 33416 16176 33468 16182
rect 33416 16118 33468 16124
rect 33324 16108 33376 16114
rect 33324 16050 33376 16056
rect 32950 15804 33258 15813
rect 32950 15802 32956 15804
rect 33012 15802 33036 15804
rect 33092 15802 33116 15804
rect 33172 15802 33196 15804
rect 33252 15802 33258 15804
rect 33012 15750 33014 15802
rect 33194 15750 33196 15802
rect 32950 15748 32956 15750
rect 33012 15748 33036 15750
rect 33092 15748 33116 15750
rect 33172 15748 33196 15750
rect 33252 15748 33258 15750
rect 32950 15739 33258 15748
rect 32950 14716 33258 14725
rect 32950 14714 32956 14716
rect 33012 14714 33036 14716
rect 33092 14714 33116 14716
rect 33172 14714 33196 14716
rect 33252 14714 33258 14716
rect 33012 14662 33014 14714
rect 33194 14662 33196 14714
rect 32950 14660 32956 14662
rect 33012 14660 33036 14662
rect 33092 14660 33116 14662
rect 33172 14660 33196 14662
rect 33252 14660 33258 14662
rect 32950 14651 33258 14660
rect 32864 14544 32916 14550
rect 32864 14486 32916 14492
rect 33336 14362 33364 16050
rect 33416 15904 33468 15910
rect 33416 15846 33468 15852
rect 33428 14414 33456 15846
rect 33520 15570 33548 19858
rect 33796 19786 33824 22918
rect 33888 22710 33916 22918
rect 33980 22710 34008 23258
rect 33876 22704 33928 22710
rect 33968 22704 34020 22710
rect 33876 22646 33928 22652
rect 33966 22672 33968 22681
rect 34020 22672 34022 22681
rect 33966 22607 34022 22616
rect 34164 22098 34192 24074
rect 34428 23792 34480 23798
rect 34428 23734 34480 23740
rect 34336 23656 34388 23662
rect 34336 23598 34388 23604
rect 34348 22574 34376 23598
rect 34440 23050 34468 23734
rect 34428 23044 34480 23050
rect 34428 22986 34480 22992
rect 34440 22710 34468 22986
rect 34808 22982 34836 24686
rect 34886 24647 34942 24656
rect 34796 22976 34848 22982
rect 34796 22918 34848 22924
rect 34900 22817 34928 24647
rect 34980 23520 35032 23526
rect 34980 23462 35032 23468
rect 34992 23254 35020 23462
rect 35084 23322 35112 26200
rect 35440 24812 35492 24818
rect 35440 24754 35492 24760
rect 35348 24268 35400 24274
rect 35348 24210 35400 24216
rect 35256 24064 35308 24070
rect 35254 24032 35256 24041
rect 35308 24032 35310 24041
rect 35254 23967 35310 23976
rect 35360 23798 35388 24210
rect 35452 24070 35480 24754
rect 35532 24268 35584 24274
rect 35532 24210 35584 24216
rect 35440 24064 35492 24070
rect 35440 24006 35492 24012
rect 35348 23792 35400 23798
rect 35348 23734 35400 23740
rect 35544 23497 35572 24210
rect 35530 23488 35586 23497
rect 35530 23423 35586 23432
rect 35728 23361 35756 26200
rect 36084 24200 36136 24206
rect 36084 24142 36136 24148
rect 35992 24064 36044 24070
rect 35992 24006 36044 24012
rect 35808 23724 35860 23730
rect 35808 23666 35860 23672
rect 35714 23352 35770 23361
rect 35072 23316 35124 23322
rect 35714 23287 35770 23296
rect 35072 23258 35124 23264
rect 34980 23248 35032 23254
rect 34980 23190 35032 23196
rect 35072 23180 35124 23186
rect 35124 23140 35756 23168
rect 35072 23122 35124 23128
rect 34980 22976 35032 22982
rect 34980 22918 35032 22924
rect 35256 22976 35308 22982
rect 35256 22918 35308 22924
rect 34886 22808 34942 22817
rect 34886 22743 34942 22752
rect 34428 22704 34480 22710
rect 34428 22646 34480 22652
rect 34336 22568 34388 22574
rect 34242 22536 34298 22545
rect 34336 22510 34388 22516
rect 34242 22471 34298 22480
rect 34152 22092 34204 22098
rect 34152 22034 34204 22040
rect 34060 21004 34112 21010
rect 34060 20946 34112 20952
rect 34072 20602 34100 20946
rect 34256 20806 34284 22471
rect 34348 22166 34376 22510
rect 34440 22166 34468 22646
rect 34336 22160 34388 22166
rect 34336 22102 34388 22108
rect 34428 22160 34480 22166
rect 34428 22102 34480 22108
rect 34428 22024 34480 22030
rect 34428 21966 34480 21972
rect 34336 21344 34388 21350
rect 34336 21286 34388 21292
rect 34348 21078 34376 21286
rect 34336 21072 34388 21078
rect 34336 21014 34388 21020
rect 34244 20800 34296 20806
rect 34164 20760 34244 20788
rect 34060 20596 34112 20602
rect 34060 20538 34112 20544
rect 33784 19780 33836 19786
rect 33784 19722 33836 19728
rect 33968 19508 34020 19514
rect 33968 19450 34020 19456
rect 33980 19417 34008 19450
rect 33966 19408 34022 19417
rect 33966 19343 34022 19352
rect 33968 18964 34020 18970
rect 33704 18924 33968 18952
rect 33704 18630 33732 18924
rect 33968 18906 34020 18912
rect 34164 18834 34192 20760
rect 34244 20742 34296 20748
rect 34440 20641 34468 21966
rect 34794 21720 34850 21729
rect 34900 21690 34928 22743
rect 34794 21655 34850 21664
rect 34888 21684 34940 21690
rect 34808 21554 34836 21655
rect 34888 21626 34940 21632
rect 34796 21548 34848 21554
rect 34796 21490 34848 21496
rect 34808 21457 34836 21490
rect 34794 21448 34850 21457
rect 34794 21383 34850 21392
rect 34520 21344 34572 21350
rect 34520 21286 34572 21292
rect 34532 21146 34560 21286
rect 34520 21140 34572 21146
rect 34520 21082 34572 21088
rect 34704 20800 34756 20806
rect 34704 20742 34756 20748
rect 34426 20632 34482 20641
rect 34610 20632 34666 20641
rect 34426 20567 34482 20576
rect 34532 20590 34610 20618
rect 34428 20528 34480 20534
rect 34532 20516 34560 20590
rect 34716 20602 34744 20742
rect 34610 20567 34666 20576
rect 34704 20596 34756 20602
rect 34704 20538 34756 20544
rect 34480 20488 34560 20516
rect 34612 20528 34664 20534
rect 34428 20470 34480 20476
rect 34612 20470 34664 20476
rect 34624 20058 34652 20470
rect 34612 20052 34664 20058
rect 34612 19994 34664 20000
rect 34518 19816 34574 19825
rect 34518 19751 34574 19760
rect 34336 19712 34388 19718
rect 34336 19654 34388 19660
rect 34244 19372 34296 19378
rect 34244 19314 34296 19320
rect 34152 18828 34204 18834
rect 34152 18770 34204 18776
rect 34256 18630 34284 19314
rect 34348 19122 34376 19654
rect 34428 19508 34480 19514
rect 34532 19496 34560 19751
rect 34480 19468 34560 19496
rect 34428 19450 34480 19456
rect 34348 19094 34468 19122
rect 34336 18964 34388 18970
rect 34336 18906 34388 18912
rect 33692 18624 33744 18630
rect 34152 18624 34204 18630
rect 33692 18566 33744 18572
rect 34150 18592 34152 18601
rect 34244 18624 34296 18630
rect 34204 18592 34206 18601
rect 34244 18566 34296 18572
rect 34150 18527 34206 18536
rect 33876 18216 33928 18222
rect 33876 18158 33928 18164
rect 33888 17134 33916 18158
rect 34152 17876 34204 17882
rect 34152 17818 34204 17824
rect 34164 17270 34192 17818
rect 34152 17264 34204 17270
rect 34152 17206 34204 17212
rect 33876 17128 33928 17134
rect 33876 17070 33928 17076
rect 33968 16992 34020 16998
rect 33968 16934 34020 16940
rect 33980 16250 34008 16934
rect 34164 16726 34192 17206
rect 34152 16720 34204 16726
rect 34152 16662 34204 16668
rect 34060 16516 34112 16522
rect 34060 16458 34112 16464
rect 33968 16244 34020 16250
rect 33968 16186 34020 16192
rect 33508 15564 33560 15570
rect 33508 15506 33560 15512
rect 33876 15360 33928 15366
rect 33876 15302 33928 15308
rect 33888 15162 33916 15302
rect 33876 15156 33928 15162
rect 33876 15098 33928 15104
rect 34072 14958 34100 16458
rect 34164 15706 34192 16662
rect 34152 15700 34204 15706
rect 34152 15642 34204 15648
rect 34152 15564 34204 15570
rect 34152 15506 34204 15512
rect 33876 14952 33928 14958
rect 33876 14894 33928 14900
rect 33968 14952 34020 14958
rect 33968 14894 34020 14900
rect 34060 14952 34112 14958
rect 34060 14894 34112 14900
rect 33244 14334 33364 14362
rect 33416 14408 33468 14414
rect 33416 14350 33468 14356
rect 33600 14340 33652 14346
rect 33244 14278 33272 14334
rect 33600 14282 33652 14288
rect 33232 14272 33284 14278
rect 33232 14214 33284 14220
rect 32864 14000 32916 14006
rect 32864 13942 32916 13948
rect 32772 13524 32824 13530
rect 32772 13466 32824 13472
rect 32876 13394 32904 13942
rect 33324 13728 33376 13734
rect 33324 13670 33376 13676
rect 32950 13628 33258 13637
rect 32950 13626 32956 13628
rect 33012 13626 33036 13628
rect 33092 13626 33116 13628
rect 33172 13626 33196 13628
rect 33252 13626 33258 13628
rect 33012 13574 33014 13626
rect 33194 13574 33196 13626
rect 32950 13572 32956 13574
rect 33012 13572 33036 13574
rect 33092 13572 33116 13574
rect 33172 13572 33196 13574
rect 33252 13572 33258 13574
rect 32950 13563 33258 13572
rect 33336 13530 33364 13670
rect 33324 13524 33376 13530
rect 33324 13466 33376 13472
rect 32772 13388 32824 13394
rect 32772 13330 32824 13336
rect 32864 13388 32916 13394
rect 32864 13330 32916 13336
rect 32784 12986 32812 13330
rect 33612 13326 33640 14282
rect 33690 13832 33746 13841
rect 33888 13802 33916 14894
rect 33980 14618 34008 14894
rect 33968 14612 34020 14618
rect 33968 14554 34020 14560
rect 33690 13767 33746 13776
rect 33876 13796 33928 13802
rect 33704 13734 33732 13767
rect 33876 13738 33928 13744
rect 33692 13728 33744 13734
rect 33692 13670 33744 13676
rect 33692 13456 33744 13462
rect 33692 13398 33744 13404
rect 33324 13320 33376 13326
rect 33600 13320 33652 13326
rect 33324 13262 33376 13268
rect 33428 13280 33600 13308
rect 32772 12980 32824 12986
rect 32772 12922 32824 12928
rect 33336 12646 33364 13262
rect 33324 12640 33376 12646
rect 33324 12582 33376 12588
rect 32950 12540 33258 12549
rect 32950 12538 32956 12540
rect 33012 12538 33036 12540
rect 33092 12538 33116 12540
rect 33172 12538 33196 12540
rect 33252 12538 33258 12540
rect 33012 12486 33014 12538
rect 33194 12486 33196 12538
rect 32950 12484 32956 12486
rect 33012 12484 33036 12486
rect 33092 12484 33116 12486
rect 33172 12484 33196 12486
rect 33252 12484 33258 12486
rect 32950 12475 33258 12484
rect 33324 12096 33376 12102
rect 33324 12038 33376 12044
rect 32864 11688 32916 11694
rect 32784 11648 32864 11676
rect 32784 11218 32812 11648
rect 32864 11630 32916 11636
rect 32950 11452 33258 11461
rect 32950 11450 32956 11452
rect 33012 11450 33036 11452
rect 33092 11450 33116 11452
rect 33172 11450 33196 11452
rect 33252 11450 33258 11452
rect 33012 11398 33014 11450
rect 33194 11398 33196 11450
rect 32950 11396 32956 11398
rect 33012 11396 33036 11398
rect 33092 11396 33116 11398
rect 33172 11396 33196 11398
rect 33252 11396 33258 11398
rect 32950 11387 33258 11396
rect 32772 11212 32824 11218
rect 32772 11154 32824 11160
rect 32680 10668 32732 10674
rect 32680 10610 32732 10616
rect 32692 10130 32720 10610
rect 32680 10124 32732 10130
rect 32680 10066 32732 10072
rect 32680 9920 32732 9926
rect 32600 9880 32680 9908
rect 32680 9862 32732 9868
rect 32680 9716 32732 9722
rect 32680 9658 32732 9664
rect 32586 9480 32642 9489
rect 32586 9415 32642 9424
rect 32312 9104 32364 9110
rect 31942 9072 31998 9081
rect 32312 9046 32364 9052
rect 31942 9007 31998 9016
rect 30932 8492 30984 8498
rect 30932 8434 30984 8440
rect 31668 8492 31720 8498
rect 31668 8434 31720 8440
rect 30944 7546 30972 8434
rect 31484 8424 31536 8430
rect 31484 8366 31536 8372
rect 32220 8424 32272 8430
rect 32220 8366 32272 8372
rect 31496 7954 31524 8366
rect 32232 7954 32260 8366
rect 32324 8362 32352 9046
rect 32600 9042 32628 9415
rect 32692 9178 32720 9658
rect 32680 9172 32732 9178
rect 32680 9114 32732 9120
rect 32588 9036 32640 9042
rect 32588 8978 32640 8984
rect 32692 8974 32720 9114
rect 32680 8968 32732 8974
rect 32680 8910 32732 8916
rect 32588 8900 32640 8906
rect 32588 8842 32640 8848
rect 32600 8566 32628 8842
rect 32692 8566 32720 8910
rect 32588 8560 32640 8566
rect 32588 8502 32640 8508
rect 32680 8560 32732 8566
rect 32680 8502 32732 8508
rect 32680 8424 32732 8430
rect 32784 8412 32812 11154
rect 33232 11076 33284 11082
rect 33336 11064 33364 12038
rect 33428 11676 33456 13280
rect 33600 13262 33652 13268
rect 33508 12776 33560 12782
rect 33508 12718 33560 12724
rect 33520 11744 33548 12718
rect 33704 11898 33732 13398
rect 33876 13252 33928 13258
rect 33876 13194 33928 13200
rect 33784 12980 33836 12986
rect 33784 12922 33836 12928
rect 33692 11892 33744 11898
rect 33692 11834 33744 11840
rect 33520 11716 33732 11744
rect 33428 11648 33640 11676
rect 33416 11552 33468 11558
rect 33416 11494 33468 11500
rect 33428 11354 33456 11494
rect 33416 11348 33468 11354
rect 33416 11290 33468 11296
rect 33284 11036 33364 11064
rect 33232 11018 33284 11024
rect 32956 11008 33008 11014
rect 32956 10950 33008 10956
rect 32968 10810 32996 10950
rect 33336 10810 33364 11036
rect 32956 10804 33008 10810
rect 32956 10746 33008 10752
rect 33324 10804 33376 10810
rect 33324 10746 33376 10752
rect 32864 10464 32916 10470
rect 32864 10406 32916 10412
rect 32876 10146 32904 10406
rect 32950 10364 33258 10373
rect 32950 10362 32956 10364
rect 33012 10362 33036 10364
rect 33092 10362 33116 10364
rect 33172 10362 33196 10364
rect 33252 10362 33258 10364
rect 33012 10310 33014 10362
rect 33194 10310 33196 10362
rect 32950 10308 32956 10310
rect 33012 10308 33036 10310
rect 33092 10308 33116 10310
rect 33172 10308 33196 10310
rect 33252 10308 33258 10310
rect 32950 10299 33258 10308
rect 33048 10192 33100 10198
rect 32876 10140 33048 10146
rect 32876 10134 33100 10140
rect 32876 10118 33088 10134
rect 33232 10124 33284 10130
rect 33232 10066 33284 10072
rect 33140 9988 33192 9994
rect 33140 9930 33192 9936
rect 33152 9874 33180 9930
rect 32732 8384 32812 8412
rect 32876 9846 33180 9874
rect 32680 8366 32732 8372
rect 32312 8356 32364 8362
rect 32312 8298 32364 8304
rect 32772 8016 32824 8022
rect 32772 7958 32824 7964
rect 31484 7948 31536 7954
rect 31484 7890 31536 7896
rect 32220 7948 32272 7954
rect 32220 7890 32272 7896
rect 31392 7744 31444 7750
rect 31392 7686 31444 7692
rect 31404 7546 31432 7686
rect 30932 7540 30984 7546
rect 30932 7482 30984 7488
rect 31392 7540 31444 7546
rect 31392 7482 31444 7488
rect 30748 6112 30800 6118
rect 30748 6054 30800 6060
rect 31496 5302 31524 7890
rect 32784 7750 32812 7958
rect 32876 7818 32904 9846
rect 33244 9761 33272 10066
rect 33230 9752 33286 9761
rect 33336 9722 33364 10746
rect 33612 10418 33640 11648
rect 33704 10713 33732 11716
rect 33796 11150 33824 12922
rect 33888 12374 33916 13194
rect 34060 12980 34112 12986
rect 34060 12922 34112 12928
rect 34072 12850 34100 12922
rect 34060 12844 34112 12850
rect 34060 12786 34112 12792
rect 33876 12368 33928 12374
rect 33876 12310 33928 12316
rect 34060 12300 34112 12306
rect 34060 12242 34112 12248
rect 34072 11218 34100 12242
rect 34164 11218 34192 15506
rect 34060 11212 34112 11218
rect 34060 11154 34112 11160
rect 34152 11212 34204 11218
rect 34152 11154 34204 11160
rect 33784 11144 33836 11150
rect 33784 11086 33836 11092
rect 33690 10704 33746 10713
rect 33690 10639 33746 10648
rect 33874 10704 33930 10713
rect 33874 10639 33930 10648
rect 33612 10390 33824 10418
rect 33230 9687 33286 9696
rect 33324 9716 33376 9722
rect 33324 9658 33376 9664
rect 32950 9276 33258 9285
rect 32950 9274 32956 9276
rect 33012 9274 33036 9276
rect 33092 9274 33116 9276
rect 33172 9274 33196 9276
rect 33252 9274 33258 9276
rect 33012 9222 33014 9274
rect 33194 9222 33196 9274
rect 32950 9220 32956 9222
rect 33012 9220 33036 9222
rect 33092 9220 33116 9222
rect 33172 9220 33196 9222
rect 33252 9220 33258 9222
rect 32950 9211 33258 9220
rect 33046 9072 33102 9081
rect 33046 9007 33102 9016
rect 33060 8430 33088 9007
rect 33796 8838 33824 10390
rect 33888 8974 33916 10639
rect 34072 10130 34100 11154
rect 34060 10124 34112 10130
rect 34060 10066 34112 10072
rect 34072 9654 34100 10066
rect 34164 9654 34192 11154
rect 34256 10713 34284 18566
rect 34348 18222 34376 18906
rect 34440 18358 34468 19094
rect 34532 18970 34560 19468
rect 34624 19378 34652 19994
rect 34992 19854 35020 22918
rect 35072 22092 35124 22098
rect 35072 22034 35124 22040
rect 35084 21690 35112 22034
rect 35164 21888 35216 21894
rect 35164 21830 35216 21836
rect 35072 21684 35124 21690
rect 35072 21626 35124 21632
rect 35072 20868 35124 20874
rect 35072 20810 35124 20816
rect 35084 20330 35112 20810
rect 35072 20324 35124 20330
rect 35072 20266 35124 20272
rect 34980 19848 35032 19854
rect 34980 19790 35032 19796
rect 35072 19780 35124 19786
rect 35072 19722 35124 19728
rect 34612 19372 34664 19378
rect 34612 19314 34664 19320
rect 34520 18964 34572 18970
rect 34520 18906 34572 18912
rect 34428 18352 34480 18358
rect 34428 18294 34480 18300
rect 34336 18216 34388 18222
rect 34336 18158 34388 18164
rect 34440 18057 34468 18294
rect 34426 18048 34482 18057
rect 34426 17983 34482 17992
rect 34624 17898 34652 19314
rect 34704 18624 34756 18630
rect 34704 18566 34756 18572
rect 34348 17870 34652 17898
rect 34348 16017 34376 17870
rect 34612 17808 34664 17814
rect 34612 17750 34664 17756
rect 34624 17270 34652 17750
rect 34612 17264 34664 17270
rect 34612 17206 34664 17212
rect 34624 16794 34652 17206
rect 34612 16788 34664 16794
rect 34612 16730 34664 16736
rect 34428 16652 34480 16658
rect 34428 16594 34480 16600
rect 34334 16008 34390 16017
rect 34334 15943 34390 15952
rect 34440 15473 34468 16594
rect 34624 16590 34652 16730
rect 34520 16584 34572 16590
rect 34520 16526 34572 16532
rect 34612 16584 34664 16590
rect 34612 16526 34664 16532
rect 34532 16454 34560 16526
rect 34520 16448 34572 16454
rect 34520 16390 34572 16396
rect 34520 16244 34572 16250
rect 34520 16186 34572 16192
rect 34532 15502 34560 16186
rect 34520 15496 34572 15502
rect 34426 15464 34482 15473
rect 34520 15438 34572 15444
rect 34426 15399 34482 15408
rect 34624 15314 34652 16526
rect 34532 15286 34652 15314
rect 34336 14000 34388 14006
rect 34336 13942 34388 13948
rect 34348 13258 34376 13942
rect 34532 13784 34560 15286
rect 34716 15162 34744 18566
rect 34886 18048 34942 18057
rect 34886 17983 34942 17992
rect 34900 17882 34928 17983
rect 34888 17876 34940 17882
rect 34888 17818 34940 17824
rect 34980 17876 35032 17882
rect 34980 17818 35032 17824
rect 34888 17536 34940 17542
rect 34888 17478 34940 17484
rect 34900 17338 34928 17478
rect 34888 17332 34940 17338
rect 34888 17274 34940 17280
rect 34888 17128 34940 17134
rect 34888 17070 34940 17076
rect 34900 16046 34928 17070
rect 34992 16454 35020 17818
rect 34980 16448 35032 16454
rect 34980 16390 35032 16396
rect 34796 16040 34848 16046
rect 34796 15982 34848 15988
rect 34888 16040 34940 16046
rect 34888 15982 34940 15988
rect 34704 15156 34756 15162
rect 34704 15098 34756 15104
rect 34612 14952 34664 14958
rect 34612 14894 34664 14900
rect 34624 14278 34652 14894
rect 34612 14272 34664 14278
rect 34612 14214 34664 14220
rect 34440 13756 34560 13784
rect 34336 13252 34388 13258
rect 34336 13194 34388 13200
rect 34348 12646 34376 13194
rect 34440 12986 34468 13756
rect 34428 12980 34480 12986
rect 34428 12922 34480 12928
rect 34520 12708 34572 12714
rect 34520 12650 34572 12656
rect 34336 12640 34388 12646
rect 34336 12582 34388 12588
rect 34348 12102 34376 12582
rect 34426 12200 34482 12209
rect 34426 12135 34482 12144
rect 34336 12096 34388 12102
rect 34336 12038 34388 12044
rect 34440 11914 34468 12135
rect 34348 11886 34468 11914
rect 34242 10704 34298 10713
rect 34242 10639 34298 10648
rect 34060 9648 34112 9654
rect 34060 9590 34112 9596
rect 34152 9648 34204 9654
rect 34152 9590 34204 9596
rect 34060 9036 34112 9042
rect 34060 8978 34112 8984
rect 33876 8968 33928 8974
rect 33876 8910 33928 8916
rect 33784 8832 33836 8838
rect 33784 8774 33836 8780
rect 33048 8424 33100 8430
rect 33048 8366 33100 8372
rect 33600 8356 33652 8362
rect 33600 8298 33652 8304
rect 33612 8242 33640 8298
rect 33428 8214 33640 8242
rect 32950 8188 33258 8197
rect 32950 8186 32956 8188
rect 33012 8186 33036 8188
rect 33092 8186 33116 8188
rect 33172 8186 33196 8188
rect 33252 8186 33258 8188
rect 33012 8134 33014 8186
rect 33194 8134 33196 8186
rect 32950 8132 32956 8134
rect 33012 8132 33036 8134
rect 33092 8132 33116 8134
rect 33172 8132 33196 8134
rect 33252 8132 33258 8134
rect 32950 8123 33258 8132
rect 33428 8022 33456 8214
rect 33416 8016 33468 8022
rect 33416 7958 33468 7964
rect 32864 7812 32916 7818
rect 32864 7754 32916 7760
rect 32772 7744 32824 7750
rect 32772 7686 32824 7692
rect 32784 7206 32812 7686
rect 32772 7200 32824 7206
rect 32772 7142 32824 7148
rect 32950 7100 33258 7109
rect 32950 7098 32956 7100
rect 33012 7098 33036 7100
rect 33092 7098 33116 7100
rect 33172 7098 33196 7100
rect 33252 7098 33258 7100
rect 33012 7046 33014 7098
rect 33194 7046 33196 7098
rect 32950 7044 32956 7046
rect 33012 7044 33036 7046
rect 33092 7044 33116 7046
rect 33172 7044 33196 7046
rect 33252 7044 33258 7046
rect 32950 7035 33258 7044
rect 33796 6866 33824 8774
rect 34072 8634 34100 8978
rect 34164 8974 34192 9590
rect 34152 8968 34204 8974
rect 34152 8910 34204 8916
rect 34060 8628 34112 8634
rect 34060 8570 34112 8576
rect 33968 8288 34020 8294
rect 33968 8230 34020 8236
rect 33980 8090 34008 8230
rect 33968 8084 34020 8090
rect 33968 8026 34020 8032
rect 34348 7410 34376 11886
rect 34428 10260 34480 10266
rect 34428 10202 34480 10208
rect 34440 8498 34468 10202
rect 34532 8974 34560 12650
rect 34624 9625 34652 14214
rect 34808 13190 34836 15982
rect 34900 15502 34928 15982
rect 34888 15496 34940 15502
rect 34888 15438 34940 15444
rect 34900 14482 34928 15438
rect 35084 15144 35112 19722
rect 35176 17882 35204 21830
rect 35268 20874 35296 22918
rect 35348 22432 35400 22438
rect 35532 22432 35584 22438
rect 35438 22400 35494 22409
rect 35400 22380 35438 22386
rect 35348 22374 35438 22380
rect 35360 22358 35438 22374
rect 35532 22374 35584 22380
rect 35438 22335 35494 22344
rect 35256 20868 35308 20874
rect 35256 20810 35308 20816
rect 35268 20398 35296 20810
rect 35256 20392 35308 20398
rect 35256 20334 35308 20340
rect 35256 20256 35308 20262
rect 35256 20198 35308 20204
rect 35268 19310 35296 20198
rect 35452 19786 35480 22335
rect 35544 21894 35572 22374
rect 35728 22166 35756 23140
rect 35820 23050 35848 23666
rect 35900 23520 35952 23526
rect 35900 23462 35952 23468
rect 35912 23225 35940 23462
rect 35898 23216 35954 23225
rect 35898 23151 35954 23160
rect 35808 23044 35860 23050
rect 35808 22986 35860 22992
rect 35716 22160 35768 22166
rect 35622 22128 35678 22137
rect 35716 22102 35768 22108
rect 35622 22063 35624 22072
rect 35676 22063 35678 22072
rect 35624 22034 35676 22040
rect 35532 21888 35584 21894
rect 35532 21830 35584 21836
rect 35544 20398 35572 21830
rect 35728 21010 35756 22102
rect 35820 21010 35848 22986
rect 36004 22778 36032 24006
rect 36096 22778 36124 24142
rect 36176 24064 36228 24070
rect 36176 24006 36228 24012
rect 35992 22772 36044 22778
rect 35992 22714 36044 22720
rect 36084 22772 36136 22778
rect 36084 22714 36136 22720
rect 35992 22636 36044 22642
rect 35992 22578 36044 22584
rect 35900 21684 35952 21690
rect 35900 21626 35952 21632
rect 35912 21185 35940 21626
rect 35898 21176 35954 21185
rect 35898 21111 35954 21120
rect 35716 21004 35768 21010
rect 35716 20946 35768 20952
rect 35808 21004 35860 21010
rect 35808 20946 35860 20952
rect 35532 20392 35584 20398
rect 35532 20334 35584 20340
rect 35532 19916 35584 19922
rect 35532 19858 35584 19864
rect 35440 19780 35492 19786
rect 35440 19722 35492 19728
rect 35256 19304 35308 19310
rect 35254 19272 35256 19281
rect 35308 19272 35310 19281
rect 35254 19207 35310 19216
rect 35268 18034 35296 19207
rect 35348 18692 35400 18698
rect 35348 18634 35400 18640
rect 35360 18222 35388 18634
rect 35348 18216 35400 18222
rect 35348 18158 35400 18164
rect 35268 18006 35388 18034
rect 35164 17876 35216 17882
rect 35164 17818 35216 17824
rect 35164 17740 35216 17746
rect 35216 17700 35296 17728
rect 35164 17682 35216 17688
rect 35268 17542 35296 17700
rect 35256 17536 35308 17542
rect 35256 17478 35308 17484
rect 35164 16244 35216 16250
rect 35164 16186 35216 16192
rect 34992 15116 35112 15144
rect 34888 14476 34940 14482
rect 34888 14418 34940 14424
rect 34992 13938 35020 15116
rect 35176 14346 35204 16186
rect 35164 14340 35216 14346
rect 35164 14282 35216 14288
rect 34980 13932 35032 13938
rect 34980 13874 35032 13880
rect 35176 13818 35204 14282
rect 34900 13790 35204 13818
rect 34796 13184 34848 13190
rect 34796 13126 34848 13132
rect 34900 13002 34928 13790
rect 35072 13388 35124 13394
rect 35072 13330 35124 13336
rect 34716 12974 34928 13002
rect 34716 12442 34744 12974
rect 34888 12912 34940 12918
rect 34888 12854 34940 12860
rect 34704 12436 34756 12442
rect 34704 12378 34756 12384
rect 34796 12300 34848 12306
rect 34796 12242 34848 12248
rect 34808 11898 34836 12242
rect 34900 12238 34928 12854
rect 35084 12288 35112 13330
rect 35164 12844 35216 12850
rect 35268 12832 35296 17478
rect 35360 17270 35388 18006
rect 35544 17728 35572 19858
rect 35624 19780 35676 19786
rect 35624 19722 35676 19728
rect 35636 19514 35664 19722
rect 35624 19508 35676 19514
rect 35624 19450 35676 19456
rect 35622 18592 35678 18601
rect 35622 18527 35678 18536
rect 35452 17700 35572 17728
rect 35452 17542 35480 17700
rect 35636 17660 35664 18527
rect 35728 18358 35756 20946
rect 35820 20874 35848 20946
rect 35808 20868 35860 20874
rect 35808 20810 35860 20816
rect 35808 20256 35860 20262
rect 35808 20198 35860 20204
rect 35820 20058 35848 20198
rect 35808 20052 35860 20058
rect 35808 19994 35860 20000
rect 35808 19712 35860 19718
rect 35808 19654 35860 19660
rect 35716 18352 35768 18358
rect 35716 18294 35768 18300
rect 35728 17746 35756 18294
rect 35716 17740 35768 17746
rect 35716 17682 35768 17688
rect 35544 17632 35664 17660
rect 35440 17536 35492 17542
rect 35440 17478 35492 17484
rect 35348 17264 35400 17270
rect 35348 17206 35400 17212
rect 35440 16176 35492 16182
rect 35440 16118 35492 16124
rect 35348 14952 35400 14958
rect 35348 14894 35400 14900
rect 35360 14618 35388 14894
rect 35348 14612 35400 14618
rect 35348 14554 35400 14560
rect 35348 13796 35400 13802
rect 35348 13738 35400 13744
rect 35360 13394 35388 13738
rect 35348 13388 35400 13394
rect 35348 13330 35400 13336
rect 35346 13288 35402 13297
rect 35346 13223 35348 13232
rect 35400 13223 35402 13232
rect 35348 13194 35400 13200
rect 35216 12804 35296 12832
rect 35164 12786 35216 12792
rect 35176 12434 35204 12786
rect 35176 12406 35388 12434
rect 35084 12260 35296 12288
rect 34888 12232 34940 12238
rect 34888 12174 34940 12180
rect 35072 12164 35124 12170
rect 35072 12106 35124 12112
rect 34796 11892 34848 11898
rect 34796 11834 34848 11840
rect 34610 9616 34666 9625
rect 34610 9551 34666 9560
rect 34520 8968 34572 8974
rect 34520 8910 34572 8916
rect 34428 8492 34480 8498
rect 34428 8434 34480 8440
rect 34808 7954 34836 11834
rect 35084 11694 35112 12106
rect 35072 11688 35124 11694
rect 35072 11630 35124 11636
rect 34980 11348 35032 11354
rect 34980 11290 35032 11296
rect 34992 8906 35020 11290
rect 35084 10810 35112 11630
rect 35072 10804 35124 10810
rect 35072 10746 35124 10752
rect 35268 10690 35296 12260
rect 35360 11898 35388 12406
rect 35348 11892 35400 11898
rect 35348 11834 35400 11840
rect 35348 10736 35400 10742
rect 35268 10684 35348 10690
rect 35268 10678 35400 10684
rect 35268 10662 35388 10678
rect 35164 10532 35216 10538
rect 35164 10474 35216 10480
rect 35176 10266 35204 10474
rect 35164 10260 35216 10266
rect 35164 10202 35216 10208
rect 35268 10130 35296 10662
rect 35348 10464 35400 10470
rect 35348 10406 35400 10412
rect 35360 10266 35388 10406
rect 35348 10260 35400 10266
rect 35348 10202 35400 10208
rect 35256 10124 35308 10130
rect 35256 10066 35308 10072
rect 35268 9450 35296 10066
rect 35256 9444 35308 9450
rect 35256 9386 35308 9392
rect 34980 8900 35032 8906
rect 34980 8842 35032 8848
rect 34888 8832 34940 8838
rect 34888 8774 34940 8780
rect 35256 8832 35308 8838
rect 35256 8774 35308 8780
rect 34900 8566 34928 8774
rect 34888 8560 34940 8566
rect 34888 8502 34940 8508
rect 35268 8022 35296 8774
rect 35256 8016 35308 8022
rect 35256 7958 35308 7964
rect 34796 7948 34848 7954
rect 34796 7890 34848 7896
rect 34336 7404 34388 7410
rect 34336 7346 34388 7352
rect 33784 6860 33836 6866
rect 33784 6802 33836 6808
rect 32950 6012 33258 6021
rect 32950 6010 32956 6012
rect 33012 6010 33036 6012
rect 33092 6010 33116 6012
rect 33172 6010 33196 6012
rect 33252 6010 33258 6012
rect 33012 5958 33014 6010
rect 33194 5958 33196 6010
rect 32950 5956 32956 5958
rect 33012 5956 33036 5958
rect 33092 5956 33116 5958
rect 33172 5956 33196 5958
rect 33252 5956 33258 5958
rect 32950 5947 33258 5956
rect 32772 5704 32824 5710
rect 32772 5646 32824 5652
rect 31484 5296 31536 5302
rect 31484 5238 31536 5244
rect 32784 4554 32812 5646
rect 32950 4924 33258 4933
rect 32950 4922 32956 4924
rect 33012 4922 33036 4924
rect 33092 4922 33116 4924
rect 33172 4922 33196 4924
rect 33252 4922 33258 4924
rect 33012 4870 33014 4922
rect 33194 4870 33196 4922
rect 32950 4868 32956 4870
rect 33012 4868 33036 4870
rect 33092 4868 33116 4870
rect 33172 4868 33196 4870
rect 33252 4868 33258 4870
rect 32950 4859 33258 4868
rect 32772 4548 32824 4554
rect 32772 4490 32824 4496
rect 32864 4480 32916 4486
rect 32864 4422 32916 4428
rect 29644 2984 29696 2990
rect 29644 2926 29696 2932
rect 30656 2984 30708 2990
rect 30656 2926 30708 2932
rect 27896 2848 27948 2854
rect 27816 2808 27896 2836
rect 27896 2790 27948 2796
rect 32876 2650 32904 4422
rect 34428 4004 34480 4010
rect 34428 3946 34480 3952
rect 32950 3836 33258 3845
rect 32950 3834 32956 3836
rect 33012 3834 33036 3836
rect 33092 3834 33116 3836
rect 33172 3834 33196 3836
rect 33252 3834 33258 3836
rect 33012 3782 33014 3834
rect 33194 3782 33196 3834
rect 32950 3780 32956 3782
rect 33012 3780 33036 3782
rect 33092 3780 33116 3782
rect 33172 3780 33196 3782
rect 33252 3780 33258 3782
rect 32950 3771 33258 3780
rect 32950 2748 33258 2757
rect 32950 2746 32956 2748
rect 33012 2746 33036 2748
rect 33092 2746 33116 2748
rect 33172 2746 33196 2748
rect 33252 2746 33258 2748
rect 33012 2694 33014 2746
rect 33194 2694 33196 2746
rect 32950 2692 32956 2694
rect 33012 2692 33036 2694
rect 33092 2692 33116 2694
rect 33172 2692 33196 2694
rect 33252 2692 33258 2694
rect 32950 2683 33258 2692
rect 34440 2650 34468 3946
rect 35452 3398 35480 16118
rect 35544 12986 35572 17632
rect 35624 17264 35676 17270
rect 35624 17206 35676 17212
rect 35532 12980 35584 12986
rect 35532 12922 35584 12928
rect 35636 12782 35664 17206
rect 35728 16658 35756 17682
rect 35716 16652 35768 16658
rect 35716 16594 35768 16600
rect 35714 16008 35770 16017
rect 35714 15943 35770 15952
rect 35728 14521 35756 15943
rect 35820 15314 35848 19654
rect 35898 19544 35954 19553
rect 35898 19479 35900 19488
rect 35952 19479 35954 19488
rect 35900 19450 35952 19456
rect 35900 19304 35952 19310
rect 35900 19246 35952 19252
rect 35912 19174 35940 19246
rect 35900 19168 35952 19174
rect 35900 19110 35952 19116
rect 36004 18834 36032 22578
rect 36084 22024 36136 22030
rect 36084 21966 36136 21972
rect 36096 19378 36124 21966
rect 36188 21894 36216 24006
rect 36360 23656 36412 23662
rect 36360 23598 36412 23604
rect 36452 23656 36504 23662
rect 36452 23598 36504 23604
rect 36372 21962 36400 23598
rect 36464 22953 36492 23598
rect 36740 23225 36768 26302
rect 37002 26200 37058 27000
rect 37646 26330 37702 27000
rect 38290 26330 38346 27000
rect 38934 26330 38990 27000
rect 39578 26330 39634 27000
rect 40132 26376 40184 26382
rect 37646 26302 37872 26330
rect 37646 26200 37702 26302
rect 37016 23769 37044 26200
rect 37372 24268 37424 24274
rect 37372 24210 37424 24216
rect 37002 23760 37058 23769
rect 37002 23695 37058 23704
rect 37280 23520 37332 23526
rect 37280 23462 37332 23468
rect 37292 23322 37320 23462
rect 37280 23316 37332 23322
rect 37280 23258 37332 23264
rect 36726 23216 36782 23225
rect 36726 23151 36782 23160
rect 37280 23180 37332 23186
rect 37280 23122 37332 23128
rect 36450 22944 36506 22953
rect 36450 22879 36506 22888
rect 37292 22642 37320 23122
rect 36820 22636 36872 22642
rect 36820 22578 36872 22584
rect 37280 22636 37332 22642
rect 37280 22578 37332 22584
rect 36636 22024 36688 22030
rect 36636 21966 36688 21972
rect 36360 21956 36412 21962
rect 36360 21898 36412 21904
rect 36176 21888 36228 21894
rect 36176 21830 36228 21836
rect 36648 21622 36676 21966
rect 36452 21616 36504 21622
rect 36452 21558 36504 21564
rect 36636 21616 36688 21622
rect 36636 21558 36688 21564
rect 36176 21480 36228 21486
rect 36176 21422 36228 21428
rect 36188 20806 36216 21422
rect 36360 21412 36412 21418
rect 36360 21354 36412 21360
rect 36176 20800 36228 20806
rect 36176 20742 36228 20748
rect 36176 19916 36228 19922
rect 36176 19858 36228 19864
rect 36084 19372 36136 19378
rect 36084 19314 36136 19320
rect 36188 19258 36216 19858
rect 36372 19378 36400 21354
rect 36268 19372 36320 19378
rect 36268 19314 36320 19320
rect 36360 19372 36412 19378
rect 36360 19314 36412 19320
rect 36096 19230 36216 19258
rect 35992 18828 36044 18834
rect 35992 18770 36044 18776
rect 35992 18284 36044 18290
rect 35992 18226 36044 18232
rect 35898 18048 35954 18057
rect 35898 17983 35954 17992
rect 35912 17542 35940 17983
rect 35900 17536 35952 17542
rect 35900 17478 35952 17484
rect 35912 16590 35940 17478
rect 35900 16584 35952 16590
rect 35900 16526 35952 16532
rect 35820 15286 35940 15314
rect 35912 15026 35940 15286
rect 35900 15020 35952 15026
rect 35900 14962 35952 14968
rect 35714 14512 35770 14521
rect 35714 14447 35770 14456
rect 36004 13530 36032 18226
rect 36096 17202 36124 19230
rect 36176 19168 36228 19174
rect 36176 19110 36228 19116
rect 36188 18426 36216 19110
rect 36176 18420 36228 18426
rect 36176 18362 36228 18368
rect 36188 17746 36216 18362
rect 36280 18086 36308 19314
rect 36360 19236 36412 19242
rect 36360 19178 36412 19184
rect 36268 18080 36320 18086
rect 36268 18022 36320 18028
rect 36176 17740 36228 17746
rect 36176 17682 36228 17688
rect 36176 17536 36228 17542
rect 36176 17478 36228 17484
rect 36084 17196 36136 17202
rect 36084 17138 36136 17144
rect 36084 15360 36136 15366
rect 36084 15302 36136 15308
rect 35992 13524 36044 13530
rect 35992 13466 36044 13472
rect 35992 13184 36044 13190
rect 35992 13126 36044 13132
rect 35808 12980 35860 12986
rect 35808 12922 35860 12928
rect 35820 12889 35848 12922
rect 35806 12880 35862 12889
rect 35806 12815 35862 12824
rect 35624 12776 35676 12782
rect 35624 12718 35676 12724
rect 35806 12744 35862 12753
rect 35806 12679 35862 12688
rect 35820 12306 35848 12679
rect 35808 12300 35860 12306
rect 35808 12242 35860 12248
rect 35716 11212 35768 11218
rect 35716 11154 35768 11160
rect 35728 10810 35756 11154
rect 35716 10804 35768 10810
rect 35716 10746 35768 10752
rect 35532 10668 35584 10674
rect 35532 10610 35584 10616
rect 35716 10668 35768 10674
rect 35716 10610 35768 10616
rect 35544 9654 35572 10610
rect 35532 9648 35584 9654
rect 35584 9608 35664 9636
rect 35532 9590 35584 9596
rect 35532 9376 35584 9382
rect 35532 9318 35584 9324
rect 35544 9042 35572 9318
rect 35532 9036 35584 9042
rect 35532 8978 35584 8984
rect 35636 8634 35664 9608
rect 35728 9110 35756 10610
rect 35900 10600 35952 10606
rect 35900 10542 35952 10548
rect 35808 9920 35860 9926
rect 35808 9862 35860 9868
rect 35820 9722 35848 9862
rect 35808 9716 35860 9722
rect 35808 9658 35860 9664
rect 35806 9616 35862 9625
rect 35806 9551 35862 9560
rect 35716 9104 35768 9110
rect 35716 9046 35768 9052
rect 35820 8906 35848 9551
rect 35912 9178 35940 10542
rect 35900 9172 35952 9178
rect 35900 9114 35952 9120
rect 35808 8900 35860 8906
rect 35808 8842 35860 8848
rect 35624 8628 35676 8634
rect 35624 8570 35676 8576
rect 35808 5840 35860 5846
rect 35808 5782 35860 5788
rect 35820 4826 35848 5782
rect 35808 4820 35860 4826
rect 35808 4762 35860 4768
rect 35440 3392 35492 3398
rect 35440 3334 35492 3340
rect 36004 2774 36032 13126
rect 36096 12986 36124 15302
rect 36188 15026 36216 17478
rect 36268 17196 36320 17202
rect 36268 17138 36320 17144
rect 36280 16726 36308 17138
rect 36268 16720 36320 16726
rect 36268 16662 36320 16668
rect 36372 16522 36400 19178
rect 36464 17270 36492 21558
rect 36728 21548 36780 21554
rect 36728 21490 36780 21496
rect 36636 21480 36688 21486
rect 36636 21422 36688 21428
rect 36648 20806 36676 21422
rect 36636 20800 36688 20806
rect 36636 20742 36688 20748
rect 36648 20641 36676 20742
rect 36634 20632 36690 20641
rect 36634 20567 36690 20576
rect 36636 20392 36688 20398
rect 36636 20334 36688 20340
rect 36542 19544 36598 19553
rect 36542 19479 36598 19488
rect 36556 19446 36584 19479
rect 36544 19440 36596 19446
rect 36544 19382 36596 19388
rect 36648 18154 36676 20334
rect 36636 18148 36688 18154
rect 36636 18090 36688 18096
rect 36544 17740 36596 17746
rect 36544 17682 36596 17688
rect 36452 17264 36504 17270
rect 36452 17206 36504 17212
rect 36556 17134 36584 17682
rect 36740 17626 36768 21490
rect 36832 18952 36860 22578
rect 37188 22228 37240 22234
rect 37188 22170 37240 22176
rect 37200 22001 37228 22170
rect 37292 22098 37320 22578
rect 37280 22092 37332 22098
rect 37280 22034 37332 22040
rect 37186 21992 37242 22001
rect 37186 21927 37242 21936
rect 37280 21956 37332 21962
rect 37280 21898 37332 21904
rect 37292 21350 37320 21898
rect 37280 21344 37332 21350
rect 37280 21286 37332 21292
rect 37292 21010 37320 21286
rect 37004 21004 37056 21010
rect 37004 20946 37056 20952
rect 37280 21004 37332 21010
rect 37280 20946 37332 20952
rect 36910 19272 36966 19281
rect 36910 19207 36912 19216
rect 36964 19207 36966 19216
rect 36912 19178 36964 19184
rect 36912 18964 36964 18970
rect 36832 18924 36912 18952
rect 36912 18906 36964 18912
rect 37016 18766 37044 20946
rect 37094 20768 37150 20777
rect 37094 20703 37150 20712
rect 37108 19990 37136 20703
rect 37384 20534 37412 24210
rect 37740 24132 37792 24138
rect 37740 24074 37792 24080
rect 37648 24064 37700 24070
rect 37646 24032 37648 24041
rect 37700 24032 37702 24041
rect 37646 23967 37702 23976
rect 37556 23792 37608 23798
rect 37556 23734 37608 23740
rect 37464 23724 37516 23730
rect 37464 23666 37516 23672
rect 37476 22506 37504 23666
rect 37568 23322 37596 23734
rect 37660 23594 37688 23967
rect 37752 23798 37780 24074
rect 37740 23792 37792 23798
rect 37740 23734 37792 23740
rect 37648 23588 37700 23594
rect 37648 23530 37700 23536
rect 37556 23316 37608 23322
rect 37556 23258 37608 23264
rect 37464 22500 37516 22506
rect 37464 22442 37516 22448
rect 37568 22234 37596 23258
rect 37844 23168 37872 26302
rect 38290 26302 38608 26330
rect 38290 26200 38346 26302
rect 37924 24812 37976 24818
rect 37924 24754 37976 24760
rect 37936 24274 37964 24754
rect 37924 24268 37976 24274
rect 37924 24210 37976 24216
rect 38292 24268 38344 24274
rect 38292 24210 38344 24216
rect 37950 23964 38258 23973
rect 37950 23962 37956 23964
rect 38012 23962 38036 23964
rect 38092 23962 38116 23964
rect 38172 23962 38196 23964
rect 38252 23962 38258 23964
rect 38012 23910 38014 23962
rect 38194 23910 38196 23962
rect 37950 23908 37956 23910
rect 38012 23908 38036 23910
rect 38092 23908 38116 23910
rect 38172 23908 38196 23910
rect 38252 23908 38258 23910
rect 37950 23899 38258 23908
rect 37660 23140 37872 23168
rect 37660 22420 37688 23140
rect 37832 23044 37884 23050
rect 37832 22986 37884 22992
rect 37844 22710 37872 22986
rect 37950 22876 38258 22885
rect 37950 22874 37956 22876
rect 38012 22874 38036 22876
rect 38092 22874 38116 22876
rect 38172 22874 38196 22876
rect 38252 22874 38258 22876
rect 38012 22822 38014 22874
rect 38194 22822 38196 22874
rect 37950 22820 37956 22822
rect 38012 22820 38036 22822
rect 38092 22820 38116 22822
rect 38172 22820 38196 22822
rect 38252 22820 38258 22822
rect 37950 22811 38258 22820
rect 37832 22704 37884 22710
rect 37832 22646 37884 22652
rect 37844 22574 37872 22646
rect 37740 22568 37792 22574
rect 37738 22536 37740 22545
rect 37832 22568 37884 22574
rect 37792 22536 37794 22545
rect 37832 22510 37884 22516
rect 37738 22471 37794 22480
rect 37740 22432 37792 22438
rect 37660 22392 37740 22420
rect 37740 22374 37792 22380
rect 37556 22228 37608 22234
rect 37556 22170 37608 22176
rect 38304 22098 38332 24210
rect 38474 23896 38530 23905
rect 38474 23831 38530 23840
rect 38384 23792 38436 23798
rect 38384 23734 38436 23740
rect 38396 23526 38424 23734
rect 38488 23594 38516 23831
rect 38476 23588 38528 23594
rect 38476 23530 38528 23536
rect 38384 23520 38436 23526
rect 38384 23462 38436 23468
rect 38580 22778 38608 26302
rect 38934 26302 39252 26330
rect 38934 26200 38990 26302
rect 38660 24744 38712 24750
rect 38660 24686 38712 24692
rect 38672 23526 38700 24686
rect 39120 24336 39172 24342
rect 39120 24278 39172 24284
rect 38936 24200 38988 24206
rect 38936 24142 38988 24148
rect 38660 23520 38712 23526
rect 38660 23462 38712 23468
rect 38842 23488 38898 23497
rect 38842 23423 38898 23432
rect 38856 23186 38884 23423
rect 38844 23180 38896 23186
rect 38844 23122 38896 23128
rect 38844 22976 38896 22982
rect 38844 22918 38896 22924
rect 38568 22772 38620 22778
rect 38568 22714 38620 22720
rect 38856 22166 38884 22918
rect 38844 22160 38896 22166
rect 38844 22102 38896 22108
rect 37648 22092 37700 22098
rect 38292 22092 38344 22098
rect 37700 22052 37780 22080
rect 37648 22034 37700 22040
rect 37752 21486 37780 22052
rect 38292 22034 38344 22040
rect 37950 21788 38258 21797
rect 37950 21786 37956 21788
rect 38012 21786 38036 21788
rect 38092 21786 38116 21788
rect 38172 21786 38196 21788
rect 38252 21786 38258 21788
rect 38012 21734 38014 21786
rect 38194 21734 38196 21786
rect 37950 21732 37956 21734
rect 38012 21732 38036 21734
rect 38092 21732 38116 21734
rect 38172 21732 38196 21734
rect 38252 21732 38258 21734
rect 37950 21723 38258 21732
rect 38304 21486 38332 22034
rect 38844 21956 38896 21962
rect 38844 21898 38896 21904
rect 38568 21888 38620 21894
rect 38568 21830 38620 21836
rect 38384 21616 38436 21622
rect 38384 21558 38436 21564
rect 38396 21486 38424 21558
rect 37740 21480 37792 21486
rect 37740 21422 37792 21428
rect 38292 21480 38344 21486
rect 38292 21422 38344 21428
rect 38384 21480 38436 21486
rect 38384 21422 38436 21428
rect 37464 21412 37516 21418
rect 37464 21354 37516 21360
rect 37372 20528 37424 20534
rect 37372 20470 37424 20476
rect 37188 20460 37240 20466
rect 37188 20402 37240 20408
rect 37096 19984 37148 19990
rect 37096 19926 37148 19932
rect 37004 18760 37056 18766
rect 37004 18702 37056 18708
rect 36740 17598 36952 17626
rect 36820 17536 36872 17542
rect 36820 17478 36872 17484
rect 36544 17128 36596 17134
rect 36544 17070 36596 17076
rect 36636 17128 36688 17134
rect 36636 17070 36688 17076
rect 36726 17096 36782 17105
rect 36544 16992 36596 16998
rect 36544 16934 36596 16940
rect 36360 16516 36412 16522
rect 36360 16458 36412 16464
rect 36452 16516 36504 16522
rect 36452 16458 36504 16464
rect 36372 15570 36400 16458
rect 36464 16114 36492 16458
rect 36556 16454 36584 16934
rect 36544 16448 36596 16454
rect 36544 16390 36596 16396
rect 36452 16108 36504 16114
rect 36452 16050 36504 16056
rect 36360 15564 36412 15570
rect 36360 15506 36412 15512
rect 36464 15434 36492 16050
rect 36452 15428 36504 15434
rect 36452 15370 36504 15376
rect 36464 15026 36492 15370
rect 36556 15366 36584 16390
rect 36544 15360 36596 15366
rect 36544 15302 36596 15308
rect 36176 15020 36228 15026
rect 36176 14962 36228 14968
rect 36452 15020 36504 15026
rect 36452 14962 36504 14968
rect 36464 14346 36492 14962
rect 36544 14952 36596 14958
rect 36544 14894 36596 14900
rect 36452 14340 36504 14346
rect 36452 14282 36504 14288
rect 36464 14074 36492 14282
rect 36452 14068 36504 14074
rect 36452 14010 36504 14016
rect 36176 13864 36228 13870
rect 36176 13806 36228 13812
rect 36084 12980 36136 12986
rect 36084 12922 36136 12928
rect 36082 12880 36138 12889
rect 36082 12815 36138 12824
rect 36096 12646 36124 12815
rect 36084 12640 36136 12646
rect 36084 12582 36136 12588
rect 36084 11892 36136 11898
rect 36084 11834 36136 11840
rect 36096 11082 36124 11834
rect 36188 11354 36216 13806
rect 36360 13252 36412 13258
rect 36360 13194 36412 13200
rect 36372 12434 36400 13194
rect 36452 13184 36504 13190
rect 36452 13126 36504 13132
rect 36464 12918 36492 13126
rect 36452 12912 36504 12918
rect 36452 12854 36504 12860
rect 36280 12406 36400 12434
rect 36176 11348 36228 11354
rect 36176 11290 36228 11296
rect 36084 11076 36136 11082
rect 36084 11018 36136 11024
rect 36280 8362 36308 12406
rect 36556 12102 36584 14894
rect 36648 14618 36676 17070
rect 36726 17031 36782 17040
rect 36740 16658 36768 17031
rect 36728 16652 36780 16658
rect 36728 16594 36780 16600
rect 36728 16448 36780 16454
rect 36728 16390 36780 16396
rect 36740 14822 36768 16390
rect 36832 16046 36860 17478
rect 36924 16590 36952 17598
rect 37200 17066 37228 20402
rect 37280 20052 37332 20058
rect 37280 19994 37332 20000
rect 37292 18086 37320 19994
rect 37372 19916 37424 19922
rect 37372 19858 37424 19864
rect 37384 19242 37412 19858
rect 37372 19236 37424 19242
rect 37372 19178 37424 19184
rect 37476 19174 37504 21354
rect 37648 20936 37700 20942
rect 37752 20890 37780 21422
rect 38304 21010 38332 21422
rect 38292 21004 38344 21010
rect 38292 20946 38344 20952
rect 37700 20884 37780 20890
rect 37648 20878 37780 20884
rect 37660 20862 37780 20878
rect 37752 20398 37780 20862
rect 38292 20800 38344 20806
rect 38292 20742 38344 20748
rect 37950 20700 38258 20709
rect 37950 20698 37956 20700
rect 38012 20698 38036 20700
rect 38092 20698 38116 20700
rect 38172 20698 38196 20700
rect 38252 20698 38258 20700
rect 38012 20646 38014 20698
rect 38194 20646 38196 20698
rect 37950 20644 37956 20646
rect 38012 20644 38036 20646
rect 38092 20644 38116 20646
rect 38172 20644 38196 20646
rect 38252 20644 38258 20646
rect 37950 20635 38258 20644
rect 38304 20534 38332 20742
rect 38292 20528 38344 20534
rect 38292 20470 38344 20476
rect 38580 20398 38608 21830
rect 38856 21622 38884 21898
rect 38844 21616 38896 21622
rect 38844 21558 38896 21564
rect 38856 21026 38884 21558
rect 38672 20998 38884 21026
rect 38672 20874 38700 20998
rect 38660 20868 38712 20874
rect 38660 20810 38712 20816
rect 38672 20534 38700 20810
rect 38660 20528 38712 20534
rect 38712 20488 38792 20516
rect 38660 20470 38712 20476
rect 37556 20392 37608 20398
rect 37556 20334 37608 20340
rect 37740 20392 37792 20398
rect 37740 20334 37792 20340
rect 38568 20392 38620 20398
rect 38568 20334 38620 20340
rect 37464 19168 37516 19174
rect 37464 19110 37516 19116
rect 37464 18896 37516 18902
rect 37464 18838 37516 18844
rect 37476 18290 37504 18838
rect 37568 18834 37596 20334
rect 37648 19916 37700 19922
rect 37648 19858 37700 19864
rect 37556 18828 37608 18834
rect 37556 18770 37608 18776
rect 37372 18284 37424 18290
rect 37372 18226 37424 18232
rect 37464 18284 37516 18290
rect 37464 18226 37516 18232
rect 37280 18080 37332 18086
rect 37280 18022 37332 18028
rect 37188 17060 37240 17066
rect 37188 17002 37240 17008
rect 37004 16720 37056 16726
rect 37004 16662 37056 16668
rect 36912 16584 36964 16590
rect 36912 16526 36964 16532
rect 36924 16250 36952 16526
rect 37016 16522 37044 16662
rect 37004 16516 37056 16522
rect 37004 16458 37056 16464
rect 36912 16244 36964 16250
rect 36912 16186 36964 16192
rect 36820 16040 36872 16046
rect 36820 15982 36872 15988
rect 37280 16040 37332 16046
rect 37280 15982 37332 15988
rect 36832 15706 36860 15982
rect 36820 15700 36872 15706
rect 36820 15642 36872 15648
rect 37004 15700 37056 15706
rect 37004 15642 37056 15648
rect 37016 14958 37044 15642
rect 37096 15360 37148 15366
rect 37096 15302 37148 15308
rect 37004 14952 37056 14958
rect 37004 14894 37056 14900
rect 36728 14816 36780 14822
rect 36728 14758 36780 14764
rect 36636 14612 36688 14618
rect 36636 14554 36688 14560
rect 36648 13870 36676 14554
rect 36636 13864 36688 13870
rect 36636 13806 36688 13812
rect 36648 13258 36676 13806
rect 37108 13394 37136 15302
rect 37292 15162 37320 15982
rect 37384 15910 37412 18226
rect 37476 17678 37504 18226
rect 37464 17672 37516 17678
rect 37464 17614 37516 17620
rect 37476 16726 37504 17614
rect 37660 17082 37688 19858
rect 37752 19378 37780 20334
rect 38660 20256 38712 20262
rect 38660 20198 38712 20204
rect 38200 19984 38252 19990
rect 38200 19926 38252 19932
rect 38212 19718 38240 19926
rect 38672 19718 38700 20198
rect 38764 19922 38792 20488
rect 38752 19916 38804 19922
rect 38752 19858 38804 19864
rect 37832 19712 37884 19718
rect 37832 19654 37884 19660
rect 38200 19712 38252 19718
rect 38200 19654 38252 19660
rect 38660 19712 38712 19718
rect 38660 19654 38712 19660
rect 37740 19372 37792 19378
rect 37740 19314 37792 19320
rect 37844 18306 37872 19654
rect 37950 19612 38258 19621
rect 37950 19610 37956 19612
rect 38012 19610 38036 19612
rect 38092 19610 38116 19612
rect 38172 19610 38196 19612
rect 38252 19610 38258 19612
rect 38012 19558 38014 19610
rect 38194 19558 38196 19610
rect 37950 19556 37956 19558
rect 38012 19556 38036 19558
rect 38092 19556 38116 19558
rect 38172 19556 38196 19558
rect 38252 19556 38258 19558
rect 37950 19547 38258 19556
rect 38382 19544 38438 19553
rect 37924 19508 37976 19514
rect 38382 19479 38384 19488
rect 37924 19450 37976 19456
rect 38436 19479 38438 19488
rect 38384 19450 38436 19456
rect 37936 19242 37964 19450
rect 38476 19440 38528 19446
rect 38476 19382 38528 19388
rect 38200 19304 38252 19310
rect 38198 19272 38200 19281
rect 38252 19272 38254 19281
rect 37924 19236 37976 19242
rect 38198 19207 38254 19216
rect 37924 19178 37976 19184
rect 38212 18970 38240 19207
rect 38292 19168 38344 19174
rect 38292 19110 38344 19116
rect 38200 18964 38252 18970
rect 38200 18906 38252 18912
rect 38014 18728 38070 18737
rect 38014 18663 38070 18672
rect 38028 18630 38056 18663
rect 38016 18624 38068 18630
rect 38016 18566 38068 18572
rect 37950 18524 38258 18533
rect 37950 18522 37956 18524
rect 38012 18522 38036 18524
rect 38092 18522 38116 18524
rect 38172 18522 38196 18524
rect 38252 18522 38258 18524
rect 38012 18470 38014 18522
rect 38194 18470 38196 18522
rect 37950 18468 37956 18470
rect 38012 18468 38036 18470
rect 38092 18468 38116 18470
rect 38172 18468 38196 18470
rect 38252 18468 38258 18470
rect 37950 18459 38258 18468
rect 37752 18278 37872 18306
rect 37752 17270 37780 18278
rect 38304 18222 38332 19110
rect 38384 18760 38436 18766
rect 38384 18702 38436 18708
rect 38396 18358 38424 18702
rect 38384 18352 38436 18358
rect 38384 18294 38436 18300
rect 37832 18216 37884 18222
rect 37832 18158 37884 18164
rect 38292 18216 38344 18222
rect 38292 18158 38344 18164
rect 37740 17264 37792 17270
rect 37740 17206 37792 17212
rect 37568 17054 37688 17082
rect 37740 17060 37792 17066
rect 37464 16720 37516 16726
rect 37464 16662 37516 16668
rect 37464 16584 37516 16590
rect 37464 16526 37516 16532
rect 37476 16182 37504 16526
rect 37464 16176 37516 16182
rect 37464 16118 37516 16124
rect 37372 15904 37424 15910
rect 37372 15846 37424 15852
rect 37476 15502 37504 16118
rect 37464 15496 37516 15502
rect 37464 15438 37516 15444
rect 37372 15428 37424 15434
rect 37372 15370 37424 15376
rect 37280 15156 37332 15162
rect 37280 15098 37332 15104
rect 37188 15088 37240 15094
rect 37188 15030 37240 15036
rect 37200 14929 37228 15030
rect 37186 14920 37242 14929
rect 37186 14855 37242 14864
rect 37280 14884 37332 14890
rect 37280 14826 37332 14832
rect 37096 13388 37148 13394
rect 37096 13330 37148 13336
rect 36636 13252 36688 13258
rect 36636 13194 36688 13200
rect 36820 12980 36872 12986
rect 36820 12922 36872 12928
rect 36728 12912 36780 12918
rect 36728 12854 36780 12860
rect 36740 12170 36768 12854
rect 36832 12186 36860 12922
rect 37292 12238 37320 14826
rect 37384 13530 37412 15370
rect 37476 15026 37504 15438
rect 37464 15020 37516 15026
rect 37464 14962 37516 14968
rect 37476 14482 37504 14962
rect 37568 14822 37596 17054
rect 37740 17002 37792 17008
rect 37648 16992 37700 16998
rect 37648 16934 37700 16940
rect 37556 14816 37608 14822
rect 37556 14758 37608 14764
rect 37464 14476 37516 14482
rect 37464 14418 37516 14424
rect 37568 14362 37596 14758
rect 37476 14346 37596 14362
rect 37464 14340 37596 14346
rect 37516 14334 37596 14340
rect 37464 14282 37516 14288
rect 37556 14272 37608 14278
rect 37556 14214 37608 14220
rect 37568 14090 37596 14214
rect 37476 14062 37596 14090
rect 37372 13524 37424 13530
rect 37372 13466 37424 13472
rect 37372 13184 37424 13190
rect 37372 13126 37424 13132
rect 37384 12850 37412 13126
rect 37372 12844 37424 12850
rect 37372 12786 37424 12792
rect 37372 12708 37424 12714
rect 37372 12650 37424 12656
rect 37280 12232 37332 12238
rect 36728 12164 36780 12170
rect 36832 12158 37044 12186
rect 37280 12174 37332 12180
rect 36728 12106 36780 12112
rect 36544 12096 36596 12102
rect 36544 12038 36596 12044
rect 36740 11830 36768 12106
rect 36820 12096 36872 12102
rect 36820 12038 36872 12044
rect 36728 11824 36780 11830
rect 36728 11766 36780 11772
rect 36636 11688 36688 11694
rect 36636 11630 36688 11636
rect 36648 10470 36676 11630
rect 36740 11082 36768 11766
rect 36832 11626 36860 12038
rect 36912 11756 36964 11762
rect 36912 11698 36964 11704
rect 36820 11620 36872 11626
rect 36820 11562 36872 11568
rect 36728 11076 36780 11082
rect 36728 11018 36780 11024
rect 36740 10742 36768 11018
rect 36924 10810 36952 11698
rect 36912 10804 36964 10810
rect 36912 10746 36964 10752
rect 36728 10736 36780 10742
rect 36728 10678 36780 10684
rect 36636 10464 36688 10470
rect 36636 10406 36688 10412
rect 36648 10266 36676 10406
rect 36740 10266 36768 10678
rect 36636 10260 36688 10266
rect 36636 10202 36688 10208
rect 36728 10260 36780 10266
rect 36728 10202 36780 10208
rect 36740 9994 36768 10202
rect 36728 9988 36780 9994
rect 36728 9930 36780 9936
rect 36268 8356 36320 8362
rect 36268 8298 36320 8304
rect 36452 6248 36504 6254
rect 36452 6190 36504 6196
rect 36464 3534 36492 6190
rect 37016 4690 37044 12158
rect 37384 11830 37412 12650
rect 37476 12306 37504 14062
rect 37660 14006 37688 16934
rect 37752 16590 37780 17002
rect 37740 16584 37792 16590
rect 37740 16526 37792 16532
rect 37740 15972 37792 15978
rect 37740 15914 37792 15920
rect 37752 14482 37780 15914
rect 37844 15706 37872 18158
rect 37950 17436 38258 17445
rect 37950 17434 37956 17436
rect 38012 17434 38036 17436
rect 38092 17434 38116 17436
rect 38172 17434 38196 17436
rect 38252 17434 38258 17436
rect 38012 17382 38014 17434
rect 38194 17382 38196 17434
rect 37950 17380 37956 17382
rect 38012 17380 38036 17382
rect 38092 17380 38116 17382
rect 38172 17380 38196 17382
rect 38252 17380 38258 17382
rect 37950 17371 38258 17380
rect 38304 17134 38332 18158
rect 38488 17746 38516 19382
rect 38764 18902 38792 19858
rect 38948 19417 38976 24142
rect 39132 21078 39160 24278
rect 39224 23254 39252 26302
rect 39578 26302 39896 26330
rect 40132 26318 40184 26324
rect 39578 26200 39634 26302
rect 39672 24608 39724 24614
rect 39672 24550 39724 24556
rect 39304 23656 39356 23662
rect 39304 23598 39356 23604
rect 39396 23656 39448 23662
rect 39396 23598 39448 23604
rect 39212 23248 39264 23254
rect 39212 23190 39264 23196
rect 39316 22094 39344 23598
rect 39408 23089 39436 23598
rect 39394 23080 39450 23089
rect 39394 23015 39450 23024
rect 39408 22137 39436 23015
rect 39580 22976 39632 22982
rect 39580 22918 39632 22924
rect 39592 22710 39620 22918
rect 39580 22704 39632 22710
rect 39580 22646 39632 22652
rect 39488 22636 39540 22642
rect 39488 22578 39540 22584
rect 39500 22438 39528 22578
rect 39488 22432 39540 22438
rect 39488 22374 39540 22380
rect 39224 22066 39344 22094
rect 39394 22128 39450 22137
rect 39120 21072 39172 21078
rect 39120 21014 39172 21020
rect 39224 20505 39252 22066
rect 39394 22063 39450 22072
rect 39592 21962 39620 22646
rect 39684 22438 39712 24550
rect 39868 22438 39896 26302
rect 40040 24676 40092 24682
rect 40040 24618 40092 24624
rect 40052 24018 40080 24618
rect 40144 24206 40172 26318
rect 40222 26200 40278 27000
rect 42154 26200 42210 27000
rect 42798 26200 42854 27000
rect 43442 26200 43498 27000
rect 44086 26200 44142 27000
rect 44730 26200 44786 27000
rect 45374 26200 45430 27000
rect 46018 26200 46074 27000
rect 46662 26330 46718 27000
rect 46662 26302 46888 26330
rect 46662 26200 46718 26302
rect 40132 24200 40184 24206
rect 40132 24142 40184 24148
rect 40052 23990 40172 24018
rect 40144 23730 40172 23990
rect 40040 23724 40092 23730
rect 40040 23666 40092 23672
rect 40132 23724 40184 23730
rect 40132 23666 40184 23672
rect 40052 23322 40080 23666
rect 40236 23322 40264 26200
rect 40408 25084 40460 25090
rect 40408 25026 40460 25032
rect 40316 24404 40368 24410
rect 40316 24346 40368 24352
rect 40040 23316 40092 23322
rect 40040 23258 40092 23264
rect 40224 23316 40276 23322
rect 40224 23258 40276 23264
rect 40040 22636 40092 22642
rect 40040 22578 40092 22584
rect 39672 22432 39724 22438
rect 39672 22374 39724 22380
rect 39856 22432 39908 22438
rect 39856 22374 39908 22380
rect 40052 22234 40080 22578
rect 40132 22568 40184 22574
rect 40132 22510 40184 22516
rect 40040 22228 40092 22234
rect 40040 22170 40092 22176
rect 39580 21956 39632 21962
rect 39580 21898 39632 21904
rect 40040 21888 40092 21894
rect 40040 21830 40092 21836
rect 40052 21690 40080 21830
rect 40144 21690 40172 22510
rect 40328 22094 40356 24346
rect 40420 23662 40448 25026
rect 40500 24812 40552 24818
rect 40500 24754 40552 24760
rect 40512 24410 40540 24754
rect 40682 24440 40738 24449
rect 40500 24404 40552 24410
rect 40682 24375 40738 24384
rect 40868 24404 40920 24410
rect 40500 24346 40552 24352
rect 40696 24274 40724 24375
rect 40868 24346 40920 24352
rect 40684 24268 40736 24274
rect 40684 24210 40736 24216
rect 40500 24064 40552 24070
rect 40500 24006 40552 24012
rect 40408 23656 40460 23662
rect 40408 23598 40460 23604
rect 40408 22976 40460 22982
rect 40408 22918 40460 22924
rect 40236 22066 40356 22094
rect 40040 21684 40092 21690
rect 40040 21626 40092 21632
rect 40132 21684 40184 21690
rect 40132 21626 40184 21632
rect 39856 21616 39908 21622
rect 39856 21558 39908 21564
rect 39868 21350 39896 21558
rect 40040 21412 40092 21418
rect 40040 21354 40092 21360
rect 39764 21344 39816 21350
rect 39764 21286 39816 21292
rect 39856 21344 39908 21350
rect 39856 21286 39908 21292
rect 39776 21078 39804 21286
rect 39764 21072 39816 21078
rect 39764 21014 39816 21020
rect 39210 20496 39266 20505
rect 39210 20431 39266 20440
rect 39028 20324 39080 20330
rect 39028 20266 39080 20272
rect 38934 19408 38990 19417
rect 38934 19343 38990 19352
rect 38752 18896 38804 18902
rect 38752 18838 38804 18844
rect 38568 18828 38620 18834
rect 38568 18770 38620 18776
rect 38476 17740 38528 17746
rect 38476 17682 38528 17688
rect 38384 17536 38436 17542
rect 38384 17478 38436 17484
rect 38292 17128 38344 17134
rect 38292 17070 38344 17076
rect 38292 16992 38344 16998
rect 38292 16934 38344 16940
rect 38304 16522 38332 16934
rect 38292 16516 38344 16522
rect 38292 16458 38344 16464
rect 37950 16348 38258 16357
rect 37950 16346 37956 16348
rect 38012 16346 38036 16348
rect 38092 16346 38116 16348
rect 38172 16346 38196 16348
rect 38252 16346 38258 16348
rect 38012 16294 38014 16346
rect 38194 16294 38196 16346
rect 37950 16292 37956 16294
rect 38012 16292 38036 16294
rect 38092 16292 38116 16294
rect 38172 16292 38196 16294
rect 38252 16292 38258 16294
rect 37950 16283 38258 16292
rect 37832 15700 37884 15706
rect 37832 15642 37884 15648
rect 37950 15260 38258 15269
rect 37950 15258 37956 15260
rect 38012 15258 38036 15260
rect 38092 15258 38116 15260
rect 38172 15258 38196 15260
rect 38252 15258 38258 15260
rect 38012 15206 38014 15258
rect 38194 15206 38196 15258
rect 37950 15204 37956 15206
rect 38012 15204 38036 15206
rect 38092 15204 38116 15206
rect 38172 15204 38196 15206
rect 38252 15204 38258 15206
rect 37950 15195 38258 15204
rect 38304 15144 38332 16458
rect 38396 16454 38424 17478
rect 38476 17128 38528 17134
rect 38474 17096 38476 17105
rect 38528 17096 38530 17105
rect 38474 17031 38530 17040
rect 38474 16552 38530 16561
rect 38474 16487 38530 16496
rect 38384 16448 38436 16454
rect 38384 16390 38436 16396
rect 38120 15116 38332 15144
rect 37832 15088 37884 15094
rect 37832 15030 37884 15036
rect 37740 14476 37792 14482
rect 37740 14418 37792 14424
rect 37844 14346 37872 15030
rect 38120 14618 38148 15116
rect 38488 14958 38516 16487
rect 38580 16436 38608 18770
rect 39040 18193 39068 20266
rect 39212 20256 39264 20262
rect 39212 20198 39264 20204
rect 39224 19310 39252 20198
rect 39764 19984 39816 19990
rect 39764 19926 39816 19932
rect 39488 19916 39540 19922
rect 39488 19858 39540 19864
rect 39500 19446 39528 19858
rect 39488 19440 39540 19446
rect 39488 19382 39540 19388
rect 39212 19304 39264 19310
rect 39212 19246 39264 19252
rect 39224 18426 39252 19246
rect 39500 19242 39528 19382
rect 39488 19236 39540 19242
rect 39488 19178 39540 19184
rect 39776 19174 39804 19926
rect 39868 19718 39896 21286
rect 40052 21162 40080 21354
rect 39960 21146 40080 21162
rect 40236 21146 40264 22066
rect 40420 21690 40448 22918
rect 40408 21684 40460 21690
rect 40408 21626 40460 21632
rect 40512 21418 40540 24006
rect 40776 23792 40828 23798
rect 40604 23740 40776 23746
rect 40604 23734 40828 23740
rect 40604 23730 40816 23734
rect 40592 23724 40816 23730
rect 40644 23718 40816 23724
rect 40592 23666 40644 23672
rect 40880 23610 40908 24346
rect 40958 24304 41014 24313
rect 40958 24239 40960 24248
rect 41012 24239 41014 24248
rect 40960 24210 41012 24216
rect 42168 24206 42196 26200
rect 42800 25016 42852 25022
rect 42800 24958 42852 24964
rect 41328 24200 41380 24206
rect 41328 24142 41380 24148
rect 42156 24200 42208 24206
rect 42156 24142 42208 24148
rect 40604 23582 40908 23610
rect 40500 21412 40552 21418
rect 40500 21354 40552 21360
rect 40314 21176 40370 21185
rect 39948 21140 40080 21146
rect 40000 21134 40080 21140
rect 40224 21140 40276 21146
rect 39948 21082 40000 21088
rect 40314 21111 40316 21120
rect 40224 21082 40276 21088
rect 40368 21111 40370 21120
rect 40316 21082 40368 21088
rect 40604 20602 40632 23582
rect 40868 23316 40920 23322
rect 40868 23258 40920 23264
rect 40880 22574 40908 23258
rect 41236 23044 41288 23050
rect 41236 22986 41288 22992
rect 41248 22778 41276 22986
rect 41236 22772 41288 22778
rect 41236 22714 41288 22720
rect 40868 22568 40920 22574
rect 40774 22536 40830 22545
rect 40868 22510 40920 22516
rect 40774 22471 40830 22480
rect 40788 22166 40816 22471
rect 40960 22432 41012 22438
rect 40960 22374 41012 22380
rect 40776 22160 40828 22166
rect 40776 22102 40828 22108
rect 40684 21888 40736 21894
rect 40684 21830 40736 21836
rect 40592 20596 40644 20602
rect 40592 20538 40644 20544
rect 40500 20392 40552 20398
rect 40500 20334 40552 20340
rect 39948 20256 40000 20262
rect 39948 20198 40000 20204
rect 39856 19712 39908 19718
rect 39856 19654 39908 19660
rect 39764 19168 39816 19174
rect 39764 19110 39816 19116
rect 39764 18692 39816 18698
rect 39764 18634 39816 18640
rect 39776 18426 39804 18634
rect 39212 18420 39264 18426
rect 39212 18362 39264 18368
rect 39764 18420 39816 18426
rect 39764 18362 39816 18368
rect 39026 18184 39082 18193
rect 39026 18119 39082 18128
rect 39856 17808 39908 17814
rect 39578 17776 39634 17785
rect 39856 17750 39908 17756
rect 39578 17711 39634 17720
rect 38660 16448 38712 16454
rect 38580 16408 38660 16436
rect 38580 16182 38608 16408
rect 38660 16390 38712 16396
rect 38568 16176 38620 16182
rect 38568 16118 38620 16124
rect 38568 15156 38620 15162
rect 38568 15098 38620 15104
rect 38476 14952 38528 14958
rect 38580 14929 38608 15098
rect 38936 14952 38988 14958
rect 38476 14894 38528 14900
rect 38566 14920 38622 14929
rect 38936 14894 38988 14900
rect 38566 14855 38622 14864
rect 38948 14618 38976 14894
rect 38108 14612 38160 14618
rect 38108 14554 38160 14560
rect 38384 14612 38436 14618
rect 38384 14554 38436 14560
rect 38936 14612 38988 14618
rect 38936 14554 38988 14560
rect 37832 14340 37884 14346
rect 37832 14282 37884 14288
rect 37556 14000 37608 14006
rect 37556 13942 37608 13948
rect 37648 14000 37700 14006
rect 37648 13942 37700 13948
rect 37568 12730 37596 13942
rect 37740 13796 37792 13802
rect 37740 13738 37792 13744
rect 37752 13190 37780 13738
rect 37844 13530 37872 14282
rect 37950 14172 38258 14181
rect 37950 14170 37956 14172
rect 38012 14170 38036 14172
rect 38092 14170 38116 14172
rect 38172 14170 38196 14172
rect 38252 14170 38258 14172
rect 38012 14118 38014 14170
rect 38194 14118 38196 14170
rect 37950 14116 37956 14118
rect 38012 14116 38036 14118
rect 38092 14116 38116 14118
rect 38172 14116 38196 14118
rect 38252 14116 38258 14118
rect 37950 14107 38258 14116
rect 38396 13734 38424 14554
rect 39592 14414 39620 17711
rect 39764 16516 39816 16522
rect 39764 16458 39816 16464
rect 39776 16182 39804 16458
rect 39764 16176 39816 16182
rect 39764 16118 39816 16124
rect 39776 15434 39804 16118
rect 39764 15428 39816 15434
rect 39764 15370 39816 15376
rect 39776 14618 39804 15370
rect 39868 15026 39896 17750
rect 39960 17746 39988 20198
rect 40406 19952 40462 19961
rect 40406 19887 40462 19896
rect 40132 19780 40184 19786
rect 40132 19722 40184 19728
rect 40040 19712 40092 19718
rect 40040 19654 40092 19660
rect 40052 18426 40080 19654
rect 40144 19514 40172 19722
rect 40420 19514 40448 19887
rect 40132 19508 40184 19514
rect 40132 19450 40184 19456
rect 40408 19508 40460 19514
rect 40408 19450 40460 19456
rect 40132 19372 40184 19378
rect 40132 19314 40184 19320
rect 40144 18873 40172 19314
rect 40224 19236 40276 19242
rect 40224 19178 40276 19184
rect 40130 18864 40186 18873
rect 40130 18799 40186 18808
rect 40040 18420 40092 18426
rect 40040 18362 40092 18368
rect 40236 18358 40264 19178
rect 40406 19136 40462 19145
rect 40406 19071 40462 19080
rect 40224 18352 40276 18358
rect 40224 18294 40276 18300
rect 39948 17740 40000 17746
rect 39948 17682 40000 17688
rect 40132 17332 40184 17338
rect 40132 17274 40184 17280
rect 40224 17332 40276 17338
rect 40224 17274 40276 17280
rect 40040 16448 40092 16454
rect 40040 16390 40092 16396
rect 40052 16250 40080 16390
rect 40040 16244 40092 16250
rect 40040 16186 40092 16192
rect 40144 15162 40172 17274
rect 40236 16658 40264 17274
rect 40420 17066 40448 19071
rect 40512 18952 40540 20334
rect 40592 19916 40644 19922
rect 40592 19858 40644 19864
rect 40604 19281 40632 19858
rect 40590 19272 40646 19281
rect 40590 19207 40646 19216
rect 40512 18924 40632 18952
rect 40604 18630 40632 18924
rect 40500 18624 40552 18630
rect 40500 18566 40552 18572
rect 40592 18624 40644 18630
rect 40592 18566 40644 18572
rect 40512 17814 40540 18566
rect 40500 17808 40552 17814
rect 40500 17750 40552 17756
rect 40604 17134 40632 18566
rect 40696 18329 40724 21830
rect 40788 21486 40816 22102
rect 40868 21548 40920 21554
rect 40868 21490 40920 21496
rect 40776 21480 40828 21486
rect 40776 21422 40828 21428
rect 40880 21049 40908 21490
rect 40866 21040 40922 21049
rect 40866 20975 40922 20984
rect 40972 20913 41000 22374
rect 41340 22137 41368 24142
rect 41788 24132 41840 24138
rect 41788 24074 41840 24080
rect 42248 24132 42300 24138
rect 42248 24074 42300 24080
rect 41800 23662 41828 24074
rect 41972 24064 42024 24070
rect 41972 24006 42024 24012
rect 42156 24064 42208 24070
rect 42156 24006 42208 24012
rect 41788 23656 41840 23662
rect 41788 23598 41840 23604
rect 41604 23520 41656 23526
rect 41604 23462 41656 23468
rect 41420 23180 41472 23186
rect 41420 23122 41472 23128
rect 41432 22710 41460 23122
rect 41420 22704 41472 22710
rect 41420 22646 41472 22652
rect 41326 22128 41382 22137
rect 41326 22063 41382 22072
rect 41432 21962 41460 22646
rect 41512 22432 41564 22438
rect 41512 22374 41564 22380
rect 41420 21956 41472 21962
rect 41420 21898 41472 21904
rect 41236 21616 41288 21622
rect 41236 21558 41288 21564
rect 41052 21140 41104 21146
rect 41052 21082 41104 21088
rect 40958 20904 41014 20913
rect 40958 20839 41014 20848
rect 41064 19922 41092 21082
rect 41248 19990 41276 21558
rect 41418 21448 41474 21457
rect 41418 21383 41420 21392
rect 41472 21383 41474 21392
rect 41420 21354 41472 21360
rect 41524 21321 41552 22374
rect 41616 22098 41644 23462
rect 41984 22778 42012 24006
rect 42168 23730 42196 24006
rect 42260 23905 42288 24074
rect 42246 23896 42302 23905
rect 42246 23831 42302 23840
rect 42156 23724 42208 23730
rect 42156 23666 42208 23672
rect 42260 23526 42288 23831
rect 42432 23792 42484 23798
rect 42432 23734 42484 23740
rect 42444 23594 42472 23734
rect 42812 23730 42840 24958
rect 42950 24508 43258 24517
rect 42950 24506 42956 24508
rect 43012 24506 43036 24508
rect 43092 24506 43116 24508
rect 43172 24506 43196 24508
rect 43252 24506 43258 24508
rect 43012 24454 43014 24506
rect 43194 24454 43196 24506
rect 42950 24452 42956 24454
rect 43012 24452 43036 24454
rect 43092 24452 43116 24454
rect 43172 24452 43196 24454
rect 43252 24452 43258 24454
rect 42950 24443 43258 24452
rect 43996 24064 44048 24070
rect 43996 24006 44048 24012
rect 42800 23724 42852 23730
rect 42800 23666 42852 23672
rect 42616 23656 42668 23662
rect 42616 23598 42668 23604
rect 43904 23656 43956 23662
rect 43904 23598 43956 23604
rect 42432 23588 42484 23594
rect 42432 23530 42484 23536
rect 42248 23520 42300 23526
rect 42248 23462 42300 23468
rect 42064 23044 42116 23050
rect 42064 22986 42116 22992
rect 41972 22772 42024 22778
rect 41972 22714 42024 22720
rect 42076 22710 42104 22986
rect 42156 22976 42208 22982
rect 42156 22918 42208 22924
rect 42168 22817 42196 22918
rect 42154 22808 42210 22817
rect 42154 22743 42210 22752
rect 42248 22772 42300 22778
rect 42064 22704 42116 22710
rect 42064 22646 42116 22652
rect 41696 22636 41748 22642
rect 41696 22578 41748 22584
rect 41708 22234 41736 22578
rect 42168 22438 42196 22743
rect 42248 22714 42300 22720
rect 42260 22642 42288 22714
rect 42248 22636 42300 22642
rect 42248 22578 42300 22584
rect 42156 22432 42208 22438
rect 42156 22374 42208 22380
rect 41696 22228 41748 22234
rect 41696 22170 41748 22176
rect 41604 22092 41656 22098
rect 41604 22034 41656 22040
rect 41708 22001 41736 22170
rect 41878 22128 41934 22137
rect 41934 22072 42012 22094
rect 41878 22066 42012 22072
rect 41878 22063 41934 22066
rect 41984 22030 42012 22066
rect 42064 22092 42116 22098
rect 42064 22034 42116 22040
rect 41972 22024 42024 22030
rect 41694 21992 41750 22001
rect 41972 21966 42024 21972
rect 41694 21927 41750 21936
rect 41788 21956 41840 21962
rect 41788 21898 41840 21904
rect 41800 21842 41828 21898
rect 42076 21842 42104 22034
rect 41800 21814 42104 21842
rect 41788 21616 41840 21622
rect 41788 21558 41840 21564
rect 41800 21486 41828 21558
rect 41788 21480 41840 21486
rect 41788 21422 41840 21428
rect 41510 21312 41566 21321
rect 41510 21247 41566 21256
rect 42168 21078 42196 22374
rect 42260 21690 42288 22578
rect 42444 22166 42472 23530
rect 42628 23361 42656 23598
rect 42950 23420 43258 23429
rect 42950 23418 42956 23420
rect 43012 23418 43036 23420
rect 43092 23418 43116 23420
rect 43172 23418 43196 23420
rect 43252 23418 43258 23420
rect 43012 23366 43014 23418
rect 43194 23366 43196 23418
rect 42950 23364 42956 23366
rect 43012 23364 43036 23366
rect 43092 23364 43116 23366
rect 43172 23364 43196 23366
rect 43252 23364 43258 23366
rect 42614 23352 42670 23361
rect 42950 23355 43258 23364
rect 42614 23287 42670 23296
rect 42800 23316 42852 23322
rect 42628 22982 42656 23287
rect 42800 23258 42852 23264
rect 42616 22976 42668 22982
rect 42616 22918 42668 22924
rect 42812 22642 42840 23258
rect 43916 23254 43944 23598
rect 43904 23248 43956 23254
rect 43902 23216 43904 23225
rect 43956 23216 43958 23225
rect 43902 23151 43958 23160
rect 44008 23118 44036 24006
rect 44100 23118 44128 26200
rect 44272 24948 44324 24954
rect 44272 24890 44324 24896
rect 44180 23860 44232 23866
rect 44180 23802 44232 23808
rect 42892 23112 42944 23118
rect 43996 23112 44048 23118
rect 42892 23054 42944 23060
rect 43534 23080 43590 23089
rect 42904 22778 42932 23054
rect 43996 23054 44048 23060
rect 44088 23112 44140 23118
rect 44088 23054 44140 23060
rect 43534 23015 43536 23024
rect 43588 23015 43590 23024
rect 43536 22986 43588 22992
rect 43996 22976 44048 22982
rect 43996 22918 44048 22924
rect 42892 22772 42944 22778
rect 42892 22714 42944 22720
rect 43720 22704 43772 22710
rect 43720 22646 43772 22652
rect 42800 22636 42852 22642
rect 42800 22578 42852 22584
rect 42614 22536 42670 22545
rect 42812 22522 42840 22578
rect 42614 22471 42616 22480
rect 42668 22471 42670 22480
rect 42720 22494 42840 22522
rect 43352 22568 43404 22574
rect 43352 22510 43404 22516
rect 42616 22442 42668 22448
rect 42720 22234 42748 22494
rect 42800 22432 42852 22438
rect 42800 22374 42852 22380
rect 42708 22228 42760 22234
rect 42708 22170 42760 22176
rect 42432 22160 42484 22166
rect 42432 22102 42484 22108
rect 42248 21684 42300 21690
rect 42248 21626 42300 21632
rect 42812 21593 42840 22374
rect 42950 22332 43258 22341
rect 42950 22330 42956 22332
rect 43012 22330 43036 22332
rect 43092 22330 43116 22332
rect 43172 22330 43196 22332
rect 43252 22330 43258 22332
rect 43012 22278 43014 22330
rect 43194 22278 43196 22330
rect 42950 22276 42956 22278
rect 43012 22276 43036 22278
rect 43092 22276 43116 22278
rect 43172 22276 43196 22278
rect 43252 22276 43258 22278
rect 42950 22267 43258 22276
rect 43364 22234 43392 22510
rect 43732 22234 43760 22646
rect 43904 22432 43956 22438
rect 43904 22374 43956 22380
rect 43352 22228 43404 22234
rect 43352 22170 43404 22176
rect 43720 22228 43772 22234
rect 43720 22170 43772 22176
rect 42892 21684 42944 21690
rect 42892 21626 42944 21632
rect 42798 21584 42854 21593
rect 42798 21519 42854 21528
rect 42904 21486 42932 21626
rect 42892 21480 42944 21486
rect 42892 21422 42944 21428
rect 42950 21244 43258 21253
rect 42950 21242 42956 21244
rect 43012 21242 43036 21244
rect 43092 21242 43116 21244
rect 43172 21242 43196 21244
rect 43252 21242 43258 21244
rect 43012 21190 43014 21242
rect 43194 21190 43196 21242
rect 42950 21188 42956 21190
rect 43012 21188 43036 21190
rect 43092 21188 43116 21190
rect 43172 21188 43196 21190
rect 43252 21188 43258 21190
rect 42950 21179 43258 21188
rect 42156 21072 42208 21078
rect 42156 21014 42208 21020
rect 42168 20874 42196 21014
rect 41420 20868 41472 20874
rect 41420 20810 41472 20816
rect 42156 20868 42208 20874
rect 42156 20810 42208 20816
rect 41432 20754 41460 20810
rect 41340 20726 41460 20754
rect 41340 20330 41368 20726
rect 41328 20324 41380 20330
rect 41328 20266 41380 20272
rect 42950 20156 43258 20165
rect 42950 20154 42956 20156
rect 43012 20154 43036 20156
rect 43092 20154 43116 20156
rect 43172 20154 43196 20156
rect 43252 20154 43258 20156
rect 43012 20102 43014 20154
rect 43194 20102 43196 20154
rect 42950 20100 42956 20102
rect 43012 20100 43036 20102
rect 43092 20100 43116 20102
rect 43172 20100 43196 20102
rect 43252 20100 43258 20102
rect 42950 20091 43258 20100
rect 41236 19984 41288 19990
rect 41236 19926 41288 19932
rect 41052 19916 41104 19922
rect 41052 19858 41104 19864
rect 41064 19786 41092 19858
rect 43916 19854 43944 22374
rect 44008 21690 44036 22918
rect 44192 22506 44220 23802
rect 44284 23730 44312 24890
rect 44546 24712 44602 24721
rect 44546 24647 44602 24656
rect 44272 23724 44324 23730
rect 44272 23666 44324 23672
rect 44560 22778 44588 24647
rect 44744 24206 44772 26200
rect 45388 24290 45416 26200
rect 45388 24262 45600 24290
rect 45572 24206 45600 24262
rect 44640 24200 44692 24206
rect 44640 24142 44692 24148
rect 44732 24200 44784 24206
rect 44732 24142 44784 24148
rect 45284 24200 45336 24206
rect 45284 24142 45336 24148
rect 45560 24200 45612 24206
rect 45560 24142 45612 24148
rect 44652 23322 44680 24142
rect 45296 23866 45324 24142
rect 46032 24138 46060 26200
rect 46662 25120 46718 25129
rect 46662 25055 46718 25064
rect 46570 24712 46626 24721
rect 46570 24647 46626 24656
rect 46020 24132 46072 24138
rect 46020 24074 46072 24080
rect 46112 24064 46164 24070
rect 46112 24006 46164 24012
rect 46204 24064 46256 24070
rect 46204 24006 46256 24012
rect 45284 23860 45336 23866
rect 45284 23802 45336 23808
rect 45374 23760 45430 23769
rect 45374 23695 45376 23704
rect 45428 23695 45430 23704
rect 45376 23666 45428 23672
rect 45190 23624 45246 23633
rect 45388 23610 45416 23666
rect 45388 23582 45508 23610
rect 45190 23559 45192 23568
rect 45244 23559 45246 23568
rect 45192 23530 45244 23536
rect 45376 23520 45428 23526
rect 45376 23462 45428 23468
rect 44640 23316 44692 23322
rect 44640 23258 44692 23264
rect 44548 22772 44600 22778
rect 44548 22714 44600 22720
rect 44180 22500 44232 22506
rect 44180 22442 44232 22448
rect 45388 21962 45416 23462
rect 45480 23322 45508 23582
rect 45468 23316 45520 23322
rect 45468 23258 45520 23264
rect 45376 21956 45428 21962
rect 45376 21898 45428 21904
rect 43996 21684 44048 21690
rect 43996 21626 44048 21632
rect 43904 19848 43956 19854
rect 43904 19790 43956 19796
rect 41052 19780 41104 19786
rect 41052 19722 41104 19728
rect 45284 19712 45336 19718
rect 45284 19654 45336 19660
rect 45296 19378 45324 19654
rect 41236 19372 41288 19378
rect 41236 19314 41288 19320
rect 45284 19372 45336 19378
rect 45284 19314 45336 19320
rect 41144 19304 41196 19310
rect 41144 19246 41196 19252
rect 41156 19174 41184 19246
rect 41144 19168 41196 19174
rect 41144 19110 41196 19116
rect 40682 18320 40738 18329
rect 40682 18255 40738 18264
rect 41052 17740 41104 17746
rect 41052 17682 41104 17688
rect 40592 17128 40644 17134
rect 40592 17070 40644 17076
rect 40408 17060 40460 17066
rect 40408 17002 40460 17008
rect 40224 16652 40276 16658
rect 40420 16640 40448 17002
rect 41064 16998 41092 17682
rect 41156 17270 41184 19110
rect 41144 17264 41196 17270
rect 41144 17206 41196 17212
rect 41052 16992 41104 16998
rect 41052 16934 41104 16940
rect 41156 16658 41184 17206
rect 41248 16726 41276 19314
rect 41604 19168 41656 19174
rect 41604 19110 41656 19116
rect 41616 18698 41644 19110
rect 42950 19068 43258 19077
rect 42950 19066 42956 19068
rect 43012 19066 43036 19068
rect 43092 19066 43116 19068
rect 43172 19066 43196 19068
rect 43252 19066 43258 19068
rect 43012 19014 43014 19066
rect 43194 19014 43196 19066
rect 42950 19012 42956 19014
rect 43012 19012 43036 19014
rect 43092 19012 43116 19014
rect 43172 19012 43196 19014
rect 43252 19012 43258 19014
rect 42950 19003 43258 19012
rect 42708 18896 42760 18902
rect 42708 18838 42760 18844
rect 41604 18692 41656 18698
rect 41604 18634 41656 18640
rect 42720 17241 42748 18838
rect 42950 17980 43258 17989
rect 42950 17978 42956 17980
rect 43012 17978 43036 17980
rect 43092 17978 43116 17980
rect 43172 17978 43196 17980
rect 43252 17978 43258 17980
rect 43012 17926 43014 17978
rect 43194 17926 43196 17978
rect 42950 17924 42956 17926
rect 43012 17924 43036 17926
rect 43092 17924 43116 17926
rect 43172 17924 43196 17926
rect 43252 17924 43258 17926
rect 42950 17915 43258 17924
rect 42706 17232 42762 17241
rect 42706 17167 42762 17176
rect 41328 17060 41380 17066
rect 41328 17002 41380 17008
rect 41340 16726 41368 17002
rect 42950 16892 43258 16901
rect 42950 16890 42956 16892
rect 43012 16890 43036 16892
rect 43092 16890 43116 16892
rect 43172 16890 43196 16892
rect 43252 16890 43258 16892
rect 43012 16838 43014 16890
rect 43194 16838 43196 16890
rect 42950 16836 42956 16838
rect 43012 16836 43036 16838
rect 43092 16836 43116 16838
rect 43172 16836 43196 16838
rect 43252 16836 43258 16838
rect 42950 16827 43258 16836
rect 46124 16726 46152 24006
rect 46216 21418 46244 24006
rect 46480 23656 46532 23662
rect 46480 23598 46532 23604
rect 46492 23186 46520 23598
rect 46480 23180 46532 23186
rect 46480 23122 46532 23128
rect 46584 22030 46612 24647
rect 46676 22642 46704 25055
rect 46756 24132 46808 24138
rect 46756 24074 46808 24080
rect 46768 23730 46796 24074
rect 46860 23798 46888 26302
rect 47306 26200 47362 27000
rect 47950 26200 48006 27000
rect 48594 26200 48650 27000
rect 49238 26200 49294 27000
rect 47320 24206 47348 26200
rect 47582 24304 47638 24313
rect 47492 24268 47544 24274
rect 47582 24239 47638 24248
rect 47492 24210 47544 24216
rect 47308 24200 47360 24206
rect 47308 24142 47360 24148
rect 46940 24064 46992 24070
rect 46940 24006 46992 24012
rect 46848 23792 46900 23798
rect 46848 23734 46900 23740
rect 46756 23724 46808 23730
rect 46756 23666 46808 23672
rect 46664 22636 46716 22642
rect 46664 22578 46716 22584
rect 46572 22024 46624 22030
rect 46572 21966 46624 21972
rect 46204 21412 46256 21418
rect 46204 21354 46256 21360
rect 46952 19553 46980 24006
rect 47124 23520 47176 23526
rect 47124 23462 47176 23468
rect 47136 22817 47164 23462
rect 47122 22808 47178 22817
rect 47320 22778 47348 24142
rect 47122 22743 47178 22752
rect 47308 22772 47360 22778
rect 47308 22714 47360 22720
rect 47504 21690 47532 24210
rect 47596 22642 47624 24239
rect 47964 24154 47992 26200
rect 48226 25528 48282 25537
rect 48226 25463 48282 25472
rect 48240 24274 48268 25463
rect 48320 24880 48372 24886
rect 48320 24822 48372 24828
rect 48228 24268 48280 24274
rect 48228 24210 48280 24216
rect 47872 24126 47992 24154
rect 47872 23730 47900 24126
rect 47950 23964 48258 23973
rect 47950 23962 47956 23964
rect 48012 23962 48036 23964
rect 48092 23962 48116 23964
rect 48172 23962 48196 23964
rect 48252 23962 48258 23964
rect 48012 23910 48014 23962
rect 48194 23910 48196 23962
rect 47950 23908 47956 23910
rect 48012 23908 48036 23910
rect 48092 23908 48116 23910
rect 48172 23908 48196 23910
rect 48252 23908 48258 23910
rect 47950 23899 48258 23908
rect 47860 23724 47912 23730
rect 47780 23684 47860 23712
rect 47780 23322 47808 23684
rect 47860 23666 47912 23672
rect 47858 23488 47914 23497
rect 47858 23423 47914 23432
rect 47768 23316 47820 23322
rect 47768 23258 47820 23264
rect 47676 23248 47728 23254
rect 47676 23190 47728 23196
rect 47584 22636 47636 22642
rect 47584 22578 47636 22584
rect 47688 21894 47716 23190
rect 47872 23118 47900 23423
rect 48332 23202 48360 24822
rect 48410 23896 48466 23905
rect 48410 23831 48466 23840
rect 48424 23662 48452 23831
rect 48608 23730 48636 26200
rect 48780 24200 48832 24206
rect 48778 24168 48780 24177
rect 48832 24168 48834 24177
rect 48778 24103 48834 24112
rect 48596 23724 48648 23730
rect 48596 23666 48648 23672
rect 48412 23656 48464 23662
rect 48412 23598 48464 23604
rect 48332 23174 48452 23202
rect 47860 23112 47912 23118
rect 48320 23112 48372 23118
rect 47860 23054 47912 23060
rect 48318 23080 48320 23089
rect 48372 23080 48374 23089
rect 47872 22778 47900 23054
rect 48318 23015 48374 23024
rect 47950 22876 48258 22885
rect 47950 22874 47956 22876
rect 48012 22874 48036 22876
rect 48092 22874 48116 22876
rect 48172 22874 48196 22876
rect 48252 22874 48258 22876
rect 48012 22822 48014 22874
rect 48194 22822 48196 22874
rect 47950 22820 47956 22822
rect 48012 22820 48036 22822
rect 48092 22820 48116 22822
rect 48172 22820 48196 22822
rect 48252 22820 48258 22822
rect 47950 22811 48258 22820
rect 48424 22778 48452 23174
rect 48608 23050 48636 23666
rect 49148 23520 49200 23526
rect 49148 23462 49200 23468
rect 48596 23044 48648 23050
rect 48596 22986 48648 22992
rect 48504 22976 48556 22982
rect 48504 22918 48556 22924
rect 47860 22772 47912 22778
rect 47860 22714 47912 22720
rect 48412 22772 48464 22778
rect 48412 22714 48464 22720
rect 48516 22094 48544 22918
rect 49056 22636 49108 22642
rect 49056 22578 49108 22584
rect 48596 22432 48648 22438
rect 48596 22374 48648 22380
rect 48332 22066 48544 22094
rect 47860 22024 47912 22030
rect 47860 21966 47912 21972
rect 47676 21888 47728 21894
rect 47676 21830 47728 21836
rect 47768 21888 47820 21894
rect 47768 21830 47820 21836
rect 47492 21684 47544 21690
rect 47492 21626 47544 21632
rect 47780 21622 47808 21830
rect 47768 21616 47820 21622
rect 47768 21558 47820 21564
rect 47872 21554 47900 21966
rect 47950 21788 48258 21797
rect 47950 21786 47956 21788
rect 48012 21786 48036 21788
rect 48092 21786 48116 21788
rect 48172 21786 48196 21788
rect 48252 21786 48258 21788
rect 48012 21734 48014 21786
rect 48194 21734 48196 21786
rect 47950 21732 47956 21734
rect 48012 21732 48036 21734
rect 48092 21732 48116 21734
rect 48172 21732 48196 21734
rect 48252 21732 48258 21734
rect 47950 21723 48258 21732
rect 47860 21548 47912 21554
rect 47860 21490 47912 21496
rect 47950 20700 48258 20709
rect 47950 20698 47956 20700
rect 48012 20698 48036 20700
rect 48092 20698 48116 20700
rect 48172 20698 48196 20700
rect 48252 20698 48258 20700
rect 48012 20646 48014 20698
rect 48194 20646 48196 20698
rect 47950 20644 47956 20646
rect 48012 20644 48036 20646
rect 48092 20644 48116 20646
rect 48172 20644 48196 20646
rect 48252 20644 48258 20646
rect 47950 20635 48258 20644
rect 48332 20369 48360 22066
rect 48412 21888 48464 21894
rect 48412 21830 48464 21836
rect 48504 21888 48556 21894
rect 48504 21830 48556 21836
rect 48424 20942 48452 21830
rect 48412 20936 48464 20942
rect 48412 20878 48464 20884
rect 48318 20360 48374 20369
rect 48318 20295 48374 20304
rect 48412 20256 48464 20262
rect 48412 20198 48464 20204
rect 47950 19612 48258 19621
rect 47950 19610 47956 19612
rect 48012 19610 48036 19612
rect 48092 19610 48116 19612
rect 48172 19610 48196 19612
rect 48252 19610 48258 19612
rect 48012 19558 48014 19610
rect 48194 19558 48196 19610
rect 47950 19556 47956 19558
rect 48012 19556 48036 19558
rect 48092 19556 48116 19558
rect 48172 19556 48196 19558
rect 48252 19556 48258 19558
rect 46938 19544 46994 19553
rect 47950 19547 48258 19556
rect 46938 19479 46994 19488
rect 48424 19446 48452 20198
rect 48516 19825 48544 21830
rect 48608 20058 48636 22374
rect 49068 22273 49096 22578
rect 49054 22264 49110 22273
rect 49054 22199 49110 22208
rect 48780 22024 48832 22030
rect 48780 21966 48832 21972
rect 48792 21865 48820 21966
rect 48778 21856 48834 21865
rect 48778 21791 48834 21800
rect 48792 21690 48820 21791
rect 49068 21690 49096 22199
rect 49160 21962 49188 23462
rect 49252 23186 49280 26200
rect 49240 23180 49292 23186
rect 49240 23122 49292 23128
rect 49332 23112 49384 23118
rect 49332 23054 49384 23060
rect 49240 22976 49292 22982
rect 49240 22918 49292 22924
rect 49252 22098 49280 22918
rect 49344 22681 49372 23054
rect 49330 22672 49386 22681
rect 49330 22607 49386 22616
rect 49344 22234 49372 22607
rect 49332 22228 49384 22234
rect 49332 22170 49384 22176
rect 49240 22092 49292 22098
rect 49240 22034 49292 22040
rect 49148 21956 49200 21962
rect 49148 21898 49200 21904
rect 48780 21684 48832 21690
rect 48780 21626 48832 21632
rect 49056 21684 49108 21690
rect 49056 21626 49108 21632
rect 49056 21548 49108 21554
rect 49056 21490 49108 21496
rect 49068 21049 49096 21490
rect 49160 21457 49188 21898
rect 49146 21448 49202 21457
rect 49146 21383 49202 21392
rect 49240 21344 49292 21350
rect 49240 21286 49292 21292
rect 49054 21040 49110 21049
rect 49054 20975 49110 20984
rect 49056 20936 49108 20942
rect 49056 20878 49108 20884
rect 48964 20800 49016 20806
rect 48964 20742 49016 20748
rect 48976 20482 49004 20742
rect 49068 20641 49096 20878
rect 49054 20632 49110 20641
rect 49054 20567 49110 20576
rect 48976 20466 49096 20482
rect 48780 20460 48832 20466
rect 48976 20460 49108 20466
rect 48976 20454 49056 20460
rect 48780 20402 48832 20408
rect 49056 20402 49108 20408
rect 48792 20233 48820 20402
rect 48778 20224 48834 20233
rect 48778 20159 48834 20168
rect 48792 20058 48820 20159
rect 48596 20052 48648 20058
rect 48596 19994 48648 20000
rect 48780 20052 48832 20058
rect 48780 19994 48832 20000
rect 49068 19825 49096 20402
rect 48502 19816 48558 19825
rect 48502 19751 48558 19760
rect 49054 19816 49110 19825
rect 49054 19751 49110 19760
rect 49252 19514 49280 21286
rect 49332 19780 49384 19786
rect 49332 19722 49384 19728
rect 49240 19508 49292 19514
rect 49240 19450 49292 19456
rect 48412 19440 48464 19446
rect 49344 19417 49372 19722
rect 48412 19382 48464 19388
rect 49330 19408 49386 19417
rect 49148 19372 49200 19378
rect 49330 19343 49386 19352
rect 49148 19314 49200 19320
rect 49056 19168 49108 19174
rect 49056 19110 49108 19116
rect 49068 18850 49096 19110
rect 49160 19009 49188 19314
rect 49146 19000 49202 19009
rect 49146 18935 49202 18944
rect 49068 18822 49188 18850
rect 49160 18766 49188 18822
rect 48780 18760 48832 18766
rect 48780 18702 48832 18708
rect 49148 18760 49200 18766
rect 49148 18702 49200 18708
rect 48412 18624 48464 18630
rect 48792 18601 48820 18702
rect 48412 18566 48464 18572
rect 48778 18592 48834 18601
rect 47950 18524 48258 18533
rect 47950 18522 47956 18524
rect 48012 18522 48036 18524
rect 48092 18522 48116 18524
rect 48172 18522 48196 18524
rect 48252 18522 48258 18524
rect 48012 18470 48014 18522
rect 48194 18470 48196 18522
rect 47950 18468 47956 18470
rect 48012 18468 48036 18470
rect 48092 18468 48116 18470
rect 48172 18468 48196 18470
rect 48252 18468 48258 18470
rect 47950 18459 48258 18468
rect 48424 18290 48452 18566
rect 48778 18527 48834 18536
rect 48792 18426 48820 18527
rect 48780 18420 48832 18426
rect 48780 18362 48832 18368
rect 48412 18284 48464 18290
rect 48412 18226 48464 18232
rect 49056 18284 49108 18290
rect 49056 18226 49108 18232
rect 48320 18080 48372 18086
rect 48320 18022 48372 18028
rect 47950 17436 48258 17445
rect 47950 17434 47956 17436
rect 48012 17434 48036 17436
rect 48092 17434 48116 17436
rect 48172 17434 48196 17436
rect 48252 17434 48258 17436
rect 48012 17382 48014 17434
rect 48194 17382 48196 17434
rect 47950 17380 47956 17382
rect 48012 17380 48036 17382
rect 48092 17380 48116 17382
rect 48172 17380 48196 17382
rect 48252 17380 48258 17382
rect 47950 17371 48258 17380
rect 48332 17338 48360 18022
rect 48596 17876 48648 17882
rect 48596 17818 48648 17824
rect 48412 17604 48464 17610
rect 48412 17546 48464 17552
rect 48504 17604 48556 17610
rect 48504 17546 48556 17552
rect 48424 17338 48452 17546
rect 48320 17332 48372 17338
rect 48320 17274 48372 17280
rect 48412 17332 48464 17338
rect 48412 17274 48464 17280
rect 48516 16794 48544 17546
rect 48608 17338 48636 17818
rect 49068 17785 49096 18226
rect 49160 18193 49188 18702
rect 49146 18184 49202 18193
rect 49146 18119 49202 18128
rect 49054 17776 49110 17785
rect 49054 17711 49110 17720
rect 49056 17672 49108 17678
rect 49056 17614 49108 17620
rect 49068 17377 49096 17614
rect 49148 17536 49200 17542
rect 49148 17478 49200 17484
rect 49054 17368 49110 17377
rect 48596 17332 48648 17338
rect 49160 17354 49188 17478
rect 49160 17326 49280 17354
rect 49054 17303 49110 17312
rect 48596 17274 48648 17280
rect 49252 17202 49280 17326
rect 48780 17196 48832 17202
rect 48780 17138 48832 17144
rect 49240 17196 49292 17202
rect 49240 17138 49292 17144
rect 48792 16969 48820 17138
rect 48778 16960 48834 16969
rect 48778 16895 48834 16904
rect 48792 16794 48820 16895
rect 48504 16788 48556 16794
rect 48504 16730 48556 16736
rect 48780 16788 48832 16794
rect 48780 16730 48832 16736
rect 41236 16720 41288 16726
rect 41236 16662 41288 16668
rect 41328 16720 41380 16726
rect 41328 16662 41380 16668
rect 46112 16720 46164 16726
rect 46112 16662 46164 16668
rect 40500 16652 40552 16658
rect 40420 16612 40500 16640
rect 40224 16594 40276 16600
rect 40500 16594 40552 16600
rect 40592 16652 40644 16658
rect 40592 16594 40644 16600
rect 41144 16652 41196 16658
rect 41144 16594 41196 16600
rect 40604 16046 40632 16594
rect 41604 16584 41656 16590
rect 41604 16526 41656 16532
rect 49148 16584 49200 16590
rect 49252 16561 49280 17138
rect 49148 16526 49200 16532
rect 49238 16552 49294 16561
rect 41328 16448 41380 16454
rect 41328 16390 41380 16396
rect 41340 16182 41368 16390
rect 41328 16176 41380 16182
rect 41328 16118 41380 16124
rect 40316 16040 40368 16046
rect 40316 15982 40368 15988
rect 40592 16040 40644 16046
rect 40592 15982 40644 15988
rect 41052 16040 41104 16046
rect 41052 15982 41104 15988
rect 40328 15570 40356 15982
rect 40316 15564 40368 15570
rect 40316 15506 40368 15512
rect 41064 15366 41092 15982
rect 41340 15434 41368 16118
rect 41616 15910 41644 16526
rect 48780 16448 48832 16454
rect 48780 16390 48832 16396
rect 47950 16348 48258 16357
rect 47950 16346 47956 16348
rect 48012 16346 48036 16348
rect 48092 16346 48116 16348
rect 48172 16346 48196 16348
rect 48252 16346 48258 16348
rect 48012 16294 48014 16346
rect 48194 16294 48196 16346
rect 47950 16292 47956 16294
rect 48012 16292 48036 16294
rect 48092 16292 48116 16294
rect 48172 16292 48196 16294
rect 48252 16292 48258 16294
rect 47950 16283 48258 16292
rect 48792 16153 48820 16390
rect 49160 16153 49188 16526
rect 49238 16487 49294 16496
rect 48778 16144 48834 16153
rect 48688 16108 48740 16114
rect 49146 16144 49202 16153
rect 48778 16079 48834 16088
rect 49056 16108 49108 16114
rect 48688 16050 48740 16056
rect 49146 16079 49202 16088
rect 49056 16050 49108 16056
rect 41604 15904 41656 15910
rect 41604 15846 41656 15852
rect 41616 15706 41644 15846
rect 42950 15804 43258 15813
rect 42950 15802 42956 15804
rect 43012 15802 43036 15804
rect 43092 15802 43116 15804
rect 43172 15802 43196 15804
rect 43252 15802 43258 15804
rect 43012 15750 43014 15802
rect 43194 15750 43196 15802
rect 42950 15748 42956 15750
rect 43012 15748 43036 15750
rect 43092 15748 43116 15750
rect 43172 15748 43196 15750
rect 43252 15748 43258 15750
rect 42950 15739 43258 15748
rect 48700 15706 48728 16050
rect 49068 15745 49096 16050
rect 49238 16008 49294 16017
rect 49238 15943 49240 15952
rect 49292 15943 49294 15952
rect 49240 15914 49292 15920
rect 49054 15736 49110 15745
rect 41604 15700 41656 15706
rect 41604 15642 41656 15648
rect 48688 15700 48740 15706
rect 49054 15671 49110 15680
rect 48688 15642 48740 15648
rect 49332 15496 49384 15502
rect 49332 15438 49384 15444
rect 41328 15428 41380 15434
rect 41328 15370 41380 15376
rect 41052 15360 41104 15366
rect 49344 15337 49372 15438
rect 41052 15302 41104 15308
rect 49330 15328 49386 15337
rect 47950 15260 48258 15269
rect 49330 15263 49386 15272
rect 47950 15258 47956 15260
rect 48012 15258 48036 15260
rect 48092 15258 48116 15260
rect 48172 15258 48196 15260
rect 48252 15258 48258 15260
rect 48012 15206 48014 15258
rect 48194 15206 48196 15258
rect 47950 15204 47956 15206
rect 48012 15204 48036 15206
rect 48092 15204 48116 15206
rect 48172 15204 48196 15206
rect 48252 15204 48258 15206
rect 47950 15195 48258 15204
rect 40132 15156 40184 15162
rect 40132 15098 40184 15104
rect 40316 15156 40368 15162
rect 40316 15098 40368 15104
rect 39856 15020 39908 15026
rect 39856 14962 39908 14968
rect 40328 14890 40356 15098
rect 48412 15088 48464 15094
rect 48412 15030 48464 15036
rect 49238 15056 49294 15065
rect 40316 14884 40368 14890
rect 40316 14826 40368 14832
rect 45836 14816 45888 14822
rect 45836 14758 45888 14764
rect 42950 14716 43258 14725
rect 42950 14714 42956 14716
rect 43012 14714 43036 14716
rect 43092 14714 43116 14716
rect 43172 14714 43196 14716
rect 43252 14714 43258 14716
rect 43012 14662 43014 14714
rect 43194 14662 43196 14714
rect 42950 14660 42956 14662
rect 43012 14660 43036 14662
rect 43092 14660 43116 14662
rect 43172 14660 43196 14662
rect 43252 14660 43258 14662
rect 42950 14651 43258 14660
rect 39764 14612 39816 14618
rect 39764 14554 39816 14560
rect 39580 14408 39632 14414
rect 39580 14350 39632 14356
rect 39304 14272 39356 14278
rect 39304 14214 39356 14220
rect 39316 14006 39344 14214
rect 39304 14000 39356 14006
rect 39304 13942 39356 13948
rect 39776 13938 39804 14554
rect 39946 14376 40002 14385
rect 39946 14311 40002 14320
rect 39396 13932 39448 13938
rect 39396 13874 39448 13880
rect 39764 13932 39816 13938
rect 39764 13874 39816 13880
rect 38384 13728 38436 13734
rect 38384 13670 38436 13676
rect 37832 13524 37884 13530
rect 37832 13466 37884 13472
rect 38752 13524 38804 13530
rect 38752 13466 38804 13472
rect 37844 13326 37872 13466
rect 37832 13320 37884 13326
rect 37832 13262 37884 13268
rect 37740 13184 37792 13190
rect 37740 13126 37792 13132
rect 37752 12918 37780 13126
rect 37844 12986 37872 13262
rect 37950 13084 38258 13093
rect 37950 13082 37956 13084
rect 38012 13082 38036 13084
rect 38092 13082 38116 13084
rect 38172 13082 38196 13084
rect 38252 13082 38258 13084
rect 38012 13030 38014 13082
rect 38194 13030 38196 13082
rect 37950 13028 37956 13030
rect 38012 13028 38036 13030
rect 38092 13028 38116 13030
rect 38172 13028 38196 13030
rect 38252 13028 38258 13030
rect 37950 13019 38258 13028
rect 37832 12980 37884 12986
rect 37832 12922 37884 12928
rect 38764 12918 38792 13466
rect 37740 12912 37792 12918
rect 37740 12854 37792 12860
rect 38752 12912 38804 12918
rect 38752 12854 38804 12860
rect 37568 12702 37872 12730
rect 37648 12436 37700 12442
rect 37648 12378 37700 12384
rect 37660 12306 37688 12378
rect 37464 12300 37516 12306
rect 37464 12242 37516 12248
rect 37648 12300 37700 12306
rect 37648 12242 37700 12248
rect 37740 12300 37792 12306
rect 37740 12242 37792 12248
rect 37464 12096 37516 12102
rect 37464 12038 37516 12044
rect 37372 11824 37424 11830
rect 37372 11766 37424 11772
rect 37372 11552 37424 11558
rect 37372 11494 37424 11500
rect 37384 11082 37412 11494
rect 37372 11076 37424 11082
rect 37372 11018 37424 11024
rect 37476 11014 37504 12038
rect 37752 11898 37780 12242
rect 37844 11898 37872 12702
rect 39408 12434 39436 13874
rect 39960 12918 39988 14311
rect 41512 14068 41564 14074
rect 41512 14010 41564 14016
rect 41524 13326 41552 14010
rect 45848 13938 45876 14758
rect 48320 14272 48372 14278
rect 48320 14214 48372 14220
rect 47950 14172 48258 14181
rect 47950 14170 47956 14172
rect 48012 14170 48036 14172
rect 48092 14170 48116 14172
rect 48172 14170 48196 14172
rect 48252 14170 48258 14172
rect 48012 14118 48014 14170
rect 48194 14118 48196 14170
rect 47950 14116 47956 14118
rect 48012 14116 48036 14118
rect 48092 14116 48116 14118
rect 48172 14116 48196 14118
rect 48252 14116 48258 14118
rect 47950 14107 48258 14116
rect 47032 14068 47084 14074
rect 47032 14010 47084 14016
rect 45836 13932 45888 13938
rect 45836 13874 45888 13880
rect 46480 13864 46532 13870
rect 46480 13806 46532 13812
rect 42950 13628 43258 13637
rect 42950 13626 42956 13628
rect 43012 13626 43036 13628
rect 43092 13626 43116 13628
rect 43172 13626 43196 13628
rect 43252 13626 43258 13628
rect 43012 13574 43014 13626
rect 43194 13574 43196 13626
rect 42950 13572 42956 13574
rect 43012 13572 43036 13574
rect 43092 13572 43116 13574
rect 43172 13572 43196 13574
rect 43252 13572 43258 13574
rect 42950 13563 43258 13572
rect 46492 13326 46520 13806
rect 41512 13320 41564 13326
rect 41512 13262 41564 13268
rect 46480 13320 46532 13326
rect 46480 13262 46532 13268
rect 46112 13184 46164 13190
rect 46112 13126 46164 13132
rect 39948 12912 40000 12918
rect 39948 12854 40000 12860
rect 46124 12850 46152 13126
rect 47044 12850 47072 14010
rect 48332 13954 48360 14214
rect 48424 14074 48452 15030
rect 49056 15020 49108 15026
rect 49238 14991 49294 15000
rect 49056 14962 49108 14968
rect 49068 14929 49096 14962
rect 49054 14920 49110 14929
rect 49054 14855 49110 14864
rect 49146 14512 49202 14521
rect 49146 14447 49202 14456
rect 49160 14414 49188 14447
rect 49148 14408 49200 14414
rect 49148 14350 49200 14356
rect 49146 14104 49202 14113
rect 48412 14068 48464 14074
rect 49252 14074 49280 14991
rect 49146 14039 49202 14048
rect 49240 14068 49292 14074
rect 48412 14010 48464 14016
rect 49160 14006 49188 14039
rect 49240 14010 49292 14016
rect 48240 13938 48360 13954
rect 49148 14000 49200 14006
rect 49148 13942 49200 13948
rect 48228 13932 48360 13938
rect 48280 13926 48360 13932
rect 48228 13874 48280 13880
rect 48240 13705 48268 13874
rect 48226 13696 48282 13705
rect 48226 13631 48282 13640
rect 49146 13288 49202 13297
rect 49146 13223 49148 13232
rect 49200 13223 49202 13232
rect 49148 13194 49200 13200
rect 47950 13084 48258 13093
rect 47950 13082 47956 13084
rect 48012 13082 48036 13084
rect 48092 13082 48116 13084
rect 48172 13082 48196 13084
rect 48252 13082 48258 13084
rect 48012 13030 48014 13082
rect 48194 13030 48196 13082
rect 47950 13028 47956 13030
rect 48012 13028 48036 13030
rect 48092 13028 48116 13030
rect 48172 13028 48196 13030
rect 48252 13028 48258 13030
rect 47950 13019 48258 13028
rect 49146 12880 49202 12889
rect 46112 12844 46164 12850
rect 46112 12786 46164 12792
rect 47032 12844 47084 12850
rect 49146 12815 49148 12824
rect 47032 12786 47084 12792
rect 49200 12815 49202 12824
rect 49148 12786 49200 12792
rect 47032 12708 47084 12714
rect 47032 12650 47084 12656
rect 39488 12640 39540 12646
rect 39488 12582 39540 12588
rect 39316 12406 39436 12434
rect 39316 12170 39344 12406
rect 39304 12164 39356 12170
rect 39304 12106 39356 12112
rect 38660 12096 38712 12102
rect 38660 12038 38712 12044
rect 37950 11996 38258 12005
rect 37950 11994 37956 11996
rect 38012 11994 38036 11996
rect 38092 11994 38116 11996
rect 38172 11994 38196 11996
rect 38252 11994 38258 11996
rect 38012 11942 38014 11994
rect 38194 11942 38196 11994
rect 37950 11940 37956 11942
rect 38012 11940 38036 11942
rect 38092 11940 38116 11942
rect 38172 11940 38196 11942
rect 38252 11940 38258 11942
rect 37950 11931 38258 11940
rect 38672 11898 38700 12038
rect 37740 11892 37792 11898
rect 37740 11834 37792 11840
rect 37832 11892 37884 11898
rect 37832 11834 37884 11840
rect 38660 11892 38712 11898
rect 38660 11834 38712 11840
rect 39028 11756 39080 11762
rect 39028 11698 39080 11704
rect 37464 11008 37516 11014
rect 37464 10950 37516 10956
rect 37950 10908 38258 10917
rect 37950 10906 37956 10908
rect 38012 10906 38036 10908
rect 38092 10906 38116 10908
rect 38172 10906 38196 10908
rect 38252 10906 38258 10908
rect 38012 10854 38014 10906
rect 38194 10854 38196 10906
rect 37950 10852 37956 10854
rect 38012 10852 38036 10854
rect 38092 10852 38116 10854
rect 38172 10852 38196 10854
rect 38252 10852 38258 10854
rect 37950 10843 38258 10852
rect 38566 10160 38622 10169
rect 38566 10095 38622 10104
rect 38580 9994 38608 10095
rect 38568 9988 38620 9994
rect 38568 9930 38620 9936
rect 38384 9920 38436 9926
rect 38384 9862 38436 9868
rect 37950 9820 38258 9829
rect 37950 9818 37956 9820
rect 38012 9818 38036 9820
rect 38092 9818 38116 9820
rect 38172 9818 38196 9820
rect 38252 9818 38258 9820
rect 38012 9766 38014 9818
rect 38194 9766 38196 9818
rect 37950 9764 37956 9766
rect 38012 9764 38036 9766
rect 38092 9764 38116 9766
rect 38172 9764 38196 9766
rect 38252 9764 38258 9766
rect 37950 9755 38258 9764
rect 38396 9722 38424 9862
rect 38384 9716 38436 9722
rect 38384 9658 38436 9664
rect 37950 8732 38258 8741
rect 37950 8730 37956 8732
rect 38012 8730 38036 8732
rect 38092 8730 38116 8732
rect 38172 8730 38196 8732
rect 38252 8730 38258 8732
rect 38012 8678 38014 8730
rect 38194 8678 38196 8730
rect 37950 8676 37956 8678
rect 38012 8676 38036 8678
rect 38092 8676 38116 8678
rect 38172 8676 38196 8678
rect 38252 8676 38258 8678
rect 37950 8667 38258 8676
rect 38752 8424 38804 8430
rect 38752 8366 38804 8372
rect 38764 7818 38792 8366
rect 39040 7886 39068 11698
rect 39316 11354 39344 12106
rect 39500 11354 39528 12582
rect 42950 12540 43258 12549
rect 42950 12538 42956 12540
rect 43012 12538 43036 12540
rect 43092 12538 43116 12540
rect 43172 12538 43196 12540
rect 43252 12538 43258 12540
rect 43012 12486 43014 12538
rect 43194 12486 43196 12538
rect 42950 12484 42956 12486
rect 43012 12484 43036 12486
rect 43092 12484 43116 12486
rect 43172 12484 43196 12486
rect 43252 12484 43258 12486
rect 42950 12475 43258 12484
rect 43352 12164 43404 12170
rect 43352 12106 43404 12112
rect 40776 12096 40828 12102
rect 40776 12038 40828 12044
rect 40788 11830 40816 12038
rect 40776 11824 40828 11830
rect 40776 11766 40828 11772
rect 39948 11756 40000 11762
rect 39948 11698 40000 11704
rect 39304 11348 39356 11354
rect 39304 11290 39356 11296
rect 39488 11348 39540 11354
rect 39488 11290 39540 11296
rect 39500 11150 39528 11290
rect 39488 11144 39540 11150
rect 39960 11121 39988 11698
rect 40224 11552 40276 11558
rect 40224 11494 40276 11500
rect 40236 11150 40264 11494
rect 42950 11452 43258 11461
rect 42950 11450 42956 11452
rect 43012 11450 43036 11452
rect 43092 11450 43116 11452
rect 43172 11450 43196 11452
rect 43252 11450 43258 11452
rect 43012 11398 43014 11450
rect 43194 11398 43196 11450
rect 42950 11396 42956 11398
rect 43012 11396 43036 11398
rect 43092 11396 43116 11398
rect 43172 11396 43196 11398
rect 43252 11396 43258 11398
rect 42950 11387 43258 11396
rect 41604 11348 41656 11354
rect 41604 11290 41656 11296
rect 40224 11144 40276 11150
rect 39488 11086 39540 11092
rect 39946 11112 40002 11121
rect 40224 11086 40276 11092
rect 39946 11047 40002 11056
rect 39762 10704 39818 10713
rect 39762 10639 39764 10648
rect 39816 10639 39818 10648
rect 39764 10610 39816 10616
rect 41616 10062 41644 11290
rect 42950 10364 43258 10373
rect 42950 10362 42956 10364
rect 43012 10362 43036 10364
rect 43092 10362 43116 10364
rect 43172 10362 43196 10364
rect 43252 10362 43258 10364
rect 43012 10310 43014 10362
rect 43194 10310 43196 10362
rect 42950 10308 42956 10310
rect 43012 10308 43036 10310
rect 43092 10308 43116 10310
rect 43172 10308 43196 10310
rect 43252 10308 43258 10310
rect 42950 10299 43258 10308
rect 41604 10056 41656 10062
rect 41604 9998 41656 10004
rect 43364 9586 43392 12106
rect 45928 12096 45980 12102
rect 45928 12038 45980 12044
rect 45940 11762 45968 12038
rect 45928 11756 45980 11762
rect 45928 11698 45980 11704
rect 43720 11620 43772 11626
rect 43720 11562 43772 11568
rect 46296 11620 46348 11626
rect 46296 11562 46348 11568
rect 43352 9580 43404 9586
rect 43352 9522 43404 9528
rect 42950 9276 43258 9285
rect 42950 9274 42956 9276
rect 43012 9274 43036 9276
rect 43092 9274 43116 9276
rect 43172 9274 43196 9276
rect 43252 9274 43258 9276
rect 43012 9222 43014 9274
rect 43194 9222 43196 9274
rect 42950 9220 42956 9222
rect 43012 9220 43036 9222
rect 43092 9220 43116 9222
rect 43172 9220 43196 9222
rect 43252 9220 43258 9222
rect 42950 9211 43258 9220
rect 43628 9172 43680 9178
rect 43628 9114 43680 9120
rect 39580 8832 39632 8838
rect 39580 8774 39632 8780
rect 39592 8566 39620 8774
rect 40224 8628 40276 8634
rect 40224 8570 40276 8576
rect 39580 8560 39632 8566
rect 39580 8502 39632 8508
rect 40132 8356 40184 8362
rect 40132 8298 40184 8304
rect 39028 7880 39080 7886
rect 39028 7822 39080 7828
rect 38752 7812 38804 7818
rect 38752 7754 38804 7760
rect 40040 7812 40092 7818
rect 40040 7754 40092 7760
rect 38660 7744 38712 7750
rect 38660 7686 38712 7692
rect 37950 7644 38258 7653
rect 37950 7642 37956 7644
rect 38012 7642 38036 7644
rect 38092 7642 38116 7644
rect 38172 7642 38196 7644
rect 38252 7642 38258 7644
rect 38012 7590 38014 7642
rect 38194 7590 38196 7642
rect 37950 7588 37956 7590
rect 38012 7588 38036 7590
rect 38092 7588 38116 7590
rect 38172 7588 38196 7590
rect 38252 7588 38258 7590
rect 37950 7579 38258 7588
rect 38672 7546 38700 7686
rect 38660 7540 38712 7546
rect 38660 7482 38712 7488
rect 37372 7200 37424 7206
rect 37372 7142 37424 7148
rect 37924 7200 37976 7206
rect 37924 7142 37976 7148
rect 37280 6180 37332 6186
rect 37280 6122 37332 6128
rect 37004 4684 37056 4690
rect 37004 4626 37056 4632
rect 37292 4146 37320 6122
rect 37384 5234 37412 7142
rect 37936 6934 37964 7142
rect 37924 6928 37976 6934
rect 37924 6870 37976 6876
rect 40052 6798 40080 7754
rect 40144 7478 40172 8298
rect 40132 7472 40184 7478
rect 40132 7414 40184 7420
rect 40132 6860 40184 6866
rect 40132 6802 40184 6808
rect 40040 6792 40092 6798
rect 40040 6734 40092 6740
rect 37950 6556 38258 6565
rect 37950 6554 37956 6556
rect 38012 6554 38036 6556
rect 38092 6554 38116 6556
rect 38172 6554 38196 6556
rect 38252 6554 38258 6556
rect 38012 6502 38014 6554
rect 38194 6502 38196 6554
rect 37950 6500 37956 6502
rect 38012 6500 38036 6502
rect 38092 6500 38116 6502
rect 38172 6500 38196 6502
rect 38252 6500 38258 6502
rect 37950 6491 38258 6500
rect 37648 6112 37700 6118
rect 37648 6054 37700 6060
rect 37660 5914 37688 6054
rect 37648 5908 37700 5914
rect 37648 5850 37700 5856
rect 37950 5468 38258 5477
rect 37950 5466 37956 5468
rect 38012 5466 38036 5468
rect 38092 5466 38116 5468
rect 38172 5466 38196 5468
rect 38252 5466 38258 5468
rect 38012 5414 38014 5466
rect 38194 5414 38196 5466
rect 37950 5412 37956 5414
rect 38012 5412 38036 5414
rect 38092 5412 38116 5414
rect 38172 5412 38196 5414
rect 38252 5412 38258 5414
rect 37950 5403 38258 5412
rect 37372 5228 37424 5234
rect 37372 5170 37424 5176
rect 37832 5024 37884 5030
rect 37832 4966 37884 4972
rect 37844 4758 37872 4966
rect 40144 4826 40172 6802
rect 40236 6390 40264 8570
rect 42950 8188 43258 8197
rect 42950 8186 42956 8188
rect 43012 8186 43036 8188
rect 43092 8186 43116 8188
rect 43172 8186 43196 8188
rect 43252 8186 43258 8188
rect 43012 8134 43014 8186
rect 43194 8134 43196 8186
rect 42950 8132 42956 8134
rect 43012 8132 43036 8134
rect 43092 8132 43116 8134
rect 43172 8132 43196 8134
rect 43252 8132 43258 8134
rect 42950 8123 43258 8132
rect 42950 7100 43258 7109
rect 42950 7098 42956 7100
rect 43012 7098 43036 7100
rect 43092 7098 43116 7100
rect 43172 7098 43196 7100
rect 43252 7098 43258 7100
rect 43012 7046 43014 7098
rect 43194 7046 43196 7098
rect 42950 7044 42956 7046
rect 43012 7044 43036 7046
rect 43092 7044 43116 7046
rect 43172 7044 43196 7046
rect 43252 7044 43258 7046
rect 42950 7035 43258 7044
rect 43640 6914 43668 9114
rect 43732 8974 43760 11562
rect 45744 11076 45796 11082
rect 45744 11018 45796 11024
rect 45756 10062 45784 11018
rect 46308 10062 46336 11562
rect 47044 11150 47072 12650
rect 47952 12640 48004 12646
rect 47952 12582 48004 12588
rect 47964 12238 47992 12582
rect 49146 12472 49202 12481
rect 49146 12407 49202 12416
rect 49160 12306 49188 12407
rect 49148 12300 49200 12306
rect 49148 12242 49200 12248
rect 47952 12232 48004 12238
rect 47952 12174 48004 12180
rect 49146 12064 49202 12073
rect 47950 11996 48258 12005
rect 49146 11999 49202 12008
rect 47950 11994 47956 11996
rect 48012 11994 48036 11996
rect 48092 11994 48116 11996
rect 48172 11994 48196 11996
rect 48252 11994 48258 11996
rect 48012 11942 48014 11994
rect 48194 11942 48196 11994
rect 47950 11940 47956 11942
rect 48012 11940 48036 11942
rect 48092 11940 48116 11942
rect 48172 11940 48196 11942
rect 48252 11940 48258 11942
rect 47950 11931 48258 11940
rect 49160 11830 49188 11999
rect 49148 11824 49200 11830
rect 49148 11766 49200 11772
rect 49146 11656 49202 11665
rect 49146 11591 49202 11600
rect 49160 11218 49188 11591
rect 49238 11248 49294 11257
rect 49148 11212 49200 11218
rect 49238 11183 49294 11192
rect 49148 11154 49200 11160
rect 47032 11144 47084 11150
rect 47032 11086 47084 11092
rect 46940 11076 46992 11082
rect 46940 11018 46992 11024
rect 46952 10674 46980 11018
rect 47950 10908 48258 10917
rect 47950 10906 47956 10908
rect 48012 10906 48036 10908
rect 48092 10906 48116 10908
rect 48172 10906 48196 10908
rect 48252 10906 48258 10908
rect 48012 10854 48014 10906
rect 48194 10854 48196 10906
rect 47950 10852 47956 10854
rect 48012 10852 48036 10854
rect 48092 10852 48116 10854
rect 48172 10852 48196 10854
rect 48252 10852 48258 10854
rect 47950 10843 48258 10852
rect 49146 10840 49202 10849
rect 49146 10775 49202 10784
rect 46940 10668 46992 10674
rect 46940 10610 46992 10616
rect 46940 10532 46992 10538
rect 46940 10474 46992 10480
rect 45744 10056 45796 10062
rect 45744 9998 45796 10004
rect 46296 10056 46348 10062
rect 46296 9998 46348 10004
rect 46020 9988 46072 9994
rect 46020 9930 46072 9936
rect 45836 9920 45888 9926
rect 45836 9862 45888 9868
rect 43720 8968 43772 8974
rect 43720 8910 43772 8916
rect 45848 8498 45876 9862
rect 46032 8498 46060 9930
rect 45836 8492 45888 8498
rect 45836 8434 45888 8440
rect 46020 8492 46072 8498
rect 46020 8434 46072 8440
rect 46848 8424 46900 8430
rect 46848 8366 46900 8372
rect 46860 7993 46888 8366
rect 46846 7984 46902 7993
rect 46846 7919 46902 7928
rect 46952 7886 46980 10474
rect 49160 10130 49188 10775
rect 49252 10742 49280 11183
rect 49240 10736 49292 10742
rect 49240 10678 49292 10684
rect 49330 10432 49386 10441
rect 49330 10367 49386 10376
rect 49148 10124 49200 10130
rect 49148 10066 49200 10072
rect 49238 10024 49294 10033
rect 47308 9988 47360 9994
rect 49238 9959 49294 9968
rect 47308 9930 47360 9936
rect 47032 9716 47084 9722
rect 47032 9658 47084 9664
rect 46940 7880 46992 7886
rect 46940 7822 46992 7828
rect 46940 7540 46992 7546
rect 46940 7482 46992 7488
rect 45836 7200 45888 7206
rect 45836 7142 45888 7148
rect 43640 6886 43760 6914
rect 40224 6384 40276 6390
rect 40224 6326 40276 6332
rect 42950 6012 43258 6021
rect 42950 6010 42956 6012
rect 43012 6010 43036 6012
rect 43092 6010 43116 6012
rect 43172 6010 43196 6012
rect 43252 6010 43258 6012
rect 43012 5958 43014 6010
rect 43194 5958 43196 6010
rect 42950 5956 42956 5958
rect 43012 5956 43036 5958
rect 43092 5956 43116 5958
rect 43172 5956 43196 5958
rect 43252 5956 43258 5958
rect 42950 5947 43258 5956
rect 43732 5710 43760 6886
rect 43720 5704 43772 5710
rect 43720 5646 43772 5652
rect 45744 5636 45796 5642
rect 45744 5578 45796 5584
rect 40408 5092 40460 5098
rect 40408 5034 40460 5040
rect 40132 4820 40184 4826
rect 40132 4762 40184 4768
rect 37832 4752 37884 4758
rect 37832 4694 37884 4700
rect 39764 4548 39816 4554
rect 39764 4490 39816 4496
rect 37372 4480 37424 4486
rect 37372 4422 37424 4428
rect 37384 4282 37412 4422
rect 37950 4380 38258 4389
rect 37950 4378 37956 4380
rect 38012 4378 38036 4380
rect 38092 4378 38116 4380
rect 38172 4378 38196 4380
rect 38252 4378 38258 4380
rect 38012 4326 38014 4378
rect 38194 4326 38196 4378
rect 37950 4324 37956 4326
rect 38012 4324 38036 4326
rect 38092 4324 38116 4326
rect 38172 4324 38196 4326
rect 38252 4324 38258 4326
rect 37950 4315 38258 4324
rect 37372 4276 37424 4282
rect 37372 4218 37424 4224
rect 37280 4140 37332 4146
rect 37280 4082 37332 4088
rect 39212 4140 39264 4146
rect 39212 4082 39264 4088
rect 36452 3528 36504 3534
rect 36452 3470 36504 3476
rect 37950 3292 38258 3301
rect 37950 3290 37956 3292
rect 38012 3290 38036 3292
rect 38092 3290 38116 3292
rect 38172 3290 38196 3292
rect 38252 3290 38258 3292
rect 38012 3238 38014 3290
rect 38194 3238 38196 3290
rect 37950 3236 37956 3238
rect 38012 3236 38036 3238
rect 38092 3236 38116 3238
rect 38172 3236 38196 3238
rect 38252 3236 38258 3238
rect 37950 3227 38258 3236
rect 37740 3188 37792 3194
rect 37740 3130 37792 3136
rect 35912 2746 36032 2774
rect 27528 2644 27580 2650
rect 27528 2586 27580 2592
rect 32864 2644 32916 2650
rect 32864 2586 32916 2592
rect 34428 2644 34480 2650
rect 34428 2586 34480 2592
rect 35912 2582 35940 2746
rect 35900 2576 35952 2582
rect 35900 2518 35952 2524
rect 37752 2514 37780 3130
rect 38292 2916 38344 2922
rect 38292 2858 38344 2864
rect 37740 2508 37792 2514
rect 37740 2450 37792 2456
rect 38304 2446 38332 2858
rect 27160 2440 27212 2446
rect 29000 2440 29052 2446
rect 27160 2382 27212 2388
rect 28920 2388 29000 2394
rect 28920 2382 29052 2388
rect 30748 2440 30800 2446
rect 30748 2382 30800 2388
rect 33140 2440 33192 2446
rect 33140 2382 33192 2388
rect 34980 2440 35032 2446
rect 34980 2382 35032 2388
rect 38292 2440 38344 2446
rect 38292 2382 38344 2388
rect 28920 2366 29040 2382
rect 27950 2204 28258 2213
rect 27950 2202 27956 2204
rect 28012 2202 28036 2204
rect 28092 2202 28116 2204
rect 28172 2202 28196 2204
rect 28252 2202 28258 2204
rect 28012 2150 28014 2202
rect 28194 2150 28196 2202
rect 27950 2148 27956 2150
rect 28012 2148 28036 2150
rect 28092 2148 28116 2150
rect 28172 2148 28196 2150
rect 28252 2148 28258 2150
rect 27950 2139 28258 2148
rect 28644 870 28764 898
rect 28644 800 28672 870
rect 18156 734 18460 762
rect 20166 0 20222 800
rect 22282 0 22338 800
rect 24398 0 24454 800
rect 26514 0 26570 800
rect 28630 0 28686 800
rect 28736 762 28764 870
rect 28920 762 28948 2366
rect 30760 800 30788 2382
rect 33152 1578 33180 2382
rect 32876 1550 33180 1578
rect 32876 800 32904 1550
rect 34992 800 35020 2382
rect 37096 2304 37148 2310
rect 37096 2246 37148 2252
rect 37108 800 37136 2246
rect 37950 2204 38258 2213
rect 37950 2202 37956 2204
rect 38012 2202 38036 2204
rect 38092 2202 38116 2204
rect 38172 2202 38196 2204
rect 38252 2202 38258 2204
rect 38012 2150 38014 2202
rect 38194 2150 38196 2202
rect 37950 2148 37956 2150
rect 38012 2148 38036 2150
rect 38092 2148 38116 2150
rect 38172 2148 38196 2150
rect 38252 2148 38258 2150
rect 37950 2139 38258 2148
rect 39224 800 39252 4082
rect 39776 3058 39804 4490
rect 40420 3670 40448 5034
rect 42950 4924 43258 4933
rect 42950 4922 42956 4924
rect 43012 4922 43036 4924
rect 43092 4922 43116 4924
rect 43172 4922 43196 4924
rect 43252 4922 43258 4924
rect 43012 4870 43014 4922
rect 43194 4870 43196 4922
rect 42950 4868 42956 4870
rect 43012 4868 43036 4870
rect 43092 4868 43116 4870
rect 43172 4868 43196 4870
rect 43252 4868 43258 4870
rect 42950 4859 43258 4868
rect 45652 4276 45704 4282
rect 45652 4218 45704 4224
rect 42950 3836 43258 3845
rect 42950 3834 42956 3836
rect 43012 3834 43036 3836
rect 43092 3834 43116 3836
rect 43172 3834 43196 3836
rect 43252 3834 43258 3836
rect 43012 3782 43014 3834
rect 43194 3782 43196 3834
rect 42950 3780 42956 3782
rect 43012 3780 43036 3782
rect 43092 3780 43116 3782
rect 43172 3780 43196 3782
rect 43252 3780 43258 3782
rect 42950 3771 43258 3780
rect 40408 3664 40460 3670
rect 40408 3606 40460 3612
rect 45560 3528 45612 3534
rect 45560 3470 45612 3476
rect 39764 3052 39816 3058
rect 39764 2994 39816 3000
rect 42950 2748 43258 2757
rect 42950 2746 42956 2748
rect 43012 2746 43036 2748
rect 43092 2746 43116 2748
rect 43172 2746 43196 2748
rect 43252 2746 43258 2748
rect 43012 2694 43014 2746
rect 43194 2694 43196 2746
rect 42950 2692 42956 2694
rect 43012 2692 43036 2694
rect 43092 2692 43116 2694
rect 43172 2692 43196 2694
rect 43252 2692 43258 2694
rect 42950 2683 43258 2692
rect 41328 2508 41380 2514
rect 41328 2450 41380 2456
rect 41340 800 41368 2450
rect 43444 2304 43496 2310
rect 43444 2246 43496 2252
rect 43456 800 43484 2246
rect 45572 800 45600 3470
rect 45664 2446 45692 4218
rect 45756 3058 45784 5578
rect 45848 5234 45876 7142
rect 45836 5228 45888 5234
rect 45836 5170 45888 5176
rect 46952 4622 46980 7482
rect 47044 7410 47072 9658
rect 47320 9625 47348 9930
rect 47950 9820 48258 9829
rect 47950 9818 47956 9820
rect 48012 9818 48036 9820
rect 48092 9818 48116 9820
rect 48172 9818 48196 9820
rect 48252 9818 48258 9820
rect 48012 9766 48014 9818
rect 48194 9766 48196 9818
rect 47950 9764 47956 9766
rect 48012 9764 48036 9766
rect 48092 9764 48116 9766
rect 48172 9764 48196 9766
rect 48252 9764 48258 9766
rect 47950 9755 48258 9764
rect 47306 9616 47362 9625
rect 47306 9551 47362 9560
rect 49146 9208 49202 9217
rect 49146 9143 49202 9152
rect 47492 8900 47544 8906
rect 47492 8842 47544 8848
rect 47032 7404 47084 7410
rect 47032 7346 47084 7352
rect 47032 6928 47084 6934
rect 47032 6870 47084 6876
rect 46940 4616 46992 4622
rect 46940 4558 46992 4564
rect 47044 4146 47072 6870
rect 47504 6322 47532 8842
rect 47950 8732 48258 8741
rect 47950 8730 47956 8732
rect 48012 8730 48036 8732
rect 48092 8730 48116 8732
rect 48172 8730 48196 8732
rect 48252 8730 48258 8732
rect 48012 8678 48014 8730
rect 48194 8678 48196 8730
rect 47950 8676 47956 8678
rect 48012 8676 48036 8678
rect 48092 8676 48116 8678
rect 48172 8676 48196 8678
rect 48252 8676 48258 8678
rect 47950 8667 48258 8676
rect 47676 8628 47728 8634
rect 47676 8570 47728 8576
rect 47492 6316 47544 6322
rect 47492 6258 47544 6264
rect 47124 6180 47176 6186
rect 47124 6122 47176 6128
rect 45836 4140 45888 4146
rect 45836 4082 45888 4088
rect 47032 4140 47084 4146
rect 47032 4082 47084 4088
rect 45848 3602 45876 4082
rect 46664 4072 46716 4078
rect 46664 4014 46716 4020
rect 45836 3596 45888 3602
rect 45836 3538 45888 3544
rect 45744 3052 45796 3058
rect 45744 2994 45796 3000
rect 45652 2440 45704 2446
rect 45652 2382 45704 2388
rect 46676 1465 46704 4014
rect 47136 3534 47164 6122
rect 47308 5908 47360 5914
rect 47308 5850 47360 5856
rect 47216 4752 47268 4758
rect 47216 4694 47268 4700
rect 47124 3528 47176 3534
rect 47124 3470 47176 3476
rect 46756 2984 46808 2990
rect 46756 2926 46808 2932
rect 46848 2984 46900 2990
rect 46848 2926 46900 2932
rect 46768 1873 46796 2926
rect 46860 2689 46888 2926
rect 46846 2680 46902 2689
rect 46846 2615 46902 2624
rect 47228 2446 47256 4694
rect 47320 3058 47348 5850
rect 47688 5710 47716 8570
rect 49160 8566 49188 9143
rect 49252 9042 49280 9959
rect 49344 9654 49372 10367
rect 49332 9648 49384 9654
rect 49332 9590 49384 9596
rect 49240 9036 49292 9042
rect 49240 8978 49292 8984
rect 49238 8800 49294 8809
rect 49238 8735 49294 8744
rect 49148 8560 49200 8566
rect 49148 8502 49200 8508
rect 47860 8356 47912 8362
rect 47860 8298 47912 8304
rect 47768 7268 47820 7274
rect 47768 7210 47820 7216
rect 47676 5704 47728 5710
rect 47676 5646 47728 5652
rect 47780 5234 47808 7210
rect 47872 6798 47900 8298
rect 49252 7954 49280 8735
rect 49330 8392 49386 8401
rect 49330 8327 49386 8336
rect 49240 7948 49292 7954
rect 49240 7890 49292 7896
rect 47950 7644 48258 7653
rect 47950 7642 47956 7644
rect 48012 7642 48036 7644
rect 48092 7642 48116 7644
rect 48172 7642 48196 7644
rect 48252 7642 48258 7644
rect 48012 7590 48014 7642
rect 48194 7590 48196 7642
rect 47950 7588 47956 7590
rect 48012 7588 48036 7590
rect 48092 7588 48116 7590
rect 48172 7588 48196 7590
rect 48252 7588 48258 7590
rect 47950 7579 48258 7588
rect 49146 7576 49202 7585
rect 49146 7511 49202 7520
rect 49160 6866 49188 7511
rect 49344 7478 49372 8327
rect 49332 7472 49384 7478
rect 49332 7414 49384 7420
rect 49238 7168 49294 7177
rect 49238 7103 49294 7112
rect 49148 6860 49200 6866
rect 49148 6802 49200 6808
rect 47860 6792 47912 6798
rect 47860 6734 47912 6740
rect 48872 6724 48924 6730
rect 48872 6666 48924 6672
rect 47950 6556 48258 6565
rect 47950 6554 47956 6556
rect 48012 6554 48036 6556
rect 48092 6554 48116 6556
rect 48172 6554 48196 6556
rect 48252 6554 48258 6556
rect 48012 6502 48014 6554
rect 48194 6502 48196 6554
rect 47950 6500 47956 6502
rect 48012 6500 48036 6502
rect 48092 6500 48116 6502
rect 48172 6500 48196 6502
rect 48252 6500 48258 6502
rect 47950 6491 48258 6500
rect 48884 6361 48912 6666
rect 49252 6390 49280 7103
rect 49422 6760 49478 6769
rect 49422 6695 49478 6704
rect 49240 6384 49292 6390
rect 48870 6352 48926 6361
rect 49240 6326 49292 6332
rect 48870 6287 48926 6296
rect 49146 5944 49202 5953
rect 49146 5879 49202 5888
rect 47950 5468 48258 5477
rect 47950 5466 47956 5468
rect 48012 5466 48036 5468
rect 48092 5466 48116 5468
rect 48172 5466 48196 5468
rect 48252 5466 48258 5468
rect 48012 5414 48014 5466
rect 48194 5414 48196 5466
rect 47950 5412 47956 5414
rect 48012 5412 48036 5414
rect 48092 5412 48116 5414
rect 48172 5412 48196 5414
rect 48252 5412 48258 5414
rect 47950 5403 48258 5412
rect 49160 5302 49188 5879
rect 49436 5778 49464 6695
rect 49424 5772 49476 5778
rect 49424 5714 49476 5720
rect 49422 5536 49478 5545
rect 49422 5471 49478 5480
rect 49148 5296 49200 5302
rect 49148 5238 49200 5244
rect 47768 5228 47820 5234
rect 47768 5170 47820 5176
rect 48320 5160 48372 5166
rect 48320 5102 48372 5108
rect 49330 5128 49386 5137
rect 48332 4729 48360 5102
rect 49330 5063 49386 5072
rect 48318 4720 48374 4729
rect 48318 4655 48374 4664
rect 47676 4548 47728 4554
rect 47676 4490 47728 4496
rect 47688 3942 47716 4490
rect 47950 4380 48258 4389
rect 47950 4378 47956 4380
rect 48012 4378 48036 4380
rect 48092 4378 48116 4380
rect 48172 4378 48196 4380
rect 48252 4378 48258 4380
rect 48012 4326 48014 4378
rect 48194 4326 48196 4378
rect 47950 4324 47956 4326
rect 48012 4324 48036 4326
rect 48092 4324 48116 4326
rect 48172 4324 48196 4326
rect 48252 4324 48258 4326
rect 47950 4315 48258 4324
rect 49146 4312 49202 4321
rect 49146 4247 49202 4256
rect 47676 3936 47728 3942
rect 47676 3878 47728 3884
rect 47308 3052 47360 3058
rect 47308 2994 47360 3000
rect 47216 2440 47268 2446
rect 47216 2382 47268 2388
rect 46754 1864 46810 1873
rect 46754 1799 46810 1808
rect 46662 1456 46718 1465
rect 46662 1391 46718 1400
rect 47688 800 47716 3878
rect 49160 3602 49188 4247
rect 49344 4146 49372 5063
rect 49436 4690 49464 5471
rect 49424 4684 49476 4690
rect 49424 4626 49476 4632
rect 49792 4480 49844 4486
rect 49792 4422 49844 4428
rect 49332 4140 49384 4146
rect 49332 4082 49384 4088
rect 49238 3904 49294 3913
rect 49238 3839 49294 3848
rect 49148 3596 49200 3602
rect 49148 3538 49200 3544
rect 49146 3496 49202 3505
rect 48688 3460 48740 3466
rect 49146 3431 49202 3440
rect 48688 3402 48740 3408
rect 47950 3292 48258 3301
rect 47950 3290 47956 3292
rect 48012 3290 48036 3292
rect 48092 3290 48116 3292
rect 48172 3290 48196 3292
rect 48252 3290 48258 3292
rect 48012 3238 48014 3290
rect 48194 3238 48196 3290
rect 47950 3236 47956 3238
rect 48012 3236 48036 3238
rect 48092 3236 48116 3238
rect 48172 3236 48196 3238
rect 48252 3236 48258 3238
rect 47950 3227 48258 3236
rect 48700 3097 48728 3402
rect 48686 3088 48742 3097
rect 48686 3023 48742 3032
rect 49160 2514 49188 3431
rect 49252 3126 49280 3839
rect 49240 3120 49292 3126
rect 49240 3062 49292 3068
rect 49148 2508 49200 2514
rect 49148 2450 49200 2456
rect 48504 2372 48556 2378
rect 48504 2314 48556 2320
rect 48516 2281 48544 2314
rect 48502 2272 48558 2281
rect 47950 2204 48258 2213
rect 48502 2207 48558 2216
rect 47950 2202 47956 2204
rect 48012 2202 48036 2204
rect 48092 2202 48116 2204
rect 48172 2202 48196 2204
rect 48252 2202 48258 2204
rect 48012 2150 48014 2202
rect 48194 2150 48196 2202
rect 47950 2148 47956 2150
rect 48012 2148 48036 2150
rect 48092 2148 48116 2150
rect 48172 2148 48196 2150
rect 48252 2148 48258 2150
rect 47950 2139 48258 2148
rect 49804 800 49832 4422
rect 28736 734 28948 762
rect 30746 0 30802 800
rect 32862 0 32918 800
rect 34978 0 35034 800
rect 37094 0 37150 800
rect 39210 0 39266 800
rect 41326 0 41382 800
rect 43442 0 43498 800
rect 45558 0 45614 800
rect 47674 0 47730 800
rect 49790 0 49846 800
<< via2 >>
rect 2778 24404 2834 24440
rect 2778 24384 2780 24404
rect 2780 24384 2832 24404
rect 2832 24384 2834 24404
rect 1306 20712 1362 20768
rect 3422 25608 3478 25664
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 4066 25200 4122 25256
rect 3882 24792 3938 24848
rect 3790 23976 3846 24032
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 2686 21528 2742 21584
rect 2778 21120 2834 21176
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 2686 19488 2742 19544
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 3330 19896 3386 19952
rect 2778 18808 2834 18864
rect 1950 18672 2006 18728
rect 2962 19216 3018 19272
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 2870 18264 2926 18320
rect 4066 23588 4122 23624
rect 4066 23568 4068 23588
rect 4068 23568 4120 23588
rect 4120 23568 4122 23588
rect 4066 23160 4122 23216
rect 3974 22752 4030 22808
rect 4066 22480 4122 22536
rect 3882 21936 3938 21992
rect 3882 20340 3884 20360
rect 3884 20340 3936 20360
rect 3936 20340 3938 20360
rect 3882 20304 3938 20340
rect 2686 17856 2742 17912
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 2778 17448 2834 17504
rect 1214 17040 1270 17096
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 1306 16632 1362 16688
rect 1306 16224 1362 16280
rect 5906 21392 5962 21448
rect 7378 24248 7434 24304
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 1306 15816 1362 15872
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 1306 15408 1362 15464
rect 1306 15000 1362 15056
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 1306 14592 1362 14648
rect 1306 14184 1362 14240
rect 2778 13776 2834 13832
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 3514 13368 3570 13424
rect 1306 12960 1362 13016
rect 1214 12552 1270 12608
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 1214 12144 1270 12200
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 8758 21392 8814 21448
rect 11334 21392 11390 21448
rect 11334 20984 11390 21040
rect 10966 19760 11022 19816
rect 9770 16496 9826 16552
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 10506 16632 10562 16688
rect 10690 17176 10746 17232
rect 11150 18128 11206 18184
rect 10506 15272 10562 15328
rect 10322 14456 10378 14512
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 1306 11736 1362 11792
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 1306 11328 1362 11384
rect 1766 11056 1822 11112
rect 1582 10920 1638 10976
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 1306 10512 1362 10568
rect 1214 10104 1270 10160
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 1306 9716 1362 9752
rect 1306 9696 1308 9716
rect 1308 9696 1360 9716
rect 1360 9696 1362 9716
rect 1766 9444 1822 9480
rect 1766 9424 1768 9444
rect 1768 9424 1820 9444
rect 1820 9424 1822 9444
rect 1306 9288 1362 9344
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 1306 8900 1362 8936
rect 1306 8880 1308 8900
rect 1308 8880 1360 8900
rect 1360 8880 1362 8900
rect 1214 8472 1270 8528
rect 1398 8084 1454 8120
rect 1398 8064 1400 8084
rect 1400 8064 1452 8084
rect 1452 8064 1454 8084
rect 1306 7656 1362 7712
rect 1306 7248 1362 7304
rect 1214 6840 1270 6896
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 12070 18808 12126 18864
rect 11794 17040 11850 17096
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 13358 19896 13414 19952
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 13634 19760 13690 19816
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 11886 15952 11942 16008
rect 11518 13812 11520 13832
rect 11520 13812 11572 13832
rect 11572 13812 11574 13832
rect 11518 13776 11574 13812
rect 12438 15408 12494 15464
rect 12438 15272 12494 15328
rect 12346 14900 12348 14920
rect 12348 14900 12400 14920
rect 12400 14900 12402 14920
rect 12346 14864 12402 14900
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 14094 19352 14150 19408
rect 14462 22516 14464 22536
rect 14464 22516 14516 22536
rect 14516 22516 14518 22536
rect 14462 22480 14518 22516
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 1306 6432 1362 6488
rect 1306 6024 1362 6080
rect 1306 5652 1308 5672
rect 1308 5652 1360 5672
rect 1360 5652 1362 5672
rect 1306 5616 1362 5652
rect 1306 4820 1362 4856
rect 1306 4800 1308 4820
rect 1308 4800 1360 4820
rect 1360 4800 1362 4820
rect 1306 4392 1362 4448
rect 1398 3984 1454 4040
rect 1306 3576 1362 3632
rect 1122 3440 1178 3496
rect 1306 3188 1362 3224
rect 1306 3168 1308 3188
rect 1308 3168 1360 3188
rect 1360 3168 1362 3188
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 2778 5208 2834 5264
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 5354 3984 5410 4040
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 1306 2760 1362 2816
rect 1306 2388 1308 2408
rect 1308 2388 1360 2408
rect 1360 2388 1362 2408
rect 1306 2352 1362 2388
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 1214 1944 1270 2000
rect 1306 1536 1362 1592
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 13358 11464 13414 11520
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 14278 17312 14334 17368
rect 14278 16088 14334 16144
rect 14554 16496 14610 16552
rect 14370 15000 14426 15056
rect 15106 19352 15162 19408
rect 15014 18264 15070 18320
rect 14922 18128 14978 18184
rect 14646 15544 14702 15600
rect 14186 14356 14188 14376
rect 14188 14356 14240 14376
rect 14240 14356 14242 14376
rect 14186 14320 14242 14356
rect 14554 13640 14610 13696
rect 14278 13504 14334 13560
rect 13542 11328 13598 11384
rect 13634 10668 13690 10704
rect 13634 10648 13636 10668
rect 13636 10648 13688 10668
rect 13688 10648 13690 10668
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 13082 10104 13138 10160
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 14370 11464 14426 11520
rect 16210 21936 16266 21992
rect 15382 19372 15438 19408
rect 15382 19352 15384 19372
rect 15384 19352 15436 19372
rect 15436 19352 15438 19372
rect 15382 18148 15438 18184
rect 15382 18128 15384 18148
rect 15384 18128 15436 18148
rect 15436 18128 15438 18148
rect 15382 17312 15438 17368
rect 14830 15988 14832 16008
rect 14832 15988 14884 16008
rect 14884 15988 14886 16008
rect 14830 15952 14886 15988
rect 15014 15000 15070 15056
rect 15658 16496 15714 16552
rect 15014 11736 15070 11792
rect 14738 11092 14740 11112
rect 14740 11092 14792 11112
rect 14792 11092 14794 11112
rect 14738 11056 14794 11092
rect 14186 9016 14242 9072
rect 15566 15408 15622 15464
rect 16670 21528 16726 21584
rect 16578 21140 16634 21176
rect 16578 21120 16580 21140
rect 16580 21120 16632 21140
rect 16632 21120 16634 21140
rect 17130 21120 17186 21176
rect 16762 20340 16764 20360
rect 16764 20340 16816 20360
rect 16816 20340 16818 20360
rect 16762 20304 16818 20340
rect 16210 18672 16266 18728
rect 15934 16632 15990 16688
rect 16118 16652 16174 16688
rect 16118 16632 16120 16652
rect 16120 16632 16172 16652
rect 16172 16632 16174 16652
rect 15842 15988 15844 16008
rect 15844 15988 15896 16008
rect 15896 15988 15898 16008
rect 15842 15952 15898 15988
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 18418 22072 18474 22128
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 17406 18708 17408 18728
rect 17408 18708 17460 18728
rect 17460 18708 17462 18728
rect 17406 18672 17462 18708
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 18694 22072 18750 22128
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 19338 23976 19394 24032
rect 18878 21936 18934 21992
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 17498 16940 17500 16960
rect 17500 16940 17552 16960
rect 17552 16940 17554 16960
rect 15198 11600 15254 11656
rect 16578 15000 16634 15056
rect 16486 13812 16488 13832
rect 16488 13812 16540 13832
rect 16540 13812 16542 13832
rect 16486 13776 16542 13812
rect 16210 12844 16266 12880
rect 16210 12824 16212 12844
rect 16212 12824 16264 12844
rect 16264 12824 16266 12844
rect 16210 12688 16266 12744
rect 15658 11600 15714 11656
rect 16118 11736 16174 11792
rect 16486 12144 16542 12200
rect 16946 15816 17002 15872
rect 17314 15564 17370 15600
rect 17314 15544 17316 15564
rect 17316 15544 17368 15564
rect 17368 15544 17370 15564
rect 17498 16904 17554 16940
rect 17590 15000 17646 15056
rect 16946 13504 17002 13560
rect 16670 11348 16726 11384
rect 16670 11328 16672 11348
rect 16672 11328 16724 11348
rect 16724 11328 16726 11348
rect 16578 9968 16634 10024
rect 16854 11056 16910 11112
rect 17130 12280 17186 12336
rect 17314 12144 17370 12200
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18510 13776 18566 13832
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18234 11500 18236 11520
rect 18236 11500 18288 11520
rect 18288 11500 18290 11520
rect 17682 11192 17738 11248
rect 18234 11464 18290 11500
rect 18418 11192 18474 11248
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 19338 21664 19394 21720
rect 19246 20984 19302 21040
rect 21178 22072 21234 22128
rect 21270 21800 21326 21856
rect 19706 20848 19762 20904
rect 19982 20576 20038 20632
rect 19338 19624 19394 19680
rect 19430 18808 19486 18864
rect 18878 18692 18934 18728
rect 18878 18672 18880 18692
rect 18880 18672 18932 18692
rect 18932 18672 18934 18692
rect 19062 18264 19118 18320
rect 19338 18400 19394 18456
rect 19798 18672 19854 18728
rect 19062 13776 19118 13832
rect 21086 20984 21142 21040
rect 20350 19488 20406 19544
rect 19706 16632 19762 16688
rect 19246 13232 19302 13288
rect 18602 11056 18658 11112
rect 19798 16088 19854 16144
rect 21638 22072 21694 22128
rect 21546 20984 21602 21040
rect 21270 18536 21326 18592
rect 19982 14184 20038 14240
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 20534 15136 20590 15192
rect 21178 16904 21234 16960
rect 20994 16496 21050 16552
rect 20074 12688 20130 12744
rect 19890 11772 19892 11792
rect 19892 11772 19944 11792
rect 19944 11772 19946 11792
rect 19890 11736 19946 11772
rect 21914 20576 21970 20632
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 22742 21936 22798 21992
rect 23202 21800 23258 21856
rect 22834 21528 22890 21584
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 21822 19896 21878 19952
rect 21638 17720 21694 17776
rect 23478 21120 23534 21176
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 23386 20032 23442 20088
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 22466 16496 22522 16552
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 24030 22480 24086 22536
rect 24674 23432 24730 23488
rect 24674 23044 24730 23080
rect 24674 23024 24676 23044
rect 24676 23024 24728 23044
rect 24728 23024 24730 23044
rect 24858 20984 24914 21040
rect 24122 20168 24178 20224
rect 23570 16632 23626 16688
rect 21638 15000 21694 15056
rect 21822 14456 21878 14512
rect 21730 14320 21786 14376
rect 20810 11076 20866 11112
rect 20810 11056 20812 11076
rect 20812 11056 20864 11076
rect 20864 11056 20866 11076
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 21638 12688 21694 12744
rect 21270 9968 21326 10024
rect 22650 12960 22706 13016
rect 23294 16088 23350 16144
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 22098 12144 22154 12200
rect 22650 12416 22706 12472
rect 23110 12980 23166 13016
rect 23110 12960 23112 12980
rect 23112 12960 23164 12980
rect 23164 12960 23166 12980
rect 23018 12688 23074 12744
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 22558 12144 22614 12200
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 22006 11056 22062 11112
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 22466 9968 22522 10024
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 23846 11056 23902 11112
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 24122 11056 24178 11112
rect 25134 22092 25190 22128
rect 25134 22072 25136 22092
rect 25136 22072 25188 22092
rect 25188 22072 25190 22092
rect 25226 21428 25228 21448
rect 25228 21428 25280 21448
rect 25280 21428 25282 21448
rect 25226 21392 25282 21428
rect 25318 20576 25374 20632
rect 25962 24248 26018 24304
rect 26146 24112 26202 24168
rect 25594 22480 25650 22536
rect 25318 19488 25374 19544
rect 25042 18692 25098 18728
rect 25042 18672 25044 18692
rect 25044 18672 25096 18692
rect 25096 18672 25098 18692
rect 25134 18284 25190 18320
rect 25134 18264 25136 18284
rect 25136 18264 25188 18284
rect 25188 18264 25190 18284
rect 25042 18128 25098 18184
rect 25410 17176 25466 17232
rect 24398 14320 24454 14376
rect 24582 14220 24584 14240
rect 24584 14220 24636 14240
rect 24636 14220 24638 14240
rect 24582 14184 24638 14220
rect 26330 23432 26386 23488
rect 27342 24012 27344 24032
rect 27344 24012 27396 24032
rect 27396 24012 27398 24032
rect 27342 23976 27398 24012
rect 27956 23962 28012 23964
rect 28036 23962 28092 23964
rect 28116 23962 28172 23964
rect 28196 23962 28252 23964
rect 27956 23910 28002 23962
rect 28002 23910 28012 23962
rect 28036 23910 28066 23962
rect 28066 23910 28078 23962
rect 28078 23910 28092 23962
rect 28116 23910 28130 23962
rect 28130 23910 28142 23962
rect 28142 23910 28172 23962
rect 28196 23910 28206 23962
rect 28206 23910 28252 23962
rect 27956 23908 28012 23910
rect 28036 23908 28092 23910
rect 28116 23908 28172 23910
rect 28196 23908 28252 23910
rect 25778 21956 25834 21992
rect 25778 21936 25780 21956
rect 25780 21936 25832 21956
rect 25832 21936 25834 21956
rect 25870 19896 25926 19952
rect 26146 21392 26202 21448
rect 26054 19760 26110 19816
rect 26146 19488 26202 19544
rect 26054 19080 26110 19136
rect 25870 18808 25926 18864
rect 25962 18264 26018 18320
rect 25594 16088 25650 16144
rect 24490 12824 24546 12880
rect 25410 11736 25466 11792
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 26698 21140 26754 21176
rect 26698 21120 26700 21140
rect 26700 21120 26752 21140
rect 26752 21120 26754 21140
rect 26882 20984 26938 21040
rect 26606 19352 26662 19408
rect 26422 18536 26478 18592
rect 26330 18128 26386 18184
rect 26514 17584 26570 17640
rect 26790 19624 26846 19680
rect 26698 17040 26754 17096
rect 27250 22092 27306 22128
rect 27250 22072 27252 22092
rect 27252 22072 27304 22092
rect 27304 22072 27306 22092
rect 27956 22874 28012 22876
rect 28036 22874 28092 22876
rect 28116 22874 28172 22876
rect 28196 22874 28252 22876
rect 27956 22822 28002 22874
rect 28002 22822 28012 22874
rect 28036 22822 28066 22874
rect 28066 22822 28078 22874
rect 28078 22822 28092 22874
rect 28116 22822 28130 22874
rect 28130 22822 28142 22874
rect 28142 22822 28172 22874
rect 28196 22822 28206 22874
rect 28206 22822 28252 22874
rect 27956 22820 28012 22822
rect 28036 22820 28092 22822
rect 28116 22820 28172 22822
rect 28196 22820 28252 22822
rect 27956 21786 28012 21788
rect 28036 21786 28092 21788
rect 28116 21786 28172 21788
rect 28196 21786 28252 21788
rect 27956 21734 28002 21786
rect 28002 21734 28012 21786
rect 28036 21734 28066 21786
rect 28066 21734 28078 21786
rect 28078 21734 28092 21786
rect 28116 21734 28130 21786
rect 28130 21734 28142 21786
rect 28142 21734 28172 21786
rect 28196 21734 28206 21786
rect 28206 21734 28252 21786
rect 27956 21732 28012 21734
rect 28036 21732 28092 21734
rect 28116 21732 28172 21734
rect 28196 21732 28252 21734
rect 27434 21392 27490 21448
rect 27342 21120 27398 21176
rect 26974 18672 27030 18728
rect 27066 18400 27122 18456
rect 27250 18164 27252 18184
rect 27252 18164 27304 18184
rect 27304 18164 27306 18184
rect 27250 18128 27306 18164
rect 27066 17992 27122 18048
rect 27066 16904 27122 16960
rect 26146 15816 26202 15872
rect 26330 14864 26386 14920
rect 25870 12708 25926 12744
rect 25870 12688 25872 12708
rect 25872 12688 25924 12708
rect 25924 12688 25926 12708
rect 25594 9016 25650 9072
rect 26238 12960 26294 13016
rect 27250 16632 27306 16688
rect 27710 19624 27766 19680
rect 27618 17856 27674 17912
rect 28814 21548 28870 21584
rect 28814 21528 28816 21548
rect 28816 21528 28868 21548
rect 28868 21528 28870 21548
rect 28446 20712 28502 20768
rect 28722 20748 28724 20768
rect 28724 20748 28776 20768
rect 28776 20748 28778 20768
rect 27956 20698 28012 20700
rect 28036 20698 28092 20700
rect 28116 20698 28172 20700
rect 28196 20698 28252 20700
rect 27956 20646 28002 20698
rect 28002 20646 28012 20698
rect 28036 20646 28066 20698
rect 28066 20646 28078 20698
rect 28078 20646 28092 20698
rect 28116 20646 28130 20698
rect 28130 20646 28142 20698
rect 28142 20646 28172 20698
rect 28196 20646 28206 20698
rect 28206 20646 28252 20698
rect 27956 20644 28012 20646
rect 28036 20644 28092 20646
rect 28116 20644 28172 20646
rect 28196 20644 28252 20646
rect 27956 19610 28012 19612
rect 28036 19610 28092 19612
rect 28116 19610 28172 19612
rect 28196 19610 28252 19612
rect 27956 19558 28002 19610
rect 28002 19558 28012 19610
rect 28036 19558 28066 19610
rect 28066 19558 28078 19610
rect 28078 19558 28092 19610
rect 28116 19558 28130 19610
rect 28130 19558 28142 19610
rect 28142 19558 28172 19610
rect 28196 19558 28206 19610
rect 28206 19558 28252 19610
rect 27956 19556 28012 19558
rect 28036 19556 28092 19558
rect 28116 19556 28172 19558
rect 28196 19556 28252 19558
rect 28722 20712 28778 20748
rect 28814 20168 28870 20224
rect 28538 19624 28594 19680
rect 28814 19488 28870 19544
rect 27956 18522 28012 18524
rect 28036 18522 28092 18524
rect 28116 18522 28172 18524
rect 28196 18522 28252 18524
rect 27956 18470 28002 18522
rect 28002 18470 28012 18522
rect 28036 18470 28066 18522
rect 28066 18470 28078 18522
rect 28078 18470 28092 18522
rect 28116 18470 28130 18522
rect 28130 18470 28142 18522
rect 28142 18470 28172 18522
rect 28196 18470 28206 18522
rect 28206 18470 28252 18522
rect 27956 18468 28012 18470
rect 28036 18468 28092 18470
rect 28116 18468 28172 18470
rect 28196 18468 28252 18470
rect 27802 17856 27858 17912
rect 27956 17434 28012 17436
rect 28036 17434 28092 17436
rect 28116 17434 28172 17436
rect 28196 17434 28252 17436
rect 27956 17382 28002 17434
rect 28002 17382 28012 17434
rect 28036 17382 28066 17434
rect 28066 17382 28078 17434
rect 28078 17382 28092 17434
rect 28116 17382 28130 17434
rect 28130 17382 28142 17434
rect 28142 17382 28172 17434
rect 28196 17382 28206 17434
rect 28206 17382 28252 17434
rect 27956 17380 28012 17382
rect 28036 17380 28092 17382
rect 28116 17380 28172 17382
rect 28196 17380 28252 17382
rect 28262 17176 28318 17232
rect 27710 16904 27766 16960
rect 27342 15952 27398 16008
rect 26974 15408 27030 15464
rect 27956 16346 28012 16348
rect 28036 16346 28092 16348
rect 28116 16346 28172 16348
rect 28196 16346 28252 16348
rect 27956 16294 28002 16346
rect 28002 16294 28012 16346
rect 28036 16294 28066 16346
rect 28066 16294 28078 16346
rect 28078 16294 28092 16346
rect 28116 16294 28130 16346
rect 28130 16294 28142 16346
rect 28142 16294 28172 16346
rect 28196 16294 28206 16346
rect 28206 16294 28252 16346
rect 27956 16292 28012 16294
rect 28036 16292 28092 16294
rect 28116 16292 28172 16294
rect 28196 16292 28252 16294
rect 27066 15020 27122 15056
rect 27066 15000 27068 15020
rect 27068 15000 27120 15020
rect 27120 15000 27122 15020
rect 26790 10104 26846 10160
rect 26146 9580 26202 9616
rect 26146 9560 26148 9580
rect 26148 9560 26200 9580
rect 26200 9560 26202 9580
rect 25410 4020 25412 4040
rect 25412 4020 25464 4040
rect 25464 4020 25466 4040
rect 25410 3984 25466 4020
rect 27956 15258 28012 15260
rect 28036 15258 28092 15260
rect 28116 15258 28172 15260
rect 28196 15258 28252 15260
rect 27956 15206 28002 15258
rect 28002 15206 28012 15258
rect 28036 15206 28066 15258
rect 28066 15206 28078 15258
rect 28078 15206 28092 15258
rect 28116 15206 28130 15258
rect 28130 15206 28142 15258
rect 28142 15206 28172 15258
rect 28196 15206 28206 15258
rect 28206 15206 28252 15258
rect 27956 15204 28012 15206
rect 28036 15204 28092 15206
rect 28116 15204 28172 15206
rect 28196 15204 28252 15206
rect 27526 15136 27582 15192
rect 28630 19080 28686 19136
rect 28998 18944 29054 19000
rect 28538 17856 28594 17912
rect 28262 14320 28318 14376
rect 28630 16788 28686 16824
rect 28630 16768 28632 16788
rect 28632 16768 28684 16788
rect 28684 16768 28686 16788
rect 27956 14170 28012 14172
rect 28036 14170 28092 14172
rect 28116 14170 28172 14172
rect 28196 14170 28252 14172
rect 27956 14118 28002 14170
rect 28002 14118 28012 14170
rect 28036 14118 28066 14170
rect 28066 14118 28078 14170
rect 28078 14118 28092 14170
rect 28116 14118 28130 14170
rect 28130 14118 28142 14170
rect 28142 14118 28172 14170
rect 28196 14118 28206 14170
rect 28206 14118 28252 14170
rect 27956 14116 28012 14118
rect 28036 14116 28092 14118
rect 28116 14116 28172 14118
rect 28196 14116 28252 14118
rect 27956 13082 28012 13084
rect 28036 13082 28092 13084
rect 28116 13082 28172 13084
rect 28196 13082 28252 13084
rect 27956 13030 28002 13082
rect 28002 13030 28012 13082
rect 28036 13030 28066 13082
rect 28066 13030 28078 13082
rect 28078 13030 28092 13082
rect 28116 13030 28130 13082
rect 28130 13030 28142 13082
rect 28142 13030 28172 13082
rect 28196 13030 28206 13082
rect 28206 13030 28252 13082
rect 27956 13028 28012 13030
rect 28036 13028 28092 13030
rect 28116 13028 28172 13030
rect 28196 13028 28252 13030
rect 27956 11994 28012 11996
rect 28036 11994 28092 11996
rect 28116 11994 28172 11996
rect 28196 11994 28252 11996
rect 27956 11942 28002 11994
rect 28002 11942 28012 11994
rect 28036 11942 28066 11994
rect 28066 11942 28078 11994
rect 28078 11942 28092 11994
rect 28116 11942 28130 11994
rect 28130 11942 28142 11994
rect 28142 11942 28172 11994
rect 28196 11942 28206 11994
rect 28206 11942 28252 11994
rect 27956 11940 28012 11942
rect 28036 11940 28092 11942
rect 28116 11940 28172 11942
rect 28196 11940 28252 11942
rect 27956 10906 28012 10908
rect 28036 10906 28092 10908
rect 28116 10906 28172 10908
rect 28196 10906 28252 10908
rect 27956 10854 28002 10906
rect 28002 10854 28012 10906
rect 28036 10854 28066 10906
rect 28066 10854 28078 10906
rect 28078 10854 28092 10906
rect 28116 10854 28130 10906
rect 28130 10854 28142 10906
rect 28142 10854 28172 10906
rect 28196 10854 28206 10906
rect 28206 10854 28252 10906
rect 27956 10852 28012 10854
rect 28036 10852 28092 10854
rect 28116 10852 28172 10854
rect 28196 10852 28252 10854
rect 27526 10104 27582 10160
rect 27956 9818 28012 9820
rect 28036 9818 28092 9820
rect 28116 9818 28172 9820
rect 28196 9818 28252 9820
rect 27956 9766 28002 9818
rect 28002 9766 28012 9818
rect 28036 9766 28066 9818
rect 28066 9766 28078 9818
rect 28078 9766 28092 9818
rect 28116 9766 28130 9818
rect 28130 9766 28142 9818
rect 28142 9766 28172 9818
rect 28196 9766 28206 9818
rect 28206 9766 28252 9818
rect 27956 9764 28012 9766
rect 28036 9764 28092 9766
rect 28116 9764 28172 9766
rect 28196 9764 28252 9766
rect 27956 8730 28012 8732
rect 28036 8730 28092 8732
rect 28116 8730 28172 8732
rect 28196 8730 28252 8732
rect 27956 8678 28002 8730
rect 28002 8678 28012 8730
rect 28036 8678 28066 8730
rect 28066 8678 28078 8730
rect 28078 8678 28092 8730
rect 28116 8678 28130 8730
rect 28130 8678 28142 8730
rect 28142 8678 28172 8730
rect 28196 8678 28206 8730
rect 28206 8678 28252 8730
rect 27956 8676 28012 8678
rect 28036 8676 28092 8678
rect 28116 8676 28172 8678
rect 28196 8676 28252 8678
rect 27956 7642 28012 7644
rect 28036 7642 28092 7644
rect 28116 7642 28172 7644
rect 28196 7642 28252 7644
rect 27956 7590 28002 7642
rect 28002 7590 28012 7642
rect 28036 7590 28066 7642
rect 28066 7590 28078 7642
rect 28078 7590 28092 7642
rect 28116 7590 28130 7642
rect 28130 7590 28142 7642
rect 28142 7590 28172 7642
rect 28196 7590 28206 7642
rect 28206 7590 28252 7642
rect 27956 7588 28012 7590
rect 28036 7588 28092 7590
rect 28116 7588 28172 7590
rect 28196 7588 28252 7590
rect 27956 6554 28012 6556
rect 28036 6554 28092 6556
rect 28116 6554 28172 6556
rect 28196 6554 28252 6556
rect 27956 6502 28002 6554
rect 28002 6502 28012 6554
rect 28036 6502 28066 6554
rect 28066 6502 28078 6554
rect 28078 6502 28092 6554
rect 28116 6502 28130 6554
rect 28130 6502 28142 6554
rect 28142 6502 28172 6554
rect 28196 6502 28206 6554
rect 28206 6502 28252 6554
rect 27956 6500 28012 6502
rect 28036 6500 28092 6502
rect 28116 6500 28172 6502
rect 28196 6500 28252 6502
rect 28998 18420 29054 18456
rect 28998 18400 29000 18420
rect 29000 18400 29052 18420
rect 29052 18400 29054 18420
rect 28722 14320 28778 14376
rect 29274 19624 29330 19680
rect 29182 19252 29184 19272
rect 29184 19252 29236 19272
rect 29236 19252 29238 19272
rect 29182 19216 29238 19252
rect 30102 24384 30158 24440
rect 30010 24248 30066 24304
rect 30194 23180 30250 23216
rect 30194 23160 30196 23180
rect 30196 23160 30248 23180
rect 30248 23160 30250 23180
rect 30010 22072 30066 22128
rect 29642 21392 29698 21448
rect 29366 18400 29422 18456
rect 29734 20848 29790 20904
rect 29642 18672 29698 18728
rect 29550 18128 29606 18184
rect 28538 11056 28594 11112
rect 29274 16652 29330 16688
rect 29274 16632 29276 16652
rect 29276 16632 29328 16652
rect 29328 16632 29330 16652
rect 30746 22772 30802 22808
rect 30746 22752 30748 22772
rect 30748 22752 30800 22772
rect 30800 22752 30802 22772
rect 30010 20304 30066 20360
rect 30010 18808 30066 18864
rect 29090 10920 29146 10976
rect 28630 9016 28686 9072
rect 29550 15544 29606 15600
rect 29734 14048 29790 14104
rect 29550 12860 29552 12880
rect 29552 12860 29604 12880
rect 29604 12860 29606 12880
rect 29550 12824 29606 12860
rect 30654 21664 30710 21720
rect 30194 20712 30250 20768
rect 30194 18128 30250 18184
rect 30010 16632 30066 16688
rect 30470 18672 30526 18728
rect 30838 21120 30894 21176
rect 30838 20460 30894 20496
rect 30838 20440 30840 20460
rect 30840 20440 30892 20460
rect 30892 20440 30894 20460
rect 31022 23568 31078 23624
rect 31206 21564 31208 21584
rect 31208 21564 31260 21584
rect 31260 21564 31262 21584
rect 31206 21528 31262 21564
rect 30654 18944 30710 19000
rect 30654 17584 30710 17640
rect 30470 15544 30526 15600
rect 27956 5466 28012 5468
rect 28036 5466 28092 5468
rect 28116 5466 28172 5468
rect 28196 5466 28252 5468
rect 27956 5414 28002 5466
rect 28002 5414 28012 5466
rect 28036 5414 28066 5466
rect 28066 5414 28078 5466
rect 28078 5414 28092 5466
rect 28116 5414 28130 5466
rect 28130 5414 28142 5466
rect 28142 5414 28172 5466
rect 28196 5414 28206 5466
rect 28206 5414 28252 5466
rect 27956 5412 28012 5414
rect 28036 5412 28092 5414
rect 28116 5412 28172 5414
rect 28196 5412 28252 5414
rect 27956 4378 28012 4380
rect 28036 4378 28092 4380
rect 28116 4378 28172 4380
rect 28196 4378 28252 4380
rect 27956 4326 28002 4378
rect 28002 4326 28012 4378
rect 28036 4326 28066 4378
rect 28066 4326 28078 4378
rect 28078 4326 28092 4378
rect 28116 4326 28130 4378
rect 28130 4326 28142 4378
rect 28142 4326 28172 4378
rect 28196 4326 28206 4378
rect 28206 4326 28252 4378
rect 27956 4324 28012 4326
rect 28036 4324 28092 4326
rect 28116 4324 28172 4326
rect 28196 4324 28252 4326
rect 26054 3440 26110 3496
rect 27956 3290 28012 3292
rect 28036 3290 28092 3292
rect 28116 3290 28172 3292
rect 28196 3290 28252 3292
rect 27956 3238 28002 3290
rect 28002 3238 28012 3290
rect 28036 3238 28066 3290
rect 28066 3238 28078 3290
rect 28078 3238 28092 3290
rect 28116 3238 28130 3290
rect 28130 3238 28142 3290
rect 28142 3238 28172 3290
rect 28196 3238 28206 3290
rect 28206 3238 28252 3290
rect 27956 3236 28012 3238
rect 28036 3236 28092 3238
rect 28116 3236 28172 3238
rect 28196 3236 28252 3238
rect 30194 11076 30250 11112
rect 30194 11056 30196 11076
rect 30196 11056 30248 11076
rect 30248 11056 30250 11076
rect 30378 12144 30434 12200
rect 32402 24404 32458 24440
rect 32402 24384 32404 24404
rect 32404 24384 32456 24404
rect 32456 24384 32458 24404
rect 31482 23024 31538 23080
rect 31482 22616 31538 22672
rect 31390 22072 31446 22128
rect 32956 24506 33012 24508
rect 33036 24506 33092 24508
rect 33116 24506 33172 24508
rect 33196 24506 33252 24508
rect 32956 24454 33002 24506
rect 33002 24454 33012 24506
rect 33036 24454 33066 24506
rect 33066 24454 33078 24506
rect 33078 24454 33092 24506
rect 33116 24454 33130 24506
rect 33130 24454 33142 24506
rect 33142 24454 33172 24506
rect 33196 24454 33206 24506
rect 33206 24454 33252 24506
rect 32956 24452 33012 24454
rect 33036 24452 33092 24454
rect 33116 24452 33172 24454
rect 33196 24452 33252 24454
rect 32586 22888 32642 22944
rect 32956 23418 33012 23420
rect 33036 23418 33092 23420
rect 33116 23418 33172 23420
rect 33196 23418 33252 23420
rect 32956 23366 33002 23418
rect 33002 23366 33012 23418
rect 33036 23366 33066 23418
rect 33066 23366 33078 23418
rect 33078 23366 33092 23418
rect 33116 23366 33130 23418
rect 33130 23366 33142 23418
rect 33142 23366 33172 23418
rect 33196 23366 33206 23418
rect 33206 23366 33252 23418
rect 32956 23364 33012 23366
rect 33036 23364 33092 23366
rect 33116 23364 33172 23366
rect 33196 23364 33252 23366
rect 32956 22330 33012 22332
rect 33036 22330 33092 22332
rect 33116 22330 33172 22332
rect 33196 22330 33252 22332
rect 32956 22278 33002 22330
rect 33002 22278 33012 22330
rect 33036 22278 33066 22330
rect 33066 22278 33078 22330
rect 33078 22278 33092 22330
rect 33116 22278 33130 22330
rect 33130 22278 33142 22330
rect 33142 22278 33172 22330
rect 33196 22278 33206 22330
rect 33206 22278 33252 22330
rect 32956 22276 33012 22278
rect 33036 22276 33092 22278
rect 33116 22276 33172 22278
rect 33196 22276 33252 22278
rect 33782 24384 33838 24440
rect 33966 23432 34022 23488
rect 33046 21972 33048 21992
rect 33048 21972 33100 21992
rect 33100 21972 33102 21992
rect 33046 21936 33102 21972
rect 32494 20984 32550 21040
rect 32402 20848 32458 20904
rect 31850 20324 31906 20360
rect 31850 20304 31852 20324
rect 31852 20304 31904 20324
rect 31904 20304 31906 20324
rect 31114 14068 31170 14104
rect 31114 14048 31116 14068
rect 31116 14048 31168 14068
rect 31168 14048 31170 14068
rect 31206 11636 31208 11656
rect 31208 11636 31260 11656
rect 31260 11636 31262 11656
rect 31206 11600 31262 11636
rect 32034 16632 32090 16688
rect 32956 21242 33012 21244
rect 33036 21242 33092 21244
rect 33116 21242 33172 21244
rect 33196 21242 33252 21244
rect 32956 21190 33002 21242
rect 33002 21190 33012 21242
rect 33036 21190 33066 21242
rect 33066 21190 33078 21242
rect 33078 21190 33092 21242
rect 33116 21190 33130 21242
rect 33130 21190 33142 21242
rect 33142 21190 33172 21242
rect 33196 21190 33206 21242
rect 33206 21190 33252 21242
rect 32956 21188 33012 21190
rect 33036 21188 33092 21190
rect 33116 21188 33172 21190
rect 33196 21188 33252 21190
rect 32956 20154 33012 20156
rect 33036 20154 33092 20156
rect 33116 20154 33172 20156
rect 33196 20154 33252 20156
rect 32956 20102 33002 20154
rect 33002 20102 33012 20154
rect 33036 20102 33066 20154
rect 33066 20102 33078 20154
rect 33078 20102 33092 20154
rect 33116 20102 33130 20154
rect 33130 20102 33142 20154
rect 33142 20102 33172 20154
rect 33196 20102 33206 20154
rect 33206 20102 33252 20154
rect 32956 20100 33012 20102
rect 33036 20100 33092 20102
rect 33116 20100 33172 20102
rect 33196 20100 33252 20102
rect 32494 15816 32550 15872
rect 32218 13796 32274 13832
rect 32218 13776 32220 13796
rect 32220 13776 32272 13796
rect 32272 13776 32274 13796
rect 32034 11600 32090 11656
rect 31482 9716 31538 9752
rect 31482 9696 31484 9716
rect 31484 9696 31536 9716
rect 31536 9696 31538 9716
rect 32956 19066 33012 19068
rect 33036 19066 33092 19068
rect 33116 19066 33172 19068
rect 33196 19066 33252 19068
rect 32956 19014 33002 19066
rect 33002 19014 33012 19066
rect 33036 19014 33066 19066
rect 33066 19014 33078 19066
rect 33078 19014 33092 19066
rect 33116 19014 33130 19066
rect 33130 19014 33142 19066
rect 33142 19014 33172 19066
rect 33196 19014 33206 19066
rect 33206 19014 33252 19066
rect 32956 19012 33012 19014
rect 33036 19012 33092 19014
rect 33116 19012 33172 19014
rect 33196 19012 33252 19014
rect 32954 18572 32956 18592
rect 32956 18572 33008 18592
rect 33008 18572 33010 18592
rect 32954 18536 33010 18572
rect 32956 17978 33012 17980
rect 33036 17978 33092 17980
rect 33116 17978 33172 17980
rect 33196 17978 33252 17980
rect 32956 17926 33002 17978
rect 33002 17926 33012 17978
rect 33036 17926 33066 17978
rect 33066 17926 33078 17978
rect 33078 17926 33092 17978
rect 33116 17926 33130 17978
rect 33130 17926 33142 17978
rect 33142 17926 33172 17978
rect 33196 17926 33206 17978
rect 33206 17926 33252 17978
rect 32956 17924 33012 17926
rect 33036 17924 33092 17926
rect 33116 17924 33172 17926
rect 33196 17924 33252 17926
rect 33690 21548 33746 21584
rect 33690 21528 33692 21548
rect 33692 21528 33744 21548
rect 33744 21528 33746 21548
rect 33598 21256 33654 21312
rect 32956 16890 33012 16892
rect 33036 16890 33092 16892
rect 33116 16890 33172 16892
rect 33196 16890 33252 16892
rect 32956 16838 33002 16890
rect 33002 16838 33012 16890
rect 33036 16838 33066 16890
rect 33066 16838 33078 16890
rect 33078 16838 33092 16890
rect 33116 16838 33130 16890
rect 33130 16838 33142 16890
rect 33142 16838 33172 16890
rect 33196 16838 33206 16890
rect 33206 16838 33252 16890
rect 32956 16836 33012 16838
rect 33036 16836 33092 16838
rect 33116 16836 33172 16838
rect 33196 16836 33252 16838
rect 32956 15802 33012 15804
rect 33036 15802 33092 15804
rect 33116 15802 33172 15804
rect 33196 15802 33252 15804
rect 32956 15750 33002 15802
rect 33002 15750 33012 15802
rect 33036 15750 33066 15802
rect 33066 15750 33078 15802
rect 33078 15750 33092 15802
rect 33116 15750 33130 15802
rect 33130 15750 33142 15802
rect 33142 15750 33172 15802
rect 33196 15750 33206 15802
rect 33206 15750 33252 15802
rect 32956 15748 33012 15750
rect 33036 15748 33092 15750
rect 33116 15748 33172 15750
rect 33196 15748 33252 15750
rect 32956 14714 33012 14716
rect 33036 14714 33092 14716
rect 33116 14714 33172 14716
rect 33196 14714 33252 14716
rect 32956 14662 33002 14714
rect 33002 14662 33012 14714
rect 33036 14662 33066 14714
rect 33066 14662 33078 14714
rect 33078 14662 33092 14714
rect 33116 14662 33130 14714
rect 33130 14662 33142 14714
rect 33142 14662 33172 14714
rect 33196 14662 33206 14714
rect 33206 14662 33252 14714
rect 32956 14660 33012 14662
rect 33036 14660 33092 14662
rect 33116 14660 33172 14662
rect 33196 14660 33252 14662
rect 33966 22652 33968 22672
rect 33968 22652 34020 22672
rect 34020 22652 34022 22672
rect 33966 22616 34022 22652
rect 34886 24656 34942 24712
rect 35254 24012 35256 24032
rect 35256 24012 35308 24032
rect 35308 24012 35310 24032
rect 35254 23976 35310 24012
rect 35530 23432 35586 23488
rect 35714 23296 35770 23352
rect 34886 22752 34942 22808
rect 34242 22480 34298 22536
rect 33966 19352 34022 19408
rect 34794 21664 34850 21720
rect 34794 21392 34850 21448
rect 34426 20576 34482 20632
rect 34610 20576 34666 20632
rect 34518 19760 34574 19816
rect 34150 18572 34152 18592
rect 34152 18572 34204 18592
rect 34204 18572 34206 18592
rect 34150 18536 34206 18572
rect 32956 13626 33012 13628
rect 33036 13626 33092 13628
rect 33116 13626 33172 13628
rect 33196 13626 33252 13628
rect 32956 13574 33002 13626
rect 33002 13574 33012 13626
rect 33036 13574 33066 13626
rect 33066 13574 33078 13626
rect 33078 13574 33092 13626
rect 33116 13574 33130 13626
rect 33130 13574 33142 13626
rect 33142 13574 33172 13626
rect 33196 13574 33206 13626
rect 33206 13574 33252 13626
rect 32956 13572 33012 13574
rect 33036 13572 33092 13574
rect 33116 13572 33172 13574
rect 33196 13572 33252 13574
rect 33690 13776 33746 13832
rect 32956 12538 33012 12540
rect 33036 12538 33092 12540
rect 33116 12538 33172 12540
rect 33196 12538 33252 12540
rect 32956 12486 33002 12538
rect 33002 12486 33012 12538
rect 33036 12486 33066 12538
rect 33066 12486 33078 12538
rect 33078 12486 33092 12538
rect 33116 12486 33130 12538
rect 33130 12486 33142 12538
rect 33142 12486 33172 12538
rect 33196 12486 33206 12538
rect 33206 12486 33252 12538
rect 32956 12484 33012 12486
rect 33036 12484 33092 12486
rect 33116 12484 33172 12486
rect 33196 12484 33252 12486
rect 32956 11450 33012 11452
rect 33036 11450 33092 11452
rect 33116 11450 33172 11452
rect 33196 11450 33252 11452
rect 32956 11398 33002 11450
rect 33002 11398 33012 11450
rect 33036 11398 33066 11450
rect 33066 11398 33078 11450
rect 33078 11398 33092 11450
rect 33116 11398 33130 11450
rect 33130 11398 33142 11450
rect 33142 11398 33172 11450
rect 33196 11398 33206 11450
rect 33206 11398 33252 11450
rect 32956 11396 33012 11398
rect 33036 11396 33092 11398
rect 33116 11396 33172 11398
rect 33196 11396 33252 11398
rect 32586 9424 32642 9480
rect 31942 9016 31998 9072
rect 32956 10362 33012 10364
rect 33036 10362 33092 10364
rect 33116 10362 33172 10364
rect 33196 10362 33252 10364
rect 32956 10310 33002 10362
rect 33002 10310 33012 10362
rect 33036 10310 33066 10362
rect 33066 10310 33078 10362
rect 33078 10310 33092 10362
rect 33116 10310 33130 10362
rect 33130 10310 33142 10362
rect 33142 10310 33172 10362
rect 33196 10310 33206 10362
rect 33206 10310 33252 10362
rect 32956 10308 33012 10310
rect 33036 10308 33092 10310
rect 33116 10308 33172 10310
rect 33196 10308 33252 10310
rect 33230 9696 33286 9752
rect 33690 10648 33746 10704
rect 33874 10648 33930 10704
rect 32956 9274 33012 9276
rect 33036 9274 33092 9276
rect 33116 9274 33172 9276
rect 33196 9274 33252 9276
rect 32956 9222 33002 9274
rect 33002 9222 33012 9274
rect 33036 9222 33066 9274
rect 33066 9222 33078 9274
rect 33078 9222 33092 9274
rect 33116 9222 33130 9274
rect 33130 9222 33142 9274
rect 33142 9222 33172 9274
rect 33196 9222 33206 9274
rect 33206 9222 33252 9274
rect 32956 9220 33012 9222
rect 33036 9220 33092 9222
rect 33116 9220 33172 9222
rect 33196 9220 33252 9222
rect 33046 9016 33102 9072
rect 34426 17992 34482 18048
rect 34334 15952 34390 16008
rect 34426 15408 34482 15464
rect 34886 17992 34942 18048
rect 34426 12144 34482 12200
rect 34242 10648 34298 10704
rect 32956 8186 33012 8188
rect 33036 8186 33092 8188
rect 33116 8186 33172 8188
rect 33196 8186 33252 8188
rect 32956 8134 33002 8186
rect 33002 8134 33012 8186
rect 33036 8134 33066 8186
rect 33066 8134 33078 8186
rect 33078 8134 33092 8186
rect 33116 8134 33130 8186
rect 33130 8134 33142 8186
rect 33142 8134 33172 8186
rect 33196 8134 33206 8186
rect 33206 8134 33252 8186
rect 32956 8132 33012 8134
rect 33036 8132 33092 8134
rect 33116 8132 33172 8134
rect 33196 8132 33252 8134
rect 32956 7098 33012 7100
rect 33036 7098 33092 7100
rect 33116 7098 33172 7100
rect 33196 7098 33252 7100
rect 32956 7046 33002 7098
rect 33002 7046 33012 7098
rect 33036 7046 33066 7098
rect 33066 7046 33078 7098
rect 33078 7046 33092 7098
rect 33116 7046 33130 7098
rect 33130 7046 33142 7098
rect 33142 7046 33172 7098
rect 33196 7046 33206 7098
rect 33206 7046 33252 7098
rect 32956 7044 33012 7046
rect 33036 7044 33092 7046
rect 33116 7044 33172 7046
rect 33196 7044 33252 7046
rect 35438 22344 35494 22400
rect 35898 23160 35954 23216
rect 35622 22092 35678 22128
rect 35622 22072 35624 22092
rect 35624 22072 35676 22092
rect 35676 22072 35678 22092
rect 35898 21120 35954 21176
rect 35254 19252 35256 19272
rect 35256 19252 35308 19272
rect 35308 19252 35310 19272
rect 35254 19216 35310 19252
rect 35622 18536 35678 18592
rect 35346 13252 35402 13288
rect 35346 13232 35348 13252
rect 35348 13232 35400 13252
rect 35400 13232 35402 13252
rect 34610 9560 34666 9616
rect 32956 6010 33012 6012
rect 33036 6010 33092 6012
rect 33116 6010 33172 6012
rect 33196 6010 33252 6012
rect 32956 5958 33002 6010
rect 33002 5958 33012 6010
rect 33036 5958 33066 6010
rect 33066 5958 33078 6010
rect 33078 5958 33092 6010
rect 33116 5958 33130 6010
rect 33130 5958 33142 6010
rect 33142 5958 33172 6010
rect 33196 5958 33206 6010
rect 33206 5958 33252 6010
rect 32956 5956 33012 5958
rect 33036 5956 33092 5958
rect 33116 5956 33172 5958
rect 33196 5956 33252 5958
rect 32956 4922 33012 4924
rect 33036 4922 33092 4924
rect 33116 4922 33172 4924
rect 33196 4922 33252 4924
rect 32956 4870 33002 4922
rect 33002 4870 33012 4922
rect 33036 4870 33066 4922
rect 33066 4870 33078 4922
rect 33078 4870 33092 4922
rect 33116 4870 33130 4922
rect 33130 4870 33142 4922
rect 33142 4870 33172 4922
rect 33196 4870 33206 4922
rect 33206 4870 33252 4922
rect 32956 4868 33012 4870
rect 33036 4868 33092 4870
rect 33116 4868 33172 4870
rect 33196 4868 33252 4870
rect 32956 3834 33012 3836
rect 33036 3834 33092 3836
rect 33116 3834 33172 3836
rect 33196 3834 33252 3836
rect 32956 3782 33002 3834
rect 33002 3782 33012 3834
rect 33036 3782 33066 3834
rect 33066 3782 33078 3834
rect 33078 3782 33092 3834
rect 33116 3782 33130 3834
rect 33130 3782 33142 3834
rect 33142 3782 33172 3834
rect 33196 3782 33206 3834
rect 33206 3782 33252 3834
rect 32956 3780 33012 3782
rect 33036 3780 33092 3782
rect 33116 3780 33172 3782
rect 33196 3780 33252 3782
rect 32956 2746 33012 2748
rect 33036 2746 33092 2748
rect 33116 2746 33172 2748
rect 33196 2746 33252 2748
rect 32956 2694 33002 2746
rect 33002 2694 33012 2746
rect 33036 2694 33066 2746
rect 33066 2694 33078 2746
rect 33078 2694 33092 2746
rect 33116 2694 33130 2746
rect 33130 2694 33142 2746
rect 33142 2694 33172 2746
rect 33196 2694 33206 2746
rect 33206 2694 33252 2746
rect 32956 2692 33012 2694
rect 33036 2692 33092 2694
rect 33116 2692 33172 2694
rect 33196 2692 33252 2694
rect 35714 15952 35770 16008
rect 35898 19508 35954 19544
rect 35898 19488 35900 19508
rect 35900 19488 35952 19508
rect 35952 19488 35954 19508
rect 37002 23704 37058 23760
rect 36726 23160 36782 23216
rect 36450 22888 36506 22944
rect 35898 17992 35954 18048
rect 35714 14456 35770 14512
rect 35806 12824 35862 12880
rect 35806 12688 35862 12744
rect 35806 9560 35862 9616
rect 36634 20576 36690 20632
rect 36542 19488 36598 19544
rect 37186 21936 37242 21992
rect 36910 19236 36966 19272
rect 36910 19216 36912 19236
rect 36912 19216 36964 19236
rect 36964 19216 36966 19236
rect 37094 20712 37150 20768
rect 37646 24012 37648 24032
rect 37648 24012 37700 24032
rect 37700 24012 37702 24032
rect 37646 23976 37702 24012
rect 37956 23962 38012 23964
rect 38036 23962 38092 23964
rect 38116 23962 38172 23964
rect 38196 23962 38252 23964
rect 37956 23910 38002 23962
rect 38002 23910 38012 23962
rect 38036 23910 38066 23962
rect 38066 23910 38078 23962
rect 38078 23910 38092 23962
rect 38116 23910 38130 23962
rect 38130 23910 38142 23962
rect 38142 23910 38172 23962
rect 38196 23910 38206 23962
rect 38206 23910 38252 23962
rect 37956 23908 38012 23910
rect 38036 23908 38092 23910
rect 38116 23908 38172 23910
rect 38196 23908 38252 23910
rect 37956 22874 38012 22876
rect 38036 22874 38092 22876
rect 38116 22874 38172 22876
rect 38196 22874 38252 22876
rect 37956 22822 38002 22874
rect 38002 22822 38012 22874
rect 38036 22822 38066 22874
rect 38066 22822 38078 22874
rect 38078 22822 38092 22874
rect 38116 22822 38130 22874
rect 38130 22822 38142 22874
rect 38142 22822 38172 22874
rect 38196 22822 38206 22874
rect 38206 22822 38252 22874
rect 37956 22820 38012 22822
rect 38036 22820 38092 22822
rect 38116 22820 38172 22822
rect 38196 22820 38252 22822
rect 37738 22516 37740 22536
rect 37740 22516 37792 22536
rect 37792 22516 37794 22536
rect 37738 22480 37794 22516
rect 38474 23840 38530 23896
rect 38842 23432 38898 23488
rect 37956 21786 38012 21788
rect 38036 21786 38092 21788
rect 38116 21786 38172 21788
rect 38196 21786 38252 21788
rect 37956 21734 38002 21786
rect 38002 21734 38012 21786
rect 38036 21734 38066 21786
rect 38066 21734 38078 21786
rect 38078 21734 38092 21786
rect 38116 21734 38130 21786
rect 38130 21734 38142 21786
rect 38142 21734 38172 21786
rect 38196 21734 38206 21786
rect 38206 21734 38252 21786
rect 37956 21732 38012 21734
rect 38036 21732 38092 21734
rect 38116 21732 38172 21734
rect 38196 21732 38252 21734
rect 36082 12824 36138 12880
rect 36726 17040 36782 17096
rect 37956 20698 38012 20700
rect 38036 20698 38092 20700
rect 38116 20698 38172 20700
rect 38196 20698 38252 20700
rect 37956 20646 38002 20698
rect 38002 20646 38012 20698
rect 38036 20646 38066 20698
rect 38066 20646 38078 20698
rect 38078 20646 38092 20698
rect 38116 20646 38130 20698
rect 38130 20646 38142 20698
rect 38142 20646 38172 20698
rect 38196 20646 38206 20698
rect 38206 20646 38252 20698
rect 37956 20644 38012 20646
rect 38036 20644 38092 20646
rect 38116 20644 38172 20646
rect 38196 20644 38252 20646
rect 37956 19610 38012 19612
rect 38036 19610 38092 19612
rect 38116 19610 38172 19612
rect 38196 19610 38252 19612
rect 37956 19558 38002 19610
rect 38002 19558 38012 19610
rect 38036 19558 38066 19610
rect 38066 19558 38078 19610
rect 38078 19558 38092 19610
rect 38116 19558 38130 19610
rect 38130 19558 38142 19610
rect 38142 19558 38172 19610
rect 38196 19558 38206 19610
rect 38206 19558 38252 19610
rect 37956 19556 38012 19558
rect 38036 19556 38092 19558
rect 38116 19556 38172 19558
rect 38196 19556 38252 19558
rect 38382 19508 38438 19544
rect 38382 19488 38384 19508
rect 38384 19488 38436 19508
rect 38436 19488 38438 19508
rect 38198 19252 38200 19272
rect 38200 19252 38252 19272
rect 38252 19252 38254 19272
rect 38198 19216 38254 19252
rect 38014 18672 38070 18728
rect 37956 18522 38012 18524
rect 38036 18522 38092 18524
rect 38116 18522 38172 18524
rect 38196 18522 38252 18524
rect 37956 18470 38002 18522
rect 38002 18470 38012 18522
rect 38036 18470 38066 18522
rect 38066 18470 38078 18522
rect 38078 18470 38092 18522
rect 38116 18470 38130 18522
rect 38130 18470 38142 18522
rect 38142 18470 38172 18522
rect 38196 18470 38206 18522
rect 38206 18470 38252 18522
rect 37956 18468 38012 18470
rect 38036 18468 38092 18470
rect 38116 18468 38172 18470
rect 38196 18468 38252 18470
rect 37186 14864 37242 14920
rect 37956 17434 38012 17436
rect 38036 17434 38092 17436
rect 38116 17434 38172 17436
rect 38196 17434 38252 17436
rect 37956 17382 38002 17434
rect 38002 17382 38012 17434
rect 38036 17382 38066 17434
rect 38066 17382 38078 17434
rect 38078 17382 38092 17434
rect 38116 17382 38130 17434
rect 38130 17382 38142 17434
rect 38142 17382 38172 17434
rect 38196 17382 38206 17434
rect 38206 17382 38252 17434
rect 37956 17380 38012 17382
rect 38036 17380 38092 17382
rect 38116 17380 38172 17382
rect 38196 17380 38252 17382
rect 39394 23024 39450 23080
rect 39394 22072 39450 22128
rect 40682 24384 40738 24440
rect 39210 20440 39266 20496
rect 38934 19352 38990 19408
rect 37956 16346 38012 16348
rect 38036 16346 38092 16348
rect 38116 16346 38172 16348
rect 38196 16346 38252 16348
rect 37956 16294 38002 16346
rect 38002 16294 38012 16346
rect 38036 16294 38066 16346
rect 38066 16294 38078 16346
rect 38078 16294 38092 16346
rect 38116 16294 38130 16346
rect 38130 16294 38142 16346
rect 38142 16294 38172 16346
rect 38196 16294 38206 16346
rect 38206 16294 38252 16346
rect 37956 16292 38012 16294
rect 38036 16292 38092 16294
rect 38116 16292 38172 16294
rect 38196 16292 38252 16294
rect 37956 15258 38012 15260
rect 38036 15258 38092 15260
rect 38116 15258 38172 15260
rect 38196 15258 38252 15260
rect 37956 15206 38002 15258
rect 38002 15206 38012 15258
rect 38036 15206 38066 15258
rect 38066 15206 38078 15258
rect 38078 15206 38092 15258
rect 38116 15206 38130 15258
rect 38130 15206 38142 15258
rect 38142 15206 38172 15258
rect 38196 15206 38206 15258
rect 38206 15206 38252 15258
rect 37956 15204 38012 15206
rect 38036 15204 38092 15206
rect 38116 15204 38172 15206
rect 38196 15204 38252 15206
rect 38474 17076 38476 17096
rect 38476 17076 38528 17096
rect 38528 17076 38530 17096
rect 38474 17040 38530 17076
rect 38474 16496 38530 16552
rect 40958 24268 41014 24304
rect 40958 24248 40960 24268
rect 40960 24248 41012 24268
rect 41012 24248 41014 24268
rect 40314 21140 40370 21176
rect 40314 21120 40316 21140
rect 40316 21120 40368 21140
rect 40368 21120 40370 21140
rect 40774 22480 40830 22536
rect 39026 18128 39082 18184
rect 39578 17720 39634 17776
rect 38566 14864 38622 14920
rect 37956 14170 38012 14172
rect 38036 14170 38092 14172
rect 38116 14170 38172 14172
rect 38196 14170 38252 14172
rect 37956 14118 38002 14170
rect 38002 14118 38012 14170
rect 38036 14118 38066 14170
rect 38066 14118 38078 14170
rect 38078 14118 38092 14170
rect 38116 14118 38130 14170
rect 38130 14118 38142 14170
rect 38142 14118 38172 14170
rect 38196 14118 38206 14170
rect 38206 14118 38252 14170
rect 37956 14116 38012 14118
rect 38036 14116 38092 14118
rect 38116 14116 38172 14118
rect 38196 14116 38252 14118
rect 40406 19896 40462 19952
rect 40130 18808 40186 18864
rect 40406 19080 40462 19136
rect 40590 19216 40646 19272
rect 40866 20984 40922 21040
rect 41326 22072 41382 22128
rect 40958 20848 41014 20904
rect 41418 21412 41474 21448
rect 41418 21392 41420 21412
rect 41420 21392 41472 21412
rect 41472 21392 41474 21412
rect 42246 23840 42302 23896
rect 42956 24506 43012 24508
rect 43036 24506 43092 24508
rect 43116 24506 43172 24508
rect 43196 24506 43252 24508
rect 42956 24454 43002 24506
rect 43002 24454 43012 24506
rect 43036 24454 43066 24506
rect 43066 24454 43078 24506
rect 43078 24454 43092 24506
rect 43116 24454 43130 24506
rect 43130 24454 43142 24506
rect 43142 24454 43172 24506
rect 43196 24454 43206 24506
rect 43206 24454 43252 24506
rect 42956 24452 43012 24454
rect 43036 24452 43092 24454
rect 43116 24452 43172 24454
rect 43196 24452 43252 24454
rect 42154 22752 42210 22808
rect 41878 22072 41934 22128
rect 41694 21936 41750 21992
rect 41510 21256 41566 21312
rect 42956 23418 43012 23420
rect 43036 23418 43092 23420
rect 43116 23418 43172 23420
rect 43196 23418 43252 23420
rect 42956 23366 43002 23418
rect 43002 23366 43012 23418
rect 43036 23366 43066 23418
rect 43066 23366 43078 23418
rect 43078 23366 43092 23418
rect 43116 23366 43130 23418
rect 43130 23366 43142 23418
rect 43142 23366 43172 23418
rect 43196 23366 43206 23418
rect 43206 23366 43252 23418
rect 42956 23364 43012 23366
rect 43036 23364 43092 23366
rect 43116 23364 43172 23366
rect 43196 23364 43252 23366
rect 42614 23296 42670 23352
rect 43902 23196 43904 23216
rect 43904 23196 43956 23216
rect 43956 23196 43958 23216
rect 43902 23160 43958 23196
rect 43534 23044 43590 23080
rect 43534 23024 43536 23044
rect 43536 23024 43588 23044
rect 43588 23024 43590 23044
rect 42614 22500 42670 22536
rect 42614 22480 42616 22500
rect 42616 22480 42668 22500
rect 42668 22480 42670 22500
rect 42956 22330 43012 22332
rect 43036 22330 43092 22332
rect 43116 22330 43172 22332
rect 43196 22330 43252 22332
rect 42956 22278 43002 22330
rect 43002 22278 43012 22330
rect 43036 22278 43066 22330
rect 43066 22278 43078 22330
rect 43078 22278 43092 22330
rect 43116 22278 43130 22330
rect 43130 22278 43142 22330
rect 43142 22278 43172 22330
rect 43196 22278 43206 22330
rect 43206 22278 43252 22330
rect 42956 22276 43012 22278
rect 43036 22276 43092 22278
rect 43116 22276 43172 22278
rect 43196 22276 43252 22278
rect 42798 21528 42854 21584
rect 42956 21242 43012 21244
rect 43036 21242 43092 21244
rect 43116 21242 43172 21244
rect 43196 21242 43252 21244
rect 42956 21190 43002 21242
rect 43002 21190 43012 21242
rect 43036 21190 43066 21242
rect 43066 21190 43078 21242
rect 43078 21190 43092 21242
rect 43116 21190 43130 21242
rect 43130 21190 43142 21242
rect 43142 21190 43172 21242
rect 43196 21190 43206 21242
rect 43206 21190 43252 21242
rect 42956 21188 43012 21190
rect 43036 21188 43092 21190
rect 43116 21188 43172 21190
rect 43196 21188 43252 21190
rect 42956 20154 43012 20156
rect 43036 20154 43092 20156
rect 43116 20154 43172 20156
rect 43196 20154 43252 20156
rect 42956 20102 43002 20154
rect 43002 20102 43012 20154
rect 43036 20102 43066 20154
rect 43066 20102 43078 20154
rect 43078 20102 43092 20154
rect 43116 20102 43130 20154
rect 43130 20102 43142 20154
rect 43142 20102 43172 20154
rect 43196 20102 43206 20154
rect 43206 20102 43252 20154
rect 42956 20100 43012 20102
rect 43036 20100 43092 20102
rect 43116 20100 43172 20102
rect 43196 20100 43252 20102
rect 44546 24656 44602 24712
rect 46662 25064 46718 25120
rect 46570 24656 46626 24712
rect 45374 23724 45430 23760
rect 45374 23704 45376 23724
rect 45376 23704 45428 23724
rect 45428 23704 45430 23724
rect 45190 23588 45246 23624
rect 45190 23568 45192 23588
rect 45192 23568 45244 23588
rect 45244 23568 45246 23588
rect 40682 18264 40738 18320
rect 42956 19066 43012 19068
rect 43036 19066 43092 19068
rect 43116 19066 43172 19068
rect 43196 19066 43252 19068
rect 42956 19014 43002 19066
rect 43002 19014 43012 19066
rect 43036 19014 43066 19066
rect 43066 19014 43078 19066
rect 43078 19014 43092 19066
rect 43116 19014 43130 19066
rect 43130 19014 43142 19066
rect 43142 19014 43172 19066
rect 43196 19014 43206 19066
rect 43206 19014 43252 19066
rect 42956 19012 43012 19014
rect 43036 19012 43092 19014
rect 43116 19012 43172 19014
rect 43196 19012 43252 19014
rect 42956 17978 43012 17980
rect 43036 17978 43092 17980
rect 43116 17978 43172 17980
rect 43196 17978 43252 17980
rect 42956 17926 43002 17978
rect 43002 17926 43012 17978
rect 43036 17926 43066 17978
rect 43066 17926 43078 17978
rect 43078 17926 43092 17978
rect 43116 17926 43130 17978
rect 43130 17926 43142 17978
rect 43142 17926 43172 17978
rect 43196 17926 43206 17978
rect 43206 17926 43252 17978
rect 42956 17924 43012 17926
rect 43036 17924 43092 17926
rect 43116 17924 43172 17926
rect 43196 17924 43252 17926
rect 42706 17176 42762 17232
rect 42956 16890 43012 16892
rect 43036 16890 43092 16892
rect 43116 16890 43172 16892
rect 43196 16890 43252 16892
rect 42956 16838 43002 16890
rect 43002 16838 43012 16890
rect 43036 16838 43066 16890
rect 43066 16838 43078 16890
rect 43078 16838 43092 16890
rect 43116 16838 43130 16890
rect 43130 16838 43142 16890
rect 43142 16838 43172 16890
rect 43196 16838 43206 16890
rect 43206 16838 43252 16890
rect 42956 16836 43012 16838
rect 43036 16836 43092 16838
rect 43116 16836 43172 16838
rect 43196 16836 43252 16838
rect 47582 24248 47638 24304
rect 47122 22752 47178 22808
rect 48226 25472 48282 25528
rect 47956 23962 48012 23964
rect 48036 23962 48092 23964
rect 48116 23962 48172 23964
rect 48196 23962 48252 23964
rect 47956 23910 48002 23962
rect 48002 23910 48012 23962
rect 48036 23910 48066 23962
rect 48066 23910 48078 23962
rect 48078 23910 48092 23962
rect 48116 23910 48130 23962
rect 48130 23910 48142 23962
rect 48142 23910 48172 23962
rect 48196 23910 48206 23962
rect 48206 23910 48252 23962
rect 47956 23908 48012 23910
rect 48036 23908 48092 23910
rect 48116 23908 48172 23910
rect 48196 23908 48252 23910
rect 47858 23432 47914 23488
rect 48410 23840 48466 23896
rect 48778 24148 48780 24168
rect 48780 24148 48832 24168
rect 48832 24148 48834 24168
rect 48778 24112 48834 24148
rect 48318 23060 48320 23080
rect 48320 23060 48372 23080
rect 48372 23060 48374 23080
rect 48318 23024 48374 23060
rect 47956 22874 48012 22876
rect 48036 22874 48092 22876
rect 48116 22874 48172 22876
rect 48196 22874 48252 22876
rect 47956 22822 48002 22874
rect 48002 22822 48012 22874
rect 48036 22822 48066 22874
rect 48066 22822 48078 22874
rect 48078 22822 48092 22874
rect 48116 22822 48130 22874
rect 48130 22822 48142 22874
rect 48142 22822 48172 22874
rect 48196 22822 48206 22874
rect 48206 22822 48252 22874
rect 47956 22820 48012 22822
rect 48036 22820 48092 22822
rect 48116 22820 48172 22822
rect 48196 22820 48252 22822
rect 47956 21786 48012 21788
rect 48036 21786 48092 21788
rect 48116 21786 48172 21788
rect 48196 21786 48252 21788
rect 47956 21734 48002 21786
rect 48002 21734 48012 21786
rect 48036 21734 48066 21786
rect 48066 21734 48078 21786
rect 48078 21734 48092 21786
rect 48116 21734 48130 21786
rect 48130 21734 48142 21786
rect 48142 21734 48172 21786
rect 48196 21734 48206 21786
rect 48206 21734 48252 21786
rect 47956 21732 48012 21734
rect 48036 21732 48092 21734
rect 48116 21732 48172 21734
rect 48196 21732 48252 21734
rect 47956 20698 48012 20700
rect 48036 20698 48092 20700
rect 48116 20698 48172 20700
rect 48196 20698 48252 20700
rect 47956 20646 48002 20698
rect 48002 20646 48012 20698
rect 48036 20646 48066 20698
rect 48066 20646 48078 20698
rect 48078 20646 48092 20698
rect 48116 20646 48130 20698
rect 48130 20646 48142 20698
rect 48142 20646 48172 20698
rect 48196 20646 48206 20698
rect 48206 20646 48252 20698
rect 47956 20644 48012 20646
rect 48036 20644 48092 20646
rect 48116 20644 48172 20646
rect 48196 20644 48252 20646
rect 48318 20304 48374 20360
rect 47956 19610 48012 19612
rect 48036 19610 48092 19612
rect 48116 19610 48172 19612
rect 48196 19610 48252 19612
rect 47956 19558 48002 19610
rect 48002 19558 48012 19610
rect 48036 19558 48066 19610
rect 48066 19558 48078 19610
rect 48078 19558 48092 19610
rect 48116 19558 48130 19610
rect 48130 19558 48142 19610
rect 48142 19558 48172 19610
rect 48196 19558 48206 19610
rect 48206 19558 48252 19610
rect 47956 19556 48012 19558
rect 48036 19556 48092 19558
rect 48116 19556 48172 19558
rect 48196 19556 48252 19558
rect 46938 19488 46994 19544
rect 49054 22208 49110 22264
rect 48778 21800 48834 21856
rect 49330 22616 49386 22672
rect 49146 21392 49202 21448
rect 49054 20984 49110 21040
rect 49054 20576 49110 20632
rect 48778 20168 48834 20224
rect 48502 19760 48558 19816
rect 49054 19760 49110 19816
rect 49330 19352 49386 19408
rect 49146 18944 49202 19000
rect 47956 18522 48012 18524
rect 48036 18522 48092 18524
rect 48116 18522 48172 18524
rect 48196 18522 48252 18524
rect 47956 18470 48002 18522
rect 48002 18470 48012 18522
rect 48036 18470 48066 18522
rect 48066 18470 48078 18522
rect 48078 18470 48092 18522
rect 48116 18470 48130 18522
rect 48130 18470 48142 18522
rect 48142 18470 48172 18522
rect 48196 18470 48206 18522
rect 48206 18470 48252 18522
rect 47956 18468 48012 18470
rect 48036 18468 48092 18470
rect 48116 18468 48172 18470
rect 48196 18468 48252 18470
rect 48778 18536 48834 18592
rect 47956 17434 48012 17436
rect 48036 17434 48092 17436
rect 48116 17434 48172 17436
rect 48196 17434 48252 17436
rect 47956 17382 48002 17434
rect 48002 17382 48012 17434
rect 48036 17382 48066 17434
rect 48066 17382 48078 17434
rect 48078 17382 48092 17434
rect 48116 17382 48130 17434
rect 48130 17382 48142 17434
rect 48142 17382 48172 17434
rect 48196 17382 48206 17434
rect 48206 17382 48252 17434
rect 47956 17380 48012 17382
rect 48036 17380 48092 17382
rect 48116 17380 48172 17382
rect 48196 17380 48252 17382
rect 49146 18128 49202 18184
rect 49054 17720 49110 17776
rect 49054 17312 49110 17368
rect 48778 16904 48834 16960
rect 47956 16346 48012 16348
rect 48036 16346 48092 16348
rect 48116 16346 48172 16348
rect 48196 16346 48252 16348
rect 47956 16294 48002 16346
rect 48002 16294 48012 16346
rect 48036 16294 48066 16346
rect 48066 16294 48078 16346
rect 48078 16294 48092 16346
rect 48116 16294 48130 16346
rect 48130 16294 48142 16346
rect 48142 16294 48172 16346
rect 48196 16294 48206 16346
rect 48206 16294 48252 16346
rect 47956 16292 48012 16294
rect 48036 16292 48092 16294
rect 48116 16292 48172 16294
rect 48196 16292 48252 16294
rect 49238 16496 49294 16552
rect 48778 16088 48834 16144
rect 49146 16088 49202 16144
rect 42956 15802 43012 15804
rect 43036 15802 43092 15804
rect 43116 15802 43172 15804
rect 43196 15802 43252 15804
rect 42956 15750 43002 15802
rect 43002 15750 43012 15802
rect 43036 15750 43066 15802
rect 43066 15750 43078 15802
rect 43078 15750 43092 15802
rect 43116 15750 43130 15802
rect 43130 15750 43142 15802
rect 43142 15750 43172 15802
rect 43196 15750 43206 15802
rect 43206 15750 43252 15802
rect 42956 15748 43012 15750
rect 43036 15748 43092 15750
rect 43116 15748 43172 15750
rect 43196 15748 43252 15750
rect 49238 15972 49294 16008
rect 49238 15952 49240 15972
rect 49240 15952 49292 15972
rect 49292 15952 49294 15972
rect 49054 15680 49110 15736
rect 49330 15272 49386 15328
rect 47956 15258 48012 15260
rect 48036 15258 48092 15260
rect 48116 15258 48172 15260
rect 48196 15258 48252 15260
rect 47956 15206 48002 15258
rect 48002 15206 48012 15258
rect 48036 15206 48066 15258
rect 48066 15206 48078 15258
rect 48078 15206 48092 15258
rect 48116 15206 48130 15258
rect 48130 15206 48142 15258
rect 48142 15206 48172 15258
rect 48196 15206 48206 15258
rect 48206 15206 48252 15258
rect 47956 15204 48012 15206
rect 48036 15204 48092 15206
rect 48116 15204 48172 15206
rect 48196 15204 48252 15206
rect 42956 14714 43012 14716
rect 43036 14714 43092 14716
rect 43116 14714 43172 14716
rect 43196 14714 43252 14716
rect 42956 14662 43002 14714
rect 43002 14662 43012 14714
rect 43036 14662 43066 14714
rect 43066 14662 43078 14714
rect 43078 14662 43092 14714
rect 43116 14662 43130 14714
rect 43130 14662 43142 14714
rect 43142 14662 43172 14714
rect 43196 14662 43206 14714
rect 43206 14662 43252 14714
rect 42956 14660 43012 14662
rect 43036 14660 43092 14662
rect 43116 14660 43172 14662
rect 43196 14660 43252 14662
rect 39946 14320 40002 14376
rect 37956 13082 38012 13084
rect 38036 13082 38092 13084
rect 38116 13082 38172 13084
rect 38196 13082 38252 13084
rect 37956 13030 38002 13082
rect 38002 13030 38012 13082
rect 38036 13030 38066 13082
rect 38066 13030 38078 13082
rect 38078 13030 38092 13082
rect 38116 13030 38130 13082
rect 38130 13030 38142 13082
rect 38142 13030 38172 13082
rect 38196 13030 38206 13082
rect 38206 13030 38252 13082
rect 37956 13028 38012 13030
rect 38036 13028 38092 13030
rect 38116 13028 38172 13030
rect 38196 13028 38252 13030
rect 47956 14170 48012 14172
rect 48036 14170 48092 14172
rect 48116 14170 48172 14172
rect 48196 14170 48252 14172
rect 47956 14118 48002 14170
rect 48002 14118 48012 14170
rect 48036 14118 48066 14170
rect 48066 14118 48078 14170
rect 48078 14118 48092 14170
rect 48116 14118 48130 14170
rect 48130 14118 48142 14170
rect 48142 14118 48172 14170
rect 48196 14118 48206 14170
rect 48206 14118 48252 14170
rect 47956 14116 48012 14118
rect 48036 14116 48092 14118
rect 48116 14116 48172 14118
rect 48196 14116 48252 14118
rect 42956 13626 43012 13628
rect 43036 13626 43092 13628
rect 43116 13626 43172 13628
rect 43196 13626 43252 13628
rect 42956 13574 43002 13626
rect 43002 13574 43012 13626
rect 43036 13574 43066 13626
rect 43066 13574 43078 13626
rect 43078 13574 43092 13626
rect 43116 13574 43130 13626
rect 43130 13574 43142 13626
rect 43142 13574 43172 13626
rect 43196 13574 43206 13626
rect 43206 13574 43252 13626
rect 42956 13572 43012 13574
rect 43036 13572 43092 13574
rect 43116 13572 43172 13574
rect 43196 13572 43252 13574
rect 49238 15000 49294 15056
rect 49054 14864 49110 14920
rect 49146 14456 49202 14512
rect 49146 14048 49202 14104
rect 48226 13640 48282 13696
rect 49146 13252 49202 13288
rect 49146 13232 49148 13252
rect 49148 13232 49200 13252
rect 49200 13232 49202 13252
rect 47956 13082 48012 13084
rect 48036 13082 48092 13084
rect 48116 13082 48172 13084
rect 48196 13082 48252 13084
rect 47956 13030 48002 13082
rect 48002 13030 48012 13082
rect 48036 13030 48066 13082
rect 48066 13030 48078 13082
rect 48078 13030 48092 13082
rect 48116 13030 48130 13082
rect 48130 13030 48142 13082
rect 48142 13030 48172 13082
rect 48196 13030 48206 13082
rect 48206 13030 48252 13082
rect 47956 13028 48012 13030
rect 48036 13028 48092 13030
rect 48116 13028 48172 13030
rect 48196 13028 48252 13030
rect 49146 12844 49202 12880
rect 49146 12824 49148 12844
rect 49148 12824 49200 12844
rect 49200 12824 49202 12844
rect 37956 11994 38012 11996
rect 38036 11994 38092 11996
rect 38116 11994 38172 11996
rect 38196 11994 38252 11996
rect 37956 11942 38002 11994
rect 38002 11942 38012 11994
rect 38036 11942 38066 11994
rect 38066 11942 38078 11994
rect 38078 11942 38092 11994
rect 38116 11942 38130 11994
rect 38130 11942 38142 11994
rect 38142 11942 38172 11994
rect 38196 11942 38206 11994
rect 38206 11942 38252 11994
rect 37956 11940 38012 11942
rect 38036 11940 38092 11942
rect 38116 11940 38172 11942
rect 38196 11940 38252 11942
rect 37956 10906 38012 10908
rect 38036 10906 38092 10908
rect 38116 10906 38172 10908
rect 38196 10906 38252 10908
rect 37956 10854 38002 10906
rect 38002 10854 38012 10906
rect 38036 10854 38066 10906
rect 38066 10854 38078 10906
rect 38078 10854 38092 10906
rect 38116 10854 38130 10906
rect 38130 10854 38142 10906
rect 38142 10854 38172 10906
rect 38196 10854 38206 10906
rect 38206 10854 38252 10906
rect 37956 10852 38012 10854
rect 38036 10852 38092 10854
rect 38116 10852 38172 10854
rect 38196 10852 38252 10854
rect 38566 10104 38622 10160
rect 37956 9818 38012 9820
rect 38036 9818 38092 9820
rect 38116 9818 38172 9820
rect 38196 9818 38252 9820
rect 37956 9766 38002 9818
rect 38002 9766 38012 9818
rect 38036 9766 38066 9818
rect 38066 9766 38078 9818
rect 38078 9766 38092 9818
rect 38116 9766 38130 9818
rect 38130 9766 38142 9818
rect 38142 9766 38172 9818
rect 38196 9766 38206 9818
rect 38206 9766 38252 9818
rect 37956 9764 38012 9766
rect 38036 9764 38092 9766
rect 38116 9764 38172 9766
rect 38196 9764 38252 9766
rect 37956 8730 38012 8732
rect 38036 8730 38092 8732
rect 38116 8730 38172 8732
rect 38196 8730 38252 8732
rect 37956 8678 38002 8730
rect 38002 8678 38012 8730
rect 38036 8678 38066 8730
rect 38066 8678 38078 8730
rect 38078 8678 38092 8730
rect 38116 8678 38130 8730
rect 38130 8678 38142 8730
rect 38142 8678 38172 8730
rect 38196 8678 38206 8730
rect 38206 8678 38252 8730
rect 37956 8676 38012 8678
rect 38036 8676 38092 8678
rect 38116 8676 38172 8678
rect 38196 8676 38252 8678
rect 42956 12538 43012 12540
rect 43036 12538 43092 12540
rect 43116 12538 43172 12540
rect 43196 12538 43252 12540
rect 42956 12486 43002 12538
rect 43002 12486 43012 12538
rect 43036 12486 43066 12538
rect 43066 12486 43078 12538
rect 43078 12486 43092 12538
rect 43116 12486 43130 12538
rect 43130 12486 43142 12538
rect 43142 12486 43172 12538
rect 43196 12486 43206 12538
rect 43206 12486 43252 12538
rect 42956 12484 43012 12486
rect 43036 12484 43092 12486
rect 43116 12484 43172 12486
rect 43196 12484 43252 12486
rect 42956 11450 43012 11452
rect 43036 11450 43092 11452
rect 43116 11450 43172 11452
rect 43196 11450 43252 11452
rect 42956 11398 43002 11450
rect 43002 11398 43012 11450
rect 43036 11398 43066 11450
rect 43066 11398 43078 11450
rect 43078 11398 43092 11450
rect 43116 11398 43130 11450
rect 43130 11398 43142 11450
rect 43142 11398 43172 11450
rect 43196 11398 43206 11450
rect 43206 11398 43252 11450
rect 42956 11396 43012 11398
rect 43036 11396 43092 11398
rect 43116 11396 43172 11398
rect 43196 11396 43252 11398
rect 39946 11056 40002 11112
rect 39762 10668 39818 10704
rect 39762 10648 39764 10668
rect 39764 10648 39816 10668
rect 39816 10648 39818 10668
rect 42956 10362 43012 10364
rect 43036 10362 43092 10364
rect 43116 10362 43172 10364
rect 43196 10362 43252 10364
rect 42956 10310 43002 10362
rect 43002 10310 43012 10362
rect 43036 10310 43066 10362
rect 43066 10310 43078 10362
rect 43078 10310 43092 10362
rect 43116 10310 43130 10362
rect 43130 10310 43142 10362
rect 43142 10310 43172 10362
rect 43196 10310 43206 10362
rect 43206 10310 43252 10362
rect 42956 10308 43012 10310
rect 43036 10308 43092 10310
rect 43116 10308 43172 10310
rect 43196 10308 43252 10310
rect 42956 9274 43012 9276
rect 43036 9274 43092 9276
rect 43116 9274 43172 9276
rect 43196 9274 43252 9276
rect 42956 9222 43002 9274
rect 43002 9222 43012 9274
rect 43036 9222 43066 9274
rect 43066 9222 43078 9274
rect 43078 9222 43092 9274
rect 43116 9222 43130 9274
rect 43130 9222 43142 9274
rect 43142 9222 43172 9274
rect 43196 9222 43206 9274
rect 43206 9222 43252 9274
rect 42956 9220 43012 9222
rect 43036 9220 43092 9222
rect 43116 9220 43172 9222
rect 43196 9220 43252 9222
rect 37956 7642 38012 7644
rect 38036 7642 38092 7644
rect 38116 7642 38172 7644
rect 38196 7642 38252 7644
rect 37956 7590 38002 7642
rect 38002 7590 38012 7642
rect 38036 7590 38066 7642
rect 38066 7590 38078 7642
rect 38078 7590 38092 7642
rect 38116 7590 38130 7642
rect 38130 7590 38142 7642
rect 38142 7590 38172 7642
rect 38196 7590 38206 7642
rect 38206 7590 38252 7642
rect 37956 7588 38012 7590
rect 38036 7588 38092 7590
rect 38116 7588 38172 7590
rect 38196 7588 38252 7590
rect 37956 6554 38012 6556
rect 38036 6554 38092 6556
rect 38116 6554 38172 6556
rect 38196 6554 38252 6556
rect 37956 6502 38002 6554
rect 38002 6502 38012 6554
rect 38036 6502 38066 6554
rect 38066 6502 38078 6554
rect 38078 6502 38092 6554
rect 38116 6502 38130 6554
rect 38130 6502 38142 6554
rect 38142 6502 38172 6554
rect 38196 6502 38206 6554
rect 38206 6502 38252 6554
rect 37956 6500 38012 6502
rect 38036 6500 38092 6502
rect 38116 6500 38172 6502
rect 38196 6500 38252 6502
rect 37956 5466 38012 5468
rect 38036 5466 38092 5468
rect 38116 5466 38172 5468
rect 38196 5466 38252 5468
rect 37956 5414 38002 5466
rect 38002 5414 38012 5466
rect 38036 5414 38066 5466
rect 38066 5414 38078 5466
rect 38078 5414 38092 5466
rect 38116 5414 38130 5466
rect 38130 5414 38142 5466
rect 38142 5414 38172 5466
rect 38196 5414 38206 5466
rect 38206 5414 38252 5466
rect 37956 5412 38012 5414
rect 38036 5412 38092 5414
rect 38116 5412 38172 5414
rect 38196 5412 38252 5414
rect 42956 8186 43012 8188
rect 43036 8186 43092 8188
rect 43116 8186 43172 8188
rect 43196 8186 43252 8188
rect 42956 8134 43002 8186
rect 43002 8134 43012 8186
rect 43036 8134 43066 8186
rect 43066 8134 43078 8186
rect 43078 8134 43092 8186
rect 43116 8134 43130 8186
rect 43130 8134 43142 8186
rect 43142 8134 43172 8186
rect 43196 8134 43206 8186
rect 43206 8134 43252 8186
rect 42956 8132 43012 8134
rect 43036 8132 43092 8134
rect 43116 8132 43172 8134
rect 43196 8132 43252 8134
rect 42956 7098 43012 7100
rect 43036 7098 43092 7100
rect 43116 7098 43172 7100
rect 43196 7098 43252 7100
rect 42956 7046 43002 7098
rect 43002 7046 43012 7098
rect 43036 7046 43066 7098
rect 43066 7046 43078 7098
rect 43078 7046 43092 7098
rect 43116 7046 43130 7098
rect 43130 7046 43142 7098
rect 43142 7046 43172 7098
rect 43196 7046 43206 7098
rect 43206 7046 43252 7098
rect 42956 7044 43012 7046
rect 43036 7044 43092 7046
rect 43116 7044 43172 7046
rect 43196 7044 43252 7046
rect 49146 12416 49202 12472
rect 49146 12008 49202 12064
rect 47956 11994 48012 11996
rect 48036 11994 48092 11996
rect 48116 11994 48172 11996
rect 48196 11994 48252 11996
rect 47956 11942 48002 11994
rect 48002 11942 48012 11994
rect 48036 11942 48066 11994
rect 48066 11942 48078 11994
rect 48078 11942 48092 11994
rect 48116 11942 48130 11994
rect 48130 11942 48142 11994
rect 48142 11942 48172 11994
rect 48196 11942 48206 11994
rect 48206 11942 48252 11994
rect 47956 11940 48012 11942
rect 48036 11940 48092 11942
rect 48116 11940 48172 11942
rect 48196 11940 48252 11942
rect 49146 11600 49202 11656
rect 49238 11192 49294 11248
rect 47956 10906 48012 10908
rect 48036 10906 48092 10908
rect 48116 10906 48172 10908
rect 48196 10906 48252 10908
rect 47956 10854 48002 10906
rect 48002 10854 48012 10906
rect 48036 10854 48066 10906
rect 48066 10854 48078 10906
rect 48078 10854 48092 10906
rect 48116 10854 48130 10906
rect 48130 10854 48142 10906
rect 48142 10854 48172 10906
rect 48196 10854 48206 10906
rect 48206 10854 48252 10906
rect 47956 10852 48012 10854
rect 48036 10852 48092 10854
rect 48116 10852 48172 10854
rect 48196 10852 48252 10854
rect 49146 10784 49202 10840
rect 46846 7928 46902 7984
rect 49330 10376 49386 10432
rect 49238 9968 49294 10024
rect 42956 6010 43012 6012
rect 43036 6010 43092 6012
rect 43116 6010 43172 6012
rect 43196 6010 43252 6012
rect 42956 5958 43002 6010
rect 43002 5958 43012 6010
rect 43036 5958 43066 6010
rect 43066 5958 43078 6010
rect 43078 5958 43092 6010
rect 43116 5958 43130 6010
rect 43130 5958 43142 6010
rect 43142 5958 43172 6010
rect 43196 5958 43206 6010
rect 43206 5958 43252 6010
rect 42956 5956 43012 5958
rect 43036 5956 43092 5958
rect 43116 5956 43172 5958
rect 43196 5956 43252 5958
rect 37956 4378 38012 4380
rect 38036 4378 38092 4380
rect 38116 4378 38172 4380
rect 38196 4378 38252 4380
rect 37956 4326 38002 4378
rect 38002 4326 38012 4378
rect 38036 4326 38066 4378
rect 38066 4326 38078 4378
rect 38078 4326 38092 4378
rect 38116 4326 38130 4378
rect 38130 4326 38142 4378
rect 38142 4326 38172 4378
rect 38196 4326 38206 4378
rect 38206 4326 38252 4378
rect 37956 4324 38012 4326
rect 38036 4324 38092 4326
rect 38116 4324 38172 4326
rect 38196 4324 38252 4326
rect 37956 3290 38012 3292
rect 38036 3290 38092 3292
rect 38116 3290 38172 3292
rect 38196 3290 38252 3292
rect 37956 3238 38002 3290
rect 38002 3238 38012 3290
rect 38036 3238 38066 3290
rect 38066 3238 38078 3290
rect 38078 3238 38092 3290
rect 38116 3238 38130 3290
rect 38130 3238 38142 3290
rect 38142 3238 38172 3290
rect 38196 3238 38206 3290
rect 38206 3238 38252 3290
rect 37956 3236 38012 3238
rect 38036 3236 38092 3238
rect 38116 3236 38172 3238
rect 38196 3236 38252 3238
rect 27956 2202 28012 2204
rect 28036 2202 28092 2204
rect 28116 2202 28172 2204
rect 28196 2202 28252 2204
rect 27956 2150 28002 2202
rect 28002 2150 28012 2202
rect 28036 2150 28066 2202
rect 28066 2150 28078 2202
rect 28078 2150 28092 2202
rect 28116 2150 28130 2202
rect 28130 2150 28142 2202
rect 28142 2150 28172 2202
rect 28196 2150 28206 2202
rect 28206 2150 28252 2202
rect 27956 2148 28012 2150
rect 28036 2148 28092 2150
rect 28116 2148 28172 2150
rect 28196 2148 28252 2150
rect 37956 2202 38012 2204
rect 38036 2202 38092 2204
rect 38116 2202 38172 2204
rect 38196 2202 38252 2204
rect 37956 2150 38002 2202
rect 38002 2150 38012 2202
rect 38036 2150 38066 2202
rect 38066 2150 38078 2202
rect 38078 2150 38092 2202
rect 38116 2150 38130 2202
rect 38130 2150 38142 2202
rect 38142 2150 38172 2202
rect 38196 2150 38206 2202
rect 38206 2150 38252 2202
rect 37956 2148 38012 2150
rect 38036 2148 38092 2150
rect 38116 2148 38172 2150
rect 38196 2148 38252 2150
rect 42956 4922 43012 4924
rect 43036 4922 43092 4924
rect 43116 4922 43172 4924
rect 43196 4922 43252 4924
rect 42956 4870 43002 4922
rect 43002 4870 43012 4922
rect 43036 4870 43066 4922
rect 43066 4870 43078 4922
rect 43078 4870 43092 4922
rect 43116 4870 43130 4922
rect 43130 4870 43142 4922
rect 43142 4870 43172 4922
rect 43196 4870 43206 4922
rect 43206 4870 43252 4922
rect 42956 4868 43012 4870
rect 43036 4868 43092 4870
rect 43116 4868 43172 4870
rect 43196 4868 43252 4870
rect 42956 3834 43012 3836
rect 43036 3834 43092 3836
rect 43116 3834 43172 3836
rect 43196 3834 43252 3836
rect 42956 3782 43002 3834
rect 43002 3782 43012 3834
rect 43036 3782 43066 3834
rect 43066 3782 43078 3834
rect 43078 3782 43092 3834
rect 43116 3782 43130 3834
rect 43130 3782 43142 3834
rect 43142 3782 43172 3834
rect 43196 3782 43206 3834
rect 43206 3782 43252 3834
rect 42956 3780 43012 3782
rect 43036 3780 43092 3782
rect 43116 3780 43172 3782
rect 43196 3780 43252 3782
rect 42956 2746 43012 2748
rect 43036 2746 43092 2748
rect 43116 2746 43172 2748
rect 43196 2746 43252 2748
rect 42956 2694 43002 2746
rect 43002 2694 43012 2746
rect 43036 2694 43066 2746
rect 43066 2694 43078 2746
rect 43078 2694 43092 2746
rect 43116 2694 43130 2746
rect 43130 2694 43142 2746
rect 43142 2694 43172 2746
rect 43196 2694 43206 2746
rect 43206 2694 43252 2746
rect 42956 2692 43012 2694
rect 43036 2692 43092 2694
rect 43116 2692 43172 2694
rect 43196 2692 43252 2694
rect 47956 9818 48012 9820
rect 48036 9818 48092 9820
rect 48116 9818 48172 9820
rect 48196 9818 48252 9820
rect 47956 9766 48002 9818
rect 48002 9766 48012 9818
rect 48036 9766 48066 9818
rect 48066 9766 48078 9818
rect 48078 9766 48092 9818
rect 48116 9766 48130 9818
rect 48130 9766 48142 9818
rect 48142 9766 48172 9818
rect 48196 9766 48206 9818
rect 48206 9766 48252 9818
rect 47956 9764 48012 9766
rect 48036 9764 48092 9766
rect 48116 9764 48172 9766
rect 48196 9764 48252 9766
rect 47306 9560 47362 9616
rect 49146 9152 49202 9208
rect 47956 8730 48012 8732
rect 48036 8730 48092 8732
rect 48116 8730 48172 8732
rect 48196 8730 48252 8732
rect 47956 8678 48002 8730
rect 48002 8678 48012 8730
rect 48036 8678 48066 8730
rect 48066 8678 48078 8730
rect 48078 8678 48092 8730
rect 48116 8678 48130 8730
rect 48130 8678 48142 8730
rect 48142 8678 48172 8730
rect 48196 8678 48206 8730
rect 48206 8678 48252 8730
rect 47956 8676 48012 8678
rect 48036 8676 48092 8678
rect 48116 8676 48172 8678
rect 48196 8676 48252 8678
rect 46846 2624 46902 2680
rect 49238 8744 49294 8800
rect 49330 8336 49386 8392
rect 47956 7642 48012 7644
rect 48036 7642 48092 7644
rect 48116 7642 48172 7644
rect 48196 7642 48252 7644
rect 47956 7590 48002 7642
rect 48002 7590 48012 7642
rect 48036 7590 48066 7642
rect 48066 7590 48078 7642
rect 48078 7590 48092 7642
rect 48116 7590 48130 7642
rect 48130 7590 48142 7642
rect 48142 7590 48172 7642
rect 48196 7590 48206 7642
rect 48206 7590 48252 7642
rect 47956 7588 48012 7590
rect 48036 7588 48092 7590
rect 48116 7588 48172 7590
rect 48196 7588 48252 7590
rect 49146 7520 49202 7576
rect 49238 7112 49294 7168
rect 47956 6554 48012 6556
rect 48036 6554 48092 6556
rect 48116 6554 48172 6556
rect 48196 6554 48252 6556
rect 47956 6502 48002 6554
rect 48002 6502 48012 6554
rect 48036 6502 48066 6554
rect 48066 6502 48078 6554
rect 48078 6502 48092 6554
rect 48116 6502 48130 6554
rect 48130 6502 48142 6554
rect 48142 6502 48172 6554
rect 48196 6502 48206 6554
rect 48206 6502 48252 6554
rect 47956 6500 48012 6502
rect 48036 6500 48092 6502
rect 48116 6500 48172 6502
rect 48196 6500 48252 6502
rect 49422 6704 49478 6760
rect 48870 6296 48926 6352
rect 49146 5888 49202 5944
rect 47956 5466 48012 5468
rect 48036 5466 48092 5468
rect 48116 5466 48172 5468
rect 48196 5466 48252 5468
rect 47956 5414 48002 5466
rect 48002 5414 48012 5466
rect 48036 5414 48066 5466
rect 48066 5414 48078 5466
rect 48078 5414 48092 5466
rect 48116 5414 48130 5466
rect 48130 5414 48142 5466
rect 48142 5414 48172 5466
rect 48196 5414 48206 5466
rect 48206 5414 48252 5466
rect 47956 5412 48012 5414
rect 48036 5412 48092 5414
rect 48116 5412 48172 5414
rect 48196 5412 48252 5414
rect 49422 5480 49478 5536
rect 49330 5072 49386 5128
rect 48318 4664 48374 4720
rect 47956 4378 48012 4380
rect 48036 4378 48092 4380
rect 48116 4378 48172 4380
rect 48196 4378 48252 4380
rect 47956 4326 48002 4378
rect 48002 4326 48012 4378
rect 48036 4326 48066 4378
rect 48066 4326 48078 4378
rect 48078 4326 48092 4378
rect 48116 4326 48130 4378
rect 48130 4326 48142 4378
rect 48142 4326 48172 4378
rect 48196 4326 48206 4378
rect 48206 4326 48252 4378
rect 47956 4324 48012 4326
rect 48036 4324 48092 4326
rect 48116 4324 48172 4326
rect 48196 4324 48252 4326
rect 49146 4256 49202 4312
rect 46754 1808 46810 1864
rect 46662 1400 46718 1456
rect 49238 3848 49294 3904
rect 49146 3440 49202 3496
rect 47956 3290 48012 3292
rect 48036 3290 48092 3292
rect 48116 3290 48172 3292
rect 48196 3290 48252 3292
rect 47956 3238 48002 3290
rect 48002 3238 48012 3290
rect 48036 3238 48066 3290
rect 48066 3238 48078 3290
rect 48078 3238 48092 3290
rect 48116 3238 48130 3290
rect 48130 3238 48142 3290
rect 48142 3238 48172 3290
rect 48196 3238 48206 3290
rect 48206 3238 48252 3290
rect 47956 3236 48012 3238
rect 48036 3236 48092 3238
rect 48116 3236 48172 3238
rect 48196 3236 48252 3238
rect 48686 3032 48742 3088
rect 48502 2216 48558 2272
rect 47956 2202 48012 2204
rect 48036 2202 48092 2204
rect 48116 2202 48172 2204
rect 48196 2202 48252 2204
rect 47956 2150 48002 2202
rect 48002 2150 48012 2202
rect 48036 2150 48066 2202
rect 48066 2150 48078 2202
rect 48078 2150 48092 2202
rect 48116 2150 48130 2202
rect 48130 2150 48142 2202
rect 48142 2150 48172 2202
rect 48196 2150 48206 2202
rect 48206 2150 48252 2202
rect 47956 2148 48012 2150
rect 48036 2148 48092 2150
rect 48116 2148 48172 2150
rect 48196 2148 48252 2150
<< metal3 >>
rect 0 25666 800 25696
rect 3417 25666 3483 25669
rect 0 25664 3483 25666
rect 0 25608 3422 25664
rect 3478 25608 3483 25664
rect 0 25606 3483 25608
rect 0 25576 800 25606
rect 3417 25603 3483 25606
rect 48221 25530 48287 25533
rect 50200 25530 51000 25560
rect 48221 25528 51000 25530
rect 48221 25472 48226 25528
rect 48282 25472 51000 25528
rect 48221 25470 51000 25472
rect 48221 25467 48287 25470
rect 50200 25440 51000 25470
rect 0 25258 800 25288
rect 4061 25258 4127 25261
rect 0 25256 4127 25258
rect 0 25200 4066 25256
rect 4122 25200 4127 25256
rect 0 25198 4127 25200
rect 0 25168 800 25198
rect 4061 25195 4127 25198
rect 46657 25122 46723 25125
rect 50200 25122 51000 25152
rect 46657 25120 51000 25122
rect 46657 25064 46662 25120
rect 46718 25064 51000 25120
rect 46657 25062 51000 25064
rect 46657 25059 46723 25062
rect 50200 25032 51000 25062
rect 0 24850 800 24880
rect 3877 24850 3943 24853
rect 0 24848 3943 24850
rect 0 24792 3882 24848
rect 3938 24792 3943 24848
rect 0 24790 3943 24792
rect 0 24760 800 24790
rect 3877 24787 3943 24790
rect 34881 24714 34947 24717
rect 44541 24714 44607 24717
rect 34881 24712 44607 24714
rect 34881 24656 34886 24712
rect 34942 24656 44546 24712
rect 44602 24656 44607 24712
rect 34881 24654 44607 24656
rect 34881 24651 34947 24654
rect 44541 24651 44607 24654
rect 46565 24714 46631 24717
rect 50200 24714 51000 24744
rect 46565 24712 51000 24714
rect 46565 24656 46570 24712
rect 46626 24656 51000 24712
rect 46565 24654 51000 24656
rect 46565 24651 46631 24654
rect 50200 24624 51000 24654
rect 2946 24512 3262 24513
rect 0 24442 800 24472
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 32946 24512 33262 24513
rect 32946 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33262 24512
rect 32946 24447 33262 24448
rect 42946 24512 43262 24513
rect 42946 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43262 24512
rect 42946 24447 43262 24448
rect 2773 24442 2839 24445
rect 0 24440 2839 24442
rect 0 24384 2778 24440
rect 2834 24384 2839 24440
rect 0 24382 2839 24384
rect 0 24352 800 24382
rect 2773 24379 2839 24382
rect 30097 24442 30163 24445
rect 32397 24442 32463 24445
rect 30097 24440 32463 24442
rect 30097 24384 30102 24440
rect 30158 24384 32402 24440
rect 32458 24384 32463 24440
rect 30097 24382 32463 24384
rect 30097 24379 30163 24382
rect 32397 24379 32463 24382
rect 33777 24442 33843 24445
rect 40677 24442 40743 24445
rect 33777 24440 40743 24442
rect 33777 24384 33782 24440
rect 33838 24384 40682 24440
rect 40738 24384 40743 24440
rect 33777 24382 40743 24384
rect 33777 24379 33843 24382
rect 40677 24379 40743 24382
rect 7373 24306 7439 24309
rect 25957 24306 26023 24309
rect 7373 24304 26023 24306
rect 7373 24248 7378 24304
rect 7434 24248 25962 24304
rect 26018 24248 26023 24304
rect 7373 24246 26023 24248
rect 7373 24243 7439 24246
rect 25957 24243 26023 24246
rect 30005 24306 30071 24309
rect 40953 24306 41019 24309
rect 30005 24304 41019 24306
rect 30005 24248 30010 24304
rect 30066 24248 40958 24304
rect 41014 24248 41019 24304
rect 30005 24246 41019 24248
rect 30005 24243 30071 24246
rect 40953 24243 41019 24246
rect 47577 24306 47643 24309
rect 50200 24306 51000 24336
rect 47577 24304 51000 24306
rect 47577 24248 47582 24304
rect 47638 24248 51000 24304
rect 47577 24246 51000 24248
rect 47577 24243 47643 24246
rect 50200 24216 51000 24246
rect 26141 24170 26207 24173
rect 48773 24170 48839 24173
rect 26141 24168 48839 24170
rect 26141 24112 26146 24168
rect 26202 24112 48778 24168
rect 48834 24112 48839 24168
rect 26141 24110 48839 24112
rect 26141 24107 26207 24110
rect 48773 24107 48839 24110
rect 0 24034 800 24064
rect 3785 24034 3851 24037
rect 0 24032 3851 24034
rect 0 23976 3790 24032
rect 3846 23976 3851 24032
rect 0 23974 3851 23976
rect 0 23944 800 23974
rect 3785 23971 3851 23974
rect 19333 24034 19399 24037
rect 27337 24034 27403 24037
rect 19333 24032 27403 24034
rect 19333 23976 19338 24032
rect 19394 23976 27342 24032
rect 27398 23976 27403 24032
rect 19333 23974 27403 23976
rect 19333 23971 19399 23974
rect 27337 23971 27403 23974
rect 28942 23972 28948 24036
rect 29012 24034 29018 24036
rect 35249 24034 35315 24037
rect 37641 24034 37707 24037
rect 29012 24032 37707 24034
rect 29012 23976 35254 24032
rect 35310 23976 37646 24032
rect 37702 23976 37707 24032
rect 29012 23974 37707 23976
rect 29012 23972 29018 23974
rect 35249 23971 35315 23974
rect 37641 23971 37707 23974
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 17946 23903 18262 23904
rect 27946 23968 28262 23969
rect 27946 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28262 23968
rect 27946 23903 28262 23904
rect 37946 23968 38262 23969
rect 37946 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38262 23968
rect 37946 23903 38262 23904
rect 47946 23968 48262 23969
rect 47946 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48262 23968
rect 47946 23903 48262 23904
rect 38469 23898 38535 23901
rect 42241 23898 42307 23901
rect 38469 23896 42307 23898
rect 38469 23840 38474 23896
rect 38530 23840 42246 23896
rect 42302 23840 42307 23896
rect 38469 23838 42307 23840
rect 38469 23835 38535 23838
rect 42241 23835 42307 23838
rect 48405 23898 48471 23901
rect 50200 23898 51000 23928
rect 48405 23896 51000 23898
rect 48405 23840 48410 23896
rect 48466 23840 51000 23896
rect 48405 23838 51000 23840
rect 48405 23835 48471 23838
rect 50200 23808 51000 23838
rect 36997 23762 37063 23765
rect 45369 23762 45435 23765
rect 36997 23760 45435 23762
rect 36997 23704 37002 23760
rect 37058 23704 45374 23760
rect 45430 23704 45435 23760
rect 36997 23702 45435 23704
rect 36997 23699 37063 23702
rect 45369 23699 45435 23702
rect 0 23626 800 23656
rect 4061 23626 4127 23629
rect 0 23624 4127 23626
rect 0 23568 4066 23624
rect 4122 23568 4127 23624
rect 0 23566 4127 23568
rect 0 23536 800 23566
rect 4061 23563 4127 23566
rect 31017 23626 31083 23629
rect 45185 23626 45251 23629
rect 31017 23624 45251 23626
rect 31017 23568 31022 23624
rect 31078 23568 45190 23624
rect 45246 23568 45251 23624
rect 31017 23566 45251 23568
rect 31017 23563 31083 23566
rect 45185 23563 45251 23566
rect 24669 23490 24735 23493
rect 26325 23490 26391 23493
rect 24669 23488 26391 23490
rect 24669 23432 24674 23488
rect 24730 23432 26330 23488
rect 26386 23432 26391 23488
rect 24669 23430 26391 23432
rect 24669 23427 24735 23430
rect 26325 23427 26391 23430
rect 33961 23490 34027 23493
rect 35525 23490 35591 23493
rect 38837 23490 38903 23493
rect 33961 23488 38903 23490
rect 33961 23432 33966 23488
rect 34022 23432 35530 23488
rect 35586 23432 38842 23488
rect 38898 23432 38903 23488
rect 33961 23430 38903 23432
rect 33961 23427 34027 23430
rect 35525 23427 35591 23430
rect 38837 23427 38903 23430
rect 47853 23490 47919 23493
rect 50200 23490 51000 23520
rect 47853 23488 51000 23490
rect 47853 23432 47858 23488
rect 47914 23432 51000 23488
rect 47853 23430 51000 23432
rect 47853 23427 47919 23430
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 32946 23424 33262 23425
rect 32946 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33262 23424
rect 32946 23359 33262 23360
rect 42946 23424 43262 23425
rect 42946 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43262 23424
rect 50200 23400 51000 23430
rect 42946 23359 43262 23360
rect 35709 23354 35775 23357
rect 42609 23354 42675 23357
rect 35709 23352 42675 23354
rect 35709 23296 35714 23352
rect 35770 23296 42614 23352
rect 42670 23296 42675 23352
rect 35709 23294 42675 23296
rect 35709 23291 35775 23294
rect 42609 23291 42675 23294
rect 0 23218 800 23248
rect 4061 23218 4127 23221
rect 0 23216 4127 23218
rect 0 23160 4066 23216
rect 4122 23160 4127 23216
rect 0 23158 4127 23160
rect 0 23128 800 23158
rect 4061 23155 4127 23158
rect 30189 23218 30255 23221
rect 35893 23218 35959 23221
rect 30189 23216 35959 23218
rect 30189 23160 30194 23216
rect 30250 23160 35898 23216
rect 35954 23160 35959 23216
rect 30189 23158 35959 23160
rect 30189 23155 30255 23158
rect 35893 23155 35959 23158
rect 36721 23218 36787 23221
rect 43897 23218 43963 23221
rect 36721 23216 43963 23218
rect 36721 23160 36726 23216
rect 36782 23160 43902 23216
rect 43958 23160 43963 23216
rect 36721 23158 43963 23160
rect 36721 23155 36787 23158
rect 43897 23155 43963 23158
rect 24669 23082 24735 23085
rect 31477 23082 31543 23085
rect 24669 23080 31543 23082
rect 24669 23024 24674 23080
rect 24730 23024 31482 23080
rect 31538 23024 31543 23080
rect 24669 23022 31543 23024
rect 24669 23019 24735 23022
rect 31477 23019 31543 23022
rect 39389 23082 39455 23085
rect 43529 23082 43595 23085
rect 39389 23080 43595 23082
rect 39389 23024 39394 23080
rect 39450 23024 43534 23080
rect 43590 23024 43595 23080
rect 39389 23022 43595 23024
rect 39389 23019 39455 23022
rect 43529 23019 43595 23022
rect 48313 23082 48379 23085
rect 50200 23082 51000 23112
rect 48313 23080 51000 23082
rect 48313 23024 48318 23080
rect 48374 23024 51000 23080
rect 48313 23022 51000 23024
rect 48313 23019 48379 23022
rect 50200 22992 51000 23022
rect 32581 22946 32647 22949
rect 36445 22946 36511 22949
rect 32581 22944 36511 22946
rect 32581 22888 32586 22944
rect 32642 22888 36450 22944
rect 36506 22888 36511 22944
rect 32581 22886 36511 22888
rect 32581 22883 32647 22886
rect 36445 22883 36511 22886
rect 7946 22880 8262 22881
rect 0 22810 800 22840
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 27946 22880 28262 22881
rect 27946 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28262 22880
rect 27946 22815 28262 22816
rect 37946 22880 38262 22881
rect 37946 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38262 22880
rect 37946 22815 38262 22816
rect 47946 22880 48262 22881
rect 47946 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48262 22880
rect 47946 22815 48262 22816
rect 3969 22810 4035 22813
rect 0 22808 4035 22810
rect 0 22752 3974 22808
rect 4030 22752 4035 22808
rect 0 22750 4035 22752
rect 0 22720 800 22750
rect 3969 22747 4035 22750
rect 30741 22810 30807 22813
rect 34881 22810 34947 22813
rect 30741 22808 34947 22810
rect 30741 22752 30746 22808
rect 30802 22752 34886 22808
rect 34942 22752 34947 22808
rect 30741 22750 34947 22752
rect 30741 22747 30807 22750
rect 34881 22747 34947 22750
rect 42149 22810 42215 22813
rect 47117 22810 47183 22813
rect 42149 22808 47183 22810
rect 42149 22752 42154 22808
rect 42210 22752 47122 22808
rect 47178 22752 47183 22808
rect 42149 22750 47183 22752
rect 42149 22747 42215 22750
rect 47117 22747 47183 22750
rect 31477 22674 31543 22677
rect 33961 22674 34027 22677
rect 31477 22672 34027 22674
rect 31477 22616 31482 22672
rect 31538 22616 33966 22672
rect 34022 22616 34027 22672
rect 31477 22614 34027 22616
rect 31477 22611 31543 22614
rect 33961 22611 34027 22614
rect 49325 22674 49391 22677
rect 50200 22674 51000 22704
rect 49325 22672 51000 22674
rect 49325 22616 49330 22672
rect 49386 22616 51000 22672
rect 49325 22614 51000 22616
rect 49325 22611 49391 22614
rect 50200 22584 51000 22614
rect 4061 22538 4127 22541
rect 2454 22536 4127 22538
rect 2454 22480 4066 22536
rect 4122 22480 4127 22536
rect 2454 22478 4127 22480
rect 0 22402 800 22432
rect 2454 22402 2514 22478
rect 4061 22475 4127 22478
rect 14457 22538 14523 22541
rect 24025 22538 24091 22541
rect 25589 22538 25655 22541
rect 14457 22536 25655 22538
rect 14457 22480 14462 22536
rect 14518 22480 24030 22536
rect 24086 22480 25594 22536
rect 25650 22480 25655 22536
rect 14457 22478 25655 22480
rect 14457 22475 14523 22478
rect 24025 22475 24091 22478
rect 25589 22475 25655 22478
rect 34237 22538 34303 22541
rect 37733 22538 37799 22541
rect 40769 22538 40835 22541
rect 42609 22538 42675 22541
rect 34237 22536 40835 22538
rect 34237 22480 34242 22536
rect 34298 22480 37738 22536
rect 37794 22480 40774 22536
rect 40830 22480 40835 22536
rect 34237 22478 40835 22480
rect 34237 22475 34303 22478
rect 37733 22475 37799 22478
rect 40769 22475 40835 22478
rect 41370 22536 42675 22538
rect 41370 22480 42614 22536
rect 42670 22480 42675 22536
rect 41370 22478 42675 22480
rect 0 22342 2514 22402
rect 35433 22402 35499 22405
rect 41370 22402 41430 22478
rect 42609 22475 42675 22478
rect 35433 22400 41430 22402
rect 35433 22344 35438 22400
rect 35494 22344 41430 22400
rect 35433 22342 41430 22344
rect 0 22312 800 22342
rect 35433 22339 35499 22342
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 22946 22271 23262 22272
rect 32946 22336 33262 22337
rect 32946 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33262 22336
rect 32946 22271 33262 22272
rect 42946 22336 43262 22337
rect 42946 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43262 22336
rect 42946 22271 43262 22272
rect 49049 22266 49115 22269
rect 50200 22266 51000 22296
rect 49049 22264 51000 22266
rect 49049 22208 49054 22264
rect 49110 22208 51000 22264
rect 49049 22206 51000 22208
rect 49049 22203 49115 22206
rect 50200 22176 51000 22206
rect 18413 22130 18479 22133
rect 18689 22130 18755 22133
rect 18413 22128 18755 22130
rect 18413 22072 18418 22128
rect 18474 22072 18694 22128
rect 18750 22072 18755 22128
rect 18413 22070 18755 22072
rect 18413 22067 18479 22070
rect 18689 22067 18755 22070
rect 21173 22130 21239 22133
rect 21633 22130 21699 22133
rect 25129 22130 25195 22133
rect 21173 22128 25195 22130
rect 21173 22072 21178 22128
rect 21234 22072 21638 22128
rect 21694 22072 25134 22128
rect 25190 22072 25195 22128
rect 21173 22070 25195 22072
rect 21173 22067 21239 22070
rect 21633 22067 21699 22070
rect 25129 22067 25195 22070
rect 27245 22130 27311 22133
rect 30005 22130 30071 22133
rect 27245 22128 30071 22130
rect 27245 22072 27250 22128
rect 27306 22072 30010 22128
rect 30066 22072 30071 22128
rect 27245 22070 30071 22072
rect 27245 22067 27311 22070
rect 30005 22067 30071 22070
rect 31385 22130 31451 22133
rect 35617 22130 35683 22133
rect 39389 22130 39455 22133
rect 31385 22128 39455 22130
rect 31385 22072 31390 22128
rect 31446 22072 35622 22128
rect 35678 22072 39394 22128
rect 39450 22072 39455 22128
rect 31385 22070 39455 22072
rect 31385 22067 31451 22070
rect 35617 22067 35683 22070
rect 39389 22067 39455 22070
rect 41321 22130 41387 22133
rect 41873 22130 41939 22133
rect 41321 22128 41939 22130
rect 41321 22072 41326 22128
rect 41382 22072 41878 22128
rect 41934 22072 41939 22128
rect 41321 22070 41939 22072
rect 41321 22067 41387 22070
rect 41873 22067 41939 22070
rect 0 21994 800 22024
rect 3877 21994 3943 21997
rect 0 21992 3943 21994
rect 0 21936 3882 21992
rect 3938 21936 3943 21992
rect 0 21934 3943 21936
rect 0 21904 800 21934
rect 3877 21931 3943 21934
rect 16205 21994 16271 21997
rect 18873 21994 18939 21997
rect 22737 21994 22803 21997
rect 16205 21992 22803 21994
rect 16205 21936 16210 21992
rect 16266 21936 18878 21992
rect 18934 21936 22742 21992
rect 22798 21936 22803 21992
rect 16205 21934 22803 21936
rect 16205 21931 16271 21934
rect 18873 21931 18939 21934
rect 22737 21931 22803 21934
rect 25773 21994 25839 21997
rect 33041 21994 33107 21997
rect 25773 21992 33107 21994
rect 25773 21936 25778 21992
rect 25834 21936 33046 21992
rect 33102 21936 33107 21992
rect 25773 21934 33107 21936
rect 25773 21931 25839 21934
rect 33041 21931 33107 21934
rect 37181 21994 37247 21997
rect 41689 21994 41755 21997
rect 37181 21992 41755 21994
rect 37181 21936 37186 21992
rect 37242 21936 41694 21992
rect 41750 21936 41755 21992
rect 37181 21934 41755 21936
rect 37181 21931 37247 21934
rect 41689 21931 41755 21934
rect 21265 21858 21331 21861
rect 23197 21858 23263 21861
rect 21265 21856 23263 21858
rect 21265 21800 21270 21856
rect 21326 21800 23202 21856
rect 23258 21800 23263 21856
rect 21265 21798 23263 21800
rect 21265 21795 21331 21798
rect 23197 21795 23263 21798
rect 48773 21858 48839 21861
rect 50200 21858 51000 21888
rect 48773 21856 51000 21858
rect 48773 21800 48778 21856
rect 48834 21800 51000 21856
rect 48773 21798 51000 21800
rect 48773 21795 48839 21798
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 27946 21792 28262 21793
rect 27946 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28262 21792
rect 27946 21727 28262 21728
rect 37946 21792 38262 21793
rect 37946 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38262 21792
rect 37946 21727 38262 21728
rect 47946 21792 48262 21793
rect 47946 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48262 21792
rect 50200 21768 51000 21798
rect 47946 21727 48262 21728
rect 19333 21722 19399 21725
rect 30649 21722 30715 21725
rect 34789 21722 34855 21725
rect 19333 21720 27860 21722
rect 19333 21664 19338 21720
rect 19394 21664 27860 21720
rect 19333 21662 27860 21664
rect 19333 21659 19399 21662
rect 0 21586 800 21616
rect 2681 21586 2747 21589
rect 0 21584 2747 21586
rect 0 21528 2686 21584
rect 2742 21528 2747 21584
rect 0 21526 2747 21528
rect 0 21496 800 21526
rect 2681 21523 2747 21526
rect 16665 21586 16731 21589
rect 22829 21586 22895 21589
rect 16665 21584 22895 21586
rect 16665 21528 16670 21584
rect 16726 21528 22834 21584
rect 22890 21528 22895 21584
rect 16665 21526 22895 21528
rect 27800 21586 27860 21662
rect 30649 21720 34855 21722
rect 30649 21664 30654 21720
rect 30710 21664 34794 21720
rect 34850 21664 34855 21720
rect 30649 21662 34855 21664
rect 30649 21659 30715 21662
rect 34789 21659 34855 21662
rect 28809 21586 28875 21589
rect 27800 21584 28875 21586
rect 27800 21528 28814 21584
rect 28870 21528 28875 21584
rect 27800 21526 28875 21528
rect 16665 21523 16731 21526
rect 22829 21523 22895 21526
rect 28809 21523 28875 21526
rect 31201 21586 31267 21589
rect 33685 21586 33751 21589
rect 42793 21586 42859 21589
rect 31201 21584 42859 21586
rect 31201 21528 31206 21584
rect 31262 21528 33690 21584
rect 33746 21528 42798 21584
rect 42854 21528 42859 21584
rect 31201 21526 42859 21528
rect 31201 21523 31267 21526
rect 33685 21523 33751 21526
rect 42793 21523 42859 21526
rect 5901 21450 5967 21453
rect 8753 21450 8819 21453
rect 5901 21448 8819 21450
rect 5901 21392 5906 21448
rect 5962 21392 8758 21448
rect 8814 21392 8819 21448
rect 5901 21390 8819 21392
rect 5901 21387 5967 21390
rect 8753 21387 8819 21390
rect 11329 21450 11395 21453
rect 25221 21450 25287 21453
rect 26141 21450 26207 21453
rect 11329 21448 26207 21450
rect 11329 21392 11334 21448
rect 11390 21392 25226 21448
rect 25282 21392 26146 21448
rect 26202 21392 26207 21448
rect 11329 21390 26207 21392
rect 11329 21387 11395 21390
rect 25221 21387 25287 21390
rect 26141 21387 26207 21390
rect 27429 21450 27495 21453
rect 29637 21450 29703 21453
rect 27429 21448 29703 21450
rect 27429 21392 27434 21448
rect 27490 21392 29642 21448
rect 29698 21392 29703 21448
rect 27429 21390 29703 21392
rect 27429 21387 27495 21390
rect 29637 21387 29703 21390
rect 34789 21450 34855 21453
rect 41413 21450 41479 21453
rect 34789 21448 41479 21450
rect 34789 21392 34794 21448
rect 34850 21392 41418 21448
rect 41474 21392 41479 21448
rect 34789 21390 41479 21392
rect 34789 21387 34855 21390
rect 41413 21387 41479 21390
rect 49141 21450 49207 21453
rect 50200 21450 51000 21480
rect 49141 21448 51000 21450
rect 49141 21392 49146 21448
rect 49202 21392 51000 21448
rect 49141 21390 51000 21392
rect 49141 21387 49207 21390
rect 50200 21360 51000 21390
rect 33593 21314 33659 21317
rect 41505 21314 41571 21317
rect 33593 21312 41571 21314
rect 33593 21256 33598 21312
rect 33654 21256 41510 21312
rect 41566 21256 41571 21312
rect 33593 21254 41571 21256
rect 33593 21251 33659 21254
rect 41505 21251 41571 21254
rect 2946 21248 3262 21249
rect 0 21178 800 21208
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 32946 21248 33262 21249
rect 32946 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33262 21248
rect 32946 21183 33262 21184
rect 42946 21248 43262 21249
rect 42946 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43262 21248
rect 42946 21183 43262 21184
rect 2773 21178 2839 21181
rect 0 21176 2839 21178
rect 0 21120 2778 21176
rect 2834 21120 2839 21176
rect 0 21118 2839 21120
rect 0 21088 800 21118
rect 2773 21115 2839 21118
rect 16573 21178 16639 21181
rect 17125 21178 17191 21181
rect 23473 21178 23539 21181
rect 26693 21178 26759 21181
rect 16573 21176 22110 21178
rect 16573 21120 16578 21176
rect 16634 21120 17130 21176
rect 17186 21120 22110 21176
rect 16573 21118 22110 21120
rect 16573 21115 16639 21118
rect 17125 21115 17191 21118
rect 11329 21042 11395 21045
rect 19241 21042 19307 21045
rect 11329 21040 19307 21042
rect 11329 20984 11334 21040
rect 11390 20984 19246 21040
rect 19302 20984 19307 21040
rect 11329 20982 19307 20984
rect 11329 20979 11395 20982
rect 19241 20979 19307 20982
rect 21081 21042 21147 21045
rect 21541 21042 21607 21045
rect 21081 21040 21607 21042
rect 21081 20984 21086 21040
rect 21142 20984 21546 21040
rect 21602 20984 21607 21040
rect 21081 20982 21607 20984
rect 22050 21042 22110 21118
rect 23473 21176 26759 21178
rect 23473 21120 23478 21176
rect 23534 21120 26698 21176
rect 26754 21120 26759 21176
rect 23473 21118 26759 21120
rect 23473 21115 23539 21118
rect 26693 21115 26759 21118
rect 27337 21178 27403 21181
rect 30833 21178 30899 21181
rect 27337 21176 30899 21178
rect 27337 21120 27342 21176
rect 27398 21120 30838 21176
rect 30894 21120 30899 21176
rect 27337 21118 30899 21120
rect 27337 21115 27403 21118
rect 30833 21115 30899 21118
rect 35893 21178 35959 21181
rect 40309 21178 40375 21181
rect 35893 21176 40375 21178
rect 35893 21120 35898 21176
rect 35954 21120 40314 21176
rect 40370 21120 40375 21176
rect 35893 21118 40375 21120
rect 35893 21115 35959 21118
rect 40309 21115 40375 21118
rect 24853 21042 24919 21045
rect 22050 21040 24919 21042
rect 22050 20984 24858 21040
rect 24914 20984 24919 21040
rect 22050 20982 24919 20984
rect 21081 20979 21147 20982
rect 21541 20979 21607 20982
rect 24853 20979 24919 20982
rect 26877 21042 26943 21045
rect 28758 21042 28764 21044
rect 26877 21040 28764 21042
rect 26877 20984 26882 21040
rect 26938 20984 28764 21040
rect 26877 20982 28764 20984
rect 26877 20979 26943 20982
rect 28758 20980 28764 20982
rect 28828 20980 28834 21044
rect 32489 21042 32555 21045
rect 40861 21042 40927 21045
rect 32489 21040 40927 21042
rect 32489 20984 32494 21040
rect 32550 20984 40866 21040
rect 40922 20984 40927 21040
rect 32489 20982 40927 20984
rect 32489 20979 32555 20982
rect 40861 20979 40927 20982
rect 49049 21042 49115 21045
rect 50200 21042 51000 21072
rect 49049 21040 51000 21042
rect 49049 20984 49054 21040
rect 49110 20984 51000 21040
rect 49049 20982 51000 20984
rect 49049 20979 49115 20982
rect 50200 20952 51000 20982
rect 19701 20906 19767 20909
rect 29729 20906 29795 20909
rect 19701 20904 29795 20906
rect 19701 20848 19706 20904
rect 19762 20848 29734 20904
rect 29790 20848 29795 20904
rect 19701 20846 29795 20848
rect 19701 20843 19767 20846
rect 29729 20843 29795 20846
rect 32397 20906 32463 20909
rect 40953 20906 41019 20909
rect 32397 20904 41019 20906
rect 32397 20848 32402 20904
rect 32458 20848 40958 20904
rect 41014 20848 41019 20904
rect 32397 20846 41019 20848
rect 32397 20843 32463 20846
rect 40953 20843 41019 20846
rect 0 20770 800 20800
rect 1301 20770 1367 20773
rect 0 20768 1367 20770
rect 0 20712 1306 20768
rect 1362 20712 1367 20768
rect 0 20710 1367 20712
rect 0 20680 800 20710
rect 1301 20707 1367 20710
rect 28441 20770 28507 20773
rect 28717 20770 28783 20773
rect 28441 20768 28783 20770
rect 28441 20712 28446 20768
rect 28502 20712 28722 20768
rect 28778 20712 28783 20768
rect 28441 20710 28783 20712
rect 28441 20707 28507 20710
rect 28717 20707 28783 20710
rect 30189 20770 30255 20773
rect 37089 20770 37155 20773
rect 30189 20768 37155 20770
rect 30189 20712 30194 20768
rect 30250 20712 37094 20768
rect 37150 20712 37155 20768
rect 30189 20710 37155 20712
rect 30189 20707 30255 20710
rect 37089 20707 37155 20710
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 17946 20639 18262 20640
rect 27946 20704 28262 20705
rect 27946 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28262 20704
rect 27946 20639 28262 20640
rect 37946 20704 38262 20705
rect 37946 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38262 20704
rect 37946 20639 38262 20640
rect 47946 20704 48262 20705
rect 47946 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48262 20704
rect 47946 20639 48262 20640
rect 19977 20634 20043 20637
rect 21909 20634 21975 20637
rect 25313 20634 25379 20637
rect 19977 20632 25379 20634
rect 19977 20576 19982 20632
rect 20038 20576 21914 20632
rect 21970 20576 25318 20632
rect 25374 20576 25379 20632
rect 19977 20574 25379 20576
rect 19977 20571 20043 20574
rect 21909 20571 21975 20574
rect 25313 20571 25379 20574
rect 28574 20572 28580 20636
rect 28644 20634 28650 20636
rect 34421 20634 34487 20637
rect 28644 20632 34487 20634
rect 28644 20576 34426 20632
rect 34482 20576 34487 20632
rect 28644 20574 34487 20576
rect 28644 20572 28650 20574
rect 34421 20571 34487 20574
rect 34605 20634 34671 20637
rect 36629 20634 36695 20637
rect 34605 20632 36695 20634
rect 34605 20576 34610 20632
rect 34666 20576 36634 20632
rect 36690 20576 36695 20632
rect 34605 20574 36695 20576
rect 34605 20571 34671 20574
rect 36629 20571 36695 20574
rect 49049 20634 49115 20637
rect 50200 20634 51000 20664
rect 49049 20632 51000 20634
rect 49049 20576 49054 20632
rect 49110 20576 51000 20632
rect 49049 20574 51000 20576
rect 49049 20571 49115 20574
rect 50200 20544 51000 20574
rect 30833 20498 30899 20501
rect 39205 20498 39271 20501
rect 30833 20496 39271 20498
rect 30833 20440 30838 20496
rect 30894 20440 39210 20496
rect 39266 20440 39271 20496
rect 30833 20438 39271 20440
rect 30833 20435 30899 20438
rect 39205 20435 39271 20438
rect 0 20362 800 20392
rect 3877 20362 3943 20365
rect 0 20360 3943 20362
rect 0 20304 3882 20360
rect 3938 20304 3943 20360
rect 0 20302 3943 20304
rect 0 20272 800 20302
rect 3877 20299 3943 20302
rect 16757 20362 16823 20365
rect 30005 20362 30071 20365
rect 16757 20360 30071 20362
rect 16757 20304 16762 20360
rect 16818 20304 30010 20360
rect 30066 20304 30071 20360
rect 16757 20302 30071 20304
rect 16757 20299 16823 20302
rect 30005 20299 30071 20302
rect 31845 20362 31911 20365
rect 48313 20362 48379 20365
rect 31845 20360 48379 20362
rect 31845 20304 31850 20360
rect 31906 20304 48318 20360
rect 48374 20304 48379 20360
rect 31845 20302 48379 20304
rect 31845 20299 31911 20302
rect 48313 20299 48379 20302
rect 24117 20226 24183 20229
rect 28390 20226 28396 20228
rect 24117 20224 28396 20226
rect 24117 20168 24122 20224
rect 24178 20168 28396 20224
rect 24117 20166 28396 20168
rect 24117 20163 24183 20166
rect 28390 20164 28396 20166
rect 28460 20164 28466 20228
rect 28809 20224 28875 20229
rect 28809 20168 28814 20224
rect 28870 20168 28875 20224
rect 28809 20163 28875 20168
rect 48773 20226 48839 20229
rect 50200 20226 51000 20256
rect 48773 20224 51000 20226
rect 48773 20168 48778 20224
rect 48834 20168 51000 20224
rect 48773 20166 51000 20168
rect 48773 20163 48839 20166
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 23381 20090 23447 20093
rect 28812 20090 28872 20163
rect 32946 20160 33262 20161
rect 32946 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33262 20160
rect 32946 20095 33262 20096
rect 42946 20160 43262 20161
rect 42946 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43262 20160
rect 50200 20136 51000 20166
rect 42946 20095 43262 20096
rect 23381 20088 28872 20090
rect 23381 20032 23386 20088
rect 23442 20032 28872 20088
rect 23381 20030 28872 20032
rect 23381 20027 23447 20030
rect 0 19954 800 19984
rect 3325 19954 3391 19957
rect 0 19952 3391 19954
rect 0 19896 3330 19952
rect 3386 19896 3391 19952
rect 0 19894 3391 19896
rect 0 19864 800 19894
rect 3325 19891 3391 19894
rect 13353 19954 13419 19957
rect 21817 19954 21883 19957
rect 25865 19954 25931 19957
rect 40401 19954 40467 19957
rect 13353 19952 40467 19954
rect 13353 19896 13358 19952
rect 13414 19896 21822 19952
rect 21878 19896 25870 19952
rect 25926 19896 40406 19952
rect 40462 19896 40467 19952
rect 13353 19894 40467 19896
rect 13353 19891 13419 19894
rect 21817 19891 21883 19894
rect 25865 19891 25931 19894
rect 40401 19891 40467 19894
rect 10961 19818 11027 19821
rect 13629 19818 13695 19821
rect 10961 19816 13695 19818
rect 10961 19760 10966 19816
rect 11022 19760 13634 19816
rect 13690 19760 13695 19816
rect 10961 19758 13695 19760
rect 10961 19755 11027 19758
rect 13629 19755 13695 19758
rect 26049 19818 26115 19821
rect 34513 19818 34579 19821
rect 48497 19818 48563 19821
rect 26049 19816 29010 19818
rect 26049 19760 26054 19816
rect 26110 19760 29010 19816
rect 26049 19758 29010 19760
rect 26049 19755 26115 19758
rect 19333 19682 19399 19685
rect 26785 19682 26851 19685
rect 27705 19682 27771 19685
rect 28533 19684 28599 19685
rect 28533 19682 28580 19684
rect 19333 19680 27771 19682
rect 19333 19624 19338 19680
rect 19394 19624 26790 19680
rect 26846 19624 27710 19680
rect 27766 19624 27771 19680
rect 19333 19622 27771 19624
rect 28488 19680 28580 19682
rect 28488 19624 28538 19680
rect 28488 19622 28580 19624
rect 19333 19619 19399 19622
rect 26785 19619 26851 19622
rect 27705 19619 27771 19622
rect 28533 19620 28580 19622
rect 28644 19620 28650 19684
rect 28950 19682 29010 19758
rect 34513 19816 48563 19818
rect 34513 19760 34518 19816
rect 34574 19760 48502 19816
rect 48558 19760 48563 19816
rect 34513 19758 48563 19760
rect 34513 19755 34579 19758
rect 48497 19755 48563 19758
rect 49049 19818 49115 19821
rect 50200 19818 51000 19848
rect 49049 19816 51000 19818
rect 49049 19760 49054 19816
rect 49110 19760 51000 19816
rect 49049 19758 51000 19760
rect 49049 19755 49115 19758
rect 50200 19728 51000 19758
rect 29269 19682 29335 19685
rect 28950 19680 35450 19682
rect 28950 19624 29274 19680
rect 29330 19624 35450 19680
rect 28950 19622 35450 19624
rect 28533 19619 28599 19620
rect 29269 19619 29335 19622
rect 7946 19616 8262 19617
rect 0 19546 800 19576
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 27946 19616 28262 19617
rect 27946 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28262 19616
rect 27946 19551 28262 19552
rect 2681 19546 2747 19549
rect 0 19544 2747 19546
rect 0 19488 2686 19544
rect 2742 19488 2747 19544
rect 0 19486 2747 19488
rect 0 19456 800 19486
rect 2681 19483 2747 19486
rect 20345 19546 20411 19549
rect 25313 19546 25379 19549
rect 26141 19546 26207 19549
rect 28809 19548 28875 19549
rect 20345 19544 26207 19546
rect 20345 19488 20350 19544
rect 20406 19488 25318 19544
rect 25374 19488 26146 19544
rect 26202 19488 26207 19544
rect 20345 19486 26207 19488
rect 20345 19483 20411 19486
rect 25313 19483 25379 19486
rect 26141 19483 26207 19486
rect 28758 19484 28764 19548
rect 28828 19546 28875 19548
rect 28828 19544 28920 19546
rect 28870 19488 28920 19544
rect 28828 19486 28920 19488
rect 28828 19484 28875 19486
rect 28809 19483 28875 19484
rect 14089 19410 14155 19413
rect 15101 19410 15167 19413
rect 14089 19408 15167 19410
rect 14089 19352 14094 19408
rect 14150 19352 15106 19408
rect 15162 19352 15167 19408
rect 14089 19350 15167 19352
rect 14089 19347 14155 19350
rect 15101 19347 15167 19350
rect 15377 19410 15443 19413
rect 26601 19410 26667 19413
rect 33961 19410 34027 19413
rect 15377 19408 34027 19410
rect 15377 19352 15382 19408
rect 15438 19352 26606 19408
rect 26662 19352 33966 19408
rect 34022 19352 34027 19408
rect 15377 19350 34027 19352
rect 35390 19410 35450 19622
rect 37946 19616 38262 19617
rect 37946 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38262 19616
rect 37946 19551 38262 19552
rect 47946 19616 48262 19617
rect 47946 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48262 19616
rect 47946 19551 48262 19552
rect 35893 19546 35959 19549
rect 36537 19546 36603 19549
rect 35893 19544 36603 19546
rect 35893 19488 35898 19544
rect 35954 19488 36542 19544
rect 36598 19488 36603 19544
rect 35893 19486 36603 19488
rect 35893 19483 35959 19486
rect 36537 19483 36603 19486
rect 38377 19546 38443 19549
rect 46933 19546 46999 19549
rect 38377 19544 46999 19546
rect 38377 19488 38382 19544
rect 38438 19488 46938 19544
rect 46994 19488 46999 19544
rect 38377 19486 46999 19488
rect 38377 19483 38443 19486
rect 46933 19483 46999 19486
rect 38929 19410 38995 19413
rect 35390 19408 38995 19410
rect 35390 19352 38934 19408
rect 38990 19352 38995 19408
rect 35390 19350 38995 19352
rect 15377 19347 15443 19350
rect 26601 19347 26667 19350
rect 33961 19347 34027 19350
rect 38929 19347 38995 19350
rect 49325 19410 49391 19413
rect 50200 19410 51000 19440
rect 49325 19408 51000 19410
rect 49325 19352 49330 19408
rect 49386 19352 51000 19408
rect 49325 19350 51000 19352
rect 49325 19347 49391 19350
rect 50200 19320 51000 19350
rect 2957 19274 3023 19277
rect 1304 19272 3023 19274
rect 1304 19216 2962 19272
rect 3018 19216 3023 19272
rect 1304 19214 3023 19216
rect 0 19138 800 19168
rect 1304 19138 1364 19214
rect 2957 19211 3023 19214
rect 28390 19212 28396 19276
rect 28460 19274 28466 19276
rect 29177 19274 29243 19277
rect 28460 19272 29243 19274
rect 28460 19216 29182 19272
rect 29238 19216 29243 19272
rect 28460 19214 29243 19216
rect 28460 19212 28466 19214
rect 29177 19211 29243 19214
rect 35249 19274 35315 19277
rect 36905 19274 36971 19277
rect 38193 19274 38259 19277
rect 40585 19274 40651 19277
rect 35249 19272 37474 19274
rect 35249 19216 35254 19272
rect 35310 19216 36910 19272
rect 36966 19216 37474 19272
rect 35249 19214 37474 19216
rect 35249 19211 35315 19214
rect 36905 19211 36971 19214
rect 0 19078 1364 19138
rect 26049 19138 26115 19141
rect 28625 19138 28691 19141
rect 26049 19136 28691 19138
rect 26049 19080 26054 19136
rect 26110 19080 28630 19136
rect 28686 19080 28691 19136
rect 26049 19078 28691 19080
rect 37414 19138 37474 19214
rect 38193 19272 40651 19274
rect 38193 19216 38198 19272
rect 38254 19216 40590 19272
rect 40646 19216 40651 19272
rect 38193 19214 40651 19216
rect 38193 19211 38259 19214
rect 40585 19211 40651 19214
rect 40401 19138 40467 19141
rect 37414 19136 40467 19138
rect 37414 19080 40406 19136
rect 40462 19080 40467 19136
rect 37414 19078 40467 19080
rect 0 19048 800 19078
rect 26049 19075 26115 19078
rect 28625 19075 28691 19078
rect 40401 19075 40467 19078
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 22946 19007 23262 19008
rect 32946 19072 33262 19073
rect 32946 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33262 19072
rect 32946 19007 33262 19008
rect 42946 19072 43262 19073
rect 42946 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43262 19072
rect 42946 19007 43262 19008
rect 28993 19002 29059 19005
rect 30649 19002 30715 19005
rect 28993 19000 30715 19002
rect 28993 18944 28998 19000
rect 29054 18944 30654 19000
rect 30710 18944 30715 19000
rect 28993 18942 30715 18944
rect 28993 18939 29059 18942
rect 30649 18939 30715 18942
rect 49141 19002 49207 19005
rect 50200 19002 51000 19032
rect 49141 19000 51000 19002
rect 49141 18944 49146 19000
rect 49202 18944 51000 19000
rect 49141 18942 51000 18944
rect 49141 18939 49207 18942
rect 50200 18912 51000 18942
rect 2773 18866 2839 18869
rect 1304 18864 2839 18866
rect 1304 18808 2778 18864
rect 2834 18808 2839 18864
rect 1304 18806 2839 18808
rect 0 18730 800 18760
rect 1304 18730 1364 18806
rect 2773 18803 2839 18806
rect 12065 18866 12131 18869
rect 19425 18866 19491 18869
rect 25865 18866 25931 18869
rect 12065 18864 25931 18866
rect 12065 18808 12070 18864
rect 12126 18808 19430 18864
rect 19486 18808 25870 18864
rect 25926 18808 25931 18864
rect 12065 18806 25931 18808
rect 12065 18803 12131 18806
rect 19425 18803 19491 18806
rect 25865 18803 25931 18806
rect 30005 18866 30071 18869
rect 40125 18866 40191 18869
rect 30005 18864 40191 18866
rect 30005 18808 30010 18864
rect 30066 18808 40130 18864
rect 40186 18808 40191 18864
rect 30005 18806 40191 18808
rect 30005 18803 30071 18806
rect 40125 18803 40191 18806
rect 0 18670 1364 18730
rect 1945 18730 2011 18733
rect 16205 18730 16271 18733
rect 1945 18728 16271 18730
rect 1945 18672 1950 18728
rect 2006 18672 16210 18728
rect 16266 18672 16271 18728
rect 1945 18670 16271 18672
rect 0 18640 800 18670
rect 1945 18667 2011 18670
rect 16205 18667 16271 18670
rect 17401 18730 17467 18733
rect 18873 18730 18939 18733
rect 17401 18728 18939 18730
rect 17401 18672 17406 18728
rect 17462 18672 18878 18728
rect 18934 18672 18939 18728
rect 17401 18670 18939 18672
rect 17401 18667 17467 18670
rect 18873 18667 18939 18670
rect 19793 18730 19859 18733
rect 25037 18730 25103 18733
rect 19793 18728 25103 18730
rect 19793 18672 19798 18728
rect 19854 18672 25042 18728
rect 25098 18672 25103 18728
rect 19793 18670 25103 18672
rect 19793 18667 19859 18670
rect 25037 18667 25103 18670
rect 26969 18730 27035 18733
rect 29637 18730 29703 18733
rect 26969 18728 29703 18730
rect 26969 18672 26974 18728
rect 27030 18672 29642 18728
rect 29698 18672 29703 18728
rect 26969 18670 29703 18672
rect 26969 18667 27035 18670
rect 29637 18667 29703 18670
rect 30465 18730 30531 18733
rect 38009 18730 38075 18733
rect 30465 18728 38075 18730
rect 30465 18672 30470 18728
rect 30526 18672 38014 18728
rect 38070 18672 38075 18728
rect 30465 18670 38075 18672
rect 30465 18667 30531 18670
rect 38009 18667 38075 18670
rect 21265 18594 21331 18597
rect 26417 18594 26483 18597
rect 21265 18592 26483 18594
rect 21265 18536 21270 18592
rect 21326 18536 26422 18592
rect 26478 18536 26483 18592
rect 21265 18534 26483 18536
rect 21265 18531 21331 18534
rect 26417 18531 26483 18534
rect 32949 18594 33015 18597
rect 34145 18594 34211 18597
rect 35617 18594 35683 18597
rect 32949 18592 35683 18594
rect 32949 18536 32954 18592
rect 33010 18536 34150 18592
rect 34206 18536 35622 18592
rect 35678 18536 35683 18592
rect 32949 18534 35683 18536
rect 32949 18531 33015 18534
rect 34145 18531 34211 18534
rect 35617 18531 35683 18534
rect 48773 18594 48839 18597
rect 50200 18594 51000 18624
rect 48773 18592 51000 18594
rect 48773 18536 48778 18592
rect 48834 18536 51000 18592
rect 48773 18534 51000 18536
rect 48773 18531 48839 18534
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 27946 18528 28262 18529
rect 27946 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28262 18528
rect 27946 18463 28262 18464
rect 37946 18528 38262 18529
rect 37946 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38262 18528
rect 37946 18463 38262 18464
rect 47946 18528 48262 18529
rect 47946 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48262 18528
rect 50200 18504 51000 18534
rect 47946 18463 48262 18464
rect 19333 18458 19399 18461
rect 27061 18458 27127 18461
rect 19333 18456 27127 18458
rect 19333 18400 19338 18456
rect 19394 18400 27066 18456
rect 27122 18400 27127 18456
rect 19333 18398 27127 18400
rect 19333 18395 19399 18398
rect 27061 18395 27127 18398
rect 28993 18458 29059 18461
rect 29361 18458 29427 18461
rect 28993 18456 29427 18458
rect 28993 18400 28998 18456
rect 29054 18400 29366 18456
rect 29422 18400 29427 18456
rect 28993 18398 29427 18400
rect 28993 18395 29059 18398
rect 29361 18395 29427 18398
rect 0 18322 800 18352
rect 2865 18322 2931 18325
rect 0 18320 2931 18322
rect 0 18264 2870 18320
rect 2926 18264 2931 18320
rect 0 18262 2931 18264
rect 0 18232 800 18262
rect 2865 18259 2931 18262
rect 15009 18322 15075 18325
rect 19057 18322 19123 18325
rect 15009 18320 19123 18322
rect 15009 18264 15014 18320
rect 15070 18264 19062 18320
rect 19118 18264 19123 18320
rect 15009 18262 19123 18264
rect 15009 18259 15075 18262
rect 19057 18259 19123 18262
rect 25129 18322 25195 18325
rect 25957 18322 26023 18325
rect 40677 18322 40743 18325
rect 25129 18320 40743 18322
rect 25129 18264 25134 18320
rect 25190 18264 25962 18320
rect 26018 18264 40682 18320
rect 40738 18264 40743 18320
rect 25129 18262 40743 18264
rect 25129 18259 25195 18262
rect 25957 18259 26023 18262
rect 40677 18259 40743 18262
rect 11145 18186 11211 18189
rect 14917 18186 14983 18189
rect 11145 18184 14983 18186
rect 11145 18128 11150 18184
rect 11206 18128 14922 18184
rect 14978 18128 14983 18184
rect 11145 18126 14983 18128
rect 11145 18123 11211 18126
rect 14917 18123 14983 18126
rect 15377 18186 15443 18189
rect 25037 18186 25103 18189
rect 26325 18186 26391 18189
rect 15377 18184 26391 18186
rect 15377 18128 15382 18184
rect 15438 18128 25042 18184
rect 25098 18128 26330 18184
rect 26386 18128 26391 18184
rect 15377 18126 26391 18128
rect 15377 18123 15443 18126
rect 25037 18123 25103 18126
rect 26325 18123 26391 18126
rect 27245 18186 27311 18189
rect 29545 18186 29611 18189
rect 30189 18186 30255 18189
rect 39021 18186 39087 18189
rect 27245 18184 30255 18186
rect 27245 18128 27250 18184
rect 27306 18128 29550 18184
rect 29606 18128 30194 18184
rect 30250 18128 30255 18184
rect 27245 18126 30255 18128
rect 27245 18123 27311 18126
rect 29545 18123 29611 18126
rect 30189 18123 30255 18126
rect 31710 18184 39087 18186
rect 31710 18128 39026 18184
rect 39082 18128 39087 18184
rect 31710 18126 39087 18128
rect 27061 18050 27127 18053
rect 31710 18050 31770 18126
rect 39021 18123 39087 18126
rect 49141 18186 49207 18189
rect 50200 18186 51000 18216
rect 49141 18184 51000 18186
rect 49141 18128 49146 18184
rect 49202 18128 51000 18184
rect 49141 18126 51000 18128
rect 49141 18123 49207 18126
rect 50200 18096 51000 18126
rect 27061 18048 31770 18050
rect 27061 17992 27066 18048
rect 27122 17992 31770 18048
rect 27061 17990 31770 17992
rect 34421 18050 34487 18053
rect 34881 18050 34947 18053
rect 35893 18050 35959 18053
rect 34421 18048 35959 18050
rect 34421 17992 34426 18048
rect 34482 17992 34886 18048
rect 34942 17992 35898 18048
rect 35954 17992 35959 18048
rect 34421 17990 35959 17992
rect 27061 17987 27127 17990
rect 34421 17987 34487 17990
rect 34881 17987 34947 17990
rect 35893 17987 35959 17990
rect 2946 17984 3262 17985
rect 0 17914 800 17944
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 32946 17984 33262 17985
rect 32946 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33262 17984
rect 32946 17919 33262 17920
rect 42946 17984 43262 17985
rect 42946 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43262 17984
rect 42946 17919 43262 17920
rect 2681 17914 2747 17917
rect 0 17912 2747 17914
rect 0 17856 2686 17912
rect 2742 17856 2747 17912
rect 0 17854 2747 17856
rect 0 17824 800 17854
rect 2681 17851 2747 17854
rect 27613 17914 27679 17917
rect 27797 17914 27863 17917
rect 28533 17914 28599 17917
rect 27613 17912 28599 17914
rect 27613 17856 27618 17912
rect 27674 17856 27802 17912
rect 27858 17856 28538 17912
rect 28594 17856 28599 17912
rect 27613 17854 28599 17856
rect 27613 17851 27679 17854
rect 27797 17851 27863 17854
rect 28533 17851 28599 17854
rect 21633 17778 21699 17781
rect 39573 17778 39639 17781
rect 21633 17776 39639 17778
rect 21633 17720 21638 17776
rect 21694 17720 39578 17776
rect 39634 17720 39639 17776
rect 21633 17718 39639 17720
rect 21633 17715 21699 17718
rect 39573 17715 39639 17718
rect 49049 17778 49115 17781
rect 50200 17778 51000 17808
rect 49049 17776 51000 17778
rect 49049 17720 49054 17776
rect 49110 17720 51000 17776
rect 49049 17718 51000 17720
rect 49049 17715 49115 17718
rect 50200 17688 51000 17718
rect 26509 17642 26575 17645
rect 30649 17642 30715 17645
rect 26509 17640 30715 17642
rect 26509 17584 26514 17640
rect 26570 17584 30654 17640
rect 30710 17584 30715 17640
rect 26509 17582 30715 17584
rect 26509 17579 26575 17582
rect 30649 17579 30715 17582
rect 0 17506 800 17536
rect 2773 17506 2839 17509
rect 0 17504 2839 17506
rect 0 17448 2778 17504
rect 2834 17448 2839 17504
rect 0 17446 2839 17448
rect 0 17416 800 17446
rect 2773 17443 2839 17446
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 17946 17375 18262 17376
rect 27946 17440 28262 17441
rect 27946 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28262 17440
rect 27946 17375 28262 17376
rect 37946 17440 38262 17441
rect 37946 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38262 17440
rect 37946 17375 38262 17376
rect 47946 17440 48262 17441
rect 47946 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48262 17440
rect 47946 17375 48262 17376
rect 14273 17370 14339 17373
rect 15377 17370 15443 17373
rect 14273 17368 15443 17370
rect 14273 17312 14278 17368
rect 14334 17312 15382 17368
rect 15438 17312 15443 17368
rect 14273 17310 15443 17312
rect 14273 17307 14339 17310
rect 15377 17307 15443 17310
rect 49049 17370 49115 17373
rect 50200 17370 51000 17400
rect 49049 17368 51000 17370
rect 49049 17312 49054 17368
rect 49110 17312 51000 17368
rect 49049 17310 51000 17312
rect 49049 17307 49115 17310
rect 50200 17280 51000 17310
rect 10685 17234 10751 17237
rect 25405 17234 25471 17237
rect 10685 17232 25471 17234
rect 10685 17176 10690 17232
rect 10746 17176 25410 17232
rect 25466 17176 25471 17232
rect 10685 17174 25471 17176
rect 10685 17171 10751 17174
rect 25405 17171 25471 17174
rect 28257 17234 28323 17237
rect 42701 17234 42767 17237
rect 28257 17232 42767 17234
rect 28257 17176 28262 17232
rect 28318 17176 42706 17232
rect 42762 17176 42767 17232
rect 28257 17174 42767 17176
rect 28257 17171 28323 17174
rect 42701 17171 42767 17174
rect 0 17098 800 17128
rect 1209 17098 1275 17101
rect 0 17096 1275 17098
rect 0 17040 1214 17096
rect 1270 17040 1275 17096
rect 0 17038 1275 17040
rect 0 17008 800 17038
rect 1209 17035 1275 17038
rect 11789 17098 11855 17101
rect 14406 17098 14412 17100
rect 11789 17096 14412 17098
rect 11789 17040 11794 17096
rect 11850 17040 14412 17096
rect 11789 17038 14412 17040
rect 11789 17035 11855 17038
rect 14406 17036 14412 17038
rect 14476 17036 14482 17100
rect 26693 17098 26759 17101
rect 36721 17098 36787 17101
rect 38469 17100 38535 17101
rect 38469 17098 38516 17100
rect 26693 17096 36787 17098
rect 26693 17040 26698 17096
rect 26754 17040 36726 17096
rect 36782 17040 36787 17096
rect 26693 17038 36787 17040
rect 38424 17096 38516 17098
rect 38424 17040 38474 17096
rect 38424 17038 38516 17040
rect 26693 17035 26759 17038
rect 36721 17035 36787 17038
rect 38469 17036 38516 17038
rect 38580 17036 38586 17100
rect 38469 17035 38535 17036
rect 17493 16962 17559 16965
rect 21173 16962 21239 16965
rect 17493 16960 21239 16962
rect 17493 16904 17498 16960
rect 17554 16904 21178 16960
rect 21234 16904 21239 16960
rect 17493 16902 21239 16904
rect 17493 16899 17559 16902
rect 21173 16899 21239 16902
rect 27061 16962 27127 16965
rect 27705 16962 27771 16965
rect 27061 16960 27771 16962
rect 27061 16904 27066 16960
rect 27122 16904 27710 16960
rect 27766 16904 27771 16960
rect 27061 16902 27771 16904
rect 27061 16899 27127 16902
rect 27705 16899 27771 16902
rect 48773 16962 48839 16965
rect 50200 16962 51000 16992
rect 48773 16960 51000 16962
rect 48773 16904 48778 16960
rect 48834 16904 51000 16960
rect 48773 16902 51000 16904
rect 48773 16899 48839 16902
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 32946 16896 33262 16897
rect 32946 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33262 16896
rect 32946 16831 33262 16832
rect 42946 16896 43262 16897
rect 42946 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43262 16896
rect 50200 16872 51000 16902
rect 42946 16831 43262 16832
rect 28625 16826 28691 16829
rect 28942 16826 28948 16828
rect 28625 16824 28948 16826
rect 28625 16768 28630 16824
rect 28686 16768 28948 16824
rect 28625 16766 28948 16768
rect 28625 16763 28691 16766
rect 28942 16764 28948 16766
rect 29012 16764 29018 16828
rect 0 16690 800 16720
rect 1301 16690 1367 16693
rect 0 16688 1367 16690
rect 0 16632 1306 16688
rect 1362 16632 1367 16688
rect 0 16630 1367 16632
rect 0 16600 800 16630
rect 1301 16627 1367 16630
rect 10501 16690 10567 16693
rect 15929 16690 15995 16693
rect 16113 16692 16179 16693
rect 10501 16688 15995 16690
rect 10501 16632 10506 16688
rect 10562 16632 15934 16688
rect 15990 16632 15995 16688
rect 10501 16630 15995 16632
rect 10501 16627 10567 16630
rect 15929 16627 15995 16630
rect 16062 16628 16068 16692
rect 16132 16690 16179 16692
rect 19701 16690 19767 16693
rect 23565 16690 23631 16693
rect 27245 16690 27311 16693
rect 16132 16688 16224 16690
rect 16174 16632 16224 16688
rect 16132 16630 16224 16632
rect 19701 16688 27311 16690
rect 19701 16632 19706 16688
rect 19762 16632 23570 16688
rect 23626 16632 27250 16688
rect 27306 16632 27311 16688
rect 19701 16630 27311 16632
rect 16132 16628 16179 16630
rect 16113 16627 16179 16628
rect 19701 16627 19767 16630
rect 23565 16627 23631 16630
rect 27245 16627 27311 16630
rect 29126 16628 29132 16692
rect 29196 16690 29202 16692
rect 29269 16690 29335 16693
rect 29196 16688 29335 16690
rect 29196 16632 29274 16688
rect 29330 16632 29335 16688
rect 29196 16630 29335 16632
rect 29196 16628 29202 16630
rect 29269 16627 29335 16630
rect 30005 16690 30071 16693
rect 32029 16690 32095 16693
rect 30005 16688 32095 16690
rect 30005 16632 30010 16688
rect 30066 16632 32034 16688
rect 32090 16632 32095 16688
rect 30005 16630 32095 16632
rect 30005 16627 30071 16630
rect 32029 16627 32095 16630
rect 9765 16554 9831 16557
rect 14549 16554 14615 16557
rect 9765 16552 14615 16554
rect 9765 16496 9770 16552
rect 9826 16496 14554 16552
rect 14610 16496 14615 16552
rect 9765 16494 14615 16496
rect 9765 16491 9831 16494
rect 14549 16491 14615 16494
rect 15653 16554 15719 16557
rect 20989 16554 21055 16557
rect 15653 16552 21055 16554
rect 15653 16496 15658 16552
rect 15714 16496 20994 16552
rect 21050 16496 21055 16552
rect 15653 16494 21055 16496
rect 15653 16491 15719 16494
rect 20989 16491 21055 16494
rect 22461 16554 22527 16557
rect 38469 16554 38535 16557
rect 22461 16552 38535 16554
rect 22461 16496 22466 16552
rect 22522 16496 38474 16552
rect 38530 16496 38535 16552
rect 22461 16494 38535 16496
rect 22461 16491 22527 16494
rect 38469 16491 38535 16494
rect 49233 16554 49299 16557
rect 50200 16554 51000 16584
rect 49233 16552 51000 16554
rect 49233 16496 49238 16552
rect 49294 16496 51000 16552
rect 49233 16494 51000 16496
rect 49233 16491 49299 16494
rect 50200 16464 51000 16494
rect 7946 16352 8262 16353
rect 0 16282 800 16312
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 27946 16352 28262 16353
rect 27946 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28262 16352
rect 27946 16287 28262 16288
rect 37946 16352 38262 16353
rect 37946 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38262 16352
rect 37946 16287 38262 16288
rect 47946 16352 48262 16353
rect 47946 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48262 16352
rect 47946 16287 48262 16288
rect 1301 16282 1367 16285
rect 0 16280 1367 16282
rect 0 16224 1306 16280
rect 1362 16224 1367 16280
rect 0 16222 1367 16224
rect 0 16192 800 16222
rect 1301 16219 1367 16222
rect 14038 16084 14044 16148
rect 14108 16146 14114 16148
rect 14273 16146 14339 16149
rect 19793 16146 19859 16149
rect 23289 16146 23355 16149
rect 14108 16144 15026 16146
rect 14108 16088 14278 16144
rect 14334 16088 15026 16144
rect 14108 16086 15026 16088
rect 14108 16084 14114 16086
rect 14273 16083 14339 16086
rect 11881 16010 11947 16013
rect 14825 16010 14891 16013
rect 11881 16008 14891 16010
rect 11881 15952 11886 16008
rect 11942 15952 14830 16008
rect 14886 15952 14891 16008
rect 11881 15950 14891 15952
rect 14966 16010 15026 16086
rect 19793 16144 23355 16146
rect 19793 16088 19798 16144
rect 19854 16088 23294 16144
rect 23350 16088 23355 16144
rect 19793 16086 23355 16088
rect 19793 16083 19859 16086
rect 23289 16083 23355 16086
rect 25589 16146 25655 16149
rect 48773 16146 48839 16149
rect 25589 16144 48839 16146
rect 25589 16088 25594 16144
rect 25650 16088 48778 16144
rect 48834 16088 48839 16144
rect 25589 16086 48839 16088
rect 25589 16083 25655 16086
rect 48773 16083 48839 16086
rect 49141 16146 49207 16149
rect 50200 16146 51000 16176
rect 49141 16144 51000 16146
rect 49141 16088 49146 16144
rect 49202 16088 51000 16144
rect 49141 16086 51000 16088
rect 49141 16083 49207 16086
rect 50200 16056 51000 16086
rect 15837 16010 15903 16013
rect 27337 16010 27403 16013
rect 34329 16010 34395 16013
rect 14966 16008 22110 16010
rect 14966 15952 15842 16008
rect 15898 15952 22110 16008
rect 14966 15950 22110 15952
rect 11881 15947 11947 15950
rect 14825 15947 14891 15950
rect 15837 15947 15903 15950
rect 0 15874 800 15904
rect 1301 15874 1367 15877
rect 16941 15876 17007 15877
rect 16941 15874 16988 15876
rect 0 15872 1367 15874
rect 0 15816 1306 15872
rect 1362 15816 1367 15872
rect 0 15814 1367 15816
rect 16896 15872 16988 15874
rect 16896 15816 16946 15872
rect 16896 15814 16988 15816
rect 0 15784 800 15814
rect 1301 15811 1367 15814
rect 16941 15812 16988 15814
rect 17052 15812 17058 15876
rect 16941 15811 17007 15812
rect 2946 15808 3262 15809
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 14641 15602 14707 15605
rect 17309 15602 17375 15605
rect 14641 15600 17375 15602
rect 14641 15544 14646 15600
rect 14702 15544 17314 15600
rect 17370 15544 17375 15600
rect 14641 15542 17375 15544
rect 22050 15602 22110 15950
rect 27337 16008 34395 16010
rect 27337 15952 27342 16008
rect 27398 15952 34334 16008
rect 34390 15952 34395 16008
rect 27337 15950 34395 15952
rect 27337 15947 27403 15950
rect 34329 15947 34395 15950
rect 35709 16010 35775 16013
rect 49233 16010 49299 16013
rect 35709 16008 49299 16010
rect 35709 15952 35714 16008
rect 35770 15952 49238 16008
rect 49294 15952 49299 16008
rect 35709 15950 49299 15952
rect 35709 15947 35775 15950
rect 49233 15947 49299 15950
rect 26141 15874 26207 15877
rect 32489 15874 32555 15877
rect 26141 15872 32555 15874
rect 26141 15816 26146 15872
rect 26202 15816 32494 15872
rect 32550 15816 32555 15872
rect 26141 15814 32555 15816
rect 26141 15811 26207 15814
rect 32489 15811 32555 15814
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 22946 15743 23262 15744
rect 32946 15808 33262 15809
rect 32946 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33262 15808
rect 32946 15743 33262 15744
rect 42946 15808 43262 15809
rect 42946 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43262 15808
rect 42946 15743 43262 15744
rect 49049 15738 49115 15741
rect 50200 15738 51000 15768
rect 49049 15736 51000 15738
rect 49049 15680 49054 15736
rect 49110 15680 51000 15736
rect 49049 15678 51000 15680
rect 49049 15675 49115 15678
rect 50200 15648 51000 15678
rect 29545 15602 29611 15605
rect 30465 15602 30531 15605
rect 22050 15600 30531 15602
rect 22050 15544 29550 15600
rect 29606 15544 30470 15600
rect 30526 15544 30531 15600
rect 22050 15542 30531 15544
rect 14641 15539 14707 15542
rect 17309 15539 17375 15542
rect 29545 15539 29611 15542
rect 30465 15539 30531 15542
rect 0 15466 800 15496
rect 1301 15466 1367 15469
rect 0 15464 1367 15466
rect 0 15408 1306 15464
rect 1362 15408 1367 15464
rect 0 15406 1367 15408
rect 0 15376 800 15406
rect 1301 15403 1367 15406
rect 12433 15466 12499 15469
rect 15561 15466 15627 15469
rect 12433 15464 15627 15466
rect 12433 15408 12438 15464
rect 12494 15408 15566 15464
rect 15622 15408 15627 15464
rect 12433 15406 15627 15408
rect 12433 15403 12499 15406
rect 15561 15403 15627 15406
rect 26969 15466 27035 15469
rect 34421 15466 34487 15469
rect 26969 15464 34487 15466
rect 26969 15408 26974 15464
rect 27030 15408 34426 15464
rect 34482 15408 34487 15464
rect 26969 15406 34487 15408
rect 26969 15403 27035 15406
rect 34421 15403 34487 15406
rect 10501 15330 10567 15333
rect 12433 15330 12499 15333
rect 10501 15328 12499 15330
rect 10501 15272 10506 15328
rect 10562 15272 12438 15328
rect 12494 15272 12499 15328
rect 10501 15270 12499 15272
rect 10501 15267 10567 15270
rect 12433 15267 12499 15270
rect 49325 15330 49391 15333
rect 50200 15330 51000 15360
rect 49325 15328 51000 15330
rect 49325 15272 49330 15328
rect 49386 15272 51000 15328
rect 49325 15270 51000 15272
rect 49325 15267 49391 15270
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 27946 15264 28262 15265
rect 27946 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28262 15264
rect 27946 15199 28262 15200
rect 37946 15264 38262 15265
rect 37946 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38262 15264
rect 37946 15199 38262 15200
rect 47946 15264 48262 15265
rect 47946 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48262 15264
rect 50200 15240 51000 15270
rect 47946 15199 48262 15200
rect 20529 15194 20595 15197
rect 27521 15194 27587 15197
rect 20529 15192 27587 15194
rect 20529 15136 20534 15192
rect 20590 15136 27526 15192
rect 27582 15136 27587 15192
rect 20529 15134 27587 15136
rect 20529 15131 20595 15134
rect 27521 15131 27587 15134
rect 0 15058 800 15088
rect 1301 15058 1367 15061
rect 0 15056 1367 15058
rect 0 15000 1306 15056
rect 1362 15000 1367 15056
rect 0 14998 1367 15000
rect 0 14968 800 14998
rect 1301 14995 1367 14998
rect 14365 15058 14431 15061
rect 15009 15058 15075 15061
rect 16573 15058 16639 15061
rect 14365 15056 16639 15058
rect 14365 15000 14370 15056
rect 14426 15000 15014 15056
rect 15070 15000 16578 15056
rect 16634 15000 16639 15056
rect 14365 14998 16639 15000
rect 14365 14995 14431 14998
rect 15009 14995 15075 14998
rect 16573 14995 16639 14998
rect 17585 15058 17651 15061
rect 21633 15058 21699 15061
rect 17585 15056 21699 15058
rect 17585 15000 17590 15056
rect 17646 15000 21638 15056
rect 21694 15000 21699 15056
rect 17585 14998 21699 15000
rect 17585 14995 17651 14998
rect 21633 14995 21699 14998
rect 27061 15058 27127 15061
rect 49233 15058 49299 15061
rect 27061 15056 49299 15058
rect 27061 15000 27066 15056
rect 27122 15000 49238 15056
rect 49294 15000 49299 15056
rect 27061 14998 49299 15000
rect 27061 14995 27127 14998
rect 49233 14995 49299 14998
rect 12341 14922 12407 14925
rect 26325 14922 26391 14925
rect 12341 14920 26391 14922
rect 12341 14864 12346 14920
rect 12402 14864 26330 14920
rect 26386 14864 26391 14920
rect 12341 14862 26391 14864
rect 12341 14859 12407 14862
rect 26325 14859 26391 14862
rect 37181 14922 37247 14925
rect 38561 14922 38627 14925
rect 37181 14920 38627 14922
rect 37181 14864 37186 14920
rect 37242 14864 38566 14920
rect 38622 14864 38627 14920
rect 37181 14862 38627 14864
rect 37181 14859 37247 14862
rect 38561 14859 38627 14862
rect 49049 14922 49115 14925
rect 50200 14922 51000 14952
rect 49049 14920 51000 14922
rect 49049 14864 49054 14920
rect 49110 14864 51000 14920
rect 49049 14862 51000 14864
rect 49049 14859 49115 14862
rect 50200 14832 51000 14862
rect 2946 14720 3262 14721
rect 0 14650 800 14680
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 32946 14720 33262 14721
rect 32946 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33262 14720
rect 32946 14655 33262 14656
rect 42946 14720 43262 14721
rect 42946 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43262 14720
rect 42946 14655 43262 14656
rect 1301 14650 1367 14653
rect 0 14648 1367 14650
rect 0 14592 1306 14648
rect 1362 14592 1367 14648
rect 0 14590 1367 14592
rect 0 14560 800 14590
rect 1301 14587 1367 14590
rect 10317 14514 10383 14517
rect 21817 14514 21883 14517
rect 35709 14514 35775 14517
rect 10317 14512 35775 14514
rect 10317 14456 10322 14512
rect 10378 14456 21822 14512
rect 21878 14456 35714 14512
rect 35770 14456 35775 14512
rect 10317 14454 35775 14456
rect 10317 14451 10383 14454
rect 21817 14451 21883 14454
rect 35709 14451 35775 14454
rect 49141 14514 49207 14517
rect 50200 14514 51000 14544
rect 49141 14512 51000 14514
rect 49141 14456 49146 14512
rect 49202 14456 51000 14512
rect 49141 14454 51000 14456
rect 49141 14451 49207 14454
rect 50200 14424 51000 14454
rect 14181 14380 14247 14381
rect 14181 14378 14228 14380
rect 14136 14376 14228 14378
rect 14136 14320 14186 14376
rect 14136 14318 14228 14320
rect 14181 14316 14228 14318
rect 14292 14316 14298 14380
rect 21725 14378 21791 14381
rect 24393 14378 24459 14381
rect 21725 14376 24459 14378
rect 21725 14320 21730 14376
rect 21786 14320 24398 14376
rect 24454 14320 24459 14376
rect 21725 14318 24459 14320
rect 14181 14315 14247 14316
rect 21725 14315 21791 14318
rect 24393 14315 24459 14318
rect 28257 14378 28323 14381
rect 28717 14378 28783 14381
rect 39941 14378 40007 14381
rect 28257 14376 40007 14378
rect 28257 14320 28262 14376
rect 28318 14320 28722 14376
rect 28778 14320 39946 14376
rect 40002 14320 40007 14376
rect 28257 14318 40007 14320
rect 28257 14315 28323 14318
rect 28717 14315 28783 14318
rect 39941 14315 40007 14318
rect 0 14242 800 14272
rect 1301 14242 1367 14245
rect 0 14240 1367 14242
rect 0 14184 1306 14240
rect 1362 14184 1367 14240
rect 0 14182 1367 14184
rect 0 14152 800 14182
rect 1301 14179 1367 14182
rect 19977 14242 20043 14245
rect 24577 14242 24643 14245
rect 19977 14240 24643 14242
rect 19977 14184 19982 14240
rect 20038 14184 24582 14240
rect 24638 14184 24643 14240
rect 19977 14182 24643 14184
rect 19977 14179 20043 14182
rect 24577 14179 24643 14182
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 17946 14111 18262 14112
rect 27946 14176 28262 14177
rect 27946 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28262 14176
rect 27946 14111 28262 14112
rect 37946 14176 38262 14177
rect 37946 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38262 14176
rect 37946 14111 38262 14112
rect 47946 14176 48262 14177
rect 47946 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48262 14176
rect 47946 14111 48262 14112
rect 29729 14106 29795 14109
rect 31109 14106 31175 14109
rect 29729 14104 31175 14106
rect 29729 14048 29734 14104
rect 29790 14048 31114 14104
rect 31170 14048 31175 14104
rect 29729 14046 31175 14048
rect 29729 14043 29795 14046
rect 31109 14043 31175 14046
rect 49141 14106 49207 14109
rect 50200 14106 51000 14136
rect 49141 14104 51000 14106
rect 49141 14048 49146 14104
rect 49202 14048 51000 14104
rect 49141 14046 51000 14048
rect 49141 14043 49207 14046
rect 50200 14016 51000 14046
rect 0 13834 800 13864
rect 2773 13834 2839 13837
rect 0 13832 2839 13834
rect 0 13776 2778 13832
rect 2834 13776 2839 13832
rect 0 13774 2839 13776
rect 0 13744 800 13774
rect 2773 13771 2839 13774
rect 11513 13834 11579 13837
rect 16481 13834 16547 13837
rect 18505 13834 18571 13837
rect 19057 13834 19123 13837
rect 11513 13832 19123 13834
rect 11513 13776 11518 13832
rect 11574 13776 16486 13832
rect 16542 13776 18510 13832
rect 18566 13776 19062 13832
rect 19118 13776 19123 13832
rect 11513 13774 19123 13776
rect 11513 13771 11579 13774
rect 16481 13771 16547 13774
rect 18505 13771 18571 13774
rect 19057 13771 19123 13774
rect 32213 13834 32279 13837
rect 33685 13834 33751 13837
rect 32213 13832 33751 13834
rect 32213 13776 32218 13832
rect 32274 13776 33690 13832
rect 33746 13776 33751 13832
rect 32213 13774 33751 13776
rect 32213 13771 32279 13774
rect 33685 13771 33751 13774
rect 14549 13698 14615 13701
rect 16062 13698 16068 13700
rect 14549 13696 16068 13698
rect 14549 13640 14554 13696
rect 14610 13640 16068 13696
rect 14549 13638 16068 13640
rect 14549 13635 14615 13638
rect 16062 13636 16068 13638
rect 16132 13636 16138 13700
rect 48221 13698 48287 13701
rect 50200 13698 51000 13728
rect 48221 13696 51000 13698
rect 48221 13640 48226 13696
rect 48282 13640 51000 13696
rect 48221 13638 51000 13640
rect 48221 13635 48287 13638
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 32946 13632 33262 13633
rect 32946 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33262 13632
rect 32946 13567 33262 13568
rect 42946 13632 43262 13633
rect 42946 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43262 13632
rect 50200 13608 51000 13638
rect 42946 13567 43262 13568
rect 14273 13562 14339 13565
rect 16941 13562 17007 13565
rect 14273 13560 17007 13562
rect 14273 13504 14278 13560
rect 14334 13504 16946 13560
rect 17002 13504 17007 13560
rect 14273 13502 17007 13504
rect 14273 13499 14339 13502
rect 16941 13499 17007 13502
rect 0 13426 800 13456
rect 3509 13426 3575 13429
rect 0 13424 3575 13426
rect 0 13368 3514 13424
rect 3570 13368 3575 13424
rect 0 13366 3575 13368
rect 0 13336 800 13366
rect 3509 13363 3575 13366
rect 19241 13290 19307 13293
rect 35341 13290 35407 13293
rect 19241 13288 35407 13290
rect 19241 13232 19246 13288
rect 19302 13232 35346 13288
rect 35402 13232 35407 13288
rect 19241 13230 35407 13232
rect 19241 13227 19307 13230
rect 35341 13227 35407 13230
rect 49141 13290 49207 13293
rect 50200 13290 51000 13320
rect 49141 13288 51000 13290
rect 49141 13232 49146 13288
rect 49202 13232 51000 13288
rect 49141 13230 51000 13232
rect 49141 13227 49207 13230
rect 50200 13200 51000 13230
rect 7946 13088 8262 13089
rect 0 13018 800 13048
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 27946 13088 28262 13089
rect 27946 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28262 13088
rect 27946 13023 28262 13024
rect 37946 13088 38262 13089
rect 37946 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38262 13088
rect 37946 13023 38262 13024
rect 47946 13088 48262 13089
rect 47946 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48262 13088
rect 47946 13023 48262 13024
rect 1301 13018 1367 13021
rect 0 13016 1367 13018
rect 0 12960 1306 13016
rect 1362 12960 1367 13016
rect 0 12958 1367 12960
rect 0 12928 800 12958
rect 1301 12955 1367 12958
rect 22645 13018 22711 13021
rect 23105 13018 23171 13021
rect 26233 13018 26299 13021
rect 22645 13016 26299 13018
rect 22645 12960 22650 13016
rect 22706 12960 23110 13016
rect 23166 12960 26238 13016
rect 26294 12960 26299 13016
rect 22645 12958 26299 12960
rect 22645 12955 22711 12958
rect 23105 12955 23171 12958
rect 26233 12955 26299 12958
rect 16205 12882 16271 12885
rect 24485 12882 24551 12885
rect 16205 12880 24551 12882
rect 16205 12824 16210 12880
rect 16266 12824 24490 12880
rect 24546 12824 24551 12880
rect 16205 12822 24551 12824
rect 16205 12819 16271 12822
rect 24485 12819 24551 12822
rect 29545 12882 29611 12885
rect 35801 12882 35867 12885
rect 36077 12882 36143 12885
rect 29545 12880 31770 12882
rect 29545 12824 29550 12880
rect 29606 12824 31770 12880
rect 29545 12822 31770 12824
rect 29545 12819 29611 12822
rect 14406 12684 14412 12748
rect 14476 12746 14482 12748
rect 16205 12746 16271 12749
rect 14476 12744 16271 12746
rect 14476 12688 16210 12744
rect 16266 12688 16271 12744
rect 14476 12686 16271 12688
rect 14476 12684 14482 12686
rect 16205 12683 16271 12686
rect 20069 12746 20135 12749
rect 21633 12746 21699 12749
rect 23013 12746 23079 12749
rect 25865 12746 25931 12749
rect 20069 12744 25931 12746
rect 20069 12688 20074 12744
rect 20130 12688 21638 12744
rect 21694 12688 23018 12744
rect 23074 12688 25870 12744
rect 25926 12688 25931 12744
rect 20069 12686 25931 12688
rect 31710 12746 31770 12822
rect 35801 12880 36143 12882
rect 35801 12824 35806 12880
rect 35862 12824 36082 12880
rect 36138 12824 36143 12880
rect 35801 12822 36143 12824
rect 35801 12819 35867 12822
rect 36077 12819 36143 12822
rect 49141 12882 49207 12885
rect 50200 12882 51000 12912
rect 49141 12880 51000 12882
rect 49141 12824 49146 12880
rect 49202 12824 51000 12880
rect 49141 12822 51000 12824
rect 49141 12819 49207 12822
rect 50200 12792 51000 12822
rect 35801 12746 35867 12749
rect 31710 12744 35867 12746
rect 31710 12688 35806 12744
rect 35862 12688 35867 12744
rect 31710 12686 35867 12688
rect 20069 12683 20135 12686
rect 21633 12683 21699 12686
rect 23013 12683 23079 12686
rect 25865 12683 25931 12686
rect 35801 12683 35867 12686
rect 0 12610 800 12640
rect 1209 12610 1275 12613
rect 0 12608 1275 12610
rect 0 12552 1214 12608
rect 1270 12552 1275 12608
rect 0 12550 1275 12552
rect 0 12520 800 12550
rect 1209 12547 1275 12550
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 22946 12479 23262 12480
rect 32946 12544 33262 12545
rect 32946 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33262 12544
rect 32946 12479 33262 12480
rect 42946 12544 43262 12545
rect 42946 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43262 12544
rect 42946 12479 43262 12480
rect 22645 12474 22711 12477
rect 22142 12472 22711 12474
rect 22142 12416 22650 12472
rect 22706 12416 22711 12472
rect 22142 12414 22711 12416
rect 17125 12338 17191 12341
rect 22142 12338 22202 12414
rect 22645 12411 22711 12414
rect 49141 12474 49207 12477
rect 50200 12474 51000 12504
rect 49141 12472 51000 12474
rect 49141 12416 49146 12472
rect 49202 12416 51000 12472
rect 49141 12414 51000 12416
rect 49141 12411 49207 12414
rect 50200 12384 51000 12414
rect 17125 12336 22202 12338
rect 17125 12280 17130 12336
rect 17186 12280 22202 12336
rect 17125 12278 22202 12280
rect 17125 12275 17191 12278
rect 0 12202 800 12232
rect 1209 12202 1275 12205
rect 0 12200 1275 12202
rect 0 12144 1214 12200
rect 1270 12144 1275 12200
rect 0 12142 1275 12144
rect 0 12112 800 12142
rect 1209 12139 1275 12142
rect 16481 12202 16547 12205
rect 17309 12202 17375 12205
rect 22093 12202 22159 12205
rect 22553 12202 22619 12205
rect 30373 12202 30439 12205
rect 34421 12202 34487 12205
rect 16481 12200 34487 12202
rect 16481 12144 16486 12200
rect 16542 12144 17314 12200
rect 17370 12144 22098 12200
rect 22154 12144 22558 12200
rect 22614 12144 30378 12200
rect 30434 12144 34426 12200
rect 34482 12144 34487 12200
rect 16481 12142 34487 12144
rect 16481 12139 16547 12142
rect 17309 12139 17375 12142
rect 22093 12139 22159 12142
rect 22553 12139 22619 12142
rect 30373 12139 30439 12142
rect 34421 12139 34487 12142
rect 49141 12066 49207 12069
rect 50200 12066 51000 12096
rect 49141 12064 51000 12066
rect 49141 12008 49146 12064
rect 49202 12008 51000 12064
rect 49141 12006 51000 12008
rect 49141 12003 49207 12006
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 27946 12000 28262 12001
rect 27946 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28262 12000
rect 27946 11935 28262 11936
rect 37946 12000 38262 12001
rect 37946 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38262 12000
rect 37946 11935 38262 11936
rect 47946 12000 48262 12001
rect 47946 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48262 12000
rect 50200 11976 51000 12006
rect 47946 11935 48262 11936
rect 0 11794 800 11824
rect 1301 11794 1367 11797
rect 0 11792 1367 11794
rect 0 11736 1306 11792
rect 1362 11736 1367 11792
rect 0 11734 1367 11736
rect 0 11704 800 11734
rect 1301 11731 1367 11734
rect 15009 11794 15075 11797
rect 16113 11794 16179 11797
rect 15009 11792 16179 11794
rect 15009 11736 15014 11792
rect 15070 11736 16118 11792
rect 16174 11736 16179 11792
rect 15009 11734 16179 11736
rect 15009 11731 15075 11734
rect 16113 11731 16179 11734
rect 19885 11794 19951 11797
rect 25405 11794 25471 11797
rect 19885 11792 25471 11794
rect 19885 11736 19890 11792
rect 19946 11736 25410 11792
rect 25466 11736 25471 11792
rect 19885 11734 25471 11736
rect 19885 11731 19951 11734
rect 25405 11731 25471 11734
rect 15193 11658 15259 11661
rect 15653 11658 15719 11661
rect 15193 11656 15719 11658
rect 15193 11600 15198 11656
rect 15254 11600 15658 11656
rect 15714 11600 15719 11656
rect 15193 11598 15719 11600
rect 15193 11595 15259 11598
rect 15653 11595 15719 11598
rect 31201 11658 31267 11661
rect 32029 11658 32095 11661
rect 31201 11656 32095 11658
rect 31201 11600 31206 11656
rect 31262 11600 32034 11656
rect 32090 11600 32095 11656
rect 31201 11598 32095 11600
rect 31201 11595 31267 11598
rect 32029 11595 32095 11598
rect 49141 11658 49207 11661
rect 50200 11658 51000 11688
rect 49141 11656 51000 11658
rect 49141 11600 49146 11656
rect 49202 11600 51000 11656
rect 49141 11598 51000 11600
rect 49141 11595 49207 11598
rect 50200 11568 51000 11598
rect 13353 11522 13419 11525
rect 14365 11522 14431 11525
rect 18229 11522 18295 11525
rect 13353 11520 18295 11522
rect 13353 11464 13358 11520
rect 13414 11464 14370 11520
rect 14426 11464 18234 11520
rect 18290 11464 18295 11520
rect 13353 11462 18295 11464
rect 13353 11459 13419 11462
rect 14365 11459 14431 11462
rect 18229 11459 18295 11462
rect 2946 11456 3262 11457
rect 0 11386 800 11416
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 32946 11456 33262 11457
rect 32946 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33262 11456
rect 32946 11391 33262 11392
rect 42946 11456 43262 11457
rect 42946 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43262 11456
rect 42946 11391 43262 11392
rect 1301 11386 1367 11389
rect 0 11384 1367 11386
rect 0 11328 1306 11384
rect 1362 11328 1367 11384
rect 0 11326 1367 11328
rect 0 11296 800 11326
rect 1301 11323 1367 11326
rect 13537 11386 13603 11389
rect 16665 11386 16731 11389
rect 13537 11384 16731 11386
rect 13537 11328 13542 11384
rect 13598 11328 16670 11384
rect 16726 11328 16731 11384
rect 13537 11326 16731 11328
rect 13537 11323 13603 11326
rect 16665 11323 16731 11326
rect 17677 11250 17743 11253
rect 18413 11250 18479 11253
rect 49233 11250 49299 11253
rect 50200 11250 51000 11280
rect 17677 11248 23858 11250
rect 17677 11192 17682 11248
rect 17738 11192 18418 11248
rect 18474 11192 23858 11248
rect 17677 11190 23858 11192
rect 17677 11187 17743 11190
rect 18413 11187 18479 11190
rect 23798 11117 23858 11190
rect 49233 11248 51000 11250
rect 49233 11192 49238 11248
rect 49294 11192 51000 11248
rect 49233 11190 51000 11192
rect 49233 11187 49299 11190
rect 50200 11160 51000 11190
rect 1761 11114 1827 11117
rect 14038 11114 14044 11116
rect 1761 11112 14044 11114
rect 1761 11056 1766 11112
rect 1822 11056 14044 11112
rect 1761 11054 14044 11056
rect 1761 11051 1827 11054
rect 14038 11052 14044 11054
rect 14108 11052 14114 11116
rect 14733 11114 14799 11117
rect 16849 11114 16915 11117
rect 18597 11114 18663 11117
rect 14733 11112 18663 11114
rect 14733 11056 14738 11112
rect 14794 11056 16854 11112
rect 16910 11056 18602 11112
rect 18658 11056 18663 11112
rect 14733 11054 18663 11056
rect 14733 11051 14799 11054
rect 16849 11051 16915 11054
rect 18597 11051 18663 11054
rect 20805 11114 20871 11117
rect 22001 11114 22067 11117
rect 20805 11112 22067 11114
rect 20805 11056 20810 11112
rect 20866 11056 22006 11112
rect 22062 11056 22067 11112
rect 20805 11054 22067 11056
rect 23798 11114 23907 11117
rect 24117 11114 24183 11117
rect 28533 11114 28599 11117
rect 23798 11112 28599 11114
rect 23798 11056 23846 11112
rect 23902 11056 24122 11112
rect 24178 11056 28538 11112
rect 28594 11056 28599 11112
rect 23798 11054 28599 11056
rect 20805 11051 20871 11054
rect 22001 11051 22067 11054
rect 23841 11051 23907 11054
rect 24117 11051 24183 11054
rect 28533 11051 28599 11054
rect 30189 11114 30255 11117
rect 39941 11114 40007 11117
rect 30189 11112 40007 11114
rect 30189 11056 30194 11112
rect 30250 11056 39946 11112
rect 40002 11056 40007 11112
rect 30189 11054 40007 11056
rect 30189 11051 30255 11054
rect 39941 11051 40007 11054
rect 0 10978 800 11008
rect 1577 10978 1643 10981
rect 0 10976 1643 10978
rect 0 10920 1582 10976
rect 1638 10920 1643 10976
rect 0 10918 1643 10920
rect 0 10888 800 10918
rect 1577 10915 1643 10918
rect 29085 10980 29151 10981
rect 29085 10976 29132 10980
rect 29196 10978 29202 10980
rect 29085 10920 29090 10976
rect 29085 10916 29132 10920
rect 29196 10918 29242 10978
rect 29196 10916 29202 10918
rect 29085 10915 29151 10916
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 17946 10847 18262 10848
rect 27946 10912 28262 10913
rect 27946 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28262 10912
rect 27946 10847 28262 10848
rect 37946 10912 38262 10913
rect 37946 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38262 10912
rect 37946 10847 38262 10848
rect 47946 10912 48262 10913
rect 47946 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48262 10912
rect 47946 10847 48262 10848
rect 49141 10842 49207 10845
rect 50200 10842 51000 10872
rect 49141 10840 51000 10842
rect 49141 10784 49146 10840
rect 49202 10784 51000 10840
rect 49141 10782 51000 10784
rect 49141 10779 49207 10782
rect 50200 10752 51000 10782
rect 13629 10706 13695 10709
rect 33685 10706 33751 10709
rect 13629 10704 33751 10706
rect 13629 10648 13634 10704
rect 13690 10648 33690 10704
rect 33746 10648 33751 10704
rect 13629 10646 33751 10648
rect 13629 10643 13695 10646
rect 33685 10643 33751 10646
rect 33869 10706 33935 10709
rect 34237 10706 34303 10709
rect 39757 10706 39823 10709
rect 33869 10704 39823 10706
rect 33869 10648 33874 10704
rect 33930 10648 34242 10704
rect 34298 10648 39762 10704
rect 39818 10648 39823 10704
rect 33869 10646 39823 10648
rect 33869 10643 33935 10646
rect 34237 10643 34303 10646
rect 39757 10643 39823 10646
rect 0 10570 800 10600
rect 1301 10570 1367 10573
rect 0 10568 1367 10570
rect 0 10512 1306 10568
rect 1362 10512 1367 10568
rect 0 10510 1367 10512
rect 0 10480 800 10510
rect 1301 10507 1367 10510
rect 49325 10434 49391 10437
rect 50200 10434 51000 10464
rect 49325 10432 51000 10434
rect 49325 10376 49330 10432
rect 49386 10376 51000 10432
rect 49325 10374 51000 10376
rect 49325 10371 49391 10374
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 32946 10368 33262 10369
rect 32946 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33262 10368
rect 32946 10303 33262 10304
rect 42946 10368 43262 10369
rect 42946 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43262 10368
rect 50200 10344 51000 10374
rect 42946 10303 43262 10304
rect 0 10162 800 10192
rect 1209 10162 1275 10165
rect 0 10160 1275 10162
rect 0 10104 1214 10160
rect 1270 10104 1275 10160
rect 0 10102 1275 10104
rect 0 10072 800 10102
rect 1209 10099 1275 10102
rect 13077 10162 13143 10165
rect 16982 10162 16988 10164
rect 13077 10160 16988 10162
rect 13077 10104 13082 10160
rect 13138 10104 16988 10160
rect 13077 10102 16988 10104
rect 13077 10099 13143 10102
rect 16982 10100 16988 10102
rect 17052 10100 17058 10164
rect 26785 10162 26851 10165
rect 27521 10162 27587 10165
rect 38561 10164 38627 10165
rect 38510 10162 38516 10164
rect 26785 10160 38516 10162
rect 38580 10160 38627 10164
rect 26785 10104 26790 10160
rect 26846 10104 27526 10160
rect 27582 10104 38516 10160
rect 38622 10104 38627 10160
rect 26785 10102 38516 10104
rect 26785 10099 26851 10102
rect 27521 10099 27587 10102
rect 38510 10100 38516 10102
rect 38580 10100 38627 10104
rect 38561 10099 38627 10100
rect 16573 10026 16639 10029
rect 21265 10026 21331 10029
rect 22461 10026 22527 10029
rect 16573 10024 22527 10026
rect 16573 9968 16578 10024
rect 16634 9968 21270 10024
rect 21326 9968 22466 10024
rect 22522 9968 22527 10024
rect 16573 9966 22527 9968
rect 16573 9963 16639 9966
rect 21265 9963 21331 9966
rect 22461 9963 22527 9966
rect 49233 10026 49299 10029
rect 50200 10026 51000 10056
rect 49233 10024 51000 10026
rect 49233 9968 49238 10024
rect 49294 9968 51000 10024
rect 49233 9966 51000 9968
rect 49233 9963 49299 9966
rect 50200 9936 51000 9966
rect 7946 9824 8262 9825
rect 0 9754 800 9784
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 27946 9824 28262 9825
rect 27946 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28262 9824
rect 27946 9759 28262 9760
rect 37946 9824 38262 9825
rect 37946 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38262 9824
rect 37946 9759 38262 9760
rect 47946 9824 48262 9825
rect 47946 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48262 9824
rect 47946 9759 48262 9760
rect 1301 9754 1367 9757
rect 0 9752 1367 9754
rect 0 9696 1306 9752
rect 1362 9696 1367 9752
rect 0 9694 1367 9696
rect 0 9664 800 9694
rect 1301 9691 1367 9694
rect 31477 9754 31543 9757
rect 33225 9754 33291 9757
rect 31477 9752 33291 9754
rect 31477 9696 31482 9752
rect 31538 9696 33230 9752
rect 33286 9696 33291 9752
rect 31477 9694 33291 9696
rect 31477 9691 31543 9694
rect 33225 9691 33291 9694
rect 26141 9618 26207 9621
rect 34605 9618 34671 9621
rect 35801 9618 35867 9621
rect 26141 9616 35867 9618
rect 26141 9560 26146 9616
rect 26202 9560 34610 9616
rect 34666 9560 35806 9616
rect 35862 9560 35867 9616
rect 26141 9558 35867 9560
rect 26141 9555 26207 9558
rect 34605 9555 34671 9558
rect 35801 9555 35867 9558
rect 47301 9618 47367 9621
rect 50200 9618 51000 9648
rect 47301 9616 51000 9618
rect 47301 9560 47306 9616
rect 47362 9560 51000 9616
rect 47301 9558 51000 9560
rect 47301 9555 47367 9558
rect 50200 9528 51000 9558
rect 1761 9482 1827 9485
rect 32581 9482 32647 9485
rect 1761 9480 32647 9482
rect 1761 9424 1766 9480
rect 1822 9424 32586 9480
rect 32642 9424 32647 9480
rect 1761 9422 32647 9424
rect 1761 9419 1827 9422
rect 32581 9419 32647 9422
rect 0 9346 800 9376
rect 1301 9346 1367 9349
rect 0 9344 1367 9346
rect 0 9288 1306 9344
rect 1362 9288 1367 9344
rect 0 9286 1367 9288
rect 0 9256 800 9286
rect 1301 9283 1367 9286
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 22946 9215 23262 9216
rect 32946 9280 33262 9281
rect 32946 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33262 9280
rect 32946 9215 33262 9216
rect 42946 9280 43262 9281
rect 42946 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43262 9280
rect 42946 9215 43262 9216
rect 49141 9210 49207 9213
rect 50200 9210 51000 9240
rect 49141 9208 51000 9210
rect 49141 9152 49146 9208
rect 49202 9152 51000 9208
rect 49141 9150 51000 9152
rect 49141 9147 49207 9150
rect 50200 9120 51000 9150
rect 14181 9076 14247 9077
rect 14181 9072 14228 9076
rect 14292 9074 14298 9076
rect 25589 9074 25655 9077
rect 14292 9072 25655 9074
rect 14181 9016 14186 9072
rect 14292 9016 25594 9072
rect 25650 9016 25655 9072
rect 14181 9012 14228 9016
rect 14292 9014 25655 9016
rect 14292 9012 14298 9014
rect 14181 9011 14247 9012
rect 25589 9011 25655 9014
rect 28625 9074 28691 9077
rect 31937 9074 32003 9077
rect 33041 9074 33107 9077
rect 28625 9072 33107 9074
rect 28625 9016 28630 9072
rect 28686 9016 31942 9072
rect 31998 9016 33046 9072
rect 33102 9016 33107 9072
rect 28625 9014 33107 9016
rect 28625 9011 28691 9014
rect 31937 9011 32003 9014
rect 33041 9011 33107 9014
rect 0 8938 800 8968
rect 1301 8938 1367 8941
rect 0 8936 1367 8938
rect 0 8880 1306 8936
rect 1362 8880 1367 8936
rect 0 8878 1367 8880
rect 0 8848 800 8878
rect 1301 8875 1367 8878
rect 49233 8802 49299 8805
rect 50200 8802 51000 8832
rect 49233 8800 51000 8802
rect 49233 8744 49238 8800
rect 49294 8744 51000 8800
rect 49233 8742 51000 8744
rect 49233 8739 49299 8742
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 27946 8736 28262 8737
rect 27946 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28262 8736
rect 27946 8671 28262 8672
rect 37946 8736 38262 8737
rect 37946 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38262 8736
rect 37946 8671 38262 8672
rect 47946 8736 48262 8737
rect 47946 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48262 8736
rect 50200 8712 51000 8742
rect 47946 8671 48262 8672
rect 0 8530 800 8560
rect 1209 8530 1275 8533
rect 0 8528 1275 8530
rect 0 8472 1214 8528
rect 1270 8472 1275 8528
rect 0 8470 1275 8472
rect 0 8440 800 8470
rect 1209 8467 1275 8470
rect 49325 8394 49391 8397
rect 50200 8394 51000 8424
rect 49325 8392 51000 8394
rect 49325 8336 49330 8392
rect 49386 8336 51000 8392
rect 49325 8334 51000 8336
rect 49325 8331 49391 8334
rect 50200 8304 51000 8334
rect 2946 8192 3262 8193
rect 0 8122 800 8152
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 32946 8192 33262 8193
rect 32946 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33262 8192
rect 32946 8127 33262 8128
rect 42946 8192 43262 8193
rect 42946 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43262 8192
rect 42946 8127 43262 8128
rect 1393 8122 1459 8125
rect 0 8120 1459 8122
rect 0 8064 1398 8120
rect 1454 8064 1459 8120
rect 0 8062 1459 8064
rect 0 8032 800 8062
rect 1393 8059 1459 8062
rect 46841 7986 46907 7989
rect 50200 7986 51000 8016
rect 46841 7984 51000 7986
rect 46841 7928 46846 7984
rect 46902 7928 51000 7984
rect 46841 7926 51000 7928
rect 46841 7923 46907 7926
rect 50200 7896 51000 7926
rect 0 7714 800 7744
rect 1301 7714 1367 7717
rect 0 7712 1367 7714
rect 0 7656 1306 7712
rect 1362 7656 1367 7712
rect 0 7654 1367 7656
rect 0 7624 800 7654
rect 1301 7651 1367 7654
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 17946 7583 18262 7584
rect 27946 7648 28262 7649
rect 27946 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28262 7648
rect 27946 7583 28262 7584
rect 37946 7648 38262 7649
rect 37946 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38262 7648
rect 37946 7583 38262 7584
rect 47946 7648 48262 7649
rect 47946 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48262 7648
rect 47946 7583 48262 7584
rect 49141 7578 49207 7581
rect 50200 7578 51000 7608
rect 49141 7576 51000 7578
rect 49141 7520 49146 7576
rect 49202 7520 51000 7576
rect 49141 7518 51000 7520
rect 49141 7515 49207 7518
rect 50200 7488 51000 7518
rect 0 7306 800 7336
rect 1301 7306 1367 7309
rect 0 7304 1367 7306
rect 0 7248 1306 7304
rect 1362 7248 1367 7304
rect 0 7246 1367 7248
rect 0 7216 800 7246
rect 1301 7243 1367 7246
rect 49233 7170 49299 7173
rect 50200 7170 51000 7200
rect 49233 7168 51000 7170
rect 49233 7112 49238 7168
rect 49294 7112 51000 7168
rect 49233 7110 51000 7112
rect 49233 7107 49299 7110
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 32946 7104 33262 7105
rect 32946 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33262 7104
rect 32946 7039 33262 7040
rect 42946 7104 43262 7105
rect 42946 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43262 7104
rect 50200 7080 51000 7110
rect 42946 7039 43262 7040
rect 0 6898 800 6928
rect 1209 6898 1275 6901
rect 0 6896 1275 6898
rect 0 6840 1214 6896
rect 1270 6840 1275 6896
rect 0 6838 1275 6840
rect 0 6808 800 6838
rect 1209 6835 1275 6838
rect 49417 6762 49483 6765
rect 50200 6762 51000 6792
rect 49417 6760 51000 6762
rect 49417 6704 49422 6760
rect 49478 6704 51000 6760
rect 49417 6702 51000 6704
rect 49417 6699 49483 6702
rect 50200 6672 51000 6702
rect 7946 6560 8262 6561
rect 0 6490 800 6520
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 27946 6560 28262 6561
rect 27946 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28262 6560
rect 27946 6495 28262 6496
rect 37946 6560 38262 6561
rect 37946 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38262 6560
rect 37946 6495 38262 6496
rect 47946 6560 48262 6561
rect 47946 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48262 6560
rect 47946 6495 48262 6496
rect 1301 6490 1367 6493
rect 0 6488 1367 6490
rect 0 6432 1306 6488
rect 1362 6432 1367 6488
rect 0 6430 1367 6432
rect 0 6400 800 6430
rect 1301 6427 1367 6430
rect 48865 6354 48931 6357
rect 50200 6354 51000 6384
rect 48865 6352 51000 6354
rect 48865 6296 48870 6352
rect 48926 6296 51000 6352
rect 48865 6294 51000 6296
rect 48865 6291 48931 6294
rect 50200 6264 51000 6294
rect 0 6082 800 6112
rect 1301 6082 1367 6085
rect 0 6080 1367 6082
rect 0 6024 1306 6080
rect 1362 6024 1367 6080
rect 0 6022 1367 6024
rect 0 5992 800 6022
rect 1301 6019 1367 6022
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 22946 5951 23262 5952
rect 32946 6016 33262 6017
rect 32946 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33262 6016
rect 32946 5951 33262 5952
rect 42946 6016 43262 6017
rect 42946 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43262 6016
rect 42946 5951 43262 5952
rect 49141 5946 49207 5949
rect 50200 5946 51000 5976
rect 49141 5944 51000 5946
rect 49141 5888 49146 5944
rect 49202 5888 51000 5944
rect 49141 5886 51000 5888
rect 49141 5883 49207 5886
rect 50200 5856 51000 5886
rect 0 5674 800 5704
rect 1301 5674 1367 5677
rect 0 5672 1367 5674
rect 0 5616 1306 5672
rect 1362 5616 1367 5672
rect 0 5614 1367 5616
rect 0 5584 800 5614
rect 1301 5611 1367 5614
rect 49417 5538 49483 5541
rect 50200 5538 51000 5568
rect 49417 5536 51000 5538
rect 49417 5480 49422 5536
rect 49478 5480 51000 5536
rect 49417 5478 51000 5480
rect 49417 5475 49483 5478
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 27946 5472 28262 5473
rect 27946 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28262 5472
rect 27946 5407 28262 5408
rect 37946 5472 38262 5473
rect 37946 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38262 5472
rect 37946 5407 38262 5408
rect 47946 5472 48262 5473
rect 47946 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48262 5472
rect 50200 5448 51000 5478
rect 47946 5407 48262 5408
rect 0 5266 800 5296
rect 2773 5266 2839 5269
rect 0 5264 2839 5266
rect 0 5208 2778 5264
rect 2834 5208 2839 5264
rect 0 5206 2839 5208
rect 0 5176 800 5206
rect 2773 5203 2839 5206
rect 49325 5130 49391 5133
rect 50200 5130 51000 5160
rect 49325 5128 51000 5130
rect 49325 5072 49330 5128
rect 49386 5072 51000 5128
rect 49325 5070 51000 5072
rect 49325 5067 49391 5070
rect 50200 5040 51000 5070
rect 2946 4928 3262 4929
rect 0 4858 800 4888
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 32946 4928 33262 4929
rect 32946 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33262 4928
rect 32946 4863 33262 4864
rect 42946 4928 43262 4929
rect 42946 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43262 4928
rect 42946 4863 43262 4864
rect 1301 4858 1367 4861
rect 0 4856 1367 4858
rect 0 4800 1306 4856
rect 1362 4800 1367 4856
rect 0 4798 1367 4800
rect 0 4768 800 4798
rect 1301 4795 1367 4798
rect 48313 4722 48379 4725
rect 50200 4722 51000 4752
rect 48313 4720 51000 4722
rect 48313 4664 48318 4720
rect 48374 4664 51000 4720
rect 48313 4662 51000 4664
rect 48313 4659 48379 4662
rect 50200 4632 51000 4662
rect 0 4450 800 4480
rect 1301 4450 1367 4453
rect 0 4448 1367 4450
rect 0 4392 1306 4448
rect 1362 4392 1367 4448
rect 0 4390 1367 4392
rect 0 4360 800 4390
rect 1301 4387 1367 4390
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 17946 4319 18262 4320
rect 27946 4384 28262 4385
rect 27946 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28262 4384
rect 27946 4319 28262 4320
rect 37946 4384 38262 4385
rect 37946 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38262 4384
rect 37946 4319 38262 4320
rect 47946 4384 48262 4385
rect 47946 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48262 4384
rect 47946 4319 48262 4320
rect 49141 4314 49207 4317
rect 50200 4314 51000 4344
rect 49141 4312 51000 4314
rect 49141 4256 49146 4312
rect 49202 4256 51000 4312
rect 49141 4254 51000 4256
rect 49141 4251 49207 4254
rect 50200 4224 51000 4254
rect 0 4042 800 4072
rect 1393 4042 1459 4045
rect 0 4040 1459 4042
rect 0 3984 1398 4040
rect 1454 3984 1459 4040
rect 0 3982 1459 3984
rect 0 3952 800 3982
rect 1393 3979 1459 3982
rect 5349 4042 5415 4045
rect 25405 4042 25471 4045
rect 5349 4040 25471 4042
rect 5349 3984 5354 4040
rect 5410 3984 25410 4040
rect 25466 3984 25471 4040
rect 5349 3982 25471 3984
rect 5349 3979 5415 3982
rect 25405 3979 25471 3982
rect 49233 3906 49299 3909
rect 50200 3906 51000 3936
rect 49233 3904 51000 3906
rect 49233 3848 49238 3904
rect 49294 3848 51000 3904
rect 49233 3846 51000 3848
rect 49233 3843 49299 3846
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 32946 3840 33262 3841
rect 32946 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33262 3840
rect 32946 3775 33262 3776
rect 42946 3840 43262 3841
rect 42946 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43262 3840
rect 50200 3816 51000 3846
rect 42946 3775 43262 3776
rect 0 3634 800 3664
rect 1301 3634 1367 3637
rect 0 3632 1367 3634
rect 0 3576 1306 3632
rect 1362 3576 1367 3632
rect 0 3574 1367 3576
rect 0 3544 800 3574
rect 1301 3571 1367 3574
rect 1117 3498 1183 3501
rect 26049 3498 26115 3501
rect 1117 3496 26115 3498
rect 1117 3440 1122 3496
rect 1178 3440 26054 3496
rect 26110 3440 26115 3496
rect 1117 3438 26115 3440
rect 1117 3435 1183 3438
rect 26049 3435 26115 3438
rect 49141 3498 49207 3501
rect 50200 3498 51000 3528
rect 49141 3496 51000 3498
rect 49141 3440 49146 3496
rect 49202 3440 51000 3496
rect 49141 3438 51000 3440
rect 49141 3435 49207 3438
rect 50200 3408 51000 3438
rect 7946 3296 8262 3297
rect 0 3226 800 3256
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 27946 3296 28262 3297
rect 27946 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28262 3296
rect 27946 3231 28262 3232
rect 37946 3296 38262 3297
rect 37946 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38262 3296
rect 37946 3231 38262 3232
rect 47946 3296 48262 3297
rect 47946 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48262 3296
rect 47946 3231 48262 3232
rect 1301 3226 1367 3229
rect 0 3224 1367 3226
rect 0 3168 1306 3224
rect 1362 3168 1367 3224
rect 0 3166 1367 3168
rect 0 3136 800 3166
rect 1301 3163 1367 3166
rect 48681 3090 48747 3093
rect 50200 3090 51000 3120
rect 48681 3088 51000 3090
rect 48681 3032 48686 3088
rect 48742 3032 51000 3088
rect 48681 3030 51000 3032
rect 48681 3027 48747 3030
rect 50200 3000 51000 3030
rect 0 2818 800 2848
rect 1301 2818 1367 2821
rect 0 2816 1367 2818
rect 0 2760 1306 2816
rect 1362 2760 1367 2816
rect 0 2758 1367 2760
rect 0 2728 800 2758
rect 1301 2755 1367 2758
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 22946 2687 23262 2688
rect 32946 2752 33262 2753
rect 32946 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33262 2752
rect 32946 2687 33262 2688
rect 42946 2752 43262 2753
rect 42946 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43262 2752
rect 42946 2687 43262 2688
rect 46841 2682 46907 2685
rect 50200 2682 51000 2712
rect 46841 2680 51000 2682
rect 46841 2624 46846 2680
rect 46902 2624 51000 2680
rect 46841 2622 51000 2624
rect 46841 2619 46907 2622
rect 50200 2592 51000 2622
rect 0 2410 800 2440
rect 1301 2410 1367 2413
rect 0 2408 1367 2410
rect 0 2352 1306 2408
rect 1362 2352 1367 2408
rect 0 2350 1367 2352
rect 0 2320 800 2350
rect 1301 2347 1367 2350
rect 48497 2274 48563 2277
rect 50200 2274 51000 2304
rect 48497 2272 51000 2274
rect 48497 2216 48502 2272
rect 48558 2216 51000 2272
rect 48497 2214 51000 2216
rect 48497 2211 48563 2214
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 27946 2208 28262 2209
rect 27946 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28262 2208
rect 27946 2143 28262 2144
rect 37946 2208 38262 2209
rect 37946 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38262 2208
rect 37946 2143 38262 2144
rect 47946 2208 48262 2209
rect 47946 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48262 2208
rect 50200 2184 51000 2214
rect 47946 2143 48262 2144
rect 0 2002 800 2032
rect 1209 2002 1275 2005
rect 0 2000 1275 2002
rect 0 1944 1214 2000
rect 1270 1944 1275 2000
rect 0 1942 1275 1944
rect 0 1912 800 1942
rect 1209 1939 1275 1942
rect 46749 1866 46815 1869
rect 50200 1866 51000 1896
rect 46749 1864 51000 1866
rect 46749 1808 46754 1864
rect 46810 1808 51000 1864
rect 46749 1806 51000 1808
rect 46749 1803 46815 1806
rect 50200 1776 51000 1806
rect 0 1594 800 1624
rect 1301 1594 1367 1597
rect 0 1592 1367 1594
rect 0 1536 1306 1592
rect 1362 1536 1367 1592
rect 0 1534 1367 1536
rect 0 1504 800 1534
rect 1301 1531 1367 1534
rect 46657 1458 46723 1461
rect 50200 1458 51000 1488
rect 46657 1456 51000 1458
rect 46657 1400 46662 1456
rect 46718 1400 51000 1456
rect 46657 1398 51000 1400
rect 46657 1395 46723 1398
rect 50200 1368 51000 1398
<< via3 >>
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 32952 24508 33016 24512
rect 32952 24452 32956 24508
rect 32956 24452 33012 24508
rect 33012 24452 33016 24508
rect 32952 24448 33016 24452
rect 33032 24508 33096 24512
rect 33032 24452 33036 24508
rect 33036 24452 33092 24508
rect 33092 24452 33096 24508
rect 33032 24448 33096 24452
rect 33112 24508 33176 24512
rect 33112 24452 33116 24508
rect 33116 24452 33172 24508
rect 33172 24452 33176 24508
rect 33112 24448 33176 24452
rect 33192 24508 33256 24512
rect 33192 24452 33196 24508
rect 33196 24452 33252 24508
rect 33252 24452 33256 24508
rect 33192 24448 33256 24452
rect 42952 24508 43016 24512
rect 42952 24452 42956 24508
rect 42956 24452 43012 24508
rect 43012 24452 43016 24508
rect 42952 24448 43016 24452
rect 43032 24508 43096 24512
rect 43032 24452 43036 24508
rect 43036 24452 43092 24508
rect 43092 24452 43096 24508
rect 43032 24448 43096 24452
rect 43112 24508 43176 24512
rect 43112 24452 43116 24508
rect 43116 24452 43172 24508
rect 43172 24452 43176 24508
rect 43112 24448 43176 24452
rect 43192 24508 43256 24512
rect 43192 24452 43196 24508
rect 43196 24452 43252 24508
rect 43252 24452 43256 24508
rect 43192 24448 43256 24452
rect 28948 23972 29012 24036
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 27952 23964 28016 23968
rect 27952 23908 27956 23964
rect 27956 23908 28012 23964
rect 28012 23908 28016 23964
rect 27952 23904 28016 23908
rect 28032 23964 28096 23968
rect 28032 23908 28036 23964
rect 28036 23908 28092 23964
rect 28092 23908 28096 23964
rect 28032 23904 28096 23908
rect 28112 23964 28176 23968
rect 28112 23908 28116 23964
rect 28116 23908 28172 23964
rect 28172 23908 28176 23964
rect 28112 23904 28176 23908
rect 28192 23964 28256 23968
rect 28192 23908 28196 23964
rect 28196 23908 28252 23964
rect 28252 23908 28256 23964
rect 28192 23904 28256 23908
rect 37952 23964 38016 23968
rect 37952 23908 37956 23964
rect 37956 23908 38012 23964
rect 38012 23908 38016 23964
rect 37952 23904 38016 23908
rect 38032 23964 38096 23968
rect 38032 23908 38036 23964
rect 38036 23908 38092 23964
rect 38092 23908 38096 23964
rect 38032 23904 38096 23908
rect 38112 23964 38176 23968
rect 38112 23908 38116 23964
rect 38116 23908 38172 23964
rect 38172 23908 38176 23964
rect 38112 23904 38176 23908
rect 38192 23964 38256 23968
rect 38192 23908 38196 23964
rect 38196 23908 38252 23964
rect 38252 23908 38256 23964
rect 38192 23904 38256 23908
rect 47952 23964 48016 23968
rect 47952 23908 47956 23964
rect 47956 23908 48012 23964
rect 48012 23908 48016 23964
rect 47952 23904 48016 23908
rect 48032 23964 48096 23968
rect 48032 23908 48036 23964
rect 48036 23908 48092 23964
rect 48092 23908 48096 23964
rect 48032 23904 48096 23908
rect 48112 23964 48176 23968
rect 48112 23908 48116 23964
rect 48116 23908 48172 23964
rect 48172 23908 48176 23964
rect 48112 23904 48176 23908
rect 48192 23964 48256 23968
rect 48192 23908 48196 23964
rect 48196 23908 48252 23964
rect 48252 23908 48256 23964
rect 48192 23904 48256 23908
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 32952 23420 33016 23424
rect 32952 23364 32956 23420
rect 32956 23364 33012 23420
rect 33012 23364 33016 23420
rect 32952 23360 33016 23364
rect 33032 23420 33096 23424
rect 33032 23364 33036 23420
rect 33036 23364 33092 23420
rect 33092 23364 33096 23420
rect 33032 23360 33096 23364
rect 33112 23420 33176 23424
rect 33112 23364 33116 23420
rect 33116 23364 33172 23420
rect 33172 23364 33176 23420
rect 33112 23360 33176 23364
rect 33192 23420 33256 23424
rect 33192 23364 33196 23420
rect 33196 23364 33252 23420
rect 33252 23364 33256 23420
rect 33192 23360 33256 23364
rect 42952 23420 43016 23424
rect 42952 23364 42956 23420
rect 42956 23364 43012 23420
rect 43012 23364 43016 23420
rect 42952 23360 43016 23364
rect 43032 23420 43096 23424
rect 43032 23364 43036 23420
rect 43036 23364 43092 23420
rect 43092 23364 43096 23420
rect 43032 23360 43096 23364
rect 43112 23420 43176 23424
rect 43112 23364 43116 23420
rect 43116 23364 43172 23420
rect 43172 23364 43176 23420
rect 43112 23360 43176 23364
rect 43192 23420 43256 23424
rect 43192 23364 43196 23420
rect 43196 23364 43252 23420
rect 43252 23364 43256 23420
rect 43192 23360 43256 23364
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 27952 22876 28016 22880
rect 27952 22820 27956 22876
rect 27956 22820 28012 22876
rect 28012 22820 28016 22876
rect 27952 22816 28016 22820
rect 28032 22876 28096 22880
rect 28032 22820 28036 22876
rect 28036 22820 28092 22876
rect 28092 22820 28096 22876
rect 28032 22816 28096 22820
rect 28112 22876 28176 22880
rect 28112 22820 28116 22876
rect 28116 22820 28172 22876
rect 28172 22820 28176 22876
rect 28112 22816 28176 22820
rect 28192 22876 28256 22880
rect 28192 22820 28196 22876
rect 28196 22820 28252 22876
rect 28252 22820 28256 22876
rect 28192 22816 28256 22820
rect 37952 22876 38016 22880
rect 37952 22820 37956 22876
rect 37956 22820 38012 22876
rect 38012 22820 38016 22876
rect 37952 22816 38016 22820
rect 38032 22876 38096 22880
rect 38032 22820 38036 22876
rect 38036 22820 38092 22876
rect 38092 22820 38096 22876
rect 38032 22816 38096 22820
rect 38112 22876 38176 22880
rect 38112 22820 38116 22876
rect 38116 22820 38172 22876
rect 38172 22820 38176 22876
rect 38112 22816 38176 22820
rect 38192 22876 38256 22880
rect 38192 22820 38196 22876
rect 38196 22820 38252 22876
rect 38252 22820 38256 22876
rect 38192 22816 38256 22820
rect 47952 22876 48016 22880
rect 47952 22820 47956 22876
rect 47956 22820 48012 22876
rect 48012 22820 48016 22876
rect 47952 22816 48016 22820
rect 48032 22876 48096 22880
rect 48032 22820 48036 22876
rect 48036 22820 48092 22876
rect 48092 22820 48096 22876
rect 48032 22816 48096 22820
rect 48112 22876 48176 22880
rect 48112 22820 48116 22876
rect 48116 22820 48172 22876
rect 48172 22820 48176 22876
rect 48112 22816 48176 22820
rect 48192 22876 48256 22880
rect 48192 22820 48196 22876
rect 48196 22820 48252 22876
rect 48252 22820 48256 22876
rect 48192 22816 48256 22820
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 32952 22332 33016 22336
rect 32952 22276 32956 22332
rect 32956 22276 33012 22332
rect 33012 22276 33016 22332
rect 32952 22272 33016 22276
rect 33032 22332 33096 22336
rect 33032 22276 33036 22332
rect 33036 22276 33092 22332
rect 33092 22276 33096 22332
rect 33032 22272 33096 22276
rect 33112 22332 33176 22336
rect 33112 22276 33116 22332
rect 33116 22276 33172 22332
rect 33172 22276 33176 22332
rect 33112 22272 33176 22276
rect 33192 22332 33256 22336
rect 33192 22276 33196 22332
rect 33196 22276 33252 22332
rect 33252 22276 33256 22332
rect 33192 22272 33256 22276
rect 42952 22332 43016 22336
rect 42952 22276 42956 22332
rect 42956 22276 43012 22332
rect 43012 22276 43016 22332
rect 42952 22272 43016 22276
rect 43032 22332 43096 22336
rect 43032 22276 43036 22332
rect 43036 22276 43092 22332
rect 43092 22276 43096 22332
rect 43032 22272 43096 22276
rect 43112 22332 43176 22336
rect 43112 22276 43116 22332
rect 43116 22276 43172 22332
rect 43172 22276 43176 22332
rect 43112 22272 43176 22276
rect 43192 22332 43256 22336
rect 43192 22276 43196 22332
rect 43196 22276 43252 22332
rect 43252 22276 43256 22332
rect 43192 22272 43256 22276
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 27952 21788 28016 21792
rect 27952 21732 27956 21788
rect 27956 21732 28012 21788
rect 28012 21732 28016 21788
rect 27952 21728 28016 21732
rect 28032 21788 28096 21792
rect 28032 21732 28036 21788
rect 28036 21732 28092 21788
rect 28092 21732 28096 21788
rect 28032 21728 28096 21732
rect 28112 21788 28176 21792
rect 28112 21732 28116 21788
rect 28116 21732 28172 21788
rect 28172 21732 28176 21788
rect 28112 21728 28176 21732
rect 28192 21788 28256 21792
rect 28192 21732 28196 21788
rect 28196 21732 28252 21788
rect 28252 21732 28256 21788
rect 28192 21728 28256 21732
rect 37952 21788 38016 21792
rect 37952 21732 37956 21788
rect 37956 21732 38012 21788
rect 38012 21732 38016 21788
rect 37952 21728 38016 21732
rect 38032 21788 38096 21792
rect 38032 21732 38036 21788
rect 38036 21732 38092 21788
rect 38092 21732 38096 21788
rect 38032 21728 38096 21732
rect 38112 21788 38176 21792
rect 38112 21732 38116 21788
rect 38116 21732 38172 21788
rect 38172 21732 38176 21788
rect 38112 21728 38176 21732
rect 38192 21788 38256 21792
rect 38192 21732 38196 21788
rect 38196 21732 38252 21788
rect 38252 21732 38256 21788
rect 38192 21728 38256 21732
rect 47952 21788 48016 21792
rect 47952 21732 47956 21788
rect 47956 21732 48012 21788
rect 48012 21732 48016 21788
rect 47952 21728 48016 21732
rect 48032 21788 48096 21792
rect 48032 21732 48036 21788
rect 48036 21732 48092 21788
rect 48092 21732 48096 21788
rect 48032 21728 48096 21732
rect 48112 21788 48176 21792
rect 48112 21732 48116 21788
rect 48116 21732 48172 21788
rect 48172 21732 48176 21788
rect 48112 21728 48176 21732
rect 48192 21788 48256 21792
rect 48192 21732 48196 21788
rect 48196 21732 48252 21788
rect 48252 21732 48256 21788
rect 48192 21728 48256 21732
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 32952 21244 33016 21248
rect 32952 21188 32956 21244
rect 32956 21188 33012 21244
rect 33012 21188 33016 21244
rect 32952 21184 33016 21188
rect 33032 21244 33096 21248
rect 33032 21188 33036 21244
rect 33036 21188 33092 21244
rect 33092 21188 33096 21244
rect 33032 21184 33096 21188
rect 33112 21244 33176 21248
rect 33112 21188 33116 21244
rect 33116 21188 33172 21244
rect 33172 21188 33176 21244
rect 33112 21184 33176 21188
rect 33192 21244 33256 21248
rect 33192 21188 33196 21244
rect 33196 21188 33252 21244
rect 33252 21188 33256 21244
rect 33192 21184 33256 21188
rect 42952 21244 43016 21248
rect 42952 21188 42956 21244
rect 42956 21188 43012 21244
rect 43012 21188 43016 21244
rect 42952 21184 43016 21188
rect 43032 21244 43096 21248
rect 43032 21188 43036 21244
rect 43036 21188 43092 21244
rect 43092 21188 43096 21244
rect 43032 21184 43096 21188
rect 43112 21244 43176 21248
rect 43112 21188 43116 21244
rect 43116 21188 43172 21244
rect 43172 21188 43176 21244
rect 43112 21184 43176 21188
rect 43192 21244 43256 21248
rect 43192 21188 43196 21244
rect 43196 21188 43252 21244
rect 43252 21188 43256 21244
rect 43192 21184 43256 21188
rect 28764 20980 28828 21044
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 27952 20700 28016 20704
rect 27952 20644 27956 20700
rect 27956 20644 28012 20700
rect 28012 20644 28016 20700
rect 27952 20640 28016 20644
rect 28032 20700 28096 20704
rect 28032 20644 28036 20700
rect 28036 20644 28092 20700
rect 28092 20644 28096 20700
rect 28032 20640 28096 20644
rect 28112 20700 28176 20704
rect 28112 20644 28116 20700
rect 28116 20644 28172 20700
rect 28172 20644 28176 20700
rect 28112 20640 28176 20644
rect 28192 20700 28256 20704
rect 28192 20644 28196 20700
rect 28196 20644 28252 20700
rect 28252 20644 28256 20700
rect 28192 20640 28256 20644
rect 37952 20700 38016 20704
rect 37952 20644 37956 20700
rect 37956 20644 38012 20700
rect 38012 20644 38016 20700
rect 37952 20640 38016 20644
rect 38032 20700 38096 20704
rect 38032 20644 38036 20700
rect 38036 20644 38092 20700
rect 38092 20644 38096 20700
rect 38032 20640 38096 20644
rect 38112 20700 38176 20704
rect 38112 20644 38116 20700
rect 38116 20644 38172 20700
rect 38172 20644 38176 20700
rect 38112 20640 38176 20644
rect 38192 20700 38256 20704
rect 38192 20644 38196 20700
rect 38196 20644 38252 20700
rect 38252 20644 38256 20700
rect 38192 20640 38256 20644
rect 47952 20700 48016 20704
rect 47952 20644 47956 20700
rect 47956 20644 48012 20700
rect 48012 20644 48016 20700
rect 47952 20640 48016 20644
rect 48032 20700 48096 20704
rect 48032 20644 48036 20700
rect 48036 20644 48092 20700
rect 48092 20644 48096 20700
rect 48032 20640 48096 20644
rect 48112 20700 48176 20704
rect 48112 20644 48116 20700
rect 48116 20644 48172 20700
rect 48172 20644 48176 20700
rect 48112 20640 48176 20644
rect 48192 20700 48256 20704
rect 48192 20644 48196 20700
rect 48196 20644 48252 20700
rect 48252 20644 48256 20700
rect 48192 20640 48256 20644
rect 28580 20572 28644 20636
rect 28396 20164 28460 20228
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 32952 20156 33016 20160
rect 32952 20100 32956 20156
rect 32956 20100 33012 20156
rect 33012 20100 33016 20156
rect 32952 20096 33016 20100
rect 33032 20156 33096 20160
rect 33032 20100 33036 20156
rect 33036 20100 33092 20156
rect 33092 20100 33096 20156
rect 33032 20096 33096 20100
rect 33112 20156 33176 20160
rect 33112 20100 33116 20156
rect 33116 20100 33172 20156
rect 33172 20100 33176 20156
rect 33112 20096 33176 20100
rect 33192 20156 33256 20160
rect 33192 20100 33196 20156
rect 33196 20100 33252 20156
rect 33252 20100 33256 20156
rect 33192 20096 33256 20100
rect 42952 20156 43016 20160
rect 42952 20100 42956 20156
rect 42956 20100 43012 20156
rect 43012 20100 43016 20156
rect 42952 20096 43016 20100
rect 43032 20156 43096 20160
rect 43032 20100 43036 20156
rect 43036 20100 43092 20156
rect 43092 20100 43096 20156
rect 43032 20096 43096 20100
rect 43112 20156 43176 20160
rect 43112 20100 43116 20156
rect 43116 20100 43172 20156
rect 43172 20100 43176 20156
rect 43112 20096 43176 20100
rect 43192 20156 43256 20160
rect 43192 20100 43196 20156
rect 43196 20100 43252 20156
rect 43252 20100 43256 20156
rect 43192 20096 43256 20100
rect 28580 19680 28644 19684
rect 28580 19624 28594 19680
rect 28594 19624 28644 19680
rect 28580 19620 28644 19624
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 27952 19612 28016 19616
rect 27952 19556 27956 19612
rect 27956 19556 28012 19612
rect 28012 19556 28016 19612
rect 27952 19552 28016 19556
rect 28032 19612 28096 19616
rect 28032 19556 28036 19612
rect 28036 19556 28092 19612
rect 28092 19556 28096 19612
rect 28032 19552 28096 19556
rect 28112 19612 28176 19616
rect 28112 19556 28116 19612
rect 28116 19556 28172 19612
rect 28172 19556 28176 19612
rect 28112 19552 28176 19556
rect 28192 19612 28256 19616
rect 28192 19556 28196 19612
rect 28196 19556 28252 19612
rect 28252 19556 28256 19612
rect 28192 19552 28256 19556
rect 28764 19544 28828 19548
rect 28764 19488 28814 19544
rect 28814 19488 28828 19544
rect 28764 19484 28828 19488
rect 37952 19612 38016 19616
rect 37952 19556 37956 19612
rect 37956 19556 38012 19612
rect 38012 19556 38016 19612
rect 37952 19552 38016 19556
rect 38032 19612 38096 19616
rect 38032 19556 38036 19612
rect 38036 19556 38092 19612
rect 38092 19556 38096 19612
rect 38032 19552 38096 19556
rect 38112 19612 38176 19616
rect 38112 19556 38116 19612
rect 38116 19556 38172 19612
rect 38172 19556 38176 19612
rect 38112 19552 38176 19556
rect 38192 19612 38256 19616
rect 38192 19556 38196 19612
rect 38196 19556 38252 19612
rect 38252 19556 38256 19612
rect 38192 19552 38256 19556
rect 47952 19612 48016 19616
rect 47952 19556 47956 19612
rect 47956 19556 48012 19612
rect 48012 19556 48016 19612
rect 47952 19552 48016 19556
rect 48032 19612 48096 19616
rect 48032 19556 48036 19612
rect 48036 19556 48092 19612
rect 48092 19556 48096 19612
rect 48032 19552 48096 19556
rect 48112 19612 48176 19616
rect 48112 19556 48116 19612
rect 48116 19556 48172 19612
rect 48172 19556 48176 19612
rect 48112 19552 48176 19556
rect 48192 19612 48256 19616
rect 48192 19556 48196 19612
rect 48196 19556 48252 19612
rect 48252 19556 48256 19612
rect 48192 19552 48256 19556
rect 28396 19212 28460 19276
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 32952 19068 33016 19072
rect 32952 19012 32956 19068
rect 32956 19012 33012 19068
rect 33012 19012 33016 19068
rect 32952 19008 33016 19012
rect 33032 19068 33096 19072
rect 33032 19012 33036 19068
rect 33036 19012 33092 19068
rect 33092 19012 33096 19068
rect 33032 19008 33096 19012
rect 33112 19068 33176 19072
rect 33112 19012 33116 19068
rect 33116 19012 33172 19068
rect 33172 19012 33176 19068
rect 33112 19008 33176 19012
rect 33192 19068 33256 19072
rect 33192 19012 33196 19068
rect 33196 19012 33252 19068
rect 33252 19012 33256 19068
rect 33192 19008 33256 19012
rect 42952 19068 43016 19072
rect 42952 19012 42956 19068
rect 42956 19012 43012 19068
rect 43012 19012 43016 19068
rect 42952 19008 43016 19012
rect 43032 19068 43096 19072
rect 43032 19012 43036 19068
rect 43036 19012 43092 19068
rect 43092 19012 43096 19068
rect 43032 19008 43096 19012
rect 43112 19068 43176 19072
rect 43112 19012 43116 19068
rect 43116 19012 43172 19068
rect 43172 19012 43176 19068
rect 43112 19008 43176 19012
rect 43192 19068 43256 19072
rect 43192 19012 43196 19068
rect 43196 19012 43252 19068
rect 43252 19012 43256 19068
rect 43192 19008 43256 19012
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 27952 18524 28016 18528
rect 27952 18468 27956 18524
rect 27956 18468 28012 18524
rect 28012 18468 28016 18524
rect 27952 18464 28016 18468
rect 28032 18524 28096 18528
rect 28032 18468 28036 18524
rect 28036 18468 28092 18524
rect 28092 18468 28096 18524
rect 28032 18464 28096 18468
rect 28112 18524 28176 18528
rect 28112 18468 28116 18524
rect 28116 18468 28172 18524
rect 28172 18468 28176 18524
rect 28112 18464 28176 18468
rect 28192 18524 28256 18528
rect 28192 18468 28196 18524
rect 28196 18468 28252 18524
rect 28252 18468 28256 18524
rect 28192 18464 28256 18468
rect 37952 18524 38016 18528
rect 37952 18468 37956 18524
rect 37956 18468 38012 18524
rect 38012 18468 38016 18524
rect 37952 18464 38016 18468
rect 38032 18524 38096 18528
rect 38032 18468 38036 18524
rect 38036 18468 38092 18524
rect 38092 18468 38096 18524
rect 38032 18464 38096 18468
rect 38112 18524 38176 18528
rect 38112 18468 38116 18524
rect 38116 18468 38172 18524
rect 38172 18468 38176 18524
rect 38112 18464 38176 18468
rect 38192 18524 38256 18528
rect 38192 18468 38196 18524
rect 38196 18468 38252 18524
rect 38252 18468 38256 18524
rect 38192 18464 38256 18468
rect 47952 18524 48016 18528
rect 47952 18468 47956 18524
rect 47956 18468 48012 18524
rect 48012 18468 48016 18524
rect 47952 18464 48016 18468
rect 48032 18524 48096 18528
rect 48032 18468 48036 18524
rect 48036 18468 48092 18524
rect 48092 18468 48096 18524
rect 48032 18464 48096 18468
rect 48112 18524 48176 18528
rect 48112 18468 48116 18524
rect 48116 18468 48172 18524
rect 48172 18468 48176 18524
rect 48112 18464 48176 18468
rect 48192 18524 48256 18528
rect 48192 18468 48196 18524
rect 48196 18468 48252 18524
rect 48252 18468 48256 18524
rect 48192 18464 48256 18468
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 32952 17980 33016 17984
rect 32952 17924 32956 17980
rect 32956 17924 33012 17980
rect 33012 17924 33016 17980
rect 32952 17920 33016 17924
rect 33032 17980 33096 17984
rect 33032 17924 33036 17980
rect 33036 17924 33092 17980
rect 33092 17924 33096 17980
rect 33032 17920 33096 17924
rect 33112 17980 33176 17984
rect 33112 17924 33116 17980
rect 33116 17924 33172 17980
rect 33172 17924 33176 17980
rect 33112 17920 33176 17924
rect 33192 17980 33256 17984
rect 33192 17924 33196 17980
rect 33196 17924 33252 17980
rect 33252 17924 33256 17980
rect 33192 17920 33256 17924
rect 42952 17980 43016 17984
rect 42952 17924 42956 17980
rect 42956 17924 43012 17980
rect 43012 17924 43016 17980
rect 42952 17920 43016 17924
rect 43032 17980 43096 17984
rect 43032 17924 43036 17980
rect 43036 17924 43092 17980
rect 43092 17924 43096 17980
rect 43032 17920 43096 17924
rect 43112 17980 43176 17984
rect 43112 17924 43116 17980
rect 43116 17924 43172 17980
rect 43172 17924 43176 17980
rect 43112 17920 43176 17924
rect 43192 17980 43256 17984
rect 43192 17924 43196 17980
rect 43196 17924 43252 17980
rect 43252 17924 43256 17980
rect 43192 17920 43256 17924
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 27952 17436 28016 17440
rect 27952 17380 27956 17436
rect 27956 17380 28012 17436
rect 28012 17380 28016 17436
rect 27952 17376 28016 17380
rect 28032 17436 28096 17440
rect 28032 17380 28036 17436
rect 28036 17380 28092 17436
rect 28092 17380 28096 17436
rect 28032 17376 28096 17380
rect 28112 17436 28176 17440
rect 28112 17380 28116 17436
rect 28116 17380 28172 17436
rect 28172 17380 28176 17436
rect 28112 17376 28176 17380
rect 28192 17436 28256 17440
rect 28192 17380 28196 17436
rect 28196 17380 28252 17436
rect 28252 17380 28256 17436
rect 28192 17376 28256 17380
rect 37952 17436 38016 17440
rect 37952 17380 37956 17436
rect 37956 17380 38012 17436
rect 38012 17380 38016 17436
rect 37952 17376 38016 17380
rect 38032 17436 38096 17440
rect 38032 17380 38036 17436
rect 38036 17380 38092 17436
rect 38092 17380 38096 17436
rect 38032 17376 38096 17380
rect 38112 17436 38176 17440
rect 38112 17380 38116 17436
rect 38116 17380 38172 17436
rect 38172 17380 38176 17436
rect 38112 17376 38176 17380
rect 38192 17436 38256 17440
rect 38192 17380 38196 17436
rect 38196 17380 38252 17436
rect 38252 17380 38256 17436
rect 38192 17376 38256 17380
rect 47952 17436 48016 17440
rect 47952 17380 47956 17436
rect 47956 17380 48012 17436
rect 48012 17380 48016 17436
rect 47952 17376 48016 17380
rect 48032 17436 48096 17440
rect 48032 17380 48036 17436
rect 48036 17380 48092 17436
rect 48092 17380 48096 17436
rect 48032 17376 48096 17380
rect 48112 17436 48176 17440
rect 48112 17380 48116 17436
rect 48116 17380 48172 17436
rect 48172 17380 48176 17436
rect 48112 17376 48176 17380
rect 48192 17436 48256 17440
rect 48192 17380 48196 17436
rect 48196 17380 48252 17436
rect 48252 17380 48256 17436
rect 48192 17376 48256 17380
rect 14412 17036 14476 17100
rect 38516 17096 38580 17100
rect 38516 17040 38530 17096
rect 38530 17040 38580 17096
rect 38516 17036 38580 17040
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 32952 16892 33016 16896
rect 32952 16836 32956 16892
rect 32956 16836 33012 16892
rect 33012 16836 33016 16892
rect 32952 16832 33016 16836
rect 33032 16892 33096 16896
rect 33032 16836 33036 16892
rect 33036 16836 33092 16892
rect 33092 16836 33096 16892
rect 33032 16832 33096 16836
rect 33112 16892 33176 16896
rect 33112 16836 33116 16892
rect 33116 16836 33172 16892
rect 33172 16836 33176 16892
rect 33112 16832 33176 16836
rect 33192 16892 33256 16896
rect 33192 16836 33196 16892
rect 33196 16836 33252 16892
rect 33252 16836 33256 16892
rect 33192 16832 33256 16836
rect 42952 16892 43016 16896
rect 42952 16836 42956 16892
rect 42956 16836 43012 16892
rect 43012 16836 43016 16892
rect 42952 16832 43016 16836
rect 43032 16892 43096 16896
rect 43032 16836 43036 16892
rect 43036 16836 43092 16892
rect 43092 16836 43096 16892
rect 43032 16832 43096 16836
rect 43112 16892 43176 16896
rect 43112 16836 43116 16892
rect 43116 16836 43172 16892
rect 43172 16836 43176 16892
rect 43112 16832 43176 16836
rect 43192 16892 43256 16896
rect 43192 16836 43196 16892
rect 43196 16836 43252 16892
rect 43252 16836 43256 16892
rect 43192 16832 43256 16836
rect 28948 16764 29012 16828
rect 16068 16688 16132 16692
rect 16068 16632 16118 16688
rect 16118 16632 16132 16688
rect 16068 16628 16132 16632
rect 29132 16628 29196 16692
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 27952 16348 28016 16352
rect 27952 16292 27956 16348
rect 27956 16292 28012 16348
rect 28012 16292 28016 16348
rect 27952 16288 28016 16292
rect 28032 16348 28096 16352
rect 28032 16292 28036 16348
rect 28036 16292 28092 16348
rect 28092 16292 28096 16348
rect 28032 16288 28096 16292
rect 28112 16348 28176 16352
rect 28112 16292 28116 16348
rect 28116 16292 28172 16348
rect 28172 16292 28176 16348
rect 28112 16288 28176 16292
rect 28192 16348 28256 16352
rect 28192 16292 28196 16348
rect 28196 16292 28252 16348
rect 28252 16292 28256 16348
rect 28192 16288 28256 16292
rect 37952 16348 38016 16352
rect 37952 16292 37956 16348
rect 37956 16292 38012 16348
rect 38012 16292 38016 16348
rect 37952 16288 38016 16292
rect 38032 16348 38096 16352
rect 38032 16292 38036 16348
rect 38036 16292 38092 16348
rect 38092 16292 38096 16348
rect 38032 16288 38096 16292
rect 38112 16348 38176 16352
rect 38112 16292 38116 16348
rect 38116 16292 38172 16348
rect 38172 16292 38176 16348
rect 38112 16288 38176 16292
rect 38192 16348 38256 16352
rect 38192 16292 38196 16348
rect 38196 16292 38252 16348
rect 38252 16292 38256 16348
rect 38192 16288 38256 16292
rect 47952 16348 48016 16352
rect 47952 16292 47956 16348
rect 47956 16292 48012 16348
rect 48012 16292 48016 16348
rect 47952 16288 48016 16292
rect 48032 16348 48096 16352
rect 48032 16292 48036 16348
rect 48036 16292 48092 16348
rect 48092 16292 48096 16348
rect 48032 16288 48096 16292
rect 48112 16348 48176 16352
rect 48112 16292 48116 16348
rect 48116 16292 48172 16348
rect 48172 16292 48176 16348
rect 48112 16288 48176 16292
rect 48192 16348 48256 16352
rect 48192 16292 48196 16348
rect 48196 16292 48252 16348
rect 48252 16292 48256 16348
rect 48192 16288 48256 16292
rect 14044 16084 14108 16148
rect 16988 15872 17052 15876
rect 16988 15816 17002 15872
rect 17002 15816 17052 15872
rect 16988 15812 17052 15816
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 32952 15804 33016 15808
rect 32952 15748 32956 15804
rect 32956 15748 33012 15804
rect 33012 15748 33016 15804
rect 32952 15744 33016 15748
rect 33032 15804 33096 15808
rect 33032 15748 33036 15804
rect 33036 15748 33092 15804
rect 33092 15748 33096 15804
rect 33032 15744 33096 15748
rect 33112 15804 33176 15808
rect 33112 15748 33116 15804
rect 33116 15748 33172 15804
rect 33172 15748 33176 15804
rect 33112 15744 33176 15748
rect 33192 15804 33256 15808
rect 33192 15748 33196 15804
rect 33196 15748 33252 15804
rect 33252 15748 33256 15804
rect 33192 15744 33256 15748
rect 42952 15804 43016 15808
rect 42952 15748 42956 15804
rect 42956 15748 43012 15804
rect 43012 15748 43016 15804
rect 42952 15744 43016 15748
rect 43032 15804 43096 15808
rect 43032 15748 43036 15804
rect 43036 15748 43092 15804
rect 43092 15748 43096 15804
rect 43032 15744 43096 15748
rect 43112 15804 43176 15808
rect 43112 15748 43116 15804
rect 43116 15748 43172 15804
rect 43172 15748 43176 15804
rect 43112 15744 43176 15748
rect 43192 15804 43256 15808
rect 43192 15748 43196 15804
rect 43196 15748 43252 15804
rect 43252 15748 43256 15804
rect 43192 15744 43256 15748
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 27952 15260 28016 15264
rect 27952 15204 27956 15260
rect 27956 15204 28012 15260
rect 28012 15204 28016 15260
rect 27952 15200 28016 15204
rect 28032 15260 28096 15264
rect 28032 15204 28036 15260
rect 28036 15204 28092 15260
rect 28092 15204 28096 15260
rect 28032 15200 28096 15204
rect 28112 15260 28176 15264
rect 28112 15204 28116 15260
rect 28116 15204 28172 15260
rect 28172 15204 28176 15260
rect 28112 15200 28176 15204
rect 28192 15260 28256 15264
rect 28192 15204 28196 15260
rect 28196 15204 28252 15260
rect 28252 15204 28256 15260
rect 28192 15200 28256 15204
rect 37952 15260 38016 15264
rect 37952 15204 37956 15260
rect 37956 15204 38012 15260
rect 38012 15204 38016 15260
rect 37952 15200 38016 15204
rect 38032 15260 38096 15264
rect 38032 15204 38036 15260
rect 38036 15204 38092 15260
rect 38092 15204 38096 15260
rect 38032 15200 38096 15204
rect 38112 15260 38176 15264
rect 38112 15204 38116 15260
rect 38116 15204 38172 15260
rect 38172 15204 38176 15260
rect 38112 15200 38176 15204
rect 38192 15260 38256 15264
rect 38192 15204 38196 15260
rect 38196 15204 38252 15260
rect 38252 15204 38256 15260
rect 38192 15200 38256 15204
rect 47952 15260 48016 15264
rect 47952 15204 47956 15260
rect 47956 15204 48012 15260
rect 48012 15204 48016 15260
rect 47952 15200 48016 15204
rect 48032 15260 48096 15264
rect 48032 15204 48036 15260
rect 48036 15204 48092 15260
rect 48092 15204 48096 15260
rect 48032 15200 48096 15204
rect 48112 15260 48176 15264
rect 48112 15204 48116 15260
rect 48116 15204 48172 15260
rect 48172 15204 48176 15260
rect 48112 15200 48176 15204
rect 48192 15260 48256 15264
rect 48192 15204 48196 15260
rect 48196 15204 48252 15260
rect 48252 15204 48256 15260
rect 48192 15200 48256 15204
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 32952 14716 33016 14720
rect 32952 14660 32956 14716
rect 32956 14660 33012 14716
rect 33012 14660 33016 14716
rect 32952 14656 33016 14660
rect 33032 14716 33096 14720
rect 33032 14660 33036 14716
rect 33036 14660 33092 14716
rect 33092 14660 33096 14716
rect 33032 14656 33096 14660
rect 33112 14716 33176 14720
rect 33112 14660 33116 14716
rect 33116 14660 33172 14716
rect 33172 14660 33176 14716
rect 33112 14656 33176 14660
rect 33192 14716 33256 14720
rect 33192 14660 33196 14716
rect 33196 14660 33252 14716
rect 33252 14660 33256 14716
rect 33192 14656 33256 14660
rect 42952 14716 43016 14720
rect 42952 14660 42956 14716
rect 42956 14660 43012 14716
rect 43012 14660 43016 14716
rect 42952 14656 43016 14660
rect 43032 14716 43096 14720
rect 43032 14660 43036 14716
rect 43036 14660 43092 14716
rect 43092 14660 43096 14716
rect 43032 14656 43096 14660
rect 43112 14716 43176 14720
rect 43112 14660 43116 14716
rect 43116 14660 43172 14716
rect 43172 14660 43176 14716
rect 43112 14656 43176 14660
rect 43192 14716 43256 14720
rect 43192 14660 43196 14716
rect 43196 14660 43252 14716
rect 43252 14660 43256 14716
rect 43192 14656 43256 14660
rect 14228 14376 14292 14380
rect 14228 14320 14242 14376
rect 14242 14320 14292 14376
rect 14228 14316 14292 14320
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 27952 14172 28016 14176
rect 27952 14116 27956 14172
rect 27956 14116 28012 14172
rect 28012 14116 28016 14172
rect 27952 14112 28016 14116
rect 28032 14172 28096 14176
rect 28032 14116 28036 14172
rect 28036 14116 28092 14172
rect 28092 14116 28096 14172
rect 28032 14112 28096 14116
rect 28112 14172 28176 14176
rect 28112 14116 28116 14172
rect 28116 14116 28172 14172
rect 28172 14116 28176 14172
rect 28112 14112 28176 14116
rect 28192 14172 28256 14176
rect 28192 14116 28196 14172
rect 28196 14116 28252 14172
rect 28252 14116 28256 14172
rect 28192 14112 28256 14116
rect 37952 14172 38016 14176
rect 37952 14116 37956 14172
rect 37956 14116 38012 14172
rect 38012 14116 38016 14172
rect 37952 14112 38016 14116
rect 38032 14172 38096 14176
rect 38032 14116 38036 14172
rect 38036 14116 38092 14172
rect 38092 14116 38096 14172
rect 38032 14112 38096 14116
rect 38112 14172 38176 14176
rect 38112 14116 38116 14172
rect 38116 14116 38172 14172
rect 38172 14116 38176 14172
rect 38112 14112 38176 14116
rect 38192 14172 38256 14176
rect 38192 14116 38196 14172
rect 38196 14116 38252 14172
rect 38252 14116 38256 14172
rect 38192 14112 38256 14116
rect 47952 14172 48016 14176
rect 47952 14116 47956 14172
rect 47956 14116 48012 14172
rect 48012 14116 48016 14172
rect 47952 14112 48016 14116
rect 48032 14172 48096 14176
rect 48032 14116 48036 14172
rect 48036 14116 48092 14172
rect 48092 14116 48096 14172
rect 48032 14112 48096 14116
rect 48112 14172 48176 14176
rect 48112 14116 48116 14172
rect 48116 14116 48172 14172
rect 48172 14116 48176 14172
rect 48112 14112 48176 14116
rect 48192 14172 48256 14176
rect 48192 14116 48196 14172
rect 48196 14116 48252 14172
rect 48252 14116 48256 14172
rect 48192 14112 48256 14116
rect 16068 13636 16132 13700
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 32952 13628 33016 13632
rect 32952 13572 32956 13628
rect 32956 13572 33012 13628
rect 33012 13572 33016 13628
rect 32952 13568 33016 13572
rect 33032 13628 33096 13632
rect 33032 13572 33036 13628
rect 33036 13572 33092 13628
rect 33092 13572 33096 13628
rect 33032 13568 33096 13572
rect 33112 13628 33176 13632
rect 33112 13572 33116 13628
rect 33116 13572 33172 13628
rect 33172 13572 33176 13628
rect 33112 13568 33176 13572
rect 33192 13628 33256 13632
rect 33192 13572 33196 13628
rect 33196 13572 33252 13628
rect 33252 13572 33256 13628
rect 33192 13568 33256 13572
rect 42952 13628 43016 13632
rect 42952 13572 42956 13628
rect 42956 13572 43012 13628
rect 43012 13572 43016 13628
rect 42952 13568 43016 13572
rect 43032 13628 43096 13632
rect 43032 13572 43036 13628
rect 43036 13572 43092 13628
rect 43092 13572 43096 13628
rect 43032 13568 43096 13572
rect 43112 13628 43176 13632
rect 43112 13572 43116 13628
rect 43116 13572 43172 13628
rect 43172 13572 43176 13628
rect 43112 13568 43176 13572
rect 43192 13628 43256 13632
rect 43192 13572 43196 13628
rect 43196 13572 43252 13628
rect 43252 13572 43256 13628
rect 43192 13568 43256 13572
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 27952 13084 28016 13088
rect 27952 13028 27956 13084
rect 27956 13028 28012 13084
rect 28012 13028 28016 13084
rect 27952 13024 28016 13028
rect 28032 13084 28096 13088
rect 28032 13028 28036 13084
rect 28036 13028 28092 13084
rect 28092 13028 28096 13084
rect 28032 13024 28096 13028
rect 28112 13084 28176 13088
rect 28112 13028 28116 13084
rect 28116 13028 28172 13084
rect 28172 13028 28176 13084
rect 28112 13024 28176 13028
rect 28192 13084 28256 13088
rect 28192 13028 28196 13084
rect 28196 13028 28252 13084
rect 28252 13028 28256 13084
rect 28192 13024 28256 13028
rect 37952 13084 38016 13088
rect 37952 13028 37956 13084
rect 37956 13028 38012 13084
rect 38012 13028 38016 13084
rect 37952 13024 38016 13028
rect 38032 13084 38096 13088
rect 38032 13028 38036 13084
rect 38036 13028 38092 13084
rect 38092 13028 38096 13084
rect 38032 13024 38096 13028
rect 38112 13084 38176 13088
rect 38112 13028 38116 13084
rect 38116 13028 38172 13084
rect 38172 13028 38176 13084
rect 38112 13024 38176 13028
rect 38192 13084 38256 13088
rect 38192 13028 38196 13084
rect 38196 13028 38252 13084
rect 38252 13028 38256 13084
rect 38192 13024 38256 13028
rect 47952 13084 48016 13088
rect 47952 13028 47956 13084
rect 47956 13028 48012 13084
rect 48012 13028 48016 13084
rect 47952 13024 48016 13028
rect 48032 13084 48096 13088
rect 48032 13028 48036 13084
rect 48036 13028 48092 13084
rect 48092 13028 48096 13084
rect 48032 13024 48096 13028
rect 48112 13084 48176 13088
rect 48112 13028 48116 13084
rect 48116 13028 48172 13084
rect 48172 13028 48176 13084
rect 48112 13024 48176 13028
rect 48192 13084 48256 13088
rect 48192 13028 48196 13084
rect 48196 13028 48252 13084
rect 48252 13028 48256 13084
rect 48192 13024 48256 13028
rect 14412 12684 14476 12748
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 32952 12540 33016 12544
rect 32952 12484 32956 12540
rect 32956 12484 33012 12540
rect 33012 12484 33016 12540
rect 32952 12480 33016 12484
rect 33032 12540 33096 12544
rect 33032 12484 33036 12540
rect 33036 12484 33092 12540
rect 33092 12484 33096 12540
rect 33032 12480 33096 12484
rect 33112 12540 33176 12544
rect 33112 12484 33116 12540
rect 33116 12484 33172 12540
rect 33172 12484 33176 12540
rect 33112 12480 33176 12484
rect 33192 12540 33256 12544
rect 33192 12484 33196 12540
rect 33196 12484 33252 12540
rect 33252 12484 33256 12540
rect 33192 12480 33256 12484
rect 42952 12540 43016 12544
rect 42952 12484 42956 12540
rect 42956 12484 43012 12540
rect 43012 12484 43016 12540
rect 42952 12480 43016 12484
rect 43032 12540 43096 12544
rect 43032 12484 43036 12540
rect 43036 12484 43092 12540
rect 43092 12484 43096 12540
rect 43032 12480 43096 12484
rect 43112 12540 43176 12544
rect 43112 12484 43116 12540
rect 43116 12484 43172 12540
rect 43172 12484 43176 12540
rect 43112 12480 43176 12484
rect 43192 12540 43256 12544
rect 43192 12484 43196 12540
rect 43196 12484 43252 12540
rect 43252 12484 43256 12540
rect 43192 12480 43256 12484
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 27952 11996 28016 12000
rect 27952 11940 27956 11996
rect 27956 11940 28012 11996
rect 28012 11940 28016 11996
rect 27952 11936 28016 11940
rect 28032 11996 28096 12000
rect 28032 11940 28036 11996
rect 28036 11940 28092 11996
rect 28092 11940 28096 11996
rect 28032 11936 28096 11940
rect 28112 11996 28176 12000
rect 28112 11940 28116 11996
rect 28116 11940 28172 11996
rect 28172 11940 28176 11996
rect 28112 11936 28176 11940
rect 28192 11996 28256 12000
rect 28192 11940 28196 11996
rect 28196 11940 28252 11996
rect 28252 11940 28256 11996
rect 28192 11936 28256 11940
rect 37952 11996 38016 12000
rect 37952 11940 37956 11996
rect 37956 11940 38012 11996
rect 38012 11940 38016 11996
rect 37952 11936 38016 11940
rect 38032 11996 38096 12000
rect 38032 11940 38036 11996
rect 38036 11940 38092 11996
rect 38092 11940 38096 11996
rect 38032 11936 38096 11940
rect 38112 11996 38176 12000
rect 38112 11940 38116 11996
rect 38116 11940 38172 11996
rect 38172 11940 38176 11996
rect 38112 11936 38176 11940
rect 38192 11996 38256 12000
rect 38192 11940 38196 11996
rect 38196 11940 38252 11996
rect 38252 11940 38256 11996
rect 38192 11936 38256 11940
rect 47952 11996 48016 12000
rect 47952 11940 47956 11996
rect 47956 11940 48012 11996
rect 48012 11940 48016 11996
rect 47952 11936 48016 11940
rect 48032 11996 48096 12000
rect 48032 11940 48036 11996
rect 48036 11940 48092 11996
rect 48092 11940 48096 11996
rect 48032 11936 48096 11940
rect 48112 11996 48176 12000
rect 48112 11940 48116 11996
rect 48116 11940 48172 11996
rect 48172 11940 48176 11996
rect 48112 11936 48176 11940
rect 48192 11996 48256 12000
rect 48192 11940 48196 11996
rect 48196 11940 48252 11996
rect 48252 11940 48256 11996
rect 48192 11936 48256 11940
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 32952 11452 33016 11456
rect 32952 11396 32956 11452
rect 32956 11396 33012 11452
rect 33012 11396 33016 11452
rect 32952 11392 33016 11396
rect 33032 11452 33096 11456
rect 33032 11396 33036 11452
rect 33036 11396 33092 11452
rect 33092 11396 33096 11452
rect 33032 11392 33096 11396
rect 33112 11452 33176 11456
rect 33112 11396 33116 11452
rect 33116 11396 33172 11452
rect 33172 11396 33176 11452
rect 33112 11392 33176 11396
rect 33192 11452 33256 11456
rect 33192 11396 33196 11452
rect 33196 11396 33252 11452
rect 33252 11396 33256 11452
rect 33192 11392 33256 11396
rect 42952 11452 43016 11456
rect 42952 11396 42956 11452
rect 42956 11396 43012 11452
rect 43012 11396 43016 11452
rect 42952 11392 43016 11396
rect 43032 11452 43096 11456
rect 43032 11396 43036 11452
rect 43036 11396 43092 11452
rect 43092 11396 43096 11452
rect 43032 11392 43096 11396
rect 43112 11452 43176 11456
rect 43112 11396 43116 11452
rect 43116 11396 43172 11452
rect 43172 11396 43176 11452
rect 43112 11392 43176 11396
rect 43192 11452 43256 11456
rect 43192 11396 43196 11452
rect 43196 11396 43252 11452
rect 43252 11396 43256 11452
rect 43192 11392 43256 11396
rect 14044 11052 14108 11116
rect 29132 10976 29196 10980
rect 29132 10920 29146 10976
rect 29146 10920 29196 10976
rect 29132 10916 29196 10920
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 27952 10908 28016 10912
rect 27952 10852 27956 10908
rect 27956 10852 28012 10908
rect 28012 10852 28016 10908
rect 27952 10848 28016 10852
rect 28032 10908 28096 10912
rect 28032 10852 28036 10908
rect 28036 10852 28092 10908
rect 28092 10852 28096 10908
rect 28032 10848 28096 10852
rect 28112 10908 28176 10912
rect 28112 10852 28116 10908
rect 28116 10852 28172 10908
rect 28172 10852 28176 10908
rect 28112 10848 28176 10852
rect 28192 10908 28256 10912
rect 28192 10852 28196 10908
rect 28196 10852 28252 10908
rect 28252 10852 28256 10908
rect 28192 10848 28256 10852
rect 37952 10908 38016 10912
rect 37952 10852 37956 10908
rect 37956 10852 38012 10908
rect 38012 10852 38016 10908
rect 37952 10848 38016 10852
rect 38032 10908 38096 10912
rect 38032 10852 38036 10908
rect 38036 10852 38092 10908
rect 38092 10852 38096 10908
rect 38032 10848 38096 10852
rect 38112 10908 38176 10912
rect 38112 10852 38116 10908
rect 38116 10852 38172 10908
rect 38172 10852 38176 10908
rect 38112 10848 38176 10852
rect 38192 10908 38256 10912
rect 38192 10852 38196 10908
rect 38196 10852 38252 10908
rect 38252 10852 38256 10908
rect 38192 10848 38256 10852
rect 47952 10908 48016 10912
rect 47952 10852 47956 10908
rect 47956 10852 48012 10908
rect 48012 10852 48016 10908
rect 47952 10848 48016 10852
rect 48032 10908 48096 10912
rect 48032 10852 48036 10908
rect 48036 10852 48092 10908
rect 48092 10852 48096 10908
rect 48032 10848 48096 10852
rect 48112 10908 48176 10912
rect 48112 10852 48116 10908
rect 48116 10852 48172 10908
rect 48172 10852 48176 10908
rect 48112 10848 48176 10852
rect 48192 10908 48256 10912
rect 48192 10852 48196 10908
rect 48196 10852 48252 10908
rect 48252 10852 48256 10908
rect 48192 10848 48256 10852
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 32952 10364 33016 10368
rect 32952 10308 32956 10364
rect 32956 10308 33012 10364
rect 33012 10308 33016 10364
rect 32952 10304 33016 10308
rect 33032 10364 33096 10368
rect 33032 10308 33036 10364
rect 33036 10308 33092 10364
rect 33092 10308 33096 10364
rect 33032 10304 33096 10308
rect 33112 10364 33176 10368
rect 33112 10308 33116 10364
rect 33116 10308 33172 10364
rect 33172 10308 33176 10364
rect 33112 10304 33176 10308
rect 33192 10364 33256 10368
rect 33192 10308 33196 10364
rect 33196 10308 33252 10364
rect 33252 10308 33256 10364
rect 33192 10304 33256 10308
rect 42952 10364 43016 10368
rect 42952 10308 42956 10364
rect 42956 10308 43012 10364
rect 43012 10308 43016 10364
rect 42952 10304 43016 10308
rect 43032 10364 43096 10368
rect 43032 10308 43036 10364
rect 43036 10308 43092 10364
rect 43092 10308 43096 10364
rect 43032 10304 43096 10308
rect 43112 10364 43176 10368
rect 43112 10308 43116 10364
rect 43116 10308 43172 10364
rect 43172 10308 43176 10364
rect 43112 10304 43176 10308
rect 43192 10364 43256 10368
rect 43192 10308 43196 10364
rect 43196 10308 43252 10364
rect 43252 10308 43256 10364
rect 43192 10304 43256 10308
rect 16988 10100 17052 10164
rect 38516 10160 38580 10164
rect 38516 10104 38566 10160
rect 38566 10104 38580 10160
rect 38516 10100 38580 10104
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 27952 9820 28016 9824
rect 27952 9764 27956 9820
rect 27956 9764 28012 9820
rect 28012 9764 28016 9820
rect 27952 9760 28016 9764
rect 28032 9820 28096 9824
rect 28032 9764 28036 9820
rect 28036 9764 28092 9820
rect 28092 9764 28096 9820
rect 28032 9760 28096 9764
rect 28112 9820 28176 9824
rect 28112 9764 28116 9820
rect 28116 9764 28172 9820
rect 28172 9764 28176 9820
rect 28112 9760 28176 9764
rect 28192 9820 28256 9824
rect 28192 9764 28196 9820
rect 28196 9764 28252 9820
rect 28252 9764 28256 9820
rect 28192 9760 28256 9764
rect 37952 9820 38016 9824
rect 37952 9764 37956 9820
rect 37956 9764 38012 9820
rect 38012 9764 38016 9820
rect 37952 9760 38016 9764
rect 38032 9820 38096 9824
rect 38032 9764 38036 9820
rect 38036 9764 38092 9820
rect 38092 9764 38096 9820
rect 38032 9760 38096 9764
rect 38112 9820 38176 9824
rect 38112 9764 38116 9820
rect 38116 9764 38172 9820
rect 38172 9764 38176 9820
rect 38112 9760 38176 9764
rect 38192 9820 38256 9824
rect 38192 9764 38196 9820
rect 38196 9764 38252 9820
rect 38252 9764 38256 9820
rect 38192 9760 38256 9764
rect 47952 9820 48016 9824
rect 47952 9764 47956 9820
rect 47956 9764 48012 9820
rect 48012 9764 48016 9820
rect 47952 9760 48016 9764
rect 48032 9820 48096 9824
rect 48032 9764 48036 9820
rect 48036 9764 48092 9820
rect 48092 9764 48096 9820
rect 48032 9760 48096 9764
rect 48112 9820 48176 9824
rect 48112 9764 48116 9820
rect 48116 9764 48172 9820
rect 48172 9764 48176 9820
rect 48112 9760 48176 9764
rect 48192 9820 48256 9824
rect 48192 9764 48196 9820
rect 48196 9764 48252 9820
rect 48252 9764 48256 9820
rect 48192 9760 48256 9764
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 32952 9276 33016 9280
rect 32952 9220 32956 9276
rect 32956 9220 33012 9276
rect 33012 9220 33016 9276
rect 32952 9216 33016 9220
rect 33032 9276 33096 9280
rect 33032 9220 33036 9276
rect 33036 9220 33092 9276
rect 33092 9220 33096 9276
rect 33032 9216 33096 9220
rect 33112 9276 33176 9280
rect 33112 9220 33116 9276
rect 33116 9220 33172 9276
rect 33172 9220 33176 9276
rect 33112 9216 33176 9220
rect 33192 9276 33256 9280
rect 33192 9220 33196 9276
rect 33196 9220 33252 9276
rect 33252 9220 33256 9276
rect 33192 9216 33256 9220
rect 42952 9276 43016 9280
rect 42952 9220 42956 9276
rect 42956 9220 43012 9276
rect 43012 9220 43016 9276
rect 42952 9216 43016 9220
rect 43032 9276 43096 9280
rect 43032 9220 43036 9276
rect 43036 9220 43092 9276
rect 43092 9220 43096 9276
rect 43032 9216 43096 9220
rect 43112 9276 43176 9280
rect 43112 9220 43116 9276
rect 43116 9220 43172 9276
rect 43172 9220 43176 9276
rect 43112 9216 43176 9220
rect 43192 9276 43256 9280
rect 43192 9220 43196 9276
rect 43196 9220 43252 9276
rect 43252 9220 43256 9276
rect 43192 9216 43256 9220
rect 14228 9072 14292 9076
rect 14228 9016 14242 9072
rect 14242 9016 14292 9072
rect 14228 9012 14292 9016
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 27952 8732 28016 8736
rect 27952 8676 27956 8732
rect 27956 8676 28012 8732
rect 28012 8676 28016 8732
rect 27952 8672 28016 8676
rect 28032 8732 28096 8736
rect 28032 8676 28036 8732
rect 28036 8676 28092 8732
rect 28092 8676 28096 8732
rect 28032 8672 28096 8676
rect 28112 8732 28176 8736
rect 28112 8676 28116 8732
rect 28116 8676 28172 8732
rect 28172 8676 28176 8732
rect 28112 8672 28176 8676
rect 28192 8732 28256 8736
rect 28192 8676 28196 8732
rect 28196 8676 28252 8732
rect 28252 8676 28256 8732
rect 28192 8672 28256 8676
rect 37952 8732 38016 8736
rect 37952 8676 37956 8732
rect 37956 8676 38012 8732
rect 38012 8676 38016 8732
rect 37952 8672 38016 8676
rect 38032 8732 38096 8736
rect 38032 8676 38036 8732
rect 38036 8676 38092 8732
rect 38092 8676 38096 8732
rect 38032 8672 38096 8676
rect 38112 8732 38176 8736
rect 38112 8676 38116 8732
rect 38116 8676 38172 8732
rect 38172 8676 38176 8732
rect 38112 8672 38176 8676
rect 38192 8732 38256 8736
rect 38192 8676 38196 8732
rect 38196 8676 38252 8732
rect 38252 8676 38256 8732
rect 38192 8672 38256 8676
rect 47952 8732 48016 8736
rect 47952 8676 47956 8732
rect 47956 8676 48012 8732
rect 48012 8676 48016 8732
rect 47952 8672 48016 8676
rect 48032 8732 48096 8736
rect 48032 8676 48036 8732
rect 48036 8676 48092 8732
rect 48092 8676 48096 8732
rect 48032 8672 48096 8676
rect 48112 8732 48176 8736
rect 48112 8676 48116 8732
rect 48116 8676 48172 8732
rect 48172 8676 48176 8732
rect 48112 8672 48176 8676
rect 48192 8732 48256 8736
rect 48192 8676 48196 8732
rect 48196 8676 48252 8732
rect 48252 8676 48256 8732
rect 48192 8672 48256 8676
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 32952 8188 33016 8192
rect 32952 8132 32956 8188
rect 32956 8132 33012 8188
rect 33012 8132 33016 8188
rect 32952 8128 33016 8132
rect 33032 8188 33096 8192
rect 33032 8132 33036 8188
rect 33036 8132 33092 8188
rect 33092 8132 33096 8188
rect 33032 8128 33096 8132
rect 33112 8188 33176 8192
rect 33112 8132 33116 8188
rect 33116 8132 33172 8188
rect 33172 8132 33176 8188
rect 33112 8128 33176 8132
rect 33192 8188 33256 8192
rect 33192 8132 33196 8188
rect 33196 8132 33252 8188
rect 33252 8132 33256 8188
rect 33192 8128 33256 8132
rect 42952 8188 43016 8192
rect 42952 8132 42956 8188
rect 42956 8132 43012 8188
rect 43012 8132 43016 8188
rect 42952 8128 43016 8132
rect 43032 8188 43096 8192
rect 43032 8132 43036 8188
rect 43036 8132 43092 8188
rect 43092 8132 43096 8188
rect 43032 8128 43096 8132
rect 43112 8188 43176 8192
rect 43112 8132 43116 8188
rect 43116 8132 43172 8188
rect 43172 8132 43176 8188
rect 43112 8128 43176 8132
rect 43192 8188 43256 8192
rect 43192 8132 43196 8188
rect 43196 8132 43252 8188
rect 43252 8132 43256 8188
rect 43192 8128 43256 8132
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 27952 7644 28016 7648
rect 27952 7588 27956 7644
rect 27956 7588 28012 7644
rect 28012 7588 28016 7644
rect 27952 7584 28016 7588
rect 28032 7644 28096 7648
rect 28032 7588 28036 7644
rect 28036 7588 28092 7644
rect 28092 7588 28096 7644
rect 28032 7584 28096 7588
rect 28112 7644 28176 7648
rect 28112 7588 28116 7644
rect 28116 7588 28172 7644
rect 28172 7588 28176 7644
rect 28112 7584 28176 7588
rect 28192 7644 28256 7648
rect 28192 7588 28196 7644
rect 28196 7588 28252 7644
rect 28252 7588 28256 7644
rect 28192 7584 28256 7588
rect 37952 7644 38016 7648
rect 37952 7588 37956 7644
rect 37956 7588 38012 7644
rect 38012 7588 38016 7644
rect 37952 7584 38016 7588
rect 38032 7644 38096 7648
rect 38032 7588 38036 7644
rect 38036 7588 38092 7644
rect 38092 7588 38096 7644
rect 38032 7584 38096 7588
rect 38112 7644 38176 7648
rect 38112 7588 38116 7644
rect 38116 7588 38172 7644
rect 38172 7588 38176 7644
rect 38112 7584 38176 7588
rect 38192 7644 38256 7648
rect 38192 7588 38196 7644
rect 38196 7588 38252 7644
rect 38252 7588 38256 7644
rect 38192 7584 38256 7588
rect 47952 7644 48016 7648
rect 47952 7588 47956 7644
rect 47956 7588 48012 7644
rect 48012 7588 48016 7644
rect 47952 7584 48016 7588
rect 48032 7644 48096 7648
rect 48032 7588 48036 7644
rect 48036 7588 48092 7644
rect 48092 7588 48096 7644
rect 48032 7584 48096 7588
rect 48112 7644 48176 7648
rect 48112 7588 48116 7644
rect 48116 7588 48172 7644
rect 48172 7588 48176 7644
rect 48112 7584 48176 7588
rect 48192 7644 48256 7648
rect 48192 7588 48196 7644
rect 48196 7588 48252 7644
rect 48252 7588 48256 7644
rect 48192 7584 48256 7588
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 32952 7100 33016 7104
rect 32952 7044 32956 7100
rect 32956 7044 33012 7100
rect 33012 7044 33016 7100
rect 32952 7040 33016 7044
rect 33032 7100 33096 7104
rect 33032 7044 33036 7100
rect 33036 7044 33092 7100
rect 33092 7044 33096 7100
rect 33032 7040 33096 7044
rect 33112 7100 33176 7104
rect 33112 7044 33116 7100
rect 33116 7044 33172 7100
rect 33172 7044 33176 7100
rect 33112 7040 33176 7044
rect 33192 7100 33256 7104
rect 33192 7044 33196 7100
rect 33196 7044 33252 7100
rect 33252 7044 33256 7100
rect 33192 7040 33256 7044
rect 42952 7100 43016 7104
rect 42952 7044 42956 7100
rect 42956 7044 43012 7100
rect 43012 7044 43016 7100
rect 42952 7040 43016 7044
rect 43032 7100 43096 7104
rect 43032 7044 43036 7100
rect 43036 7044 43092 7100
rect 43092 7044 43096 7100
rect 43032 7040 43096 7044
rect 43112 7100 43176 7104
rect 43112 7044 43116 7100
rect 43116 7044 43172 7100
rect 43172 7044 43176 7100
rect 43112 7040 43176 7044
rect 43192 7100 43256 7104
rect 43192 7044 43196 7100
rect 43196 7044 43252 7100
rect 43252 7044 43256 7100
rect 43192 7040 43256 7044
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 27952 6556 28016 6560
rect 27952 6500 27956 6556
rect 27956 6500 28012 6556
rect 28012 6500 28016 6556
rect 27952 6496 28016 6500
rect 28032 6556 28096 6560
rect 28032 6500 28036 6556
rect 28036 6500 28092 6556
rect 28092 6500 28096 6556
rect 28032 6496 28096 6500
rect 28112 6556 28176 6560
rect 28112 6500 28116 6556
rect 28116 6500 28172 6556
rect 28172 6500 28176 6556
rect 28112 6496 28176 6500
rect 28192 6556 28256 6560
rect 28192 6500 28196 6556
rect 28196 6500 28252 6556
rect 28252 6500 28256 6556
rect 28192 6496 28256 6500
rect 37952 6556 38016 6560
rect 37952 6500 37956 6556
rect 37956 6500 38012 6556
rect 38012 6500 38016 6556
rect 37952 6496 38016 6500
rect 38032 6556 38096 6560
rect 38032 6500 38036 6556
rect 38036 6500 38092 6556
rect 38092 6500 38096 6556
rect 38032 6496 38096 6500
rect 38112 6556 38176 6560
rect 38112 6500 38116 6556
rect 38116 6500 38172 6556
rect 38172 6500 38176 6556
rect 38112 6496 38176 6500
rect 38192 6556 38256 6560
rect 38192 6500 38196 6556
rect 38196 6500 38252 6556
rect 38252 6500 38256 6556
rect 38192 6496 38256 6500
rect 47952 6556 48016 6560
rect 47952 6500 47956 6556
rect 47956 6500 48012 6556
rect 48012 6500 48016 6556
rect 47952 6496 48016 6500
rect 48032 6556 48096 6560
rect 48032 6500 48036 6556
rect 48036 6500 48092 6556
rect 48092 6500 48096 6556
rect 48032 6496 48096 6500
rect 48112 6556 48176 6560
rect 48112 6500 48116 6556
rect 48116 6500 48172 6556
rect 48172 6500 48176 6556
rect 48112 6496 48176 6500
rect 48192 6556 48256 6560
rect 48192 6500 48196 6556
rect 48196 6500 48252 6556
rect 48252 6500 48256 6556
rect 48192 6496 48256 6500
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 32952 6012 33016 6016
rect 32952 5956 32956 6012
rect 32956 5956 33012 6012
rect 33012 5956 33016 6012
rect 32952 5952 33016 5956
rect 33032 6012 33096 6016
rect 33032 5956 33036 6012
rect 33036 5956 33092 6012
rect 33092 5956 33096 6012
rect 33032 5952 33096 5956
rect 33112 6012 33176 6016
rect 33112 5956 33116 6012
rect 33116 5956 33172 6012
rect 33172 5956 33176 6012
rect 33112 5952 33176 5956
rect 33192 6012 33256 6016
rect 33192 5956 33196 6012
rect 33196 5956 33252 6012
rect 33252 5956 33256 6012
rect 33192 5952 33256 5956
rect 42952 6012 43016 6016
rect 42952 5956 42956 6012
rect 42956 5956 43012 6012
rect 43012 5956 43016 6012
rect 42952 5952 43016 5956
rect 43032 6012 43096 6016
rect 43032 5956 43036 6012
rect 43036 5956 43092 6012
rect 43092 5956 43096 6012
rect 43032 5952 43096 5956
rect 43112 6012 43176 6016
rect 43112 5956 43116 6012
rect 43116 5956 43172 6012
rect 43172 5956 43176 6012
rect 43112 5952 43176 5956
rect 43192 6012 43256 6016
rect 43192 5956 43196 6012
rect 43196 5956 43252 6012
rect 43252 5956 43256 6012
rect 43192 5952 43256 5956
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 27952 5468 28016 5472
rect 27952 5412 27956 5468
rect 27956 5412 28012 5468
rect 28012 5412 28016 5468
rect 27952 5408 28016 5412
rect 28032 5468 28096 5472
rect 28032 5412 28036 5468
rect 28036 5412 28092 5468
rect 28092 5412 28096 5468
rect 28032 5408 28096 5412
rect 28112 5468 28176 5472
rect 28112 5412 28116 5468
rect 28116 5412 28172 5468
rect 28172 5412 28176 5468
rect 28112 5408 28176 5412
rect 28192 5468 28256 5472
rect 28192 5412 28196 5468
rect 28196 5412 28252 5468
rect 28252 5412 28256 5468
rect 28192 5408 28256 5412
rect 37952 5468 38016 5472
rect 37952 5412 37956 5468
rect 37956 5412 38012 5468
rect 38012 5412 38016 5468
rect 37952 5408 38016 5412
rect 38032 5468 38096 5472
rect 38032 5412 38036 5468
rect 38036 5412 38092 5468
rect 38092 5412 38096 5468
rect 38032 5408 38096 5412
rect 38112 5468 38176 5472
rect 38112 5412 38116 5468
rect 38116 5412 38172 5468
rect 38172 5412 38176 5468
rect 38112 5408 38176 5412
rect 38192 5468 38256 5472
rect 38192 5412 38196 5468
rect 38196 5412 38252 5468
rect 38252 5412 38256 5468
rect 38192 5408 38256 5412
rect 47952 5468 48016 5472
rect 47952 5412 47956 5468
rect 47956 5412 48012 5468
rect 48012 5412 48016 5468
rect 47952 5408 48016 5412
rect 48032 5468 48096 5472
rect 48032 5412 48036 5468
rect 48036 5412 48092 5468
rect 48092 5412 48096 5468
rect 48032 5408 48096 5412
rect 48112 5468 48176 5472
rect 48112 5412 48116 5468
rect 48116 5412 48172 5468
rect 48172 5412 48176 5468
rect 48112 5408 48176 5412
rect 48192 5468 48256 5472
rect 48192 5412 48196 5468
rect 48196 5412 48252 5468
rect 48252 5412 48256 5468
rect 48192 5408 48256 5412
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 32952 4924 33016 4928
rect 32952 4868 32956 4924
rect 32956 4868 33012 4924
rect 33012 4868 33016 4924
rect 32952 4864 33016 4868
rect 33032 4924 33096 4928
rect 33032 4868 33036 4924
rect 33036 4868 33092 4924
rect 33092 4868 33096 4924
rect 33032 4864 33096 4868
rect 33112 4924 33176 4928
rect 33112 4868 33116 4924
rect 33116 4868 33172 4924
rect 33172 4868 33176 4924
rect 33112 4864 33176 4868
rect 33192 4924 33256 4928
rect 33192 4868 33196 4924
rect 33196 4868 33252 4924
rect 33252 4868 33256 4924
rect 33192 4864 33256 4868
rect 42952 4924 43016 4928
rect 42952 4868 42956 4924
rect 42956 4868 43012 4924
rect 43012 4868 43016 4924
rect 42952 4864 43016 4868
rect 43032 4924 43096 4928
rect 43032 4868 43036 4924
rect 43036 4868 43092 4924
rect 43092 4868 43096 4924
rect 43032 4864 43096 4868
rect 43112 4924 43176 4928
rect 43112 4868 43116 4924
rect 43116 4868 43172 4924
rect 43172 4868 43176 4924
rect 43112 4864 43176 4868
rect 43192 4924 43256 4928
rect 43192 4868 43196 4924
rect 43196 4868 43252 4924
rect 43252 4868 43256 4924
rect 43192 4864 43256 4868
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 27952 4380 28016 4384
rect 27952 4324 27956 4380
rect 27956 4324 28012 4380
rect 28012 4324 28016 4380
rect 27952 4320 28016 4324
rect 28032 4380 28096 4384
rect 28032 4324 28036 4380
rect 28036 4324 28092 4380
rect 28092 4324 28096 4380
rect 28032 4320 28096 4324
rect 28112 4380 28176 4384
rect 28112 4324 28116 4380
rect 28116 4324 28172 4380
rect 28172 4324 28176 4380
rect 28112 4320 28176 4324
rect 28192 4380 28256 4384
rect 28192 4324 28196 4380
rect 28196 4324 28252 4380
rect 28252 4324 28256 4380
rect 28192 4320 28256 4324
rect 37952 4380 38016 4384
rect 37952 4324 37956 4380
rect 37956 4324 38012 4380
rect 38012 4324 38016 4380
rect 37952 4320 38016 4324
rect 38032 4380 38096 4384
rect 38032 4324 38036 4380
rect 38036 4324 38092 4380
rect 38092 4324 38096 4380
rect 38032 4320 38096 4324
rect 38112 4380 38176 4384
rect 38112 4324 38116 4380
rect 38116 4324 38172 4380
rect 38172 4324 38176 4380
rect 38112 4320 38176 4324
rect 38192 4380 38256 4384
rect 38192 4324 38196 4380
rect 38196 4324 38252 4380
rect 38252 4324 38256 4380
rect 38192 4320 38256 4324
rect 47952 4380 48016 4384
rect 47952 4324 47956 4380
rect 47956 4324 48012 4380
rect 48012 4324 48016 4380
rect 47952 4320 48016 4324
rect 48032 4380 48096 4384
rect 48032 4324 48036 4380
rect 48036 4324 48092 4380
rect 48092 4324 48096 4380
rect 48032 4320 48096 4324
rect 48112 4380 48176 4384
rect 48112 4324 48116 4380
rect 48116 4324 48172 4380
rect 48172 4324 48176 4380
rect 48112 4320 48176 4324
rect 48192 4380 48256 4384
rect 48192 4324 48196 4380
rect 48196 4324 48252 4380
rect 48252 4324 48256 4380
rect 48192 4320 48256 4324
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 32952 3836 33016 3840
rect 32952 3780 32956 3836
rect 32956 3780 33012 3836
rect 33012 3780 33016 3836
rect 32952 3776 33016 3780
rect 33032 3836 33096 3840
rect 33032 3780 33036 3836
rect 33036 3780 33092 3836
rect 33092 3780 33096 3836
rect 33032 3776 33096 3780
rect 33112 3836 33176 3840
rect 33112 3780 33116 3836
rect 33116 3780 33172 3836
rect 33172 3780 33176 3836
rect 33112 3776 33176 3780
rect 33192 3836 33256 3840
rect 33192 3780 33196 3836
rect 33196 3780 33252 3836
rect 33252 3780 33256 3836
rect 33192 3776 33256 3780
rect 42952 3836 43016 3840
rect 42952 3780 42956 3836
rect 42956 3780 43012 3836
rect 43012 3780 43016 3836
rect 42952 3776 43016 3780
rect 43032 3836 43096 3840
rect 43032 3780 43036 3836
rect 43036 3780 43092 3836
rect 43092 3780 43096 3836
rect 43032 3776 43096 3780
rect 43112 3836 43176 3840
rect 43112 3780 43116 3836
rect 43116 3780 43172 3836
rect 43172 3780 43176 3836
rect 43112 3776 43176 3780
rect 43192 3836 43256 3840
rect 43192 3780 43196 3836
rect 43196 3780 43252 3836
rect 43252 3780 43256 3836
rect 43192 3776 43256 3780
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 27952 3292 28016 3296
rect 27952 3236 27956 3292
rect 27956 3236 28012 3292
rect 28012 3236 28016 3292
rect 27952 3232 28016 3236
rect 28032 3292 28096 3296
rect 28032 3236 28036 3292
rect 28036 3236 28092 3292
rect 28092 3236 28096 3292
rect 28032 3232 28096 3236
rect 28112 3292 28176 3296
rect 28112 3236 28116 3292
rect 28116 3236 28172 3292
rect 28172 3236 28176 3292
rect 28112 3232 28176 3236
rect 28192 3292 28256 3296
rect 28192 3236 28196 3292
rect 28196 3236 28252 3292
rect 28252 3236 28256 3292
rect 28192 3232 28256 3236
rect 37952 3292 38016 3296
rect 37952 3236 37956 3292
rect 37956 3236 38012 3292
rect 38012 3236 38016 3292
rect 37952 3232 38016 3236
rect 38032 3292 38096 3296
rect 38032 3236 38036 3292
rect 38036 3236 38092 3292
rect 38092 3236 38096 3292
rect 38032 3232 38096 3236
rect 38112 3292 38176 3296
rect 38112 3236 38116 3292
rect 38116 3236 38172 3292
rect 38172 3236 38176 3292
rect 38112 3232 38176 3236
rect 38192 3292 38256 3296
rect 38192 3236 38196 3292
rect 38196 3236 38252 3292
rect 38252 3236 38256 3292
rect 38192 3232 38256 3236
rect 47952 3292 48016 3296
rect 47952 3236 47956 3292
rect 47956 3236 48012 3292
rect 48012 3236 48016 3292
rect 47952 3232 48016 3236
rect 48032 3292 48096 3296
rect 48032 3236 48036 3292
rect 48036 3236 48092 3292
rect 48092 3236 48096 3292
rect 48032 3232 48096 3236
rect 48112 3292 48176 3296
rect 48112 3236 48116 3292
rect 48116 3236 48172 3292
rect 48172 3236 48176 3292
rect 48112 3232 48176 3236
rect 48192 3292 48256 3296
rect 48192 3236 48196 3292
rect 48196 3236 48252 3292
rect 48252 3236 48256 3292
rect 48192 3232 48256 3236
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 32952 2748 33016 2752
rect 32952 2692 32956 2748
rect 32956 2692 33012 2748
rect 33012 2692 33016 2748
rect 32952 2688 33016 2692
rect 33032 2748 33096 2752
rect 33032 2692 33036 2748
rect 33036 2692 33092 2748
rect 33092 2692 33096 2748
rect 33032 2688 33096 2692
rect 33112 2748 33176 2752
rect 33112 2692 33116 2748
rect 33116 2692 33172 2748
rect 33172 2692 33176 2748
rect 33112 2688 33176 2692
rect 33192 2748 33256 2752
rect 33192 2692 33196 2748
rect 33196 2692 33252 2748
rect 33252 2692 33256 2748
rect 33192 2688 33256 2692
rect 42952 2748 43016 2752
rect 42952 2692 42956 2748
rect 42956 2692 43012 2748
rect 43012 2692 43016 2748
rect 42952 2688 43016 2692
rect 43032 2748 43096 2752
rect 43032 2692 43036 2748
rect 43036 2692 43092 2748
rect 43092 2692 43096 2748
rect 43032 2688 43096 2692
rect 43112 2748 43176 2752
rect 43112 2692 43116 2748
rect 43116 2692 43172 2748
rect 43172 2692 43176 2748
rect 43112 2688 43176 2692
rect 43192 2748 43256 2752
rect 43192 2692 43196 2748
rect 43196 2692 43252 2748
rect 43252 2692 43256 2748
rect 43192 2688 43256 2692
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 27952 2204 28016 2208
rect 27952 2148 27956 2204
rect 27956 2148 28012 2204
rect 28012 2148 28016 2204
rect 27952 2144 28016 2148
rect 28032 2204 28096 2208
rect 28032 2148 28036 2204
rect 28036 2148 28092 2204
rect 28092 2148 28096 2204
rect 28032 2144 28096 2148
rect 28112 2204 28176 2208
rect 28112 2148 28116 2204
rect 28116 2148 28172 2204
rect 28172 2148 28176 2204
rect 28112 2144 28176 2148
rect 28192 2204 28256 2208
rect 28192 2148 28196 2204
rect 28196 2148 28252 2204
rect 28252 2148 28256 2204
rect 28192 2144 28256 2148
rect 37952 2204 38016 2208
rect 37952 2148 37956 2204
rect 37956 2148 38012 2204
rect 38012 2148 38016 2204
rect 37952 2144 38016 2148
rect 38032 2204 38096 2208
rect 38032 2148 38036 2204
rect 38036 2148 38092 2204
rect 38092 2148 38096 2204
rect 38032 2144 38096 2148
rect 38112 2204 38176 2208
rect 38112 2148 38116 2204
rect 38116 2148 38172 2204
rect 38172 2148 38176 2204
rect 38112 2144 38176 2148
rect 38192 2204 38256 2208
rect 38192 2148 38196 2204
rect 38196 2148 38252 2204
rect 38252 2148 38256 2204
rect 38192 2144 38256 2148
rect 47952 2204 48016 2208
rect 47952 2148 47956 2204
rect 47956 2148 48012 2204
rect 48012 2148 48016 2204
rect 47952 2144 48016 2148
rect 48032 2204 48096 2208
rect 48032 2148 48036 2204
rect 48036 2148 48092 2204
rect 48092 2148 48096 2204
rect 48032 2144 48096 2148
rect 48112 2204 48176 2208
rect 48112 2148 48116 2204
rect 48116 2148 48172 2204
rect 48172 2148 48176 2204
rect 48112 2144 48176 2148
rect 48192 2204 48256 2208
rect 48192 2148 48196 2204
rect 48196 2148 48252 2204
rect 48252 2148 48256 2204
rect 48192 2144 48256 2148
<< metal4 >>
rect 2944 24512 3264 24528
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2944 23424 3264 24448
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 23968 8264 24528
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 7944 22880 8264 23904
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7944 20704 8264 21728
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7944 17440 8264 18464
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7944 14176 8264 15200
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 10912 8264 11936
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7944 8736 8264 9760
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 7648 8264 8672
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 24512 13264 24528
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 12944 23424 13264 24448
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12944 22336 13264 23360
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12944 21248 13264 22272
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12944 20160 13264 21184
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12944 19072 13264 20096
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12944 16896 13264 17920
rect 17944 23968 18264 24528
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 17944 22880 18264 23904
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17944 21792 18264 22816
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 17944 20704 18264 21728
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17944 19616 18264 20640
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17944 18528 18264 19552
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17944 17440 18264 18464
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 14411 17100 14477 17101
rect 14411 17036 14412 17100
rect 14476 17036 14477 17100
rect 14411 17035 14477 17036
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12944 15808 13264 16832
rect 14043 16148 14109 16149
rect 14043 16084 14044 16148
rect 14108 16084 14109 16148
rect 14043 16083 14109 16084
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12944 13632 13264 14656
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 14046 11117 14106 16083
rect 14227 14380 14293 14381
rect 14227 14316 14228 14380
rect 14292 14316 14293 14380
rect 14227 14315 14293 14316
rect 14043 11116 14109 11117
rect 14043 11052 14044 11116
rect 14108 11052 14109 11116
rect 14043 11051 14109 11052
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 9280 13264 10304
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12944 8192 13264 9216
rect 14230 9077 14290 14315
rect 14414 12749 14474 17035
rect 16067 16692 16133 16693
rect 16067 16628 16068 16692
rect 16132 16628 16133 16692
rect 16067 16627 16133 16628
rect 16070 13701 16130 16627
rect 17944 16352 18264 17376
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 16987 15876 17053 15877
rect 16987 15812 16988 15876
rect 17052 15812 17053 15876
rect 16987 15811 17053 15812
rect 16067 13700 16133 13701
rect 16067 13636 16068 13700
rect 16132 13636 16133 13700
rect 16067 13635 16133 13636
rect 14411 12748 14477 12749
rect 14411 12684 14412 12748
rect 14476 12684 14477 12748
rect 14411 12683 14477 12684
rect 16990 10165 17050 15811
rect 17944 15264 18264 16288
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 17944 13088 18264 14112
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17944 12000 18264 13024
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 17944 10912 18264 11936
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 16987 10164 17053 10165
rect 16987 10100 16988 10164
rect 17052 10100 17053 10164
rect 16987 10099 17053 10100
rect 17944 9824 18264 10848
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 14227 9076 14293 9077
rect 14227 9012 14228 9076
rect 14292 9012 14293 9076
rect 14227 9011 14293 9012
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12944 4928 13264 5952
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 17944 8736 18264 9760
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 17944 7648 18264 8672
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17944 6560 18264 7584
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 17944 5472 18264 6496
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 17944 3296 18264 4320
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 17944 2208 18264 3232
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 22944 24512 23264 24528
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 22944 23424 23264 24448
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 22944 22336 23264 23360
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 22944 21248 23264 22272
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22944 19072 23264 20096
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 22944 17984 23264 19008
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 22944 12544 23264 13568
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 22944 9280 23264 10304
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 22944 6016 23264 7040
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 22944 4928 23264 5952
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 22944 3840 23264 4864
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 22944 2752 23264 3776
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22944 2128 23264 2688
rect 27944 23968 28264 24528
rect 32944 24512 33264 24528
rect 32944 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33264 24512
rect 28947 24036 29013 24037
rect 28947 23972 28948 24036
rect 29012 23972 29013 24036
rect 28947 23971 29013 23972
rect 27944 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28264 23968
rect 27944 22880 28264 23904
rect 27944 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28264 22880
rect 27944 21792 28264 22816
rect 27944 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28264 21792
rect 27944 20704 28264 21728
rect 28763 21044 28829 21045
rect 28763 20980 28764 21044
rect 28828 20980 28829 21044
rect 28763 20979 28829 20980
rect 27944 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28264 20704
rect 27944 19616 28264 20640
rect 28579 20636 28645 20637
rect 28579 20572 28580 20636
rect 28644 20572 28645 20636
rect 28579 20571 28645 20572
rect 28395 20228 28461 20229
rect 28395 20164 28396 20228
rect 28460 20164 28461 20228
rect 28395 20163 28461 20164
rect 27944 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28264 19616
rect 27944 18528 28264 19552
rect 28398 19277 28458 20163
rect 28582 19685 28642 20571
rect 28579 19684 28645 19685
rect 28579 19620 28580 19684
rect 28644 19620 28645 19684
rect 28579 19619 28645 19620
rect 28766 19549 28826 20979
rect 28763 19548 28829 19549
rect 28763 19484 28764 19548
rect 28828 19484 28829 19548
rect 28763 19483 28829 19484
rect 28395 19276 28461 19277
rect 28395 19212 28396 19276
rect 28460 19212 28461 19276
rect 28395 19211 28461 19212
rect 27944 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28264 18528
rect 27944 17440 28264 18464
rect 27944 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28264 17440
rect 27944 16352 28264 17376
rect 28950 16829 29010 23971
rect 32944 23424 33264 24448
rect 32944 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33264 23424
rect 32944 22336 33264 23360
rect 32944 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33264 22336
rect 32944 21248 33264 22272
rect 32944 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33264 21248
rect 32944 20160 33264 21184
rect 32944 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33264 20160
rect 32944 19072 33264 20096
rect 32944 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33264 19072
rect 32944 17984 33264 19008
rect 32944 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33264 17984
rect 32944 16896 33264 17920
rect 32944 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33264 16896
rect 28947 16828 29013 16829
rect 28947 16764 28948 16828
rect 29012 16764 29013 16828
rect 28947 16763 29013 16764
rect 29131 16692 29197 16693
rect 29131 16628 29132 16692
rect 29196 16628 29197 16692
rect 29131 16627 29197 16628
rect 27944 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28264 16352
rect 27944 15264 28264 16288
rect 27944 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28264 15264
rect 27944 14176 28264 15200
rect 27944 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28264 14176
rect 27944 13088 28264 14112
rect 27944 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28264 13088
rect 27944 12000 28264 13024
rect 27944 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28264 12000
rect 27944 10912 28264 11936
rect 29134 10981 29194 16627
rect 32944 15808 33264 16832
rect 32944 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33264 15808
rect 32944 14720 33264 15744
rect 32944 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33264 14720
rect 32944 13632 33264 14656
rect 32944 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33264 13632
rect 32944 12544 33264 13568
rect 32944 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33264 12544
rect 32944 11456 33264 12480
rect 32944 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33264 11456
rect 29131 10980 29197 10981
rect 29131 10916 29132 10980
rect 29196 10916 29197 10980
rect 29131 10915 29197 10916
rect 27944 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28264 10912
rect 27944 9824 28264 10848
rect 27944 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28264 9824
rect 27944 8736 28264 9760
rect 27944 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28264 8736
rect 27944 7648 28264 8672
rect 27944 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28264 7648
rect 27944 6560 28264 7584
rect 27944 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28264 6560
rect 27944 5472 28264 6496
rect 27944 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28264 5472
rect 27944 4384 28264 5408
rect 27944 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28264 4384
rect 27944 3296 28264 4320
rect 27944 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28264 3296
rect 27944 2208 28264 3232
rect 27944 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28264 2208
rect 27944 2128 28264 2144
rect 32944 10368 33264 11392
rect 32944 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33264 10368
rect 32944 9280 33264 10304
rect 32944 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33264 9280
rect 32944 8192 33264 9216
rect 32944 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33264 8192
rect 32944 7104 33264 8128
rect 32944 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33264 7104
rect 32944 6016 33264 7040
rect 32944 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33264 6016
rect 32944 4928 33264 5952
rect 32944 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33264 4928
rect 32944 3840 33264 4864
rect 32944 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33264 3840
rect 32944 2752 33264 3776
rect 32944 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33264 2752
rect 32944 2128 33264 2688
rect 37944 23968 38264 24528
rect 37944 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38264 23968
rect 37944 22880 38264 23904
rect 37944 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38264 22880
rect 37944 21792 38264 22816
rect 37944 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38264 21792
rect 37944 20704 38264 21728
rect 37944 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38264 20704
rect 37944 19616 38264 20640
rect 37944 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38264 19616
rect 37944 18528 38264 19552
rect 37944 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38264 18528
rect 37944 17440 38264 18464
rect 37944 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38264 17440
rect 37944 16352 38264 17376
rect 42944 24512 43264 24528
rect 42944 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43264 24512
rect 42944 23424 43264 24448
rect 42944 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43264 23424
rect 42944 22336 43264 23360
rect 42944 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43264 22336
rect 42944 21248 43264 22272
rect 42944 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43264 21248
rect 42944 20160 43264 21184
rect 42944 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43264 20160
rect 42944 19072 43264 20096
rect 42944 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43264 19072
rect 42944 17984 43264 19008
rect 42944 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43264 17984
rect 38515 17100 38581 17101
rect 38515 17036 38516 17100
rect 38580 17036 38581 17100
rect 38515 17035 38581 17036
rect 37944 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38264 16352
rect 37944 15264 38264 16288
rect 37944 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38264 15264
rect 37944 14176 38264 15200
rect 37944 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38264 14176
rect 37944 13088 38264 14112
rect 37944 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38264 13088
rect 37944 12000 38264 13024
rect 37944 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38264 12000
rect 37944 10912 38264 11936
rect 37944 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38264 10912
rect 37944 9824 38264 10848
rect 38518 10165 38578 17035
rect 42944 16896 43264 17920
rect 42944 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43264 16896
rect 42944 15808 43264 16832
rect 42944 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43264 15808
rect 42944 14720 43264 15744
rect 42944 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43264 14720
rect 42944 13632 43264 14656
rect 42944 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43264 13632
rect 42944 12544 43264 13568
rect 42944 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43264 12544
rect 42944 11456 43264 12480
rect 42944 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43264 11456
rect 42944 10368 43264 11392
rect 42944 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43264 10368
rect 38515 10164 38581 10165
rect 38515 10100 38516 10164
rect 38580 10100 38581 10164
rect 38515 10099 38581 10100
rect 37944 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38264 9824
rect 37944 8736 38264 9760
rect 37944 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38264 8736
rect 37944 7648 38264 8672
rect 37944 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38264 7648
rect 37944 6560 38264 7584
rect 37944 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38264 6560
rect 37944 5472 38264 6496
rect 37944 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38264 5472
rect 37944 4384 38264 5408
rect 37944 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38264 4384
rect 37944 3296 38264 4320
rect 37944 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38264 3296
rect 37944 2208 38264 3232
rect 37944 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38264 2208
rect 37944 2128 38264 2144
rect 42944 9280 43264 10304
rect 42944 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43264 9280
rect 42944 8192 43264 9216
rect 42944 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43264 8192
rect 42944 7104 43264 8128
rect 42944 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43264 7104
rect 42944 6016 43264 7040
rect 42944 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43264 6016
rect 42944 4928 43264 5952
rect 42944 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43264 4928
rect 42944 3840 43264 4864
rect 42944 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43264 3840
rect 42944 2752 43264 3776
rect 42944 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43264 2752
rect 42944 2128 43264 2688
rect 47944 23968 48264 24528
rect 47944 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48264 23968
rect 47944 22880 48264 23904
rect 47944 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48264 22880
rect 47944 21792 48264 22816
rect 47944 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48264 21792
rect 47944 20704 48264 21728
rect 47944 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48264 20704
rect 47944 19616 48264 20640
rect 47944 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48264 19616
rect 47944 18528 48264 19552
rect 47944 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48264 18528
rect 47944 17440 48264 18464
rect 47944 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48264 17440
rect 47944 16352 48264 17376
rect 47944 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48264 16352
rect 47944 15264 48264 16288
rect 47944 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48264 15264
rect 47944 14176 48264 15200
rect 47944 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48264 14176
rect 47944 13088 48264 14112
rect 47944 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48264 13088
rect 47944 12000 48264 13024
rect 47944 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48264 12000
rect 47944 10912 48264 11936
rect 47944 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48264 10912
rect 47944 9824 48264 10848
rect 47944 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48264 9824
rect 47944 8736 48264 9760
rect 47944 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48264 8736
rect 47944 7648 48264 8672
rect 47944 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48264 7648
rect 47944 6560 48264 7584
rect 47944 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48264 6560
rect 47944 5472 48264 6496
rect 47944 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48264 5472
rect 47944 4384 48264 5408
rect 47944 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48264 4384
rect 47944 3296 48264 4320
rect 47944 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48264 3296
rect 47944 2208 48264 3232
rect 47944 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48264 2208
rect 47944 2128 48264 2144
use sky130_fd_sc_hd__clkbuf_2  _104_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14260 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _105_
timestamp 1676037725
transform 1 0 11040 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _106_
timestamp 1676037725
transform 1 0 9476 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _107_
timestamp 1676037725
transform 1 0 6348 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _108_
timestamp 1676037725
transform 1 0 10212 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _109_
timestamp 1676037725
transform 1 0 10856 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _110_
timestamp 1676037725
transform 1 0 14076 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _111_
timestamp 1676037725
transform 1 0 8096 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _112_
timestamp 1676037725
transform 1 0 10304 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _113_
timestamp 1676037725
transform 1 0 10856 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _114_
timestamp 1676037725
transform 1 0 11684 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _115_
timestamp 1676037725
transform 1 0 9108 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _116_
timestamp 1676037725
transform 1 0 14904 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _117_
timestamp 1676037725
transform 1 0 16008 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _118_
timestamp 1676037725
transform 1 0 11960 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _119_
timestamp 1676037725
transform 1 0 7636 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _120_
timestamp 1676037725
transform 1 0 11224 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1676037725
transform 1 0 12420 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _122_
timestamp 1676037725
transform 1 0 15272 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _123_
timestamp 1676037725
transform 1 0 7636 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _124_
timestamp 1676037725
transform 1 0 11684 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _125_
timestamp 1676037725
transform 1 0 12144 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _126_
timestamp 1676037725
transform 1 0 11776 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _127_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7820 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _128_
timestamp 1676037725
transform 1 0 5244 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _129_
timestamp 1676037725
transform 1 0 11684 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1676037725
transform 1 0 7728 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _131_
timestamp 1676037725
transform 1 0 3864 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _132_
timestamp 1676037725
transform 1 0 5704 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1676037725
transform 1 0 6624 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _134_
timestamp 1676037725
transform 1 0 36340 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _135_
timestamp 1676037725
transform 1 0 37904 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _136_
timestamp 1676037725
transform 1 0 37168 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _137_
timestamp 1676037725
transform 1 0 43608 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _138_
timestamp 1676037725
transform 1 0 38364 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _139_
timestamp 1676037725
transform 1 0 37628 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _140_
timestamp 1676037725
transform 1 0 37444 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _141_
timestamp 1676037725
transform 1 0 43884 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _142_
timestamp 1676037725
transform 1 0 38456 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _143_
timestamp 1676037725
transform 1 0 37720 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _144_
timestamp 1676037725
transform 1 0 37904 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _145_
timestamp 1676037725
transform 1 0 44804 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _146_
timestamp 1676037725
transform 1 0 38640 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _147_
timestamp 1676037725
transform 1 0 40204 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _148_
timestamp 1676037725
transform 1 0 39192 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _149_
timestamp 1676037725
transform 1 0 44068 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _150_
timestamp 1676037725
transform 1 0 40020 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _151_
timestamp 1676037725
transform 1 0 38180 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _152_
timestamp 1676037725
transform 1 0 39652 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _153_
timestamp 1676037725
transform 1 0 44252 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _154_
timestamp 1676037725
transform 1 0 40020 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _155_
timestamp 1676037725
transform 1 0 39836 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _156_
timestamp 1676037725
transform 1 0 40020 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _157_
timestamp 1676037725
transform 1 0 44988 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _158_
timestamp 1676037725
transform 1 0 45540 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _159_
timestamp 1676037725
transform 1 0 39928 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _160_
timestamp 1676037725
transform 1 0 45908 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _161_
timestamp 1676037725
transform 1 0 45908 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _162_
timestamp 1676037725
transform 1 0 45632 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _163_
timestamp 1676037725
transform 1 0 44896 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _164_
timestamp 1676037725
transform 1 0 9108 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _165_
timestamp 1676037725
transform 1 0 4048 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _166_
timestamp 1676037725
transform 1 0 5244 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _167_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4140 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _168_
timestamp 1676037725
transform 1 0 6624 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _169_
timestamp 1676037725
transform 1 0 4692 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _170_
timestamp 1676037725
transform 1 0 3404 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _171_
timestamp 1676037725
transform 1 0 2116 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _172_
timestamp 1676037725
transform 1 0 6532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _173_
timestamp 1676037725
transform 1 0 3956 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _174_
timestamp 1676037725
transform 1 0 25760 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _175_
timestamp 1676037725
transform 1 0 14260 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _176_
timestamp 1676037725
transform 1 0 11684 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _177_
timestamp 1676037725
transform 1 0 12696 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _178_
timestamp 1676037725
transform 1 0 12328 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _179_
timestamp 1676037725
transform 1 0 13064 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _180_
timestamp 1676037725
transform 1 0 14628 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _181_
timestamp 1676037725
transform 1 0 13892 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _182_
timestamp 1676037725
transform 1 0 14444 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _183_
timestamp 1676037725
transform 1 0 7268 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _184_
timestamp 1676037725
transform 1 0 23368 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _185_
timestamp 1676037725
transform 1 0 19596 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _186_
timestamp 1676037725
transform 1 0 19596 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _187_
timestamp 1676037725
transform 1 0 22540 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _188_
timestamp 1676037725
transform 1 0 21160 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _189_
timestamp 1676037725
transform 1 0 24564 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _190_
timestamp 1676037725
transform 1 0 19412 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _191_
timestamp 1676037725
transform 1 0 27140 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _192_
timestamp 1676037725
transform 1 0 21252 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _193_
timestamp 1676037725
transform 1 0 23184 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _194_
timestamp 1676037725
transform 1 0 16376 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _195_
timestamp 1676037725
transform 1 0 17388 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _196_
timestamp 1676037725
transform 1 0 18676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _197_
timestamp 1676037725
transform 1 0 19964 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _198_
timestamp 1676037725
transform 1 0 19412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _199_
timestamp 1676037725
transform 1 0 20608 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _200_
timestamp 1676037725
transform 1 0 21252 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _201_
timestamp 1676037725
transform 1 0 26404 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 15548 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1676037725
transform 1 0 13616 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1676037725
transform 1 0 10580 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1676037725
transform 1 0 9844 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A
timestamp 1676037725
transform 1 0 10396 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1676037725
transform 1 0 10488 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1676037725
transform 1 0 15088 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1676037725
transform 1 0 9936 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1676037725
transform 1 0 10304 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1676037725
transform 1 0 10028 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1676037725
transform 1 0 14720 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__A
timestamp 1676037725
transform 1 0 11592 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A
timestamp 1676037725
transform 1 0 12328 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1676037725
transform 1 0 12972 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__A
timestamp 1676037725
transform 1 0 14904 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A
timestamp 1676037725
transform 1 0 13156 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A
timestamp 1676037725
transform 1 0 11776 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__A
timestamp 1676037725
transform 1 0 12696 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__A
timestamp 1676037725
transform 1 0 14260 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__134__A
timestamp 1676037725
transform 1 0 36892 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__A
timestamp 1676037725
transform 1 0 38456 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__136__A
timestamp 1676037725
transform 1 0 36800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__138__A
timestamp 1676037725
transform 1 0 38916 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__A
timestamp 1676037725
transform 1 0 37260 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__140__A
timestamp 1676037725
transform 1 0 37996 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__A
timestamp 1676037725
transform 1 0 39008 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__A
timestamp 1676037725
transform 1 0 37352 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__A
timestamp 1676037725
transform 1 0 37536 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__146__A
timestamp 1676037725
transform 1 0 39192 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__147__A
timestamp 1676037725
transform 1 0 40756 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__148__A
timestamp 1676037725
transform 1 0 39836 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__150__A
timestamp 1676037725
transform 1 0 40572 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__A
timestamp 1676037725
transform 1 0 38732 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__A
timestamp 1676037725
transform 1 0 40204 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__154__A
timestamp 1676037725
transform 1 0 39560 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__A
timestamp 1676037725
transform 1 0 40388 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__A
timestamp 1676037725
transform 1 0 39376 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__159__A
timestamp 1676037725
transform 1 0 40480 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 20332 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16836 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 18216 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 18676 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16192 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14812 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 15640 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 15640 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 14812 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 12604 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13156 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 15180 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 12880 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 11224 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 14904 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 17020 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3__A0
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 20516 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 15824 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3__A1
timestamp 1676037725
transform 1 0 16376 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 9844 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 12328 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 21988 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 19320 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3__A0
timestamp 1676037725
transform 1 0 17664 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 16836 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 16192 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 12328 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3__A1
timestamp 1676037725
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 17480 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 16376 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 15180 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 10488 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 11592 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 16652 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3__A0
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 17940 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 13524 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 13340 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 12972 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__A1
timestamp 1676037725
transform 1 0 16744 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 23000 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 26220 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 31004 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1676037725
transform 1 0 28060 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_0_0_prog_clk_A
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_1_0_prog_clk_A
timestamp 1676037725
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_2_0_prog_clk_A
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_3_0_prog_clk_A
timestamp 1676037725
transform 1 0 22172 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_4_0_prog_clk_A
timestamp 1676037725
transform 1 0 18768 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_5_0_prog_clk_A
timestamp 1676037725
transform 1 0 18952 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_6_0_prog_clk_A
timestamp 1676037725
transform 1 0 22908 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_7_0_prog_clk_A
timestamp 1676037725
transform 1 0 24656 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_8_0_prog_clk_A
timestamp 1676037725
transform 1 0 28428 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_9_0_prog_clk_A
timestamp 1676037725
transform 1 0 28888 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_10_0_prog_clk_A
timestamp 1676037725
transform 1 0 34684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_11_0_prog_clk_A
timestamp 1676037725
transform 1 0 33672 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_12_0_prog_clk_A
timestamp 1676037725
transform 1 0 29256 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_13_0_prog_clk_A
timestamp 1676037725
transform 1 0 30360 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_14_0_prog_clk_A
timestamp 1676037725
transform 1 0 34408 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_15_0_prog_clk_A
timestamp 1676037725
transform 1 0 34408 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1676037725
transform 1 0 10120 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1676037725
transform 1 0 46644 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1676037725
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1676037725
transform 1 0 3036 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1676037725
transform 1 0 2300 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1676037725
transform 1 0 2760 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1676037725
transform 1 0 2116 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1676037725
transform 1 0 2116 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1676037725
transform 1 0 2300 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1676037725
transform 1 0 2116 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1676037725
transform 1 0 2852 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1676037725
transform 1 0 3036 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1676037725
transform 1 0 2300 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1676037725
transform 1 0 2300 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1676037725
transform 1 0 2116 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1676037725
transform 1 0 2852 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1676037725
transform 1 0 3036 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1676037725
transform 1 0 2300 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1676037725
transform 1 0 2760 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1676037725
transform 1 0 2668 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1676037725
transform 1 0 2116 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1676037725
transform 1 0 3312 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1676037725
transform 1 0 2116 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1676037725
transform 1 0 3956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1676037725
transform 1 0 2668 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1676037725
transform 1 0 2484 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1676037725
transform 1 0 2116 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1676037725
transform 1 0 2852 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1676037725
transform 1 0 3036 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1676037725
transform 1 0 2300 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1676037725
transform 1 0 2116 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1676037725
transform 1 0 2852 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1676037725
transform 1 0 48668 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1676037725
transform 1 0 48484 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1676037725
transform 1 0 48668 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1676037725
transform 1 0 48668 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1676037725
transform 1 0 48484 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1676037725
transform 1 0 48484 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1676037725
transform 1 0 48668 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1676037725
transform 1 0 48668 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1676037725
transform 1 0 48484 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1676037725
transform 1 0 48484 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1676037725
transform 1 0 49404 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1676037725
transform 1 0 48024 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1676037725
transform 1 0 48668 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1676037725
transform 1 0 48300 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1676037725
transform 1 0 47380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1676037725
transform 1 0 46000 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1676037725
transform 1 0 47932 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1676037725
transform 1 0 46368 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1676037725
transform 1 0 47748 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1676037725
transform 1 0 48024 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1676037725
transform 1 0 47564 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1676037725
transform 1 0 47840 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1676037725
transform 1 0 48484 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1676037725
transform 1 0 48668 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1676037725
transform 1 0 48760 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1676037725
transform 1 0 48668 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1676037725
transform 1 0 48484 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1676037725
transform 1 0 48668 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1676037725
transform 1 0 48668 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1676037725
transform 1 0 48484 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1676037725
transform 1 0 26680 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1676037725
transform 1 0 29532 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1676037725
transform 1 0 31648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1676037725
transform 1 0 31004 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1676037725
transform 1 0 34040 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1676037725
transform 1 0 44620 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1676037725
transform 1 0 34316 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1676037725
transform 1 0 41952 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1676037725
transform 1 0 42596 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1676037725
transform 1 0 42596 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1676037725
transform 1 0 43240 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1676037725
transform 1 0 12236 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1676037725
transform 1 0 41768 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1676037725
transform 1 0 42136 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1676037725
transform 1 0 43792 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1676037725
transform 1 0 45172 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1676037725
transform 1 0 45632 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1676037725
transform 1 0 41952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1676037725
transform 1 0 43700 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1676037725
transform 1 0 42780 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1676037725
transform 1 0 44988 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1676037725
transform 1 0 43056 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1676037725
transform 1 0 24472 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1676037725
transform 1 0 25024 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 1676037725
transform 1 0 31464 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input89_A
timestamp 1676037725
transform 1 0 25116 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input90_A
timestamp 1676037725
transform 1 0 28980 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input91_A
timestamp 1676037725
transform 1 0 28888 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input92_A
timestamp 1676037725
transform 1 0 29164 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input93_A
timestamp 1676037725
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input94_A
timestamp 1676037725
transform 1 0 31280 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input95_A
timestamp 1676037725
transform 1 0 33396 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input96_A
timestamp 1676037725
transform 1 0 35512 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input97_A
timestamp 1676037725
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input98_A
timestamp 1676037725
transform 1 0 44712 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input99_A
timestamp 1676037725
transform 1 0 43148 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input100_A
timestamp 1676037725
transform 1 0 44988 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input101_A
timestamp 1676037725
transform 1 0 47564 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input102_A
timestamp 1676037725
transform 1 0 46092 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input103_A
timestamp 1676037725
transform 1 0 47196 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input104_A
timestamp 1676037725
transform 1 0 47564 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input105_A
timestamp 1676037725
transform 1 0 47288 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input106_A
timestamp 1676037725
transform 1 0 46644 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input107_A
timestamp 1676037725
transform 1 0 46184 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input108_A
timestamp 1676037725
transform 1 0 45816 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input109_A
timestamp 1676037725
transform 1 0 45356 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input110_A
timestamp 1676037725
transform 1 0 45632 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 26588 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 24472 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25024 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 20148 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 19044 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 20608 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 22080 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 20516 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21252 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 23460 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 20700 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 23184 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 22724 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 21160 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21068 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 20792 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24288 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 25300 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 25208 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 27784 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 29072 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 27600 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 29164 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 30176 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 26680 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 29072 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 27600 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 22080 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 23920 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 31556 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 34316 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 34224 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 34224 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 36892 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 37260 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 36708 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 38456 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 39560 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 36800 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 36984 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 38640 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 35880 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 36892 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 37260 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 33304 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 34316 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 33488 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 34132 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 31740 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 28980 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 30636 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 32200 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 33304 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 34316 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 32752 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 31740 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 30176 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 29072 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 44988 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 33304 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 31832 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 34132 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 34684 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 36892 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 39284 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 36892 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 34408 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 34408 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 41032 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 41952 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 39468 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 41860 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 39468 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 39560 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 37628 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 35420 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 37628 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 41124 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 40020 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 42044 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 40940 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 41032 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 41492 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 42044 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 39836 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 40020 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 38916 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 34316 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 31740 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 27416 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 26680 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 26036 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 26588 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 25852 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 26404 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 26588 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25300 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24564 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24012 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21160 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21620 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21436 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21344 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 23828 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21896 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 12696 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 14996 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16284 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13524 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11500 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13340 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16836 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 17020 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18860 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 28152 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 25852 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 26220 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 20332 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_3.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 26404 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_3.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 27968 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_3.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 17388 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_5.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 26220 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_5.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 25852 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_5.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 19320 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 25484 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 25300 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 19412 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 18952 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 26588 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 19136 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 20516 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 25760 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 25944 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 22172 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 22356 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 25576 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 24380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 22264 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 22540 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 28980 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 25116 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 24564 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_37.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 30176 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_37.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_45.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 30176 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_left_track_53.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 24104 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 35880 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 27600 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 27600 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_2.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 33856 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_2.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 29072 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_2.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 29532 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 36984 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 30728 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 29256 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 33764 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 36432 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 36616 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 32752 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 34684 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 32936 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 30452 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 34500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 26220 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 26036 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 32292 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 26036 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 26680 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 31740 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 31832 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 25668 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 25484 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_36.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 30268 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_44.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 27784 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_right_track_52.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 35696 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 36708 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 42136 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 22724 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 28336 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 38456 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 42136 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 30728 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 31740 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_4.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 35696 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_4.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 35512 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_4.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 42228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_4.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 29716 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 42044 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 42412 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 42412 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 33672 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 34040 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 41768 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 42228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 34224 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 34408 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_10.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 37260 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_10.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 36892 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_10.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 41308 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_10.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 29256 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_12.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 41032 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_12.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 41216 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_12.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 38456 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_14.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 41584 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_14.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 34408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_16.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 41216 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_16.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 41400 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_16.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 36064 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_18.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 38824 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_18.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 39008 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_18.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 31832 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_20.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 28336 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_20.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 28520 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_20.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 24472 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_22.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 26864 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_22.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 27048 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_22.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 23644 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_24.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 27968 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_24.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 28152 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_24.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 21988 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_26.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 28428 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_26.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 28612 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_26.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 24012 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_28.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 24748 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_28.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_30.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 21344 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_30.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 23000 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_32.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16008 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_32.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_34.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16560 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_34.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16744 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_36.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_36.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 27140 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_36.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 23000 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_40.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 12788 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_42.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_42.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 17756 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_44.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 13708 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_44.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16376 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_46.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_48.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16560 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_48.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_50.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_1__0_.mux_top_track_58.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 26312 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18032 0 -1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16376 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16376 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 16836 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16836 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14260 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 14260 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 13616 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 13340 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 10764 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 9476 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 10948 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11684 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13248 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 10764 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 9108 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14444 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 15548 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2_
timestamp 1676037725
transform -1 0 16376 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3_
timestamp 1676037725
transform 1 0 20700 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4_
timestamp 1676037725
transform 1 0 15548 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15180 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 17112 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_2_
timestamp 1676037725
transform 1 0 16928 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3_
timestamp 1676037725
transform 1 0 18308 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3__254 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18676 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 15548 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_1_
timestamp 1676037725
transform 1 0 16652 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l4_in_0_
timestamp 1676037725
transform 1 0 17848 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19596 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 10396 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 12696 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2_
timestamp 1676037725
transform 1 0 19504 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3_
timestamp 1676037725
transform 1 0 16836 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4_
timestamp 1676037725
transform 1 0 17940 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_1_
timestamp 1676037725
transform 1 0 15548 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_2_
timestamp 1676037725
transform 1 0 12696 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3__255
timestamp 1676037725
transform 1 0 13524 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3_
timestamp 1676037725
transform 1 0 17112 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_0_
timestamp 1676037725
transform 1 0 13892 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_1_
timestamp 1676037725
transform 1 0 15548 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l4_in_0_
timestamp 1676037725
transform 1 0 15180 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17664 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 7728 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 7912 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 18124 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3_
timestamp 1676037725
transform 1 0 14444 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4_
timestamp 1676037725
transform 1 0 16744 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 9384 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 14260 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_2_
timestamp 1676037725
transform 1 0 14352 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3__256
timestamp 1676037725
transform 1 0 10948 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3_
timestamp 1676037725
transform 1 0 11684 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 11684 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_1_
timestamp 1676037725
transform 1 0 12328 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l4_in_0_
timestamp 1676037725
transform 1 0 12144 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 15548 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_1_
timestamp 1676037725
transform 1 0 14352 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2_
timestamp 1676037725
transform 1 0 15640 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3_
timestamp 1676037725
transform 1 0 18308 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4_
timestamp 1676037725
transform 1 0 15088 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 13156 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_1_
timestamp 1676037725
transform 1 0 15548 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_2_
timestamp 1676037725
transform 1 0 14352 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__257
timestamp 1676037725
transform 1 0 15732 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3_
timestamp 1676037725
transform 1 0 16376 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_0_
timestamp 1676037725
transform 1 0 11960 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_1_
timestamp 1676037725
transform 1 0 12972 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l4_in_0_
timestamp 1676037725
transform 1 0 11040 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14260 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27140 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23552 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22172 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21896 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14536 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 25116 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 22908 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 23276 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 20424 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20976 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 24196 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 23000 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 23552 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 18860 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 24196 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 24564 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 22264 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 27508 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 18032 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_2  cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 28888 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27140 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17940 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1676037725
transform 1 0 17848 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1676037725
transform 1 0 22448 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1676037725
transform 1 0 22540 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1676037725
transform 1 0 17756 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1676037725
transform 1 0 17940 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1676037725
transform 1 0 21988 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1676037725
transform 1 0 23276 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1676037725
transform 1 0 28796 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1676037725
transform 1 0 28244 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1676037725
transform 1 0 33304 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1676037725
transform 1 0 34040 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1676037725
transform 1 0 29900 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1676037725
transform 1 0 30728 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1676037725
transform 1 0 34592 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1676037725
transform 1 0 34868 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17
timestamp 1676037725
transform 1 0 2668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24
timestamp 1676037725
transform 1 0 3312 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1676037725
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1676037725
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1676037725
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_96
timestamp 1676037725
transform 1 0 9936 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100
timestamp 1676037725
transform 1 0 10304 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_132
timestamp 1676037725
transform 1 0 13248 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_159
timestamp 1676037725
transform 1 0 15732 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_187
timestamp 1676037725
transform 1 0 18308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1676037725
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_202
timestamp 1676037725
transform 1 0 19688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1676037725
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_225 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_247
timestamp 1676037725
transform 1 0 23828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1676037725
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_271
timestamp 1676037725
transform 1 0 26036 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_275
timestamp 1676037725
transform 1 0 26404 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1676037725
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1676037725
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_299
timestamp 1676037725
transform 1 0 28612 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 1676037725
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_311
timestamp 1676037725
transform 1 0 29716 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_326
timestamp 1676037725
transform 1 0 31096 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_330
timestamp 1676037725
transform 1 0 31464 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_337
timestamp 1676037725
transform 1 0 32108 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_345
timestamp 1676037725
transform 1 0 32844 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_349
timestamp 1676037725
transform 1 0 33212 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_353
timestamp 1676037725
transform 1 0 33580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1676037725
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_365
timestamp 1676037725
transform 1 0 34684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_372
timestamp 1676037725
transform 1 0 35328 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_376
timestamp 1676037725
transform 1 0 35696 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_388
timestamp 1676037725
transform 1 0 36800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1676037725
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_405
timestamp 1676037725
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp 1676037725
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_421
timestamp 1676037725
transform 1 0 39836 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_429
timestamp 1676037725
transform 1 0 40572 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_446
timestamp 1676037725
transform 1 0 42136 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_449
timestamp 1676037725
transform 1 0 42412 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_459
timestamp 1676037725
transform 1 0 43332 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_471
timestamp 1676037725
transform 1 0 44436 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_475
timestamp 1676037725
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_477
timestamp 1676037725
transform 1 0 44988 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_485
timestamp 1676037725
transform 1 0 45724 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_502
timestamp 1676037725
transform 1 0 47288 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_505
timestamp 1676037725
transform 1 0 47564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_525
timestamp 1676037725
transform 1 0 49404 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_9
timestamp 1676037725
transform 1 0 1932 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_19
timestamp 1676037725
transform 1 0 2852 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_31
timestamp 1676037725
transform 1 0 3956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_43
timestamp 1676037725
transform 1 0 5060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1676037725
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1676037725
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1676037725
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1676037725
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1676037725
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1676037725
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_137
timestamp 1676037725
transform 1 0 13708 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_145
timestamp 1676037725
transform 1 0 14444 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1676037725
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_171
timestamp 1676037725
transform 1 0 16836 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_180
timestamp 1676037725
transform 1 0 17664 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_184
timestamp 1676037725
transform 1 0 18032 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_201
timestamp 1676037725
transform 1 0 19596 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_208
timestamp 1676037725
transform 1 0 20240 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_215
timestamp 1676037725
transform 1 0 20884 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1676037725
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_235
timestamp 1676037725
transform 1 0 22724 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_247
timestamp 1676037725
transform 1 0 23828 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_271
timestamp 1676037725
transform 1 0 26036 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 1676037725
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_293
timestamp 1676037725
transform 1 0 28060 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_301
timestamp 1676037725
transform 1 0 28796 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_323
timestamp 1676037725
transform 1 0 30820 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_327
timestamp 1676037725
transform 1 0 31188 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1676037725
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1676037725
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1676037725
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1676037725
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1676037725
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1676037725
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1676037725
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1676037725
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1676037725
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1676037725
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1676037725
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1676037725
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1676037725
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1676037725
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_461
timestamp 1676037725
transform 1 0 43516 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_465
timestamp 1676037725
transform 1 0 43884 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_482
timestamp 1676037725
transform 1 0 45448 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_502
timestamp 1676037725
transform 1 0 47288 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_505
timestamp 1676037725
transform 1 0 47564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_525
timestamp 1676037725
transform 1 0 49404 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1676037725
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1676037725
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1676037725
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1676037725
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1676037725
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1676037725
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_165
timestamp 1676037725
transform 1 0 16284 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_170
timestamp 1676037725
transform 1 0 16744 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_182
timestamp 1676037725
transform 1 0 17848 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1676037725
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_209
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_215
timestamp 1676037725
transform 1 0 20884 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_236
timestamp 1676037725
transform 1 0 22816 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_240
timestamp 1676037725
transform 1 0 23184 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1676037725
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_276
timestamp 1676037725
transform 1 0 26496 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_288
timestamp 1676037725
transform 1 0 27600 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_300
timestamp 1676037725
transform 1 0 28704 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1676037725
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1676037725
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1676037725
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1676037725
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1676037725
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1676037725
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1676037725
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_377
timestamp 1676037725
transform 1 0 35788 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_387
timestamp 1676037725
transform 1 0 36708 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_391
timestamp 1676037725
transform 1 0 37076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_403
timestamp 1676037725
transform 1 0 38180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_415
timestamp 1676037725
transform 1 0 39284 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1676037725
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1676037725
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1676037725
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1676037725
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1676037725
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1676037725
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1676037725
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_479
timestamp 1676037725
transform 1 0 45172 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_485
timestamp 1676037725
transform 1 0 45724 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_505
timestamp 1676037725
transform 1 0 47564 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_525
timestamp 1676037725
transform 1 0 49404 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_9
timestamp 1676037725
transform 1 0 1932 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_17
timestamp 1676037725
transform 1 0 2668 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_23
timestamp 1676037725
transform 1 0 3220 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_35
timestamp 1676037725
transform 1 0 4324 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_47
timestamp 1676037725
transform 1 0 5428 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1676037725
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1676037725
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1676037725
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1676037725
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1676037725
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_229
timestamp 1676037725
transform 1 0 22172 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_233
timestamp 1676037725
transform 1 0 22540 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_240
timestamp 1676037725
transform 1 0 23184 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_247
timestamp 1676037725
transform 1 0 23828 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_272
timestamp 1676037725
transform 1 0 26128 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_304
timestamp 1676037725
transform 1 0 29072 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_316
timestamp 1676037725
transform 1 0 30176 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_328
timestamp 1676037725
transform 1 0 31280 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1676037725
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1676037725
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1676037725
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1676037725
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1676037725
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1676037725
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1676037725
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1676037725
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1676037725
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1676037725
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1676037725
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1676037725
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1676037725
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1676037725
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1676037725
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_485
timestamp 1676037725
transform 1 0 45724 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_502
timestamp 1676037725
transform 1 0 47288 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_507
timestamp 1676037725
transform 1 0 47748 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_525
timestamp 1676037725
transform 1 0 49404 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_9
timestamp 1676037725
transform 1 0 1932 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1676037725
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1676037725
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1676037725
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1676037725
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_209
timestamp 1676037725
transform 1 0 20332 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_218
timestamp 1676037725
transform 1 0 21160 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_234
timestamp 1676037725
transform 1 0 22632 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_241
timestamp 1676037725
transform 1 0 23276 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_249
timestamp 1676037725
transform 1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_282
timestamp 1676037725
transform 1 0 27048 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_294
timestamp 1676037725
transform 1 0 28152 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_306
timestamp 1676037725
transform 1 0 29256 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1676037725
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1676037725
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1676037725
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1676037725
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1676037725
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1676037725
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1676037725
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_377
timestamp 1676037725
transform 1 0 35788 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_385
timestamp 1676037725
transform 1 0 36524 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_390
timestamp 1676037725
transform 1 0 36984 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_396
timestamp 1676037725
transform 1 0 37536 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_404
timestamp 1676037725
transform 1 0 38272 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_408
timestamp 1676037725
transform 1 0 38640 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1676037725
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1676037725
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1676037725
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1676037725
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1676037725
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1676037725
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1676037725
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_491
timestamp 1676037725
transform 1 0 46276 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_497
timestamp 1676037725
transform 1 0 46828 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_505
timestamp 1676037725
transform 1 0 47564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_525
timestamp 1676037725
transform 1 0 49404 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1676037725
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1676037725
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1676037725
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1676037725
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1676037725
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_201
timestamp 1676037725
transform 1 0 19596 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_213
timestamp 1676037725
transform 1 0 20700 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_221
timestamp 1676037725
transform 1 0 21436 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1676037725
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1676037725
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1676037725
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1676037725
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1676037725
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1676037725
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1676037725
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1676037725
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1676037725
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1676037725
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1676037725
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1676037725
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1676037725
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1676037725
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1676037725
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1676037725
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_395
timestamp 1676037725
transform 1 0 37444 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_401
timestamp 1676037725
transform 1 0 37996 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_409
timestamp 1676037725
transform 1 0 38732 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_413
timestamp 1676037725
transform 1 0 39100 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_425
timestamp 1676037725
transform 1 0 40204 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_437
timestamp 1676037725
transform 1 0 41308 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_445
timestamp 1676037725
transform 1 0 42044 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1676037725
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1676037725
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1676037725
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_485
timestamp 1676037725
transform 1 0 45724 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_502
timestamp 1676037725
transform 1 0 47288 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_505
timestamp 1676037725
transform 1 0 47564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_525
timestamp 1676037725
transform 1 0 49404 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_9
timestamp 1676037725
transform 1 0 1932 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_17
timestamp 1676037725
transform 1 0 2668 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_23
timestamp 1676037725
transform 1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1676037725
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1676037725
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1676037725
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1676037725
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1676037725
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1676037725
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1676037725
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1676037725
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1676037725
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1676037725
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1676037725
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1676037725
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1676037725
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1676037725
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1676037725
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1676037725
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1676037725
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1676037725
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1676037725
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1676037725
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1676037725
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1676037725
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1676037725
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1676037725
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1676037725
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1676037725
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1676037725
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1676037725
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_457
timestamp 1676037725
transform 1 0 43148 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_461
timestamp 1676037725
transform 1 0 43516 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_466
timestamp 1676037725
transform 1 0 43976 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_474
timestamp 1676037725
transform 1 0 44712 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1676037725
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1676037725
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_501
timestamp 1676037725
transform 1 0 47196 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_525
timestamp 1676037725
transform 1 0 49404 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_9
timestamp 1676037725
transform 1 0 1932 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1676037725
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1676037725
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1676037725
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1676037725
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1676037725
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_192
timestamp 1676037725
transform 1 0 18768 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_204
timestamp 1676037725
transform 1 0 19872 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_216
timestamp 1676037725
transform 1 0 20976 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1676037725
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1676037725
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1676037725
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1676037725
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1676037725
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1676037725
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1676037725
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1676037725
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1676037725
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1676037725
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1676037725
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1676037725
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1676037725
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1676037725
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1676037725
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1676037725
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_393
timestamp 1676037725
transform 1 0 37260 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_399
timestamp 1676037725
transform 1 0 37812 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_403
timestamp 1676037725
transform 1 0 38180 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_415
timestamp 1676037725
transform 1 0 39284 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_427
timestamp 1676037725
transform 1 0 40388 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_439
timestamp 1676037725
transform 1 0 41492 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1676037725
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1676037725
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_461
timestamp 1676037725
transform 1 0 43516 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_469
timestamp 1676037725
transform 1 0 44252 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_481
timestamp 1676037725
transform 1 0 45356 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_493
timestamp 1676037725
transform 1 0 46460 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_501
timestamp 1676037725
transform 1 0 47196 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_505
timestamp 1676037725
transform 1 0 47564 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_525
timestamp 1676037725
transform 1 0 49404 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_9
timestamp 1676037725
transform 1 0 1932 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_16
timestamp 1676037725
transform 1 0 2576 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_20
timestamp 1676037725
transform 1 0 2944 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1676037725
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1676037725
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1676037725
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1676037725
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_177
timestamp 1676037725
transform 1 0 17388 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_183
timestamp 1676037725
transform 1 0 17940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1676037725
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_204
timestamp 1676037725
transform 1 0 19872 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_216
timestamp 1676037725
transform 1 0 20976 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_228
timestamp 1676037725
transform 1 0 22080 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_240
timestamp 1676037725
transform 1 0 23184 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1676037725
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1676037725
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1676037725
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1676037725
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1676037725
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1676037725
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1676037725
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1676037725
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1676037725
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1676037725
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1676037725
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1676037725
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1676037725
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1676037725
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1676037725
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1676037725
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1676037725
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1676037725
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1676037725
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1676037725
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1676037725
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1676037725
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1676037725
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1676037725
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_505
timestamp 1676037725
transform 1 0 47564 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_525
timestamp 1676037725
transform 1 0 49404 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_9
timestamp 1676037725
transform 1 0 1932 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_13
timestamp 1676037725
transform 1 0 2300 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_25
timestamp 1676037725
transform 1 0 3404 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_37
timestamp 1676037725
transform 1 0 4508 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_49
timestamp 1676037725
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1676037725
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1676037725
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1676037725
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1676037725
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1676037725
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1676037725
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_181
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_185
timestamp 1676037725
transform 1 0 18124 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_188
timestamp 1676037725
transform 1 0 18400 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1676037725
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1676037725
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_217
timestamp 1676037725
transform 1 0 21068 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_236
timestamp 1676037725
transform 1 0 22816 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_240
timestamp 1676037725
transform 1 0 23184 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_252
timestamp 1676037725
transform 1 0 24288 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_264
timestamp 1676037725
transform 1 0 25392 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_276
timestamp 1676037725
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1676037725
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1676037725
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_317
timestamp 1676037725
transform 1 0 30268 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_323
timestamp 1676037725
transform 1 0 30820 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_327
timestamp 1676037725
transform 1 0 31188 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1676037725
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_337
timestamp 1676037725
transform 1 0 32108 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_342
timestamp 1676037725
transform 1 0 32568 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_346
timestamp 1676037725
transform 1 0 32936 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_358
timestamp 1676037725
transform 1 0 34040 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_370
timestamp 1676037725
transform 1 0 35144 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_382
timestamp 1676037725
transform 1 0 36248 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_390
timestamp 1676037725
transform 1 0 36984 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_393
timestamp 1676037725
transform 1 0 37260 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_396
timestamp 1676037725
transform 1 0 37536 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_402
timestamp 1676037725
transform 1 0 38088 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_410
timestamp 1676037725
transform 1 0 38824 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_414
timestamp 1676037725
transform 1 0 39192 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_426
timestamp 1676037725
transform 1 0 40296 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_438
timestamp 1676037725
transform 1 0 41400 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_446
timestamp 1676037725
transform 1 0 42136 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1676037725
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1676037725
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_473
timestamp 1676037725
transform 1 0 44620 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_479
timestamp 1676037725
transform 1 0 45172 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_491
timestamp 1676037725
transform 1 0 46276 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1676037725
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_505
timestamp 1676037725
transform 1 0 47564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_525
timestamp 1676037725
transform 1 0 49404 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_9
timestamp 1676037725
transform 1 0 1932 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1676037725
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1676037725
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1676037725
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1676037725
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1676037725
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1676037725
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1676037725
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_153
timestamp 1676037725
transform 1 0 15180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_160
timestamp 1676037725
transform 1 0 15824 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_168
timestamp 1676037725
transform 1 0 16560 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_178
timestamp 1676037725
transform 1 0 17480 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_191
timestamp 1676037725
transform 1 0 18676 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_219
timestamp 1676037725
transform 1 0 21252 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_225
timestamp 1676037725
transform 1 0 21804 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_236
timestamp 1676037725
transform 1 0 22816 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_240
timestamp 1676037725
transform 1 0 23184 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1676037725
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1676037725
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1676037725
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1676037725
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1676037725
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1676037725
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_314
timestamp 1676037725
transform 1 0 29992 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_323
timestamp 1676037725
transform 1 0 30820 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_334
timestamp 1676037725
transform 1 0 31832 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_338
timestamp 1676037725
transform 1 0 32200 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_348
timestamp 1676037725
transform 1 0 33120 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_360
timestamp 1676037725
transform 1 0 34224 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1676037725
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1676037725
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_389
timestamp 1676037725
transform 1 0 36892 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_395
timestamp 1676037725
transform 1 0 37444 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_398
timestamp 1676037725
transform 1 0 37720 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_404
timestamp 1676037725
transform 1 0 38272 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_412
timestamp 1676037725
transform 1 0 39008 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_416
timestamp 1676037725
transform 1 0 39376 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1676037725
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1676037725
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1676037725
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1676037725
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1676037725
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1676037725
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1676037725
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1676037725
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_501
timestamp 1676037725
transform 1 0 47196 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_525
timestamp 1676037725
transform 1 0 49404 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1676037725
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1676037725
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1676037725
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1676037725
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1676037725
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1676037725
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_125
timestamp 1676037725
transform 1 0 12604 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_133
timestamp 1676037725
transform 1 0 13340 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_156
timestamp 1676037725
transform 1 0 15456 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_160
timestamp 1676037725
transform 1 0 15824 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_191
timestamp 1676037725
transform 1 0 18676 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_198
timestamp 1676037725
transform 1 0 19320 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1676037725
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_247
timestamp 1676037725
transform 1 0 23828 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_251
timestamp 1676037725
transform 1 0 24196 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_263
timestamp 1676037725
transform 1 0 25300 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_275
timestamp 1676037725
transform 1 0 26404 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1676037725
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1676037725
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_293
timestamp 1676037725
transform 1 0 28060 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_321
timestamp 1676037725
transform 1 0 30636 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_334
timestamp 1676037725
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_337
timestamp 1676037725
transform 1 0 32108 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_359
timestamp 1676037725
transform 1 0 34132 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_363
timestamp 1676037725
transform 1 0 34500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_375
timestamp 1676037725
transform 1 0 35604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_387
timestamp 1676037725
transform 1 0 36708 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1676037725
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_393
timestamp 1676037725
transform 1 0 37260 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_398
timestamp 1676037725
transform 1 0 37720 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_410
timestamp 1676037725
transform 1 0 38824 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_414
timestamp 1676037725
transform 1 0 39192 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_422
timestamp 1676037725
transform 1 0 39928 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_429
timestamp 1676037725
transform 1 0 40572 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_433
timestamp 1676037725
transform 1 0 40940 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_445
timestamp 1676037725
transform 1 0 42044 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1676037725
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_461
timestamp 1676037725
transform 1 0 43516 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_471
timestamp 1676037725
transform 1 0 44436 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_483
timestamp 1676037725
transform 1 0 45540 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_502
timestamp 1676037725
transform 1 0 47288 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_505
timestamp 1676037725
transform 1 0 47564 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_525
timestamp 1676037725
transform 1 0 49404 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_9
timestamp 1676037725
transform 1 0 1932 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_17
timestamp 1676037725
transform 1 0 2668 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_23
timestamp 1676037725
transform 1 0 3220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1676037725
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1676037725
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1676037725
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1676037725
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_146
timestamp 1676037725
transform 1 0 14536 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_151
timestamp 1676037725
transform 1 0 14996 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_162
timestamp 1676037725
transform 1 0 16008 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_186
timestamp 1676037725
transform 1 0 18216 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_190
timestamp 1676037725
transform 1 0 18584 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1676037725
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_219
timestamp 1676037725
transform 1 0 21252 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_226
timestamp 1676037725
transform 1 0 21896 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1676037725
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_259
timestamp 1676037725
transform 1 0 24932 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_269
timestamp 1676037725
transform 1 0 25852 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_281
timestamp 1676037725
transform 1 0 26956 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_289
timestamp 1676037725
transform 1 0 27692 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_292
timestamp 1676037725
transform 1 0 27968 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_303
timestamp 1676037725
transform 1 0 28980 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1676037725
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_309
timestamp 1676037725
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_314
timestamp 1676037725
transform 1 0 29992 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_318
timestamp 1676037725
transform 1 0 30360 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_342
timestamp 1676037725
transform 1 0 32568 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_348
timestamp 1676037725
transform 1 0 33120 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_359
timestamp 1676037725
transform 1 0 34132 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1676037725
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_365
timestamp 1676037725
transform 1 0 34684 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_376
timestamp 1676037725
transform 1 0 35696 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_384
timestamp 1676037725
transform 1 0 36432 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_388
timestamp 1676037725
transform 1 0 36800 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_396
timestamp 1676037725
transform 1 0 37536 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_400
timestamp 1676037725
transform 1 0 37904 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_412
timestamp 1676037725
transform 1 0 39008 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_418
timestamp 1676037725
transform 1 0 39560 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_423
timestamp 1676037725
transform 1 0 40020 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_435
timestamp 1676037725
transform 1 0 41124 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_447
timestamp 1676037725
transform 1 0 42228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_459
timestamp 1676037725
transform 1 0 43332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_471
timestamp 1676037725
transform 1 0 44436 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1676037725
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1676037725
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1676037725
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_501
timestamp 1676037725
transform 1 0 47196 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_525
timestamp 1676037725
transform 1 0 49404 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_9
timestamp 1676037725
transform 1 0 1932 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1676037725
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1676037725
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1676037725
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1676037725
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1676037725
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1676037725
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1676037725
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1676037725
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1676037725
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_119
timestamp 1676037725
transform 1 0 12052 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_129
timestamp 1676037725
transform 1 0 12972 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_156
timestamp 1676037725
transform 1 0 15456 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_194
timestamp 1676037725
transform 1 0 18952 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_218
timestamp 1676037725
transform 1 0 21160 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_228
timestamp 1676037725
transform 1 0 22080 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_239
timestamp 1676037725
transform 1 0 23092 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_263
timestamp 1676037725
transform 1 0 25300 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_276
timestamp 1676037725
transform 1 0 26496 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_281
timestamp 1676037725
transform 1 0 26956 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_307
timestamp 1676037725
transform 1 0 29348 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_331
timestamp 1676037725
transform 1 0 31556 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1676037725
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_337
timestamp 1676037725
transform 1 0 32108 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_340
timestamp 1676037725
transform 1 0 32384 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_351
timestamp 1676037725
transform 1 0 33396 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_355
timestamp 1676037725
transform 1 0 33764 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_376
timestamp 1676037725
transform 1 0 35696 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_380
timestamp 1676037725
transform 1 0 36064 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1676037725
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1676037725
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1676037725
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1676037725
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1676037725
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1676037725
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1676037725
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1676037725
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1676037725
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1676037725
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1676037725
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1676037725
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_505
timestamp 1676037725
transform 1 0 47564 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_525
timestamp 1676037725
transform 1 0 49404 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1676037725
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1676037725
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1676037725
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_121
timestamp 1676037725
transform 1 0 12236 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_124
timestamp 1676037725
transform 1 0 12512 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_135
timestamp 1676037725
transform 1 0 13524 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_163
timestamp 1676037725
transform 1 0 16100 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_170
timestamp 1676037725
transform 1 0 16744 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_181
timestamp 1676037725
transform 1 0 17756 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1676037725
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_203
timestamp 1676037725
transform 1 0 19780 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_207
timestamp 1676037725
transform 1 0 20148 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_228
timestamp 1676037725
transform 1 0 22080 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_243
timestamp 1676037725
transform 1 0 23460 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1676037725
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_275
timestamp 1676037725
transform 1 0 26404 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_279
timestamp 1676037725
transform 1 0 26772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_301
timestamp 1676037725
transform 1 0 28796 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_305
timestamp 1676037725
transform 1 0 29164 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_309
timestamp 1676037725
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_314
timestamp 1676037725
transform 1 0 29992 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_338
timestamp 1676037725
transform 1 0 32200 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_351
timestamp 1676037725
transform 1 0 33396 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_358
timestamp 1676037725
transform 1 0 34040 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_365
timestamp 1676037725
transform 1 0 34684 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_387
timestamp 1676037725
transform 1 0 36708 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_391
timestamp 1676037725
transform 1 0 37076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_407
timestamp 1676037725
transform 1 0 38548 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_411
timestamp 1676037725
transform 1 0 38916 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1676037725
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_421
timestamp 1676037725
transform 1 0 39836 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_427
timestamp 1676037725
transform 1 0 40388 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_431
timestamp 1676037725
transform 1 0 40756 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_443
timestamp 1676037725
transform 1 0 41860 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_455
timestamp 1676037725
transform 1 0 42964 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_467
timestamp 1676037725
transform 1 0 44068 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_473
timestamp 1676037725
transform 1 0 44620 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1676037725
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_505
timestamp 1676037725
transform 1 0 47564 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_525
timestamp 1676037725
transform 1 0 49404 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_9
timestamp 1676037725
transform 1 0 1932 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_17
timestamp 1676037725
transform 1 0 2668 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_23
timestamp 1676037725
transform 1 0 3220 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_35
timestamp 1676037725
transform 1 0 4324 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_47
timestamp 1676037725
transform 1 0 5428 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1676037725
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1676037725
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1676037725
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1676037725
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1676037725
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_129
timestamp 1676037725
transform 1 0 12972 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_140
timestamp 1676037725
transform 1 0 13984 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_153
timestamp 1676037725
transform 1 0 15180 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1676037725
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_172
timestamp 1676037725
transform 1 0 16928 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_183
timestamp 1676037725
transform 1 0 17940 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_196
timestamp 1676037725
transform 1 0 19136 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_209
timestamp 1676037725
transform 1 0 20332 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1676037725
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_247
timestamp 1676037725
transform 1 0 23828 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_260
timestamp 1676037725
transform 1 0 25024 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_267
timestamp 1676037725
transform 1 0 25668 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_277
timestamp 1676037725
transform 1 0 26588 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1676037725
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_292
timestamp 1676037725
transform 1 0 27968 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_296
timestamp 1676037725
transform 1 0 28336 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_299
timestamp 1676037725
transform 1 0 28612 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_312
timestamp 1676037725
transform 1 0 29808 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_325
timestamp 1676037725
transform 1 0 31004 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_332
timestamp 1676037725
transform 1 0 31648 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_337
timestamp 1676037725
transform 1 0 32108 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_348
timestamp 1676037725
transform 1 0 33120 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_352
timestamp 1676037725
transform 1 0 33488 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_376
timestamp 1676037725
transform 1 0 35696 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_389
timestamp 1676037725
transform 1 0 36892 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_395
timestamp 1676037725
transform 1 0 37444 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_407
timestamp 1676037725
transform 1 0 38548 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_423
timestamp 1676037725
transform 1 0 40020 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_427
timestamp 1676037725
transform 1 0 40388 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_439
timestamp 1676037725
transform 1 0 41492 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1676037725
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1676037725
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1676037725
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1676037725
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1676037725
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1676037725
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1676037725
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_505
timestamp 1676037725
transform 1 0 47564 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_525
timestamp 1676037725
transform 1 0 49404 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_9
timestamp 1676037725
transform 1 0 1932 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1676037725
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1676037725
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1676037725
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1676037725
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_97
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_105
timestamp 1676037725
transform 1 0 10764 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_127
timestamp 1676037725
transform 1 0 12788 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_133
timestamp 1676037725
transform 1 0 13340 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1676037725
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_153
timestamp 1676037725
transform 1 0 15180 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_166
timestamp 1676037725
transform 1 0 16376 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_179
timestamp 1676037725
transform 1 0 17572 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_192
timestamp 1676037725
transform 1 0 18768 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_201
timestamp 1676037725
transform 1 0 19596 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_206
timestamp 1676037725
transform 1 0 20056 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_230
timestamp 1676037725
transform 1 0 22264 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_237
timestamp 1676037725
transform 1 0 22908 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1676037725
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_275
timestamp 1676037725
transform 1 0 26404 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_279
timestamp 1676037725
transform 1 0 26772 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_300
timestamp 1676037725
transform 1 0 28704 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1676037725
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_320
timestamp 1676037725
transform 1 0 30544 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_324
timestamp 1676037725
transform 1 0 30912 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_346
timestamp 1676037725
transform 1 0 32936 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_361
timestamp 1676037725
transform 1 0 34316 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_367
timestamp 1676037725
transform 1 0 34868 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_375
timestamp 1676037725
transform 1 0 35604 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_399
timestamp 1676037725
transform 1 0 37812 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_406
timestamp 1676037725
transform 1 0 38456 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_410
timestamp 1676037725
transform 1 0 38824 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_421
timestamp 1676037725
transform 1 0 39836 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_427
timestamp 1676037725
transform 1 0 40388 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_434
timestamp 1676037725
transform 1 0 41032 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_446
timestamp 1676037725
transform 1 0 42136 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_458
timestamp 1676037725
transform 1 0 43240 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_470
timestamp 1676037725
transform 1 0 44344 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_477
timestamp 1676037725
transform 1 0 44988 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_487
timestamp 1676037725
transform 1 0 45908 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_499
timestamp 1676037725
transform 1 0 47012 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_507
timestamp 1676037725
transform 1 0 47748 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_525
timestamp 1676037725
transform 1 0 49404 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_9
timestamp 1676037725
transform 1 0 1932 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_16
timestamp 1676037725
transform 1 0 2576 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_20
timestamp 1676037725
transform 1 0 2944 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_32
timestamp 1676037725
transform 1 0 4048 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_44
timestamp 1676037725
transform 1 0 5152 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1676037725
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1676037725
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1676037725
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1676037725
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1676037725
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_115
timestamp 1676037725
transform 1 0 11684 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1676037725
transform 1 0 12236 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_131
timestamp 1676037725
transform 1 0 13156 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_137
timestamp 1676037725
transform 1 0 13708 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_148
timestamp 1676037725
transform 1 0 14720 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_161
timestamp 1676037725
transform 1 0 15916 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_191
timestamp 1676037725
transform 1 0 18676 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_198
timestamp 1676037725
transform 1 0 19320 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_209
timestamp 1676037725
transform 1 0 20332 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1676037725
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_231
timestamp 1676037725
transform 1 0 22356 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_244
timestamp 1676037725
transform 1 0 23552 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_268
timestamp 1676037725
transform 1 0 25760 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_273
timestamp 1676037725
transform 1 0 26220 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_278
timestamp 1676037725
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1676037725
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_292
timestamp 1676037725
transform 1 0 27968 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_296
timestamp 1676037725
transform 1 0 28336 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_318
timestamp 1676037725
transform 1 0 30360 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_331
timestamp 1676037725
transform 1 0 31556 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1676037725
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_337
timestamp 1676037725
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_348
timestamp 1676037725
transform 1 0 33120 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_361
timestamp 1676037725
transform 1 0 34316 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_369
timestamp 1676037725
transform 1 0 35052 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_390
timestamp 1676037725
transform 1 0 36984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_393
timestamp 1676037725
transform 1 0 37260 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_404
timestamp 1676037725
transform 1 0 38272 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_417
timestamp 1676037725
transform 1 0 39468 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_425
timestamp 1676037725
transform 1 0 40204 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_429
timestamp 1676037725
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1676037725
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1676037725
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1676037725
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1676037725
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_473
timestamp 1676037725
transform 1 0 44620 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_481
timestamp 1676037725
transform 1 0 45356 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_493
timestamp 1676037725
transform 1 0 46460 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_501
timestamp 1676037725
transform 1 0 47196 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_505
timestamp 1676037725
transform 1 0 47564 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_525
timestamp 1676037725
transform 1 0 49404 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_19
timestamp 1676037725
transform 1 0 2852 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1676037725
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1676037725
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1676037725
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_111
timestamp 1676037725
transform 1 0 11316 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1676037725
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_164
timestamp 1676037725
transform 1 0 16192 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_168
timestamp 1676037725
transform 1 0 16560 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_179
timestamp 1676037725
transform 1 0 17572 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1676037725
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_208
timestamp 1676037725
transform 1 0 20240 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_213
timestamp 1676037725
transform 1 0 20700 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_224
timestamp 1676037725
transform 1 0 21712 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_237
timestamp 1676037725
transform 1 0 22908 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1676037725
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_275
timestamp 1676037725
transform 1 0 26404 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_279
timestamp 1676037725
transform 1 0 26772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_290
timestamp 1676037725
transform 1 0 27784 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_294
timestamp 1676037725
transform 1 0 28152 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_306
timestamp 1676037725
transform 1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_309
timestamp 1676037725
transform 1 0 29532 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_331
timestamp 1676037725
transform 1 0 31556 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_335
timestamp 1676037725
transform 1 0 31924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_357
timestamp 1676037725
transform 1 0 33948 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1676037725
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_365
timestamp 1676037725
transform 1 0 34684 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_387
timestamp 1676037725
transform 1 0 36708 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_400
timestamp 1676037725
transform 1 0 37904 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_413
timestamp 1676037725
transform 1 0 39100 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_421
timestamp 1676037725
transform 1 0 39836 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_427
timestamp 1676037725
transform 1 0 40388 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_434
timestamp 1676037725
transform 1 0 41032 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_441
timestamp 1676037725
transform 1 0 41676 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_453
timestamp 1676037725
transform 1 0 42780 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_465
timestamp 1676037725
transform 1 0 43884 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_473
timestamp 1676037725
transform 1 0 44620 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_477
timestamp 1676037725
transform 1 0 44988 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_485
timestamp 1676037725
transform 1 0 45724 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_490
timestamp 1676037725
transform 1 0 46184 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_502
timestamp 1676037725
transform 1 0 47288 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_508
timestamp 1676037725
transform 1 0 47840 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_525
timestamp 1676037725
transform 1 0 49404 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_9
timestamp 1676037725
transform 1 0 1932 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_13
timestamp 1676037725
transform 1 0 2300 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_22
timestamp 1676037725
transform 1 0 3128 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_26
timestamp 1676037725
transform 1 0 3496 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_38
timestamp 1676037725
transform 1 0 4600 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_50
timestamp 1676037725
transform 1 0 5704 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1676037725
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1676037725
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1676037725
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_105
timestamp 1676037725
transform 1 0 10764 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_109
timestamp 1676037725
transform 1 0 11132 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_124
timestamp 1676037725
transform 1 0 12512 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_128
timestamp 1676037725
transform 1 0 12880 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_150
timestamp 1676037725
transform 1 0 14904 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_155
timestamp 1676037725
transform 1 0 15364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1676037725
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_173
timestamp 1676037725
transform 1 0 17020 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_178
timestamp 1676037725
transform 1 0 17480 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_193
timestamp 1676037725
transform 1 0 18860 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_206
timestamp 1676037725
transform 1 0 20056 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_211
timestamp 1676037725
transform 1 0 20516 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1676037725
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_230
timestamp 1676037725
transform 1 0 22264 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_243
timestamp 1676037725
transform 1 0 23460 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_267
timestamp 1676037725
transform 1 0 25668 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_275
timestamp 1676037725
transform 1 0 26404 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_281
timestamp 1676037725
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_306
timestamp 1676037725
transform 1 0 29256 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_311
timestamp 1676037725
transform 1 0 29716 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_334
timestamp 1676037725
transform 1 0 31832 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_337
timestamp 1676037725
transform 1 0 32108 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_348
timestamp 1676037725
transform 1 0 33120 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_356
timestamp 1676037725
transform 1 0 33856 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_369
timestamp 1676037725
transform 1 0 35052 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_382
timestamp 1676037725
transform 1 0 36248 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_393
timestamp 1676037725
transform 1 0 37260 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_418
timestamp 1676037725
transform 1 0 39560 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_426
timestamp 1676037725
transform 1 0 40296 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_430
timestamp 1676037725
transform 1 0 40664 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_442
timestamp 1676037725
transform 1 0 41768 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1676037725
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1676037725
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1676037725
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_485
timestamp 1676037725
transform 1 0 45724 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_490
timestamp 1676037725
transform 1 0 46184 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_502
timestamp 1676037725
transform 1 0 47288 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_505
timestamp 1676037725
transform 1 0 47564 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_525
timestamp 1676037725
transform 1 0 49404 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_21
timestamp 1676037725
transform 1 0 3036 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1676037725
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1676037725
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1676037725
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_97
timestamp 1676037725
transform 1 0 10028 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_126
timestamp 1676037725
transform 1 0 12696 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_133
timestamp 1676037725
transform 1 0 13340 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_147
timestamp 1676037725
transform 1 0 14628 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1676037725
transform 1 0 14996 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_162
timestamp 1676037725
transform 1 0 16008 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_187
timestamp 1676037725
transform 1 0 18308 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1676037725
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_200
timestamp 1676037725
transform 1 0 19504 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_211
timestamp 1676037725
transform 1 0 20516 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_224
timestamp 1676037725
transform 1 0 21712 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_237
timestamp 1676037725
transform 1 0 22908 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1676037725
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_256
timestamp 1676037725
transform 1 0 24656 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_267
timestamp 1676037725
transform 1 0 25668 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_274
timestamp 1676037725
transform 1 0 26312 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_280
timestamp 1676037725
transform 1 0 26864 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_290
timestamp 1676037725
transform 1 0 27784 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_295
timestamp 1676037725
transform 1 0 28244 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_306
timestamp 1676037725
transform 1 0 29256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_309
timestamp 1676037725
transform 1 0 29532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_320
timestamp 1676037725
transform 1 0 30544 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_324
timestamp 1676037725
transform 1 0 30912 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_346
timestamp 1676037725
transform 1 0 32936 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_359
timestamp 1676037725
transform 1 0 34132 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1676037725
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_365
timestamp 1676037725
transform 1 0 34684 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_376
timestamp 1676037725
transform 1 0 35696 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_382
timestamp 1676037725
transform 1 0 36248 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_404
timestamp 1676037725
transform 1 0 38272 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_408
timestamp 1676037725
transform 1 0 38640 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1676037725
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_433
timestamp 1676037725
transform 1 0 40940 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_440
timestamp 1676037725
transform 1 0 41584 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_452
timestamp 1676037725
transform 1 0 42688 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_464
timestamp 1676037725
transform 1 0 43792 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1676037725
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1676037725
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_501
timestamp 1676037725
transform 1 0 47196 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_525
timestamp 1676037725
transform 1 0 49404 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_21
timestamp 1676037725
transform 1 0 3036 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_29
timestamp 1676037725
transform 1 0 3772 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_33
timestamp 1676037725
transform 1 0 4140 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_45
timestamp 1676037725
transform 1 0 5244 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1676037725
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1676037725
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_93
timestamp 1676037725
transform 1 0 9660 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_97
timestamp 1676037725
transform 1 0 10028 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_105
timestamp 1676037725
transform 1 0 10764 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1676037725
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_124
timestamp 1676037725
transform 1 0 12512 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_128
timestamp 1676037725
transform 1 0 12880 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_149
timestamp 1676037725
transform 1 0 14812 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_155
timestamp 1676037725
transform 1 0 15364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1676037725
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_172
timestamp 1676037725
transform 1 0 16928 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_183
timestamp 1676037725
transform 1 0 17940 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_196
timestamp 1676037725
transform 1 0 19136 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_200
timestamp 1676037725
transform 1 0 19504 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1676037725
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_247
timestamp 1676037725
transform 1 0 23828 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_254
timestamp 1676037725
transform 1 0 24472 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1676037725
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1676037725
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_303
timestamp 1676037725
transform 1 0 28980 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_327
timestamp 1676037725
transform 1 0 31188 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_334
timestamp 1676037725
transform 1 0 31832 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_337
timestamp 1676037725
transform 1 0 32108 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_359
timestamp 1676037725
transform 1 0 34132 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_372
timestamp 1676037725
transform 1 0 35328 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_385
timestamp 1676037725
transform 1 0 36524 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_389
timestamp 1676037725
transform 1 0 36892 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_393
timestamp 1676037725
transform 1 0 37260 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_404
timestamp 1676037725
transform 1 0 38272 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_410
timestamp 1676037725
transform 1 0 38824 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_413
timestamp 1676037725
transform 1 0 39100 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_425
timestamp 1676037725
transform 1 0 40204 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_437
timestamp 1676037725
transform 1 0 41308 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_445
timestamp 1676037725
transform 1 0 42044 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1676037725
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1676037725
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_473
timestamp 1676037725
transform 1 0 44620 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_480
timestamp 1676037725
transform 1 0 45264 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_487
timestamp 1676037725
transform 1 0 45908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_499
timestamp 1676037725
transform 1 0 47012 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1676037725
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_505
timestamp 1676037725
transform 1 0 47564 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_509
timestamp 1676037725
transform 1 0 47932 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_512
timestamp 1676037725
transform 1 0 48208 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_517
timestamp 1676037725
transform 1 0 48668 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_525
timestamp 1676037725
transform 1 0 49404 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_21
timestamp 1676037725
transform 1 0 3036 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1676037725
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1676037725
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1676037725
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_95
timestamp 1676037725
transform 1 0 9844 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_103
timestamp 1676037725
transform 1 0 10580 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_107
timestamp 1676037725
transform 1 0 10948 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_112
timestamp 1676037725
transform 1 0 11408 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_125
timestamp 1676037725
transform 1 0 12604 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1676037725
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_143
timestamp 1676037725
transform 1 0 14260 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_154
timestamp 1676037725
transform 1 0 15272 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_158
timestamp 1676037725
transform 1 0 15640 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_162
timestamp 1676037725
transform 1 0 16008 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_175
timestamp 1676037725
transform 1 0 17204 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_182
timestamp 1676037725
transform 1 0 17848 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1676037725
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_209
timestamp 1676037725
transform 1 0 20332 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_215
timestamp 1676037725
transform 1 0 20884 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_238
timestamp 1676037725
transform 1 0 23000 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_242
timestamp 1676037725
transform 1 0 23368 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_245
timestamp 1676037725
transform 1 0 23644 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1676037725
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_257
timestamp 1676037725
transform 1 0 24748 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_262
timestamp 1676037725
transform 1 0 25208 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_286
timestamp 1676037725
transform 1 0 27416 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_299
timestamp 1676037725
transform 1 0 28612 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_306
timestamp 1676037725
transform 1 0 29256 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_309
timestamp 1676037725
transform 1 0 29532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_320
timestamp 1676037725
transform 1 0 30544 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_333
timestamp 1676037725
transform 1 0 31740 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_346
timestamp 1676037725
transform 1 0 32936 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_359
timestamp 1676037725
transform 1 0 34132 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_365
timestamp 1676037725
transform 1 0 34684 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_387
timestamp 1676037725
transform 1 0 36708 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_411
timestamp 1676037725
transform 1 0 38916 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_418
timestamp 1676037725
transform 1 0 39560 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_425
timestamp 1676037725
transform 1 0 40204 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_437
timestamp 1676037725
transform 1 0 41308 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_449
timestamp 1676037725
transform 1 0 42412 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_461
timestamp 1676037725
transform 1 0 43516 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_473
timestamp 1676037725
transform 1 0 44620 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1676037725
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1676037725
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1676037725
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_513
timestamp 1676037725
transform 1 0 48300 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_519
timestamp 1676037725
transform 1 0 48852 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_525
timestamp 1676037725
transform 1 0 49404 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_21
timestamp 1676037725
transform 1 0 3036 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_33
timestamp 1676037725
transform 1 0 4140 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_45
timestamp 1676037725
transform 1 0 5244 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_53
timestamp 1676037725
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_81
timestamp 1676037725
transform 1 0 8556 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_89
timestamp 1676037725
transform 1 0 9292 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_99
timestamp 1676037725
transform 1 0 10212 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_104
timestamp 1676037725
transform 1 0 10672 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1676037725
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_115
timestamp 1676037725
transform 1 0 11684 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_126
timestamp 1676037725
transform 1 0 12696 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_130
timestamp 1676037725
transform 1 0 13064 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_153
timestamp 1676037725
transform 1 0 15180 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1676037725
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_180
timestamp 1676037725
transform 1 0 17664 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_185
timestamp 1676037725
transform 1 0 18124 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_196
timestamp 1676037725
transform 1 0 19136 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_209
timestamp 1676037725
transform 1 0 20332 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1676037725
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_229
timestamp 1676037725
transform 1 0 22172 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_246
timestamp 1676037725
transform 1 0 23736 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_259
timestamp 1676037725
transform 1 0 24932 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_267
timestamp 1676037725
transform 1 0 25668 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1676037725
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_285
timestamp 1676037725
transform 1 0 27324 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_290
timestamp 1676037725
transform 1 0 27784 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_312
timestamp 1676037725
transform 1 0 29808 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_325
timestamp 1676037725
transform 1 0 31004 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_332
timestamp 1676037725
transform 1 0 31648 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_337
timestamp 1676037725
transform 1 0 32108 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_348
timestamp 1676037725
transform 1 0 33120 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_361
timestamp 1676037725
transform 1 0 34316 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_374
timestamp 1676037725
transform 1 0 35512 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_387
timestamp 1676037725
transform 1 0 36708 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1676037725
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_393
timestamp 1676037725
transform 1 0 37260 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_415
timestamp 1676037725
transform 1 0 39284 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_428
timestamp 1676037725
transform 1 0 40480 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_435
timestamp 1676037725
transform 1 0 41124 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1676037725
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1676037725
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1676037725
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1676037725
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1676037725
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1676037725
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1676037725
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1676037725
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_519
timestamp 1676037725
transform 1 0 48852 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_525
timestamp 1676037725
transform 1 0 49404 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_21
timestamp 1676037725
transform 1 0 3036 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_61
timestamp 1676037725
transform 1 0 6716 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_73
timestamp 1676037725
transform 1 0 7820 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_81
timestamp 1676037725
transform 1 0 8556 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_97
timestamp 1676037725
transform 1 0 10028 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_125
timestamp 1676037725
transform 1 0 12604 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1676037725
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_152
timestamp 1676037725
transform 1 0 15088 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_156
timestamp 1676037725
transform 1 0 15456 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_166
timestamp 1676037725
transform 1 0 16376 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_179
timestamp 1676037725
transform 1 0 17572 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_183
timestamp 1676037725
transform 1 0 17940 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_187
timestamp 1676037725
transform 1 0 18308 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_191
timestamp 1676037725
transform 1 0 18676 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_199
timestamp 1676037725
transform 1 0 19412 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_203
timestamp 1676037725
transform 1 0 19780 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_213
timestamp 1676037725
transform 1 0 20700 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_217
timestamp 1676037725
transform 1 0 21068 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_227
timestamp 1676037725
transform 1 0 21988 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_233
timestamp 1676037725
transform 1 0 22540 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_248
timestamp 1676037725
transform 1 0 23920 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_265
timestamp 1676037725
transform 1 0 25484 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_278
timestamp 1676037725
transform 1 0 26680 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_284
timestamp 1676037725
transform 1 0 27232 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_295
timestamp 1676037725
transform 1 0 28244 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_301
timestamp 1676037725
transform 1 0 28796 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_309
timestamp 1676037725
transform 1 0 29532 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_315
timestamp 1676037725
transform 1 0 30084 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_339
timestamp 1676037725
transform 1 0 32292 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_352
timestamp 1676037725
transform 1 0 33488 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_359
timestamp 1676037725
transform 1 0 34132 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1676037725
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_365
timestamp 1676037725
transform 1 0 34684 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_387
timestamp 1676037725
transform 1 0 36708 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_394
timestamp 1676037725
transform 1 0 37352 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_418
timestamp 1676037725
transform 1 0 39560 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_421
timestamp 1676037725
transform 1 0 39836 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_443
timestamp 1676037725
transform 1 0 41860 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_447
timestamp 1676037725
transform 1 0 42228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_459
timestamp 1676037725
transform 1 0 43332 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_471
timestamp 1676037725
transform 1 0 44436 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1676037725
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1676037725
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1676037725
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1676037725
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_513
timestamp 1676037725
transform 1 0 48300 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_517
timestamp 1676037725
transform 1 0 48668 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_520
timestamp 1676037725
transform 1 0 48944 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_525
timestamp 1676037725
transform 1 0 49404 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_21
timestamp 1676037725
transform 1 0 3036 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_33
timestamp 1676037725
transform 1 0 4140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_45
timestamp 1676037725
transform 1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1676037725
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_69
timestamp 1676037725
transform 1 0 7452 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_73
timestamp 1676037725
transform 1 0 7820 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_83
timestamp 1676037725
transform 1 0 8740 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_91
timestamp 1676037725
transform 1 0 9476 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_99
timestamp 1676037725
transform 1 0 10212 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_104
timestamp 1676037725
transform 1 0 10672 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1676037725
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_116
timestamp 1676037725
transform 1 0 11776 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_127
timestamp 1676037725
transform 1 0 12788 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_140
timestamp 1676037725
transform 1 0 13984 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_153
timestamp 1676037725
transform 1 0 15180 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1676037725
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_175
timestamp 1676037725
transform 1 0 17204 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_186
timestamp 1676037725
transform 1 0 18216 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_194
timestamp 1676037725
transform 1 0 18952 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_217
timestamp 1676037725
transform 1 0 21068 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_221
timestamp 1676037725
transform 1 0 21436 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_233
timestamp 1676037725
transform 1 0 22540 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_237
timestamp 1676037725
transform 1 0 22908 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_248
timestamp 1676037725
transform 1 0 23920 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_254
timestamp 1676037725
transform 1 0 24472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_275
timestamp 1676037725
transform 1 0 26404 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1676037725
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1676037725
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_292
timestamp 1676037725
transform 1 0 27968 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_316
timestamp 1676037725
transform 1 0 30176 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_329
timestamp 1676037725
transform 1 0 31372 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1676037725
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_337
timestamp 1676037725
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_348
timestamp 1676037725
transform 1 0 33120 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_361
timestamp 1676037725
transform 1 0 34316 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_367
timestamp 1676037725
transform 1 0 34868 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_390
timestamp 1676037725
transform 1 0 36984 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_393
timestamp 1676037725
transform 1 0 37260 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_398
timestamp 1676037725
transform 1 0 37720 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_402
timestamp 1676037725
transform 1 0 38088 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_423
timestamp 1676037725
transform 1 0 40020 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_427
timestamp 1676037725
transform 1 0 40388 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_437
timestamp 1676037725
transform 1 0 41308 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1676037725
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1676037725
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1676037725
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1676037725
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1676037725
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1676037725
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1676037725
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1676037725
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1676037725
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_519
timestamp 1676037725
transform 1 0 48852 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_525
timestamp 1676037725
transform 1 0 49404 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_21
timestamp 1676037725
transform 1 0 3036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1676037725
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1676037725
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1676037725
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_65
timestamp 1676037725
transform 1 0 7084 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_71
timestamp 1676037725
transform 1 0 7636 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_81
timestamp 1676037725
transform 1 0 8556 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_93
timestamp 1676037725
transform 1 0 9660 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_98
timestamp 1676037725
transform 1 0 10120 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_104
timestamp 1676037725
transform 1 0 10672 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_117
timestamp 1676037725
transform 1 0 11868 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_121
timestamp 1676037725
transform 1 0 12236 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_125
timestamp 1676037725
transform 1 0 12604 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1676037725
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_143
timestamp 1676037725
transform 1 0 14260 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_154
timestamp 1676037725
transform 1 0 15272 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_167
timestamp 1676037725
transform 1 0 16468 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_171
timestamp 1676037725
transform 1 0 16836 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1676037725
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_202
timestamp 1676037725
transform 1 0 19688 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_209
timestamp 1676037725
transform 1 0 20332 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_213
timestamp 1676037725
transform 1 0 20700 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_236
timestamp 1676037725
transform 1 0 22816 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_240
timestamp 1676037725
transform 1 0 23184 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1676037725
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_258
timestamp 1676037725
transform 1 0 24840 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_286
timestamp 1676037725
transform 1 0 27416 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_290
timestamp 1676037725
transform 1 0 27784 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_300
timestamp 1676037725
transform 1 0 28704 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1676037725
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_320
timestamp 1676037725
transform 1 0 30544 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_333
timestamp 1676037725
transform 1 0 31740 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_337
timestamp 1676037725
transform 1 0 32108 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_358
timestamp 1676037725
transform 1 0 34040 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_365
timestamp 1676037725
transform 1 0 34684 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_378
timestamp 1676037725
transform 1 0 35880 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_391
timestamp 1676037725
transform 1 0 37076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_395
timestamp 1676037725
transform 1 0 37444 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_418
timestamp 1676037725
transform 1 0 39560 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_421
timestamp 1676037725
transform 1 0 39836 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_432
timestamp 1676037725
transform 1 0 40848 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_440
timestamp 1676037725
transform 1 0 41584 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_452
timestamp 1676037725
transform 1 0 42688 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_464
timestamp 1676037725
transform 1 0 43792 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1676037725
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1676037725
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1676037725
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_513
timestamp 1676037725
transform 1 0 48300 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_519
timestamp 1676037725
transform 1 0 48852 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_525
timestamp 1676037725
transform 1 0 49404 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_21
timestamp 1676037725
transform 1 0 3036 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_33
timestamp 1676037725
transform 1 0 4140 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_45
timestamp 1676037725
transform 1 0 5244 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_53
timestamp 1676037725
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1676037725
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1676037725
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_93
timestamp 1676037725
transform 1 0 9660 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_99
timestamp 1676037725
transform 1 0 10212 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1676037725
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_119
timestamp 1676037725
transform 1 0 12052 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_124
timestamp 1676037725
transform 1 0 12512 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_135
timestamp 1676037725
transform 1 0 13524 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_139
timestamp 1676037725
transform 1 0 13892 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_145
timestamp 1676037725
transform 1 0 14444 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_149
timestamp 1676037725
transform 1 0 14812 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_153
timestamp 1676037725
transform 1 0 15180 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1676037725
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_175
timestamp 1676037725
transform 1 0 17204 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_179
timestamp 1676037725
transform 1 0 17572 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_192
timestamp 1676037725
transform 1 0 18768 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_216
timestamp 1676037725
transform 1 0 20976 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_220
timestamp 1676037725
transform 1 0 21344 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_230
timestamp 1676037725
transform 1 0 22264 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_254
timestamp 1676037725
transform 1 0 24472 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_267
timestamp 1676037725
transform 1 0 25668 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_271
timestamp 1676037725
transform 1 0 26036 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1676037725
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_281
timestamp 1676037725
transform 1 0 26956 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_294
timestamp 1676037725
transform 1 0 28152 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_298
timestamp 1676037725
transform 1 0 28520 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_308
timestamp 1676037725
transform 1 0 29440 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_321
timestamp 1676037725
transform 1 0 30636 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_334
timestamp 1676037725
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_337
timestamp 1676037725
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_360
timestamp 1676037725
transform 1 0 34224 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_375
timestamp 1676037725
transform 1 0 35604 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_388
timestamp 1676037725
transform 1 0 36800 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_393
timestamp 1676037725
transform 1 0 37260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_404
timestamp 1676037725
transform 1 0 38272 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_408
timestamp 1676037725
transform 1 0 38640 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_431
timestamp 1676037725
transform 1 0 40756 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_435
timestamp 1676037725
transform 1 0 41124 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1676037725
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1676037725
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1676037725
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1676037725
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1676037725
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1676037725
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1676037725
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_505
timestamp 1676037725
transform 1 0 47564 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_513
timestamp 1676037725
transform 1 0 48300 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_517
timestamp 1676037725
transform 1 0 48668 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_525
timestamp 1676037725
transform 1 0 49404 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_21
timestamp 1676037725
transform 1 0 3036 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1676037725
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1676037725
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1676037725
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1676037725
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1676037725
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1676037725
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_97
timestamp 1676037725
transform 1 0 10028 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_123
timestamp 1676037725
transform 1 0 12420 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_127
timestamp 1676037725
transform 1 0 12788 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_131
timestamp 1676037725
transform 1 0 13156 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1676037725
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_163
timestamp 1676037725
transform 1 0 16100 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_168
timestamp 1676037725
transform 1 0 16560 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_179
timestamp 1676037725
transform 1 0 17572 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1676037725
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_202
timestamp 1676037725
transform 1 0 19688 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_228
timestamp 1676037725
transform 1 0 22080 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_232
timestamp 1676037725
transform 1 0 22448 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_237
timestamp 1676037725
transform 1 0 22908 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1676037725
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_264
timestamp 1676037725
transform 1 0 25392 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_271
timestamp 1676037725
transform 1 0 26036 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_277
timestamp 1676037725
transform 1 0 26588 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_281
timestamp 1676037725
transform 1 0 26956 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_302
timestamp 1676037725
transform 1 0 28888 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_311
timestamp 1676037725
transform 1 0 29716 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_324
timestamp 1676037725
transform 1 0 30912 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_337
timestamp 1676037725
transform 1 0 32108 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_341
timestamp 1676037725
transform 1 0 32476 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_353
timestamp 1676037725
transform 1 0 33580 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_357
timestamp 1676037725
transform 1 0 33948 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_365
timestamp 1676037725
transform 1 0 34684 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_370
timestamp 1676037725
transform 1 0 35144 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_375
timestamp 1676037725
transform 1 0 35604 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_397
timestamp 1676037725
transform 1 0 37628 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_410
timestamp 1676037725
transform 1 0 38824 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_418
timestamp 1676037725
transform 1 0 39560 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_421
timestamp 1676037725
transform 1 0 39836 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_427
timestamp 1676037725
transform 1 0 40388 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_437
timestamp 1676037725
transform 1 0 41308 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_449
timestamp 1676037725
transform 1 0 42412 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_461
timestamp 1676037725
transform 1 0 43516 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_473
timestamp 1676037725
transform 1 0 44620 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1676037725
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1676037725
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1676037725
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_513
timestamp 1676037725
transform 1 0 48300 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_519
timestamp 1676037725
transform 1 0 48852 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_525
timestamp 1676037725
transform 1 0 49404 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_21
timestamp 1676037725
transform 1 0 3036 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_28
timestamp 1676037725
transform 1 0 3680 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_32
timestamp 1676037725
transform 1 0 4048 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_43
timestamp 1676037725
transform 1 0 5060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1676037725
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_69
timestamp 1676037725
transform 1 0 7452 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_75
timestamp 1676037725
transform 1 0 8004 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_87
timestamp 1676037725
transform 1 0 9108 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_93
timestamp 1676037725
transform 1 0 9660 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_97
timestamp 1676037725
transform 1 0 10028 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1676037725
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_135
timestamp 1676037725
transform 1 0 13524 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_148
timestamp 1676037725
transform 1 0 14720 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_154
timestamp 1676037725
transform 1 0 15272 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_159
timestamp 1676037725
transform 1 0 15732 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1676037725
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_171
timestamp 1676037725
transform 1 0 16836 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_179
timestamp 1676037725
transform 1 0 17572 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_192
timestamp 1676037725
transform 1 0 18768 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_196
timestamp 1676037725
transform 1 0 19136 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_200
timestamp 1676037725
transform 1 0 19504 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1676037725
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_237
timestamp 1676037725
transform 1 0 22908 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_252
timestamp 1676037725
transform 1 0 24288 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_265
timestamp 1676037725
transform 1 0 25484 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1676037725
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1676037725
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_292
timestamp 1676037725
transform 1 0 27968 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_305
timestamp 1676037725
transform 1 0 29164 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_313
timestamp 1676037725
transform 1 0 29900 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_324
timestamp 1676037725
transform 1 0 30912 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_331
timestamp 1676037725
transform 1 0 31556 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1676037725
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_337
timestamp 1676037725
transform 1 0 32108 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_348
timestamp 1676037725
transform 1 0 33120 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_352
timestamp 1676037725
transform 1 0 33488 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_373
timestamp 1676037725
transform 1 0 35420 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_377
timestamp 1676037725
transform 1 0 35788 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_387
timestamp 1676037725
transform 1 0 36708 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1676037725
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_393
timestamp 1676037725
transform 1 0 37260 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_399
timestamp 1676037725
transform 1 0 37812 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_421
timestamp 1676037725
transform 1 0 39836 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_425
timestamp 1676037725
transform 1 0 40204 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_436
timestamp 1676037725
transform 1 0 41216 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1676037725
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1676037725
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1676037725
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1676037725
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1676037725
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1676037725
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_505
timestamp 1676037725
transform 1 0 47564 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_513
timestamp 1676037725
transform 1 0 48300 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_519
timestamp 1676037725
transform 1 0 48852 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_525
timestamp 1676037725
transform 1 0 49404 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_21
timestamp 1676037725
transform 1 0 3036 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1676037725
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_47
timestamp 1676037725
transform 1 0 5428 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_59
timestamp 1676037725
transform 1 0 6532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_71
timestamp 1676037725
transform 1 0 7636 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_75
timestamp 1676037725
transform 1 0 8004 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_80
timestamp 1676037725
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_108
timestamp 1676037725
transform 1 0 11040 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_112
timestamp 1676037725
transform 1 0 11408 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_115
timestamp 1676037725
transform 1 0 11684 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_120
timestamp 1676037725
transform 1 0 12144 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_133
timestamp 1676037725
transform 1 0 13340 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_137
timestamp 1676037725
transform 1 0 13708 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_163
timestamp 1676037725
transform 1 0 16100 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_167
timestamp 1676037725
transform 1 0 16468 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_170
timestamp 1676037725
transform 1 0 16744 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_181
timestamp 1676037725
transform 1 0 17756 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1676037725
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_199
timestamp 1676037725
transform 1 0 19412 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_203
timestamp 1676037725
transform 1 0 19780 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_213
timestamp 1676037725
transform 1 0 20700 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_226
timestamp 1676037725
transform 1 0 21896 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1676037725
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_264
timestamp 1676037725
transform 1 0 25392 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_288
timestamp 1676037725
transform 1 0 27600 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_298
timestamp 1676037725
transform 1 0 28520 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_302
timestamp 1676037725
transform 1 0 28888 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_306
timestamp 1676037725
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_309
timestamp 1676037725
transform 1 0 29532 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_320
timestamp 1676037725
transform 1 0 30544 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_324
timestamp 1676037725
transform 1 0 30912 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_339
timestamp 1676037725
transform 1 0 32292 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_352
timestamp 1676037725
transform 1 0 33488 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_365
timestamp 1676037725
transform 1 0 34684 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_371
timestamp 1676037725
transform 1 0 35236 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_395
timestamp 1676037725
transform 1 0 37444 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_399
timestamp 1676037725
transform 1 0 37812 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_410
timestamp 1676037725
transform 1 0 38824 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_418
timestamp 1676037725
transform 1 0 39560 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_421
timestamp 1676037725
transform 1 0 39836 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_443
timestamp 1676037725
transform 1 0 41860 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_447
timestamp 1676037725
transform 1 0 42228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_459
timestamp 1676037725
transform 1 0 43332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_471
timestamp 1676037725
transform 1 0 44436 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1676037725
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1676037725
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1676037725
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1676037725
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_513
timestamp 1676037725
transform 1 0 48300 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_517
timestamp 1676037725
transform 1 0 48668 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_525
timestamp 1676037725
transform 1 0 49404 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_21
timestamp 1676037725
transform 1 0 3036 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_41
timestamp 1676037725
transform 1 0 4876 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_49
timestamp 1676037725
transform 1 0 5612 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1676037725
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1676037725
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1676037725
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_96
timestamp 1676037725
transform 1 0 9936 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_103
timestamp 1676037725
transform 1 0 10580 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1676037725
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_116
timestamp 1676037725
transform 1 0 11776 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_122
timestamp 1676037725
transform 1 0 12328 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_146
timestamp 1676037725
transform 1 0 14536 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_152
timestamp 1676037725
transform 1 0 15088 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_158
timestamp 1676037725
transform 1 0 15640 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1676037725
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_180
timestamp 1676037725
transform 1 0 17664 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_207
timestamp 1676037725
transform 1 0 20148 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_211
timestamp 1676037725
transform 1 0 20516 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1676037725
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_238
timestamp 1676037725
transform 1 0 23000 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_242
timestamp 1676037725
transform 1 0 23368 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_263
timestamp 1676037725
transform 1 0 25300 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_267
timestamp 1676037725
transform 1 0 25668 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_277
timestamp 1676037725
transform 1 0 26588 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_281
timestamp 1676037725
transform 1 0 26956 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_293
timestamp 1676037725
transform 1 0 28060 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_306
timestamp 1676037725
transform 1 0 29256 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_310
timestamp 1676037725
transform 1 0 29624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_314
timestamp 1676037725
transform 1 0 29992 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_320
timestamp 1676037725
transform 1 0 30544 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_333
timestamp 1676037725
transform 1 0 31740 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_337
timestamp 1676037725
transform 1 0 32108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_348
timestamp 1676037725
transform 1 0 33120 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_361
timestamp 1676037725
transform 1 0 34316 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_374
timestamp 1676037725
transform 1 0 35512 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_387
timestamp 1676037725
transform 1 0 36708 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1676037725
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_395
timestamp 1676037725
transform 1 0 37444 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_399
timestamp 1676037725
transform 1 0 37812 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_420
timestamp 1676037725
transform 1 0 39744 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_433
timestamp 1676037725
transform 1 0 40940 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_439
timestamp 1676037725
transform 1 0 41492 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1676037725
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1676037725
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1676037725
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1676037725
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1676037725
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1676037725
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1676037725
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_505
timestamp 1676037725
transform 1 0 47564 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_513
timestamp 1676037725
transform 1 0 48300 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_519
timestamp 1676037725
transform 1 0 48852 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_525
timestamp 1676037725
transform 1 0 49404 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_21
timestamp 1676037725
transform 1 0 3036 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1676037725
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_47
timestamp 1676037725
transform 1 0 5428 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_67
timestamp 1676037725
transform 1 0 7268 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_71
timestamp 1676037725
transform 1 0 7636 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_75
timestamp 1676037725
transform 1 0 8004 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1676037725
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_93
timestamp 1676037725
transform 1 0 9660 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_99
timestamp 1676037725
transform 1 0 10212 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_106
timestamp 1676037725
transform 1 0 10856 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_114
timestamp 1676037725
transform 1 0 11592 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1676037725
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_146
timestamp 1676037725
transform 1 0 14536 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_154
timestamp 1676037725
transform 1 0 15272 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_167
timestamp 1676037725
transform 1 0 16468 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_180
timestamp 1676037725
transform 1 0 17664 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_184
timestamp 1676037725
transform 1 0 18032 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1676037725
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_199
timestamp 1676037725
transform 1 0 19412 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_205
timestamp 1676037725
transform 1 0 19964 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_209
timestamp 1676037725
transform 1 0 20332 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_231
timestamp 1676037725
transform 1 0 22356 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_239
timestamp 1676037725
transform 1 0 23092 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1676037725
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_258
timestamp 1676037725
transform 1 0 24840 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_264
timestamp 1676037725
transform 1 0 25392 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_275
timestamp 1676037725
transform 1 0 26404 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_288
timestamp 1676037725
transform 1 0 27600 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_301
timestamp 1676037725
transform 1 0 28796 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1676037725
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1676037725
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_320
timestamp 1676037725
transform 1 0 30544 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_333
timestamp 1676037725
transform 1 0 31740 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_346
timestamp 1676037725
transform 1 0 32936 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_350
timestamp 1676037725
transform 1 0 33304 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_360
timestamp 1676037725
transform 1 0 34224 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_365
timestamp 1676037725
transform 1 0 34684 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_376
timestamp 1676037725
transform 1 0 35696 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_389
timestamp 1676037725
transform 1 0 36892 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_397
timestamp 1676037725
transform 1 0 37628 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_408
timestamp 1676037725
transform 1 0 38640 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_414
timestamp 1676037725
transform 1 0 39192 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_421
timestamp 1676037725
transform 1 0 39836 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_432
timestamp 1676037725
transform 1 0 40848 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_438
timestamp 1676037725
transform 1 0 41400 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_450
timestamp 1676037725
transform 1 0 42504 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_462
timestamp 1676037725
transform 1 0 43608 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_474
timestamp 1676037725
transform 1 0 44712 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1676037725
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1676037725
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1676037725
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_513
timestamp 1676037725
transform 1 0 48300 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_519
timestamp 1676037725
transform 1 0 48852 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_525
timestamp 1676037725
transform 1 0 49404 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_21
timestamp 1676037725
transform 1 0 3036 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_41
timestamp 1676037725
transform 1 0 4876 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_48
timestamp 1676037725
transform 1 0 5520 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_75
timestamp 1676037725
transform 1 0 8004 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_83
timestamp 1676037725
transform 1 0 8740 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_89
timestamp 1676037725
transform 1 0 9292 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_96
timestamp 1676037725
transform 1 0 9936 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_103
timestamp 1676037725
transform 1 0 10580 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1676037725
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_119
timestamp 1676037725
transform 1 0 12052 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_127
timestamp 1676037725
transform 1 0 12788 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_135
timestamp 1676037725
transform 1 0 13524 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_146
timestamp 1676037725
transform 1 0 14536 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_153
timestamp 1676037725
transform 1 0 15180 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1676037725
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_171
timestamp 1676037725
transform 1 0 16836 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_193
timestamp 1676037725
transform 1 0 18860 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_197
timestamp 1676037725
transform 1 0 19228 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_201
timestamp 1676037725
transform 1 0 19596 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1676037725
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_236
timestamp 1676037725
transform 1 0 22816 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_243
timestamp 1676037725
transform 1 0 23460 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_267
timestamp 1676037725
transform 1 0 25668 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_274
timestamp 1676037725
transform 1 0 26312 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1676037725
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_281
timestamp 1676037725
transform 1 0 26956 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_304
timestamp 1676037725
transform 1 0 29072 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_317
timestamp 1676037725
transform 1 0 30268 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_330
timestamp 1676037725
transform 1 0 31464 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1676037725
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_337
timestamp 1676037725
transform 1 0 32108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_359
timestamp 1676037725
transform 1 0 34132 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_372
timestamp 1676037725
transform 1 0 35328 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_378
timestamp 1676037725
transform 1 0 35880 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_389
timestamp 1676037725
transform 1 0 36892 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_393
timestamp 1676037725
transform 1 0 37260 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_397
timestamp 1676037725
transform 1 0 37628 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_418
timestamp 1676037725
transform 1 0 39560 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_431
timestamp 1676037725
transform 1 0 40756 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_438
timestamp 1676037725
transform 1 0 41400 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_442
timestamp 1676037725
transform 1 0 41768 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1676037725
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1676037725
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1676037725
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1676037725
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1676037725
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1676037725
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_505
timestamp 1676037725
transform 1 0 47564 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_513
timestamp 1676037725
transform 1 0 48300 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_517
timestamp 1676037725
transform 1 0 48668 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_525
timestamp 1676037725
transform 1 0 49404 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_21
timestamp 1676037725
transform 1 0 3036 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1676037725
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_47
timestamp 1676037725
transform 1 0 5428 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_67
timestamp 1676037725
transform 1 0 7268 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_76
timestamp 1676037725
transform 1 0 8096 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_91
timestamp 1676037725
transform 1 0 9476 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_98
timestamp 1676037725
transform 1 0 10120 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_105
timestamp 1676037725
transform 1 0 10764 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_112
timestamp 1676037725
transform 1 0 11408 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_120
timestamp 1676037725
transform 1 0 12144 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_124
timestamp 1676037725
transform 1 0 12512 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_130
timestamp 1676037725
transform 1 0 13064 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_134
timestamp 1676037725
transform 1 0 13432 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1676037725
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_163
timestamp 1676037725
transform 1 0 16100 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_170
timestamp 1676037725
transform 1 0 16744 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1676037725
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_199
timestamp 1676037725
transform 1 0 19412 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_214
timestamp 1676037725
transform 1 0 20792 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_238
timestamp 1676037725
transform 1 0 23000 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_246
timestamp 1676037725
transform 1 0 23736 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_258
timestamp 1676037725
transform 1 0 24840 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_262
timestamp 1676037725
transform 1 0 25208 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_265
timestamp 1676037725
transform 1 0 25484 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_276
timestamp 1676037725
transform 1 0 26496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_280
timestamp 1676037725
transform 1 0 26864 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_288
timestamp 1676037725
transform 1 0 27600 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_292
timestamp 1676037725
transform 1 0 27968 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_305
timestamp 1676037725
transform 1 0 29164 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1676037725
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_314
timestamp 1676037725
transform 1 0 29992 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_318
timestamp 1676037725
transform 1 0 30360 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_322
timestamp 1676037725
transform 1 0 30728 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_332
timestamp 1676037725
transform 1 0 31648 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_340
timestamp 1676037725
transform 1 0 32384 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_362
timestamp 1676037725
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_365
timestamp 1676037725
transform 1 0 34684 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_387
timestamp 1676037725
transform 1 0 36708 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_391
timestamp 1676037725
transform 1 0 37076 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_34_417
timestamp 1676037725
transform 1 0 39468 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_421
timestamp 1676037725
transform 1 0 39836 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_432
timestamp 1676037725
transform 1 0 40848 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_445
timestamp 1676037725
transform 1 0 42044 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_449
timestamp 1676037725
transform 1 0 42412 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_461
timestamp 1676037725
transform 1 0 43516 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_473
timestamp 1676037725
transform 1 0 44620 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1676037725
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1676037725
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1676037725
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_513
timestamp 1676037725
transform 1 0 48300 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_519
timestamp 1676037725
transform 1 0 48852 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_525
timestamp 1676037725
transform 1 0 49404 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_21
timestamp 1676037725
transform 1 0 3036 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_41
timestamp 1676037725
transform 1 0 4876 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_49
timestamp 1676037725
transform 1 0 5612 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_53
timestamp 1676037725
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_75
timestamp 1676037725
transform 1 0 8004 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_95
timestamp 1676037725
transform 1 0 9844 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_101
timestamp 1676037725
transform 1 0 10396 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1676037725
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1676037725
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_118
timestamp 1676037725
transform 1 0 11960 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_124
timestamp 1676037725
transform 1 0 12512 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_128
timestamp 1676037725
transform 1 0 12880 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_134
timestamp 1676037725
transform 1 0 13432 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_138
timestamp 1676037725
transform 1 0 13800 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_142
timestamp 1676037725
transform 1 0 14168 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1676037725
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_175
timestamp 1676037725
transform 1 0 17204 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_186
timestamp 1676037725
transform 1 0 18216 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_210
timestamp 1676037725
transform 1 0 20424 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_214
timestamp 1676037725
transform 1 0 20792 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1676037725
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_227
timestamp 1676037725
transform 1 0 21988 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_230
timestamp 1676037725
transform 1 0 22264 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_253
timestamp 1676037725
transform 1 0 24380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_266
timestamp 1676037725
transform 1 0 25576 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_272
timestamp 1676037725
transform 1 0 26128 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1676037725
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_281
timestamp 1676037725
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_292
timestamp 1676037725
transform 1 0 27968 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_305
timestamp 1676037725
transform 1 0 29164 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_318
timestamp 1676037725
transform 1 0 30360 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_331
timestamp 1676037725
transform 1 0 31556 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1676037725
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_337
timestamp 1676037725
transform 1 0 32108 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_341
timestamp 1676037725
transform 1 0 32476 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_345
timestamp 1676037725
transform 1 0 32844 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_358
timestamp 1676037725
transform 1 0 34040 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_371
timestamp 1676037725
transform 1 0 35236 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_375
timestamp 1676037725
transform 1 0 35604 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_385
timestamp 1676037725
transform 1 0 36524 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_389
timestamp 1676037725
transform 1 0 36892 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_393
timestamp 1676037725
transform 1 0 37260 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_421
timestamp 1676037725
transform 1 0 39836 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_434
timestamp 1676037725
transform 1 0 41032 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_441
timestamp 1676037725
transform 1 0 41676 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1676037725
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_453
timestamp 1676037725
transform 1 0 42780 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_465
timestamp 1676037725
transform 1 0 43884 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_477
timestamp 1676037725
transform 1 0 44988 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_489
timestamp 1676037725
transform 1 0 46092 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_501
timestamp 1676037725
transform 1 0 47196 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_505
timestamp 1676037725
transform 1 0 47564 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_512
timestamp 1676037725
transform 1 0 48208 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_519
timestamp 1676037725
transform 1 0 48852 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_525
timestamp 1676037725
transform 1 0 49404 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_21
timestamp 1676037725
transform 1 0 3036 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1676037725
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_47
timestamp 1676037725
transform 1 0 5428 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_67
timestamp 1676037725
transform 1 0 7268 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_75
timestamp 1676037725
transform 1 0 8004 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1676037725
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_85
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_103
timestamp 1676037725
transform 1 0 10580 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_107
timestamp 1676037725
transform 1 0 10948 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_118
timestamp 1676037725
transform 1 0 11960 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_125
timestamp 1676037725
transform 1 0 12604 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1676037725
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_149
timestamp 1676037725
transform 1 0 14812 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_173
timestamp 1676037725
transform 1 0 17020 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_193
timestamp 1676037725
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_215
timestamp 1676037725
transform 1 0 20884 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_219
timestamp 1676037725
transform 1 0 21252 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_230
timestamp 1676037725
transform 1 0 22264 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_243
timestamp 1676037725
transform 1 0 23460 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1676037725
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_264
timestamp 1676037725
transform 1 0 25392 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_268
timestamp 1676037725
transform 1 0 25760 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_279
timestamp 1676037725
transform 1 0 26772 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_292
timestamp 1676037725
transform 1 0 27968 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_305
timestamp 1676037725
transform 1 0 29164 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_309
timestamp 1676037725
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_314
timestamp 1676037725
transform 1 0 29992 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_318
timestamp 1676037725
transform 1 0 30360 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_322
timestamp 1676037725
transform 1 0 30728 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_343
timestamp 1676037725
transform 1 0 32660 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_356
timestamp 1676037725
transform 1 0 33856 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_360
timestamp 1676037725
transform 1 0 34224 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_365
timestamp 1676037725
transform 1 0 34684 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_376
timestamp 1676037725
transform 1 0 35696 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_389
timestamp 1676037725
transform 1 0 36892 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_414
timestamp 1676037725
transform 1 0 39192 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1676037725
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_421
timestamp 1676037725
transform 1 0 39836 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_432
timestamp 1676037725
transform 1 0 40848 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_445
timestamp 1676037725
transform 1 0 42044 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_455
timestamp 1676037725
transform 1 0 42964 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_460
timestamp 1676037725
transform 1 0 43424 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_465
timestamp 1676037725
transform 1 0 43884 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_473
timestamp 1676037725
transform 1 0 44620 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1676037725
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1676037725
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_501
timestamp 1676037725
transform 1 0 47196 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_505
timestamp 1676037725
transform 1 0 47564 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_510
timestamp 1676037725
transform 1 0 48024 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_517
timestamp 1676037725
transform 1 0 48668 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_525
timestamp 1676037725
transform 1 0 49404 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_21
timestamp 1676037725
transform 1 0 3036 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_29
timestamp 1676037725
transform 1 0 3772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_34
timestamp 1676037725
transform 1 0 4232 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1676037725
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_37_63
timestamp 1676037725
transform 1 0 6900 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_37_85
timestamp 1676037725
transform 1 0 8924 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_93
timestamp 1676037725
transform 1 0 9660 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1676037725
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_119
timestamp 1676037725
transform 1 0 12052 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_123
timestamp 1676037725
transform 1 0 12420 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_141
timestamp 1676037725
transform 1 0 14076 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_145
timestamp 1676037725
transform 1 0 14444 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_149
timestamp 1676037725
transform 1 0 14812 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1676037725
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_191
timestamp 1676037725
transform 1 0 18676 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_195
timestamp 1676037725
transform 1 0 19044 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_220
timestamp 1676037725
transform 1 0 21344 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_248
timestamp 1676037725
transform 1 0 23920 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_252
timestamp 1676037725
transform 1 0 24288 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_255
timestamp 1676037725
transform 1 0 24564 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1676037725
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_281
timestamp 1676037725
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_286
timestamp 1676037725
transform 1 0 27416 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_290
timestamp 1676037725
transform 1 0 27784 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_313
timestamp 1676037725
transform 1 0 29900 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_326
timestamp 1676037725
transform 1 0 31096 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_333
timestamp 1676037725
transform 1 0 31740 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_337
timestamp 1676037725
transform 1 0 32108 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_348
timestamp 1676037725
transform 1 0 33120 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_352
timestamp 1676037725
transform 1 0 33488 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_374
timestamp 1676037725
transform 1 0 35512 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_378
timestamp 1676037725
transform 1 0 35880 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_389
timestamp 1676037725
transform 1 0 36892 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_393
timestamp 1676037725
transform 1 0 37260 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_415
timestamp 1676037725
transform 1 0 39284 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_428
timestamp 1676037725
transform 1 0 40480 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_435
timestamp 1676037725
transform 1 0 41124 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_442
timestamp 1676037725
transform 1 0 41768 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_449
timestamp 1676037725
transform 1 0 42412 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_454
timestamp 1676037725
transform 1 0 42872 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_461
timestamp 1676037725
transform 1 0 43516 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_468
timestamp 1676037725
transform 1 0 44160 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_475
timestamp 1676037725
transform 1 0 44804 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_479
timestamp 1676037725
transform 1 0 45172 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_491
timestamp 1676037725
transform 1 0 46276 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_497
timestamp 1676037725
transform 1 0 46828 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_502
timestamp 1676037725
transform 1 0 47288 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_511
timestamp 1676037725
transform 1 0 48116 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_517
timestamp 1676037725
transform 1 0 48668 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_525
timestamp 1676037725
transform 1 0 49404 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_21
timestamp 1676037725
transform 1 0 3036 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1676037725
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_35
timestamp 1676037725
transform 1 0 4324 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_42
timestamp 1676037725
transform 1 0 4968 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_62
timestamp 1676037725
transform 1 0 6808 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1676037725
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_91
timestamp 1676037725
transform 1 0 9476 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_98
timestamp 1676037725
transform 1 0 10120 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_118
timestamp 1676037725
transform 1 0 11960 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1676037725
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_143
timestamp 1676037725
transform 1 0 14260 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_150
timestamp 1676037725
transform 1 0 14904 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_170
timestamp 1676037725
transform 1 0 16744 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1676037725
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_199
timestamp 1676037725
transform 1 0 19412 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_205
timestamp 1676037725
transform 1 0 19964 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_229
timestamp 1676037725
transform 1 0 22172 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_237
timestamp 1676037725
transform 1 0 22908 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1676037725
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_259
timestamp 1676037725
transform 1 0 24932 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_263
timestamp 1676037725
transform 1 0 25300 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_287
timestamp 1676037725
transform 1 0 27508 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_300
timestamp 1676037725
transform 1 0 28704 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_306
timestamp 1676037725
transform 1 0 29256 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_309
timestamp 1676037725
transform 1 0 29532 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_320
timestamp 1676037725
transform 1 0 30544 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_324
timestamp 1676037725
transform 1 0 30912 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_327
timestamp 1676037725
transform 1 0 31188 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_350
timestamp 1676037725
transform 1 0 33304 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_357
timestamp 1676037725
transform 1 0 33948 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1676037725
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_367
timestamp 1676037725
transform 1 0 34868 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_389
timestamp 1676037725
transform 1 0 36892 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_413
timestamp 1676037725
transform 1 0 39100 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1676037725
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_421
timestamp 1676037725
transform 1 0 39836 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_432
timestamp 1676037725
transform 1 0 40848 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_436
timestamp 1676037725
transform 1 0 41216 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_462
timestamp 1676037725
transform 1 0 43608 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_466
timestamp 1676037725
transform 1 0 43976 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_472
timestamp 1676037725
transform 1 0 44528 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_483
timestamp 1676037725
transform 1 0 45540 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_494
timestamp 1676037725
transform 1 0 46552 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_497
timestamp 1676037725
transform 1 0 46828 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_502
timestamp 1676037725
transform 1 0 47288 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_509
timestamp 1676037725
transform 1 0 47932 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_517
timestamp 1676037725
transform 1 0 48668 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_525
timestamp 1676037725
transform 1 0 49404 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_14
timestamp 1676037725
transform 1 0 2392 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_34
timestamp 1676037725
transform 1 0 4232 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1676037725
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_57
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_63
timestamp 1676037725
transform 1 0 6900 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_70
timestamp 1676037725
transform 1 0 7544 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_90
timestamp 1676037725
transform 1 0 9384 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1676037725
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_113
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_126
timestamp 1676037725
transform 1 0 12696 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_146
timestamp 1676037725
transform 1 0 14536 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1676037725
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_188
timestamp 1676037725
transform 1 0 18400 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_212
timestamp 1676037725
transform 1 0 20608 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_216
timestamp 1676037725
transform 1 0 20976 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1676037725
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_237
timestamp 1676037725
transform 1 0 22908 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_250
timestamp 1676037725
transform 1 0 24104 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_256
timestamp 1676037725
transform 1 0 24656 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1676037725
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_281
timestamp 1676037725
transform 1 0 26956 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_286
timestamp 1676037725
transform 1 0 27416 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_293
timestamp 1676037725
transform 1 0 28060 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_300
timestamp 1676037725
transform 1 0 28704 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_307
timestamp 1676037725
transform 1 0 29348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_311
timestamp 1676037725
transform 1 0 29716 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_334
timestamp 1676037725
transform 1 0 31832 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_337
timestamp 1676037725
transform 1 0 32108 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_348
timestamp 1676037725
transform 1 0 33120 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_352
timestamp 1676037725
transform 1 0 33488 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_373
timestamp 1676037725
transform 1 0 35420 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_377
timestamp 1676037725
transform 1 0 35788 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_387
timestamp 1676037725
transform 1 0 36708 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1676037725
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_393
timestamp 1676037725
transform 1 0 37260 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_404
timestamp 1676037725
transform 1 0 38272 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_408
timestamp 1676037725
transform 1 0 38640 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_419
timestamp 1676037725
transform 1 0 39652 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_426
timestamp 1676037725
transform 1 0 40296 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_440
timestamp 1676037725
transform 1 0 41584 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_449
timestamp 1676037725
transform 1 0 42412 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_461
timestamp 1676037725
transform 1 0 43516 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_475
timestamp 1676037725
transform 1 0 44804 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_482
timestamp 1676037725
transform 1 0 45448 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_486
timestamp 1676037725
transform 1 0 45816 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_492
timestamp 1676037725
transform 1 0 46368 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_500
timestamp 1676037725
transform 1 0 47104 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_507
timestamp 1676037725
transform 1 0 47748 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_514
timestamp 1676037725
transform 1 0 48392 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_522
timestamp 1676037725
transform 1 0 49128 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_9
timestamp 1676037725
transform 1 0 1932 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1676037725
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_34
timestamp 1676037725
transform 1 0 4232 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_54
timestamp 1676037725
transform 1 0 6072 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_57
timestamp 1676037725
transform 1 0 6348 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_62
timestamp 1676037725
transform 1 0 6808 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1676037725
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_90
timestamp 1676037725
transform 1 0 9384 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_110
timestamp 1676037725
transform 1 0 11224 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_113
timestamp 1676037725
transform 1 0 11500 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_118
timestamp 1676037725
transform 1 0 11960 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1676037725
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_146
timestamp 1676037725
transform 1 0 14536 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_166
timestamp 1676037725
transform 1 0 16376 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_169
timestamp 1676037725
transform 1 0 16652 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_174
timestamp 1676037725
transform 1 0 17112 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1676037725
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_202
timestamp 1676037725
transform 1 0 19688 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_222
timestamp 1676037725
transform 1 0 21528 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_225
timestamp 1676037725
transform 1 0 21804 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_243
timestamp 1676037725
transform 1 0 23460 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1676037725
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_264
timestamp 1676037725
transform 1 0 25392 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_272
timestamp 1676037725
transform 1 0 26128 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_276
timestamp 1676037725
transform 1 0 26496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_281
timestamp 1676037725
transform 1 0 26956 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_287
timestamp 1676037725
transform 1 0 27508 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_294
timestamp 1676037725
transform 1 0 28152 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_301
timestamp 1676037725
transform 1 0 28796 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1676037725
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_309
timestamp 1676037725
transform 1 0 29532 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_314
timestamp 1676037725
transform 1 0 29992 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_321
timestamp 1676037725
transform 1 0 30636 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_328
timestamp 1676037725
transform 1 0 31280 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_337
timestamp 1676037725
transform 1 0 32108 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_342
timestamp 1676037725
transform 1 0 32568 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_349
timestamp 1676037725
transform 1 0 33212 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_362
timestamp 1676037725
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_365
timestamp 1676037725
transform 1 0 34684 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_376
timestamp 1676037725
transform 1 0 35696 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_389
timestamp 1676037725
transform 1 0 36892 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_393
timestamp 1676037725
transform 1 0 37260 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_404
timestamp 1676037725
transform 1 0 38272 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_418
timestamp 1676037725
transform 1 0 39560 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_421
timestamp 1676037725
transform 1 0 39836 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_426
timestamp 1676037725
transform 1 0 40296 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_440
timestamp 1676037725
transform 1 0 41584 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_449
timestamp 1676037725
transform 1 0 42412 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_471
timestamp 1676037725
transform 1 0 44436 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1676037725
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_477
timestamp 1676037725
transform 1 0 44988 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_483
timestamp 1676037725
transform 1 0 45540 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_491
timestamp 1676037725
transform 1 0 46276 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_499
timestamp 1676037725
transform 1 0 47012 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_503
timestamp 1676037725
transform 1 0 47380 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_505
timestamp 1676037725
transform 1 0 47564 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_511
timestamp 1676037725
transform 1 0 48116 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_525
timestamp 1676037725
transform 1 0 49404 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1676037725
transform 1 0 9660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1676037725
transform 1 0 47012 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1676037725
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input4 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1564 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input5
timestamp 1676037725
transform 1 0 1564 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1676037725
transform 1 0 2300 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1676037725
transform 1 0 1564 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input8
timestamp 1676037725
transform 1 0 1564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input9
timestamp 1676037725
transform 1 0 1564 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1676037725
transform 1 0 1564 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input11
timestamp 1676037725
transform 1 0 2300 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1676037725
transform 1 0 1564 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input13
timestamp 1676037725
transform 1 0 1564 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1676037725
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1676037725
transform 1 0 1564 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input16
timestamp 1676037725
transform 1 0 2300 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input17
timestamp 1676037725
transform 1 0 1564 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input18
timestamp 1676037725
transform 1 0 1564 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1676037725
transform 1 0 2300 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input20
timestamp 1676037725
transform 1 0 1564 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input21
timestamp 1676037725
transform 1 0 1564 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1676037725
transform 1 0 2852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1676037725
transform 1 0 1564 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1676037725
transform 1 0 3404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input25
timestamp 1676037725
transform 1 0 1564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input26
timestamp 1676037725
transform 1 0 1564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1676037725
transform 1 0 1564 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input28
timestamp 1676037725
transform 1 0 2300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1676037725
transform 1 0 1564 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input30
timestamp 1676037725
transform 1 0 1564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input31
timestamp 1676037725
transform 1 0 1564 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input32
timestamp 1676037725
transform 1 0 2300 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1676037725
transform 1 0 48392 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input34
timestamp 1676037725
transform 1 0 49036 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input35
timestamp 1676037725
transform 1 0 49036 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1676037725
transform 1 0 48392 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1676037725
transform 1 0 49036 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1676037725
transform 1 0 49036 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input39
timestamp 1676037725
transform 1 0 49036 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1676037725
transform 1 0 48392 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input41
timestamp 1676037725
transform 1 0 49036 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input42
timestamp 1676037725
transform 1 0 49036 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1676037725
transform 1 0 49036 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1676037725
transform 1 0 49036 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1676037725
transform 1 0 48392 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input46
timestamp 1676037725
transform 1 0 49036 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input47
timestamp 1676037725
transform 1 0 49036 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input48
timestamp 1676037725
transform 1 0 48300 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1676037725
transform 1 0 47656 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1676037725
transform 1 0 46092 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input51
timestamp 1676037725
transform 1 0 48300 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1676037725
transform 1 0 47748 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1676037725
transform 1 0 47012 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp 1676037725
transform 1 0 48484 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1676037725
transform 1 0 49036 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input56
timestamp 1676037725
transform 1 0 49036 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1676037725
transform 1 0 49128 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input58
timestamp 1676037725
transform 1 0 49036 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input59
timestamp 1676037725
transform 1 0 49036 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1676037725
transform 1 0 49036 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1676037725
transform 1 0 48392 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input62
timestamp 1676037725
transform 1 0 49036 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1676037725
transform 1 0 26036 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1676037725
transform 1 0 29072 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1676037725
transform 1 0 31004 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1676037725
transform 1 0 32292 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1676037725
transform 1 0 32936 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1676037725
transform 1 0 40020 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1676037725
transform 1 0 33672 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1676037725
transform 1 0 40020 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1676037725
transform 1 0 41400 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1676037725
transform 1 0 41492 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input73
timestamp 1676037725
transform 1 0 40664 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input74
timestamp 1676037725
transform 1 0 11040 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input75
timestamp 1676037725
transform 1 0 38640 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input76
timestamp 1676037725
transform 1 0 40664 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input77
timestamp 1676037725
transform 1 0 42596 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input78
timestamp 1676037725
transform 1 0 43884 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1676037725
transform 1 0 45172 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1676037725
transform 1 0 40848 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1676037725
transform 1 0 43884 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1676037725
transform 1 0 42596 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1676037725
transform 1 0 44528 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1676037725
transform 1 0 43240 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input85
timestamp 1676037725
transform 1 0 11776 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input86
timestamp 1676037725
transform 1 0 21988 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1676037725
transform 1 0 24564 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 1676037725
transform 1 0 30360 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 1676037725
transform 1 0 23828 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input90
timestamp 1676037725
transform 1 0 27876 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1676037725
transform 1 0 27784 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input92
timestamp 1676037725
transform 1 0 28520 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1676037725
transform 1 0 28980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1676037725
transform 1 0 30820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 1676037725
transform 1 0 32936 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 1676037725
transform 1 0 35052 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input97
timestamp 1676037725
transform 1 0 37444 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_16  input98
timestamp 1676037725
transform 1 0 42596 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input99
timestamp 1676037725
transform 1 0 43516 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input100
timestamp 1676037725
transform 1 0 45356 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input101
timestamp 1676037725
transform 1 0 47196 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input102
timestamp 1676037725
transform 1 0 46460 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input103
timestamp 1676037725
transform 1 0 45908 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input104
timestamp 1676037725
transform 1 0 46644 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input105
timestamp 1676037725
transform 1 0 46736 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input106
timestamp 1676037725
transform 1 0 47748 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input107
timestamp 1676037725
transform 1 0 48024 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input108
timestamp 1676037725
transform 1 0 48760 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input109
timestamp 1676037725
transform 1 0 44160 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input110
timestamp 1676037725
transform 1 0 45172 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  output111 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 40664 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output112
timestamp 1676037725
transform 1 0 3404 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output113
timestamp 1676037725
transform 1 0 1564 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1676037725
transform 1 0 1564 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1676037725
transform 1 0 1564 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1676037725
transform 1 0 1564 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1676037725
transform 1 0 1564 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1676037725
transform 1 0 1564 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1676037725
transform 1 0 1564 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1676037725
transform 1 0 3404 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1676037725
transform 1 0 1564 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1676037725
transform 1 0 1564 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1676037725
transform 1 0 1564 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1676037725
transform 1 0 1564 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1676037725
transform 1 0 3956 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1676037725
transform 1 0 3956 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1676037725
transform 1 0 5796 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1676037725
transform 1 0 5796 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1676037725
transform 1 0 6532 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1676037725
transform 1 0 3956 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1676037725
transform 1 0 5796 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output132
timestamp 1676037725
transform 1 0 6532 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output133
timestamp 1676037725
transform 1 0 8372 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output134
timestamp 1676037725
transform 1 0 9108 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output135
timestamp 1676037725
transform 1 0 1564 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output136
timestamp 1676037725
transform 1 0 1564 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output137
timestamp 1676037725
transform 1 0 1564 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output138
timestamp 1676037725
transform 1 0 1564 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output139
timestamp 1676037725
transform 1 0 1564 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output140
timestamp 1676037725
transform 1 0 1564 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output141
timestamp 1676037725
transform 1 0 1564 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output142
timestamp 1676037725
transform 1 0 1564 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output143
timestamp 1676037725
transform 1 0 45816 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output144
timestamp 1676037725
transform 1 0 47932 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output145
timestamp 1676037725
transform 1 0 47932 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output146
timestamp 1676037725
transform 1 0 46092 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output147
timestamp 1676037725
transform 1 0 47932 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output148
timestamp 1676037725
transform 1 0 47932 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output149
timestamp 1676037725
transform 1 0 47932 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output150
timestamp 1676037725
transform 1 0 45816 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output151
timestamp 1676037725
transform 1 0 47932 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output152
timestamp 1676037725
transform 1 0 47932 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output153
timestamp 1676037725
transform 1 0 47932 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output154
timestamp 1676037725
transform 1 0 43976 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output155
timestamp 1676037725
transform 1 0 46092 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output156
timestamp 1676037725
transform 1 0 47932 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output157
timestamp 1676037725
transform 1 0 47932 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output158
timestamp 1676037725
transform 1 0 47932 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output159
timestamp 1676037725
transform 1 0 47932 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output160
timestamp 1676037725
transform 1 0 47932 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output161
timestamp 1676037725
transform 1 0 47932 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output162
timestamp 1676037725
transform 1 0 47932 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output163
timestamp 1676037725
transform 1 0 47932 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output164
timestamp 1676037725
transform 1 0 47932 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output165
timestamp 1676037725
transform 1 0 45816 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output166
timestamp 1676037725
transform 1 0 45816 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output167
timestamp 1676037725
transform 1 0 46092 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output168
timestamp 1676037725
transform 1 0 47932 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output169
timestamp 1676037725
transform 1 0 47932 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output170
timestamp 1676037725
transform 1 0 47932 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output171
timestamp 1676037725
transform 1 0 45816 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output172
timestamp 1676037725
transform 1 0 47932 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output173
timestamp 1676037725
transform 1 0 3956 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output174
timestamp 1676037725
transform 1 0 7176 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output175
timestamp 1676037725
transform 1 0 7912 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output176
timestamp 1676037725
transform 1 0 9752 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output177
timestamp 1676037725
transform 1 0 9752 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output178
timestamp 1676037725
transform 1 0 10488 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output179
timestamp 1676037725
transform 1 0 9752 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output180
timestamp 1676037725
transform 1 0 12604 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output181
timestamp 1676037725
transform 1 0 12328 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output182
timestamp 1676037725
transform 1 0 12328 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output183
timestamp 1676037725
transform 1 0 13064 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output184
timestamp 1676037725
transform 1 0 3404 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output185
timestamp 1676037725
transform 1 0 14904 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output186
timestamp 1676037725
transform 1 0 15272 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output187
timestamp 1676037725
transform 1 0 14904 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output188
timestamp 1676037725
transform 1 0 17388 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output189
timestamp 1676037725
transform 1 0 14904 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output190
timestamp 1676037725
transform 1 0 16928 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output191
timestamp 1676037725
transform 1 0 19412 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output192
timestamp 1676037725
transform 1 0 17480 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output193
timestamp 1676037725
transform 1 0 21988 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output194
timestamp 1676037725
transform 1 0 20056 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output195
timestamp 1676037725
transform 1 0 2024 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output196
timestamp 1676037725
transform 1 0 2760 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output197
timestamp 1676037725
transform 1 0 4600 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output198
timestamp 1676037725
transform 1 0 4600 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output199
timestamp 1676037725
transform 1 0 5336 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output200
timestamp 1676037725
transform 1 0 4600 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output201
timestamp 1676037725
transform 1 0 7452 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output202
timestamp 1676037725
transform 1 0 7176 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output203
timestamp 1676037725
transform 1 0 11776 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output204
timestamp 1676037725
transform 1 0 14260 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output205
timestamp 1676037725
transform 1 0 16836 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output206
timestamp 1676037725
transform 1 0 18124 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output207
timestamp 1676037725
transform 1 0 20056 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output208
timestamp 1676037725
transform 1 0 22356 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output209
timestamp 1676037725
transform 1 0 24564 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output210
timestamp 1676037725
transform 1 0 27140 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 49864 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 49864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 49864 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 49864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 49864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 49864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 49864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 49864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 49864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 49864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 49864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 49864 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 49864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 49864 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 49864 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 49864 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 49864 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 49864 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 49864 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 49864 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 49864 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 49864 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 49864 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 49864 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 49864 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 49864 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 49864 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 49864 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 49864 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 49864 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 49864 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 49864 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 49864 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 49864 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 49864 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 49864 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 49864 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 49864 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 49864 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 49864 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 49864 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 27140 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24564 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 22632 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22264 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20516 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 17020 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 18584 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20240 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 17112 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19136 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21988 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 19688 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21068 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20976 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 19136 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19596 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19688 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 17112 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19412 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20332 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 18768 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21988 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23828 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 23460 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 25760 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 27048 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 25576 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 27232 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 28060 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 24840 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 25668 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24840 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 21160 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22448 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 28336 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 30452 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 32292 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 32200 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 34868 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 35052 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 34868 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 36432 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 37444 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 34868 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 35144 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 35696 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 33856 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 34868 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 33764 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 29992 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 32108 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 31004 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 27968 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 29716 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 28428 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 26956 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 28796 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 30360 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 31096 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 32292 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 30728 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 29716 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 27508 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 26864 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 41492 0 1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 30820 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 29992 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 31372 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 33672 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 33580 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 35052 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 34868 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 32292 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 32476 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 37444 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 37260 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 37260 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 37996 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 37628 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 37720 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 35788 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 33580 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 35604 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 37904 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 37996 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 40020 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 38916 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 37720 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 38180 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 40020 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 37720 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 37444 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 37076 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 32292 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 29348 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 25576 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 24840 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23828 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 24564 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23920 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 24564 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24564 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23460 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22264 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21988 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19688 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19412 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19320 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20240 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21988 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20424 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16836 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13064 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 12972 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14260 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14260 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 12696 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11684 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 10580 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11960 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14260 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14536 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 15180 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16836 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17112 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30728 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 27232 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l1_in_2_
timestamp 1676037725
transform 1 0 22632 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_1.mux_l1_in_3__258
timestamp 1676037725
transform 1 0 26036 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l1_in_3_
timestamp 1676037725
transform 1 0 20884 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 25852 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l2_in_1_
timestamp 1676037725
transform 1 0 23092 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_1.mux_l3_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17204 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27140 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24564 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19872 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_3.mux_l2_in_1__211
timestamp 1676037725
transform 1 0 15456 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l2_in_1_
timestamp 1676037725
transform 1 0 16744 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_3.mux_l3_in_0_
timestamp 1676037725
transform 1 0 16836 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9936 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l1_in_0_
timestamp 1676037725
transform 1 0 25576 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24656 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_5.mux_l2_in_1__214
timestamp 1676037725
transform 1 0 19412 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l2_in_1_
timestamp 1676037725
transform 1 0 18308 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_5.mux_l3_in_0_
timestamp 1676037725
transform 1 0 17388 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10948 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27140 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24656 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l1_in_2_
timestamp 1676037725
transform 1 0 19504 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l2_in_0_
timestamp 1676037725
transform 1 0 23092 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l2_in_1_
timestamp 1676037725
transform 1 0 19688 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_7.mux_l2_in_1__216
timestamp 1676037725
transform 1 0 18676 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_7.mux_l3_in_0_
timestamp 1676037725
transform 1 0 19872 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16836 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27968 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l1_in_1_
timestamp 1676037725
transform 1 0 25760 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l1_in_2_
timestamp 1676037725
transform 1 0 20884 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_11.mux_l1_in_3__259
timestamp 1676037725
transform 1 0 21988 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l1_in_3_
timestamp 1676037725
transform 1 0 20700 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22080 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l2_in_1_
timestamp 1676037725
transform 1 0 19504 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_11.mux_l3_in_0_
timestamp 1676037725
transform 1 0 17940 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 11868 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27140 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24748 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l1_in_2_
timestamp 1676037725
transform 1 0 21160 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21436 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_13.mux_l2_in_1__260
timestamp 1676037725
transform 1 0 16468 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l2_in_1_
timestamp 1676037725
transform 1 0 18124 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_13.mux_l3_in_0_
timestamp 1676037725
transform 1 0 15640 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10580 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27876 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24564 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l1_in_2_
timestamp 1676037725
transform 1 0 21068 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l2_in_0_
timestamp 1676037725
transform 1 0 23276 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_21.mux_l2_in_1__261
timestamp 1676037725
transform 1 0 16836 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l2_in_1_
timestamp 1676037725
transform 1 0 18124 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_21.mux_l3_in_0_
timestamp 1676037725
transform 1 0 17388 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9660 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l1_in_0_
timestamp 1676037725
transform 1 0 29532 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l1_in_1_
timestamp 1676037725
transform 1 0 26772 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l1_in_2_
timestamp 1676037725
transform 1 0 24104 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l2_in_0_
timestamp 1676037725
transform 1 0 25668 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l2_in_1_
timestamp 1676037725
transform 1 0 23276 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_29.mux_l2_in_1__262
timestamp 1676037725
transform 1 0 22632 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_29.mux_l3_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 13524 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l1_in_0_
timestamp 1676037725
transform 1 0 32108 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l1_in_1_
timestamp 1676037725
transform 1 0 29716 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l2_in_0_
timestamp 1676037725
transform 1 0 28336 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_37.mux_l2_in_1__212
timestamp 1676037725
transform 1 0 23828 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l2_in_1_
timestamp 1676037725
transform 1 0 23276 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_37.mux_l3_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18400 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_45.mux_l1_in_0_
timestamp 1676037725
transform 1 0 32292 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_45.mux_l2_in_0_
timestamp 1676037725
transform 1 0 28336 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_45.mux_l2_in_1_
timestamp 1676037725
transform 1 0 28336 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_45.mux_l2_in_1__213
timestamp 1676037725
transform 1 0 27692 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_45.mux_l3_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 11132 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_53.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30268 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_53.mux_l2_in_0_
timestamp 1676037725
transform 1 0 25944 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_53.mux_l2_in_1_
timestamp 1676037725
transform 1 0 22632 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_left_track_53.mux_l2_in_1__215
timestamp 1676037725
transform 1 0 24564 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_left_track_53.mux_l3_in_0_
timestamp 1676037725
transform 1 0 19964 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 13524 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l1_in_0_
timestamp 1676037725
transform 1 0 29440 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 33304 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l1_in_2_
timestamp 1676037725
transform 1 0 27784 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 31004 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_0.mux_l2_in_1__217
timestamp 1676037725
transform 1 0 29808 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 30912 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 33488 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 39284 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 33212 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 32292 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 29716 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 35880 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_2.mux_l2_in_1__220
timestamp 1676037725
transform 1 0 33856 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 33488 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 37996 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 40848 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l1_in_0_
timestamp 1676037725
transform 1 0 34408 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l1_in_1_
timestamp 1676037725
transform 1 0 36248 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l1_in_2_
timestamp 1676037725
transform 1 0 29716 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 35972 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l2_in_1_
timestamp 1676037725
transform 1 0 35696 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_4.mux_l2_in_1__224
timestamp 1676037725
transform 1 0 31556 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_4.mux_l3_in_0_
timestamp 1676037725
transform 1 0 37444 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 41308 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l1_in_0_
timestamp 1676037725
transform 1 0 34868 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l1_in_1_
timestamp 1676037725
transform 1 0 32752 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l1_in_2_
timestamp 1676037725
transform 1 0 35420 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_6.mux_l1_in_3__227
timestamp 1676037725
transform 1 0 33764 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l1_in_3_
timestamp 1676037725
transform 1 0 32292 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l2_in_0_
timestamp 1676037725
transform 1 0 35880 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l2_in_1_
timestamp 1676037725
transform 1 0 38640 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_6.mux_l3_in_0_
timestamp 1676037725
transform 1 0 38272 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 41400 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l1_in_0_
timestamp 1676037725
transform 1 0 33396 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l1_in_1_
timestamp 1676037725
transform 1 0 32660 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l1_in_2_
timestamp 1676037725
transform 1 0 33304 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l1_in_3_
timestamp 1676037725
transform 1 0 31004 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_10.mux_l1_in_3__218
timestamp 1676037725
transform 1 0 30912 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 34500 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l2_in_1_
timestamp 1676037725
transform 1 0 36064 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_10.mux_l3_in_0_
timestamp 1676037725
transform 1 0 37444 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 40756 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l1_in_0_
timestamp 1676037725
transform 1 0 32292 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l1_in_1_
timestamp 1676037725
transform 1 0 32292 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l1_in_2_
timestamp 1676037725
transform 1 0 27140 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l2_in_0_
timestamp 1676037725
transform 1 0 33304 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l2_in_1_
timestamp 1676037725
transform 1 0 32292 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_12.mux_l2_in_1__219
timestamp 1676037725
transform 1 0 29716 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_12.mux_l3_in_0_
timestamp 1676037725
transform 1 0 37076 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 40756 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30636 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l1_in_1_
timestamp 1676037725
transform 1 0 29808 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l1_in_2_
timestamp 1676037725
transform 1 0 27140 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l2_in_0_
timestamp 1676037725
transform 1 0 30544 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_20.mux_l2_in_1__221
timestamp 1676037725
transform 1 0 28980 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l2_in_1_
timestamp 1676037725
transform 1 0 28428 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_20.mux_l3_in_0_
timestamp 1676037725
transform 1 0 33488 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 38180 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 29716 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l1_in_1_
timestamp 1676037725
transform 1 0 30176 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l1_in_2_
timestamp 1676037725
transform 1 0 25668 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l2_in_0_
timestamp 1676037725
transform 1 0 29716 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l2_in_1_
timestamp 1676037725
transform 1 0 30176 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_28.mux_l2_in_1__222
timestamp 1676037725
transform 1 0 29716 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_28.mux_l3_in_0_
timestamp 1676037725
transform 1 0 32568 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 37628 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l1_in_0_
timestamp 1676037725
transform 1 0 31280 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l1_in_1_
timestamp 1676037725
transform 1 0 32108 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l2_in_0_
timestamp 1676037725
transform 1 0 32292 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l2_in_1_
timestamp 1676037725
transform 1 0 31004 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_36.mux_l2_in_1__223
timestamp 1676037725
transform 1 0 32292 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_36.mux_l3_in_0_
timestamp 1676037725
transform 1 0 34868 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 38916 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_44.mux_l1_in_0_
timestamp 1676037725
transform 1 0 29716 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_44.mux_l1_in_1__225
timestamp 1676037725
transform 1 0 29716 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_44.mux_l1_in_1_
timestamp 1676037725
transform 1 0 28152 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_44.mux_l2_in_0_
timestamp 1676037725
transform 1 0 32568 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 37444 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_52.mux_l1_in_0_
timestamp 1676037725
transform 1 0 28612 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_52.mux_l1_in_1_
timestamp 1676037725
transform 1 0 26956 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_right_track_52.mux_l1_in_1__226
timestamp 1676037725
transform 1 0 26404 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_right_track_52.mux_l2_in_0_
timestamp 1676037725
transform 1 0 32292 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 36524 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l1_in_0_
timestamp 1676037725
transform 1 0 34868 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 38824 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l1_in_2_
timestamp 1676037725
transform 1 0 23276 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_0.mux_l1_in_3__228
timestamp 1676037725
transform 1 0 29716 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l1_in_3_
timestamp 1676037725
transform 1 0 28428 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 35880 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 28336 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 29716 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 27140 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 34868 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 40020 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 30912 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 37444 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 33028 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_2.mux_l2_in_1__234
timestamp 1676037725
transform 1 0 32568 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 32292 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 28428 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l1_in_0_
timestamp 1676037725
transform 1 0 34500 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l1_in_1_
timestamp 1676037725
transform 1 0 40020 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 35696 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_4.mux_l2_in_1__244
timestamp 1676037725
transform 1 0 31280 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l2_in_1_
timestamp 1676037725
transform 1 0 30084 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_4.mux_l3_in_0_
timestamp 1676037725
transform 1 0 30820 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 27140 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l1_in_0_
timestamp 1676037725
transform 1 0 40204 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l1_in_1_
timestamp 1676037725
transform 1 0 41216 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l1_in_2_
timestamp 1676037725
transform 1 0 32660 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l2_in_0_
timestamp 1676037725
transform 1 0 39652 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l2_in_1_
timestamp 1676037725
transform 1 0 36064 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_6.mux_l2_in_1__252
timestamp 1676037725
transform 1 0 34960 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_6.mux_l3_in_0_
timestamp 1676037725
transform 1 0 33580 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 29716 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l1_in_0_
timestamp 1676037725
transform 1 0 37444 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l1_in_1_
timestamp 1676037725
transform 1 0 41216 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l1_in_2_
timestamp 1676037725
transform 1 0 33488 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l2_in_0_
timestamp 1676037725
transform 1 0 40020 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l2_in_1_
timestamp 1676037725
transform 1 0 36064 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_8.mux_l2_in_1__253
timestamp 1676037725
transform 1 0 41124 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_8.mux_l3_in_0_
timestamp 1676037725
transform 1 0 36064 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 31464 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l1_in_0_
timestamp 1676037725
transform 1 0 34684 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l1_in_1_
timestamp 1676037725
transform 1 0 40112 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 36064 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l2_in_1_
timestamp 1676037725
transform 1 0 30912 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_10.mux_l2_in_1__229
timestamp 1676037725
transform 1 0 31372 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_10.mux_l3_in_0_
timestamp 1676037725
transform 1 0 31464 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 26404 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_12.mux_l1_in_0_
timestamp 1676037725
transform 1 0 40020 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_12.mux_l2_in_0_
timestamp 1676037725
transform 1 0 40388 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_12.mux_l2_in_1__230
timestamp 1676037725
transform 1 0 34868 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_12.mux_l2_in_1_
timestamp 1676037725
transform 1 0 37444 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_12.mux_l3_in_0_
timestamp 1676037725
transform 1 0 36064 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 29716 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_14.mux_l1_in_0_
timestamp 1676037725
transform 1 0 39928 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_14.mux_l2_in_0_
timestamp 1676037725
transform 1 0 40480 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_14.mux_l2_in_1__231
timestamp 1676037725
transform 1 0 37444 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_14.mux_l2_in_1_
timestamp 1676037725
transform 1 0 34684 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_14.mux_l3_in_0_
timestamp 1676037725
transform 1 0 37996 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 29716 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_16.mux_l1_in_0_
timestamp 1676037725
transform 1 0 40020 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_16.mux_l2_in_0_
timestamp 1676037725
transform 1 0 40480 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_16.mux_l2_in_1__232
timestamp 1676037725
transform 1 0 37076 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_16.mux_l2_in_1_
timestamp 1676037725
transform 1 0 34868 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_16.mux_l3_in_0_
timestamp 1676037725
transform 1 0 35880 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 28980 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_18.mux_l1_in_0_
timestamp 1676037725
transform 1 0 37812 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_18.mux_l2_in_0_
timestamp 1676037725
transform 1 0 39652 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_18.mux_l2_in_1_
timestamp 1676037725
transform 1 0 30728 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_18.mux_l2_in_1__233
timestamp 1676037725
transform 1 0 31372 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_18.mux_l3_in_0_
timestamp 1676037725
transform 1 0 32292 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 25760 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_20.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27324 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_20.mux_l1_in_1__235
timestamp 1676037725
transform 1 0 24932 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_20.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24840 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_20.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24840 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 23828 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_22.mux_l1_in_0_
timestamp 1676037725
transform 1 0 25852 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_22.mux_l1_in_1__236
timestamp 1676037725
transform 1 0 24196 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_22.mux_l1_in_1_
timestamp 1676037725
transform 1 0 23276 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_22.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22908 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20056 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_24.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27140 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_24.mux_l1_in_1_
timestamp 1676037725
transform 1 0 22080 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_24.mux_l1_in_1__237
timestamp 1676037725
transform 1 0 19780 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_24.mux_l2_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16100 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_26.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27416 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_26.mux_l1_in_1__238
timestamp 1676037725
transform 1 0 25392 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_26.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24196 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_26.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22080 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19412 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 22264 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_28.mux_l2_in_0__239
timestamp 1676037725
transform 1 0 22632 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_28.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14904 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_30.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_30.mux_l2_in_0__240
timestamp 1676037725
transform 1 0 17204 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_30.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 12880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_32.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_32.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16744 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_32.mux_l2_in_0__241
timestamp 1676037725
transform 1 0 19044 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 12328 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_34.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19504 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_34.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19228 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_34.mux_l2_in_0__242
timestamp 1676037725
transform 1 0 19504 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14904 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_36.mux_l1_in_0_
timestamp 1676037725
transform 1 0 25852 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_36.mux_l1_in_1__243
timestamp 1676037725
transform 1 0 21620 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_36.mux_l1_in_1_
timestamp 1676037725
transform 1 0 21988 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_36.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14260 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_40.mux_l1_in_0_
timestamp 1676037725
transform 1 0 13156 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_40.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11776 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_40.mux_l2_in_0__245
timestamp 1676037725
transform 1 0 13064 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_40.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9752 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_42.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16744 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_42.mux_l2_in_0__246
timestamp 1676037725
transform 1 0 10948 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_42.mux_l2_in_0_
timestamp 1676037725
transform 1 0 13892 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_42.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10488 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_44.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_44.mux_l2_in_0__247
timestamp 1676037725
transform 1 0 10304 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_44.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12512 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10304 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_46.mux_l1_in_0_
timestamp 1676037725
transform 1 0 11868 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_46.mux_l2_in_0__248
timestamp 1676037725
transform 1 0 9660 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_46.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10396 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9016 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_48.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_48.mux_l2_in_0_
timestamp 1676037725
transform 1 0 13708 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_48.mux_l2_in_0__249
timestamp 1676037725
transform 1 0 10488 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9200 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_50.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16928 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_50.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_50.mux_l2_in_0__250
timestamp 1676037725
transform 1 0 9844 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 8372 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_58.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_1__0_.mux_top_track_58.mux_l2_in_0__251
timestamp 1676037725
transform 1 0 9844 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_1__0_.mux_top_track_58.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_1__0_.mux_top_track_58.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9108 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1676037725
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1676037725
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1676037725
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1676037725
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1676037725
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1676037725
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1676037725
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1676037725
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1676037725
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1676037725
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1676037725
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1676037725
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1676037725
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1676037725
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1676037725
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1676037725
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 6256 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 11408 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 16560 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 21712 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 26864 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 32016 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 37168 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 42320 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 47472 0 1 23936
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 27944 2128 28264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 37944 2128 38264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 47944 2128 48264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 32944 2128 33264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 42944 2128 43264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 ccff_head
port 2 nsew signal input
flabel metal2 s 49238 26200 49294 27000 0 FreeSans 224 90 0 0 ccff_head_1
port 3 nsew signal input
flabel metal2 s 41326 0 41382 800 0 FreeSans 224 90 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal2 s 1582 26200 1638 27000 0 FreeSans 224 90 0 0 ccff_tail_0
port 5 nsew signal tristate
flabel metal3 s 0 1504 800 1624 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 6 nsew signal input
flabel metal3 s 0 5584 800 5704 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 7 nsew signal input
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 8 nsew signal input
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 9 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 10 nsew signal input
flabel metal3 s 0 7216 800 7336 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 11 nsew signal input
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 12 nsew signal input
flabel metal3 s 0 8032 800 8152 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 13 nsew signal input
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 14 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 15 nsew signal input
flabel metal3 s 0 9256 800 9376 0 FreeSans 480 0 0 0 chanx_left_in[19]
port 16 nsew signal input
flabel metal3 s 0 1912 800 2032 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 17 nsew signal input
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 chanx_left_in[20]
port 18 nsew signal input
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 chanx_left_in[21]
port 19 nsew signal input
flabel metal3 s 0 10480 800 10600 0 FreeSans 480 0 0 0 chanx_left_in[22]
port 20 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 chanx_left_in[23]
port 21 nsew signal input
flabel metal3 s 0 11296 800 11416 0 FreeSans 480 0 0 0 chanx_left_in[24]
port 22 nsew signal input
flabel metal3 s 0 11704 800 11824 0 FreeSans 480 0 0 0 chanx_left_in[25]
port 23 nsew signal input
flabel metal3 s 0 12112 800 12232 0 FreeSans 480 0 0 0 chanx_left_in[26]
port 24 nsew signal input
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 chanx_left_in[27]
port 25 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 chanx_left_in[28]
port 26 nsew signal input
flabel metal3 s 0 13336 800 13456 0 FreeSans 480 0 0 0 chanx_left_in[29]
port 27 nsew signal input
flabel metal3 s 0 2320 800 2440 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 28 nsew signal input
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 29 nsew signal input
flabel metal3 s 0 3136 800 3256 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 30 nsew signal input
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 31 nsew signal input
flabel metal3 s 0 3952 800 4072 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 32 nsew signal input
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 33 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 34 nsew signal input
flabel metal3 s 0 5176 800 5296 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 35 nsew signal input
flabel metal3 s 0 13744 800 13864 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 36 nsew signal tristate
flabel metal3 s 0 17824 800 17944 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 37 nsew signal tristate
flabel metal3 s 0 18232 800 18352 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 38 nsew signal tristate
flabel metal3 s 0 18640 800 18760 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 39 nsew signal tristate
flabel metal3 s 0 19048 800 19168 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 40 nsew signal tristate
flabel metal3 s 0 19456 800 19576 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 41 nsew signal tristate
flabel metal3 s 0 19864 800 19984 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 42 nsew signal tristate
flabel metal3 s 0 20272 800 20392 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 43 nsew signal tristate
flabel metal3 s 0 20680 800 20800 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 44 nsew signal tristate
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 45 nsew signal tristate
flabel metal3 s 0 21496 800 21616 0 FreeSans 480 0 0 0 chanx_left_out[19]
port 46 nsew signal tristate
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 47 nsew signal tristate
flabel metal3 s 0 21904 800 22024 0 FreeSans 480 0 0 0 chanx_left_out[20]
port 48 nsew signal tristate
flabel metal3 s 0 22312 800 22432 0 FreeSans 480 0 0 0 chanx_left_out[21]
port 49 nsew signal tristate
flabel metal3 s 0 22720 800 22840 0 FreeSans 480 0 0 0 chanx_left_out[22]
port 50 nsew signal tristate
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 chanx_left_out[23]
port 51 nsew signal tristate
flabel metal3 s 0 23536 800 23656 0 FreeSans 480 0 0 0 chanx_left_out[24]
port 52 nsew signal tristate
flabel metal3 s 0 23944 800 24064 0 FreeSans 480 0 0 0 chanx_left_out[25]
port 53 nsew signal tristate
flabel metal3 s 0 24352 800 24472 0 FreeSans 480 0 0 0 chanx_left_out[26]
port 54 nsew signal tristate
flabel metal3 s 0 24760 800 24880 0 FreeSans 480 0 0 0 chanx_left_out[27]
port 55 nsew signal tristate
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 chanx_left_out[28]
port 56 nsew signal tristate
flabel metal3 s 0 25576 800 25696 0 FreeSans 480 0 0 0 chanx_left_out[29]
port 57 nsew signal tristate
flabel metal3 s 0 14560 800 14680 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 58 nsew signal tristate
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 59 nsew signal tristate
flabel metal3 s 0 15376 800 15496 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 60 nsew signal tristate
flabel metal3 s 0 15784 800 15904 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 61 nsew signal tristate
flabel metal3 s 0 16192 800 16312 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 62 nsew signal tristate
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 63 nsew signal tristate
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 64 nsew signal tristate
flabel metal3 s 0 17416 800 17536 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 65 nsew signal tristate
flabel metal3 s 50200 13608 51000 13728 0 FreeSans 480 0 0 0 chanx_right_in_0[0]
port 66 nsew signal input
flabel metal3 s 50200 17688 51000 17808 0 FreeSans 480 0 0 0 chanx_right_in_0[10]
port 67 nsew signal input
flabel metal3 s 50200 18096 51000 18216 0 FreeSans 480 0 0 0 chanx_right_in_0[11]
port 68 nsew signal input
flabel metal3 s 50200 18504 51000 18624 0 FreeSans 480 0 0 0 chanx_right_in_0[12]
port 69 nsew signal input
flabel metal3 s 50200 18912 51000 19032 0 FreeSans 480 0 0 0 chanx_right_in_0[13]
port 70 nsew signal input
flabel metal3 s 50200 19320 51000 19440 0 FreeSans 480 0 0 0 chanx_right_in_0[14]
port 71 nsew signal input
flabel metal3 s 50200 19728 51000 19848 0 FreeSans 480 0 0 0 chanx_right_in_0[15]
port 72 nsew signal input
flabel metal3 s 50200 20136 51000 20256 0 FreeSans 480 0 0 0 chanx_right_in_0[16]
port 73 nsew signal input
flabel metal3 s 50200 20544 51000 20664 0 FreeSans 480 0 0 0 chanx_right_in_0[17]
port 74 nsew signal input
flabel metal3 s 50200 20952 51000 21072 0 FreeSans 480 0 0 0 chanx_right_in_0[18]
port 75 nsew signal input
flabel metal3 s 50200 21360 51000 21480 0 FreeSans 480 0 0 0 chanx_right_in_0[19]
port 76 nsew signal input
flabel metal3 s 50200 14016 51000 14136 0 FreeSans 480 0 0 0 chanx_right_in_0[1]
port 77 nsew signal input
flabel metal3 s 50200 21768 51000 21888 0 FreeSans 480 0 0 0 chanx_right_in_0[20]
port 78 nsew signal input
flabel metal3 s 50200 22176 51000 22296 0 FreeSans 480 0 0 0 chanx_right_in_0[21]
port 79 nsew signal input
flabel metal3 s 50200 22584 51000 22704 0 FreeSans 480 0 0 0 chanx_right_in_0[22]
port 80 nsew signal input
flabel metal3 s 50200 22992 51000 23112 0 FreeSans 480 0 0 0 chanx_right_in_0[23]
port 81 nsew signal input
flabel metal3 s 50200 23400 51000 23520 0 FreeSans 480 0 0 0 chanx_right_in_0[24]
port 82 nsew signal input
flabel metal3 s 50200 23808 51000 23928 0 FreeSans 480 0 0 0 chanx_right_in_0[25]
port 83 nsew signal input
flabel metal3 s 50200 24216 51000 24336 0 FreeSans 480 0 0 0 chanx_right_in_0[26]
port 84 nsew signal input
flabel metal3 s 50200 24624 51000 24744 0 FreeSans 480 0 0 0 chanx_right_in_0[27]
port 85 nsew signal input
flabel metal3 s 50200 25032 51000 25152 0 FreeSans 480 0 0 0 chanx_right_in_0[28]
port 86 nsew signal input
flabel metal3 s 50200 25440 51000 25560 0 FreeSans 480 0 0 0 chanx_right_in_0[29]
port 87 nsew signal input
flabel metal3 s 50200 14424 51000 14544 0 FreeSans 480 0 0 0 chanx_right_in_0[2]
port 88 nsew signal input
flabel metal3 s 50200 14832 51000 14952 0 FreeSans 480 0 0 0 chanx_right_in_0[3]
port 89 nsew signal input
flabel metal3 s 50200 15240 51000 15360 0 FreeSans 480 0 0 0 chanx_right_in_0[4]
port 90 nsew signal input
flabel metal3 s 50200 15648 51000 15768 0 FreeSans 480 0 0 0 chanx_right_in_0[5]
port 91 nsew signal input
flabel metal3 s 50200 16056 51000 16176 0 FreeSans 480 0 0 0 chanx_right_in_0[6]
port 92 nsew signal input
flabel metal3 s 50200 16464 51000 16584 0 FreeSans 480 0 0 0 chanx_right_in_0[7]
port 93 nsew signal input
flabel metal3 s 50200 16872 51000 16992 0 FreeSans 480 0 0 0 chanx_right_in_0[8]
port 94 nsew signal input
flabel metal3 s 50200 17280 51000 17400 0 FreeSans 480 0 0 0 chanx_right_in_0[9]
port 95 nsew signal input
flabel metal3 s 50200 1368 51000 1488 0 FreeSans 480 0 0 0 chanx_right_out_0[0]
port 96 nsew signal tristate
flabel metal3 s 50200 5448 51000 5568 0 FreeSans 480 0 0 0 chanx_right_out_0[10]
port 97 nsew signal tristate
flabel metal3 s 50200 5856 51000 5976 0 FreeSans 480 0 0 0 chanx_right_out_0[11]
port 98 nsew signal tristate
flabel metal3 s 50200 6264 51000 6384 0 FreeSans 480 0 0 0 chanx_right_out_0[12]
port 99 nsew signal tristate
flabel metal3 s 50200 6672 51000 6792 0 FreeSans 480 0 0 0 chanx_right_out_0[13]
port 100 nsew signal tristate
flabel metal3 s 50200 7080 51000 7200 0 FreeSans 480 0 0 0 chanx_right_out_0[14]
port 101 nsew signal tristate
flabel metal3 s 50200 7488 51000 7608 0 FreeSans 480 0 0 0 chanx_right_out_0[15]
port 102 nsew signal tristate
flabel metal3 s 50200 7896 51000 8016 0 FreeSans 480 0 0 0 chanx_right_out_0[16]
port 103 nsew signal tristate
flabel metal3 s 50200 8304 51000 8424 0 FreeSans 480 0 0 0 chanx_right_out_0[17]
port 104 nsew signal tristate
flabel metal3 s 50200 8712 51000 8832 0 FreeSans 480 0 0 0 chanx_right_out_0[18]
port 105 nsew signal tristate
flabel metal3 s 50200 9120 51000 9240 0 FreeSans 480 0 0 0 chanx_right_out_0[19]
port 106 nsew signal tristate
flabel metal3 s 50200 1776 51000 1896 0 FreeSans 480 0 0 0 chanx_right_out_0[1]
port 107 nsew signal tristate
flabel metal3 s 50200 9528 51000 9648 0 FreeSans 480 0 0 0 chanx_right_out_0[20]
port 108 nsew signal tristate
flabel metal3 s 50200 9936 51000 10056 0 FreeSans 480 0 0 0 chanx_right_out_0[21]
port 109 nsew signal tristate
flabel metal3 s 50200 10344 51000 10464 0 FreeSans 480 0 0 0 chanx_right_out_0[22]
port 110 nsew signal tristate
flabel metal3 s 50200 10752 51000 10872 0 FreeSans 480 0 0 0 chanx_right_out_0[23]
port 111 nsew signal tristate
flabel metal3 s 50200 11160 51000 11280 0 FreeSans 480 0 0 0 chanx_right_out_0[24]
port 112 nsew signal tristate
flabel metal3 s 50200 11568 51000 11688 0 FreeSans 480 0 0 0 chanx_right_out_0[25]
port 113 nsew signal tristate
flabel metal3 s 50200 11976 51000 12096 0 FreeSans 480 0 0 0 chanx_right_out_0[26]
port 114 nsew signal tristate
flabel metal3 s 50200 12384 51000 12504 0 FreeSans 480 0 0 0 chanx_right_out_0[27]
port 115 nsew signal tristate
flabel metal3 s 50200 12792 51000 12912 0 FreeSans 480 0 0 0 chanx_right_out_0[28]
port 116 nsew signal tristate
flabel metal3 s 50200 13200 51000 13320 0 FreeSans 480 0 0 0 chanx_right_out_0[29]
port 117 nsew signal tristate
flabel metal3 s 50200 2184 51000 2304 0 FreeSans 480 0 0 0 chanx_right_out_0[2]
port 118 nsew signal tristate
flabel metal3 s 50200 2592 51000 2712 0 FreeSans 480 0 0 0 chanx_right_out_0[3]
port 119 nsew signal tristate
flabel metal3 s 50200 3000 51000 3120 0 FreeSans 480 0 0 0 chanx_right_out_0[4]
port 120 nsew signal tristate
flabel metal3 s 50200 3408 51000 3528 0 FreeSans 480 0 0 0 chanx_right_out_0[5]
port 121 nsew signal tristate
flabel metal3 s 50200 3816 51000 3936 0 FreeSans 480 0 0 0 chanx_right_out_0[6]
port 122 nsew signal tristate
flabel metal3 s 50200 4224 51000 4344 0 FreeSans 480 0 0 0 chanx_right_out_0[7]
port 123 nsew signal tristate
flabel metal3 s 50200 4632 51000 4752 0 FreeSans 480 0 0 0 chanx_right_out_0[8]
port 124 nsew signal tristate
flabel metal3 s 50200 5040 51000 5160 0 FreeSans 480 0 0 0 chanx_right_out_0[9]
port 125 nsew signal tristate
flabel metal2 s 21546 26200 21602 27000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 126 nsew signal input
flabel metal2 s 27986 26200 28042 27000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 127 nsew signal input
flabel metal2 s 28630 26200 28686 27000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 128 nsew signal input
flabel metal2 s 29274 26200 29330 27000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 129 nsew signal input
flabel metal2 s 29918 26200 29974 27000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 130 nsew signal input
flabel metal2 s 30562 26200 30618 27000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 131 nsew signal input
flabel metal2 s 31206 26200 31262 27000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 132 nsew signal input
flabel metal2 s 31850 26200 31906 27000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 133 nsew signal input
flabel metal2 s 32494 26200 32550 27000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 134 nsew signal input
flabel metal2 s 33138 26200 33194 27000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 135 nsew signal input
flabel metal2 s 33782 26200 33838 27000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 136 nsew signal input
flabel metal2 s 22190 26200 22246 27000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 137 nsew signal input
flabel metal2 s 34426 26200 34482 27000 0 FreeSans 224 90 0 0 chany_top_in[20]
port 138 nsew signal input
flabel metal2 s 35070 26200 35126 27000 0 FreeSans 224 90 0 0 chany_top_in[21]
port 139 nsew signal input
flabel metal2 s 35714 26200 35770 27000 0 FreeSans 224 90 0 0 chany_top_in[22]
port 140 nsew signal input
flabel metal2 s 36358 26200 36414 27000 0 FreeSans 224 90 0 0 chany_top_in[23]
port 141 nsew signal input
flabel metal2 s 37002 26200 37058 27000 0 FreeSans 224 90 0 0 chany_top_in[24]
port 142 nsew signal input
flabel metal2 s 37646 26200 37702 27000 0 FreeSans 224 90 0 0 chany_top_in[25]
port 143 nsew signal input
flabel metal2 s 38290 26200 38346 27000 0 FreeSans 224 90 0 0 chany_top_in[26]
port 144 nsew signal input
flabel metal2 s 38934 26200 38990 27000 0 FreeSans 224 90 0 0 chany_top_in[27]
port 145 nsew signal input
flabel metal2 s 39578 26200 39634 27000 0 FreeSans 224 90 0 0 chany_top_in[28]
port 146 nsew signal input
flabel metal2 s 40222 26200 40278 27000 0 FreeSans 224 90 0 0 chany_top_in[29]
port 147 nsew signal input
flabel metal2 s 22834 26200 22890 27000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 148 nsew signal input
flabel metal2 s 23478 26200 23534 27000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 149 nsew signal input
flabel metal2 s 24122 26200 24178 27000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 150 nsew signal input
flabel metal2 s 24766 26200 24822 27000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 151 nsew signal input
flabel metal2 s 25410 26200 25466 27000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 152 nsew signal input
flabel metal2 s 26054 26200 26110 27000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 153 nsew signal input
flabel metal2 s 26698 26200 26754 27000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 154 nsew signal input
flabel metal2 s 27342 26200 27398 27000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 155 nsew signal input
flabel metal2 s 2226 26200 2282 27000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 156 nsew signal tristate
flabel metal2 s 8666 26200 8722 27000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 157 nsew signal tristate
flabel metal2 s 9310 26200 9366 27000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 158 nsew signal tristate
flabel metal2 s 9954 26200 10010 27000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 159 nsew signal tristate
flabel metal2 s 10598 26200 10654 27000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 160 nsew signal tristate
flabel metal2 s 11242 26200 11298 27000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 161 nsew signal tristate
flabel metal2 s 11886 26200 11942 27000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 162 nsew signal tristate
flabel metal2 s 12530 26200 12586 27000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 163 nsew signal tristate
flabel metal2 s 13174 26200 13230 27000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 164 nsew signal tristate
flabel metal2 s 13818 26200 13874 27000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 165 nsew signal tristate
flabel metal2 s 14462 26200 14518 27000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 166 nsew signal tristate
flabel metal2 s 2870 26200 2926 27000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 167 nsew signal tristate
flabel metal2 s 15106 26200 15162 27000 0 FreeSans 224 90 0 0 chany_top_out[20]
port 168 nsew signal tristate
flabel metal2 s 15750 26200 15806 27000 0 FreeSans 224 90 0 0 chany_top_out[21]
port 169 nsew signal tristate
flabel metal2 s 16394 26200 16450 27000 0 FreeSans 224 90 0 0 chany_top_out[22]
port 170 nsew signal tristate
flabel metal2 s 17038 26200 17094 27000 0 FreeSans 224 90 0 0 chany_top_out[23]
port 171 nsew signal tristate
flabel metal2 s 17682 26200 17738 27000 0 FreeSans 224 90 0 0 chany_top_out[24]
port 172 nsew signal tristate
flabel metal2 s 18326 26200 18382 27000 0 FreeSans 224 90 0 0 chany_top_out[25]
port 173 nsew signal tristate
flabel metal2 s 18970 26200 19026 27000 0 FreeSans 224 90 0 0 chany_top_out[26]
port 174 nsew signal tristate
flabel metal2 s 19614 26200 19670 27000 0 FreeSans 224 90 0 0 chany_top_out[27]
port 175 nsew signal tristate
flabel metal2 s 20258 26200 20314 27000 0 FreeSans 224 90 0 0 chany_top_out[28]
port 176 nsew signal tristate
flabel metal2 s 20902 26200 20958 27000 0 FreeSans 224 90 0 0 chany_top_out[29]
port 177 nsew signal tristate
flabel metal2 s 3514 26200 3570 27000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 178 nsew signal tristate
flabel metal2 s 4158 26200 4214 27000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 179 nsew signal tristate
flabel metal2 s 4802 26200 4858 27000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 180 nsew signal tristate
flabel metal2 s 5446 26200 5502 27000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 181 nsew signal tristate
flabel metal2 s 6090 26200 6146 27000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 182 nsew signal tristate
flabel metal2 s 6734 26200 6790 27000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 183 nsew signal tristate
flabel metal2 s 7378 26200 7434 27000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 184 nsew signal tristate
flabel metal2 s 8022 26200 8078 27000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 185 nsew signal tristate
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[0]
port 186 nsew signal tristate
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[1]
port 187 nsew signal tristate
flabel metal2 s 15934 0 15990 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[2]
port 188 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[3]
port 189 nsew signal tristate
flabel metal2 s 28630 0 28686 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[0]
port 190 nsew signal input
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[1]
port 191 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[2]
port 192 nsew signal input
flabel metal2 s 34978 0 35034 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[3]
port 193 nsew signal input
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[0]
port 194 nsew signal tristate
flabel metal2 s 22282 0 22338 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[1]
port 195 nsew signal tristate
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[2]
port 196 nsew signal tristate
flabel metal2 s 26514 0 26570 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[3]
port 197 nsew signal tristate
flabel metal2 s 37094 0 37150 800 0 FreeSans 224 90 0 0 isol_n
port 198 nsew signal input
flabel metal2 s 39210 0 39266 800 0 FreeSans 224 90 0 0 prog_clk
port 199 nsew signal input
flabel metal2 s 42154 26200 42210 27000 0 FreeSans 224 90 0 0 prog_reset_top_in
port 200 nsew signal input
flabel metal2 s 42798 26200 42854 27000 0 FreeSans 224 90 0 0 reset_top_in
port 201 nsew signal input
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 202 nsew signal input
flabel metal2 s 45558 0 45614 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
port 203 nsew signal input
flabel metal2 s 47674 0 47730 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
port 204 nsew signal input
flabel metal2 s 49790 0 49846 800 0 FreeSans 224 90 0 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
port 205 nsew signal input
flabel metal2 s 43442 26200 43498 27000 0 FreeSans 224 90 0 0 test_enable_top_in
port 206 nsew signal input
flabel metal2 s 45374 26200 45430 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
port 207 nsew signal input
flabel metal2 s 46018 26200 46074 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
port 208 nsew signal input
flabel metal2 s 46662 26200 46718 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
port 209 nsew signal input
flabel metal2 s 47306 26200 47362 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
port 210 nsew signal input
flabel metal2 s 47950 26200 48006 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
port 211 nsew signal input
flabel metal2 s 48594 26200 48650 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
port 212 nsew signal input
flabel metal2 s 44086 26200 44142 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
port 213 nsew signal input
flabel metal2 s 44730 26200 44786 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
port 214 nsew signal input
flabel metal2 s 1122 0 1178 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_0__pin_inpad_0_
port 215 nsew signal tristate
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_1__pin_inpad_0_
port 216 nsew signal tristate
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_2__pin_inpad_0_
port 217 nsew signal tristate
flabel metal2 s 7470 0 7526 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_3__pin_inpad_0_
port 218 nsew signal tristate
rlabel metal1 25484 23936 25484 23936 0 VGND
rlabel metal1 25484 24480 25484 24480 0 VPWR
rlabel metal2 21942 5644 21942 5644 0 cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal1 19826 4658 19826 4658 0 cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal2 18906 6630 18906 6630 0 cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal1 17986 6290 17986 6290 0 cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal1 20516 20978 20516 20978 0 cbx_1__0_.cbx_8__0_.ccff_head
rlabel metal2 18630 9044 18630 9044 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.ccff_tail
rlabel metal1 21298 14960 21298 14960 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\]
rlabel metal1 16698 8840 16698 8840 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\]
rlabel metal1 17112 8534 17112 8534 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[2\]
rlabel metal1 14720 9010 14720 9010 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.ccff_tail
rlabel metal1 13294 17136 13294 17136 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\]
rlabel metal2 16238 14654 16238 14654 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\]
rlabel metal1 14996 9894 14996 9894 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[2\]
rlabel metal1 12006 12104 12006 12104 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.ccff_tail
rlabel metal1 14582 14450 14582 14450 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\]
rlabel metal1 9936 12138 9936 12138 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\]
rlabel metal2 11270 11560 11270 11560 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[2\]
rlabel metal1 13754 14926 13754 14926 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\]
rlabel metal1 13340 16014 13340 16014 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\]
rlabel metal2 12558 14892 12558 14892 0 cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[2\]
rlabel metal1 15226 13362 15226 13362 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17480 7786 17480 7786 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 19550 6766 19550 6766 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 15594 13736 15594 13736 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17158 13906 17158 13906 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 17526 14450 17526 14450 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 16514 12614 16514 12614 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 15778 11186 15778 11186 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 16882 14042 16882 14042 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 17066 7922 17066 7922 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 17756 7854 17756 7854 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 18584 7718 18584 7718 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 13478 16422 13478 16422 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 15594 9690 15594 9690 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 17250 6766 17250 6766 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 13064 15470 13064 15470 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16054 13872 16054 13872 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15916 13906 15916 13906 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 13478 10030 13478 10030 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 13340 15402 13340 15402 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 15410 14042 15410 14042 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 14398 10234 14398 10234 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 16560 10778 16560 10778 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal2 15686 10234 15686 10234 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 9752 15062 9752 15062 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12558 10574 12558 10574 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal2 12834 8602 12834 8602 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 9522 15130 9522 15130 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18032 14586 18032 14586 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 14490 14926 14490 14926 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 15686 10642 15686 10642 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 11592 12954 11592 12954 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 12098 14246 12098 14246 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 14306 10778 14306 10778 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 12466 11866 12466 11866 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal2 12650 11118 12650 11118 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 13340 16150 13340 16150 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12834 14586 12834 14586 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 12926 8942 12926 8942 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 13984 16218 13984 16218 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15870 15062 15870 15062 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17158 15130 17158 15130 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 14858 11356 14858 11356 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 12834 16218 12834 16218 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 15594 15283 15594 15283 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 13938 11322 13938 11322 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 14214 14314 14214 14314 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 11776 16218 11776 16218 0 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 21252 3434 21252 3434 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.ccff_tail
rlabel metal1 20194 3060 20194 3060 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
rlabel metal1 26174 3026 26174 3026 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
rlabel metal1 27278 4182 27278 4182 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel via1 23414 3094 23414 3094 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.ccff_tail
rlabel metal1 20102 4590 20102 4590 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
rlabel metal2 21482 3740 21482 3740 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
rlabel metal1 23161 4114 23161 4114 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 27600 2958 27600 2958 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.ccff_tail
rlabel metal2 19090 4114 19090 4114 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
rlabel metal2 20838 4012 20838 4012 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
rlabel metal2 24426 4250 24426 4250 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 17250 3502 17250 3502 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
rlabel metal1 19182 6086 19182 6086 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
rlabel metal1 23828 3570 23828 3570 0 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 9798 2414 9798 2414 0 ccff_head
rlabel metal1 47242 23120 47242 23120 0 ccff_head_1
rlabel metal2 41354 1622 41354 1622 0 ccff_tail
rlabel metal2 1610 24728 1610 24728 0 ccff_tail_0
rlabel metal1 3266 2346 3266 2346 0 chanx_left_in[0]
rlabel metal1 1472 5678 1472 5678 0 chanx_left_in[10]
rlabel metal1 1472 6290 1472 6290 0 chanx_left_in[11]
rlabel metal1 1932 6766 1932 6766 0 chanx_left_in[12]
rlabel metal1 1472 6698 1472 6698 0 chanx_left_in[13]
rlabel metal1 1472 7378 1472 7378 0 chanx_left_in[14]
rlabel metal1 1472 7854 1472 7854 0 chanx_left_in[15]
rlabel metal1 1518 8398 1518 8398 0 chanx_left_in[16]
rlabel metal1 1794 8942 1794 8942 0 chanx_left_in[17]
rlabel metal1 1518 8874 1518 8874 0 chanx_left_in[18]
rlabel metal1 1472 9554 1472 9554 0 chanx_left_in[19]
rlabel metal1 1840 2346 1840 2346 0 chanx_left_in[1]
rlabel metal1 1472 10030 1472 10030 0 chanx_left_in[20]
rlabel metal1 2346 10676 2346 10676 0 chanx_left_in[21]
rlabel metal1 1472 10642 1472 10642 0 chanx_left_in[22]
rlabel metal2 1610 11033 1610 11033 0 chanx_left_in[23]
rlabel metal1 2530 11696 2530 11696 0 chanx_left_in[24]
rlabel metal1 1472 12206 1472 12206 0 chanx_left_in[25]
rlabel metal1 1426 11730 1426 11730 0 chanx_left_in[26]
rlabel metal2 1242 12699 1242 12699 0 chanx_left_in[27]
rlabel metal1 1518 12886 1518 12886 0 chanx_left_in[28]
rlabel metal2 3542 13651 3542 13651 0 chanx_left_in[29]
rlabel metal1 2208 2414 2208 2414 0 chanx_left_in[2]
rlabel metal1 1472 3026 1472 3026 0 chanx_left_in[3]
rlabel metal1 1472 3502 1472 3502 0 chanx_left_in[4]
rlabel metal1 1840 4114 1840 4114 0 chanx_left_in[5]
rlabel metal1 1564 4182 1564 4182 0 chanx_left_in[6]
rlabel metal1 1472 4590 1472 4590 0 chanx_left_in[7]
rlabel metal1 1472 5134 1472 5134 0 chanx_left_in[8]
rlabel metal1 2576 5678 2576 5678 0 chanx_left_in[9]
rlabel metal2 2806 13549 2806 13549 0 chanx_left_out[0]
rlabel metal3 1694 17884 1694 17884 0 chanx_left_out[10]
rlabel metal2 2898 18853 2898 18853 0 chanx_left_out[11]
rlabel metal3 1004 18700 1004 18700 0 chanx_left_out[12]
rlabel metal3 1004 19108 1004 19108 0 chanx_left_out[13]
rlabel metal3 1694 19516 1694 19516 0 chanx_left_out[14]
rlabel metal2 3358 20689 3358 20689 0 chanx_left_out[15]
rlabel via2 3910 20349 3910 20349 0 chanx_left_out[16]
rlabel metal3 1004 20740 1004 20740 0 chanx_left_out[17]
rlabel metal2 2852 21148 2852 21148 0 chanx_left_out[18]
rlabel metal3 1694 21556 1694 21556 0 chanx_left_out[19]
rlabel metal3 1004 14212 1004 14212 0 chanx_left_out[1]
rlabel metal2 3910 22015 3910 22015 0 chanx_left_out[20]
rlabel metal3 1579 22372 1579 22372 0 chanx_left_out[21]
rlabel metal2 4002 22457 4002 22457 0 chanx_left_out[22]
rlabel metal1 5934 20978 5934 20978 0 chanx_left_out[23]
rlabel metal1 6900 21454 6900 21454 0 chanx_left_out[24]
rlabel metal1 4140 18802 4140 18802 0 chanx_left_out[25]
rlabel metal1 6256 19890 6256 19890 0 chanx_left_out[26]
rlabel metal1 6854 20366 6854 20366 0 chanx_left_out[27]
rlabel metal2 4094 25075 4094 25075 0 chanx_left_out[28]
rlabel metal2 3450 25347 3450 25347 0 chanx_left_out[29]
rlabel metal3 1004 14620 1004 14620 0 chanx_left_out[2]
rlabel metal3 1004 15028 1004 15028 0 chanx_left_out[3]
rlabel metal3 1004 15436 1004 15436 0 chanx_left_out[4]
rlabel metal3 1004 15844 1004 15844 0 chanx_left_out[5]
rlabel metal3 1004 16252 1004 16252 0 chanx_left_out[6]
rlabel metal3 1004 16660 1004 16660 0 chanx_left_out[7]
rlabel metal3 958 17068 958 17068 0 chanx_left_out[8]
rlabel metal2 2806 17833 2806 17833 0 chanx_left_out[9]
rlabel metal1 48438 13906 48438 13906 0 chanx_right_in_0[0]
rlabel metal2 49082 18003 49082 18003 0 chanx_right_in_0[10]
rlabel metal1 49128 18734 49128 18734 0 chanx_right_in_0[11]
rlabel metal2 48806 18479 48806 18479 0 chanx_right_in_0[12]
rlabel metal2 49174 19159 49174 19159 0 chanx_right_in_0[13]
rlabel metal1 49266 19754 49266 19754 0 chanx_right_in_0[14]
rlabel metal2 49082 20111 49082 20111 0 chanx_right_in_0[15]
rlabel metal2 48806 20111 48806 20111 0 chanx_right_in_0[16]
rlabel metal2 49082 20757 49082 20757 0 chanx_right_in_0[17]
rlabel metal2 49082 21267 49082 21267 0 chanx_right_in_0[18]
rlabel metal1 49312 23494 49312 23494 0 chanx_right_in_0[19]
rlabel metal2 49174 14025 49174 14025 0 chanx_right_in_0[1]
rlabel metal2 48806 21743 48806 21743 0 chanx_right_in_0[20]
rlabel metal2 49082 22423 49082 22423 0 chanx_right_in_0[21]
rlabel metal1 49220 23086 49220 23086 0 chanx_right_in_0[22]
rlabel via2 48346 23069 48346 23069 0 chanx_right_in_0[23]
rlabel metal2 47886 23273 47886 23273 0 chanx_right_in_0[24]
rlabel metal1 46322 23664 46322 23664 0 chanx_right_in_0[25]
rlabel metal1 47748 22610 47748 22610 0 chanx_right_in_0[26]
rlabel metal3 48446 24684 48446 24684 0 chanx_right_in_0[27]
rlabel metal1 46966 22610 46966 22610 0 chanx_right_in_0[28]
rlabel metal1 48392 24242 48392 24242 0 chanx_right_in_0[29]
rlabel metal2 49174 14433 49174 14433 0 chanx_right_in_0[2]
rlabel metal2 49082 14943 49082 14943 0 chanx_right_in_0[3]
rlabel metal2 49358 15385 49358 15385 0 chanx_right_in_0[4]
rlabel metal2 49082 15895 49082 15895 0 chanx_right_in_0[5]
rlabel metal1 49128 16558 49128 16558 0 chanx_right_in_0[6]
rlabel metal1 49220 17170 49220 17170 0 chanx_right_in_0[7]
rlabel metal2 48806 16847 48806 16847 0 chanx_right_in_0[8]
rlabel metal2 49082 17493 49082 17493 0 chanx_right_in_0[9]
rlabel metal2 46690 2737 46690 2737 0 chanx_right_out_0[0]
rlabel metal1 49312 4658 49312 4658 0 chanx_right_out_0[10]
rlabel metal2 49174 5593 49174 5593 0 chanx_right_out_0[11]
rlabel metal3 49596 6324 49596 6324 0 chanx_right_out_0[12]
rlabel metal1 49312 5746 49312 5746 0 chanx_right_out_0[13]
rlabel metal1 49220 6358 49220 6358 0 chanx_right_out_0[14]
rlabel metal3 49734 7548 49734 7548 0 chanx_right_out_0[15]
rlabel metal2 46874 8177 46874 8177 0 chanx_right_out_0[16]
rlabel metal1 49266 7446 49266 7446 0 chanx_right_out_0[17]
rlabel metal1 49220 7922 49220 7922 0 chanx_right_out_0[18]
rlabel metal2 49174 8857 49174 8857 0 chanx_right_out_0[19]
rlabel metal2 46782 2397 46782 2397 0 chanx_right_out_0[1]
rlabel metal3 48814 9588 48814 9588 0 chanx_right_out_0[20]
rlabel metal1 49220 9010 49220 9010 0 chanx_right_out_0[21]
rlabel metal1 49266 9622 49266 9622 0 chanx_right_out_0[22]
rlabel metal2 49174 10455 49174 10455 0 chanx_right_out_0[23]
rlabel metal1 49220 10710 49220 10710 0 chanx_right_out_0[24]
rlabel metal2 49174 11407 49174 11407 0 chanx_right_out_0[25]
rlabel metal2 49174 11917 49174 11917 0 chanx_right_out_0[26]
rlabel metal3 49734 12444 49734 12444 0 chanx_right_out_0[27]
rlabel via2 49174 12835 49174 12835 0 chanx_right_out_0[28]
rlabel metal3 49734 13260 49734 13260 0 chanx_right_out_0[29]
rlabel metal3 49412 2244 49412 2244 0 chanx_right_out_0[2]
rlabel metal2 46874 2805 46874 2805 0 chanx_right_out_0[3]
rlabel metal3 49504 3060 49504 3060 0 chanx_right_out_0[4]
rlabel metal2 49174 2975 49174 2975 0 chanx_right_out_0[5]
rlabel metal1 49220 3094 49220 3094 0 chanx_right_out_0[6]
rlabel metal2 49174 3927 49174 3927 0 chanx_right_out_0[7]
rlabel metal1 47610 5134 47610 5134 0 chanx_right_out_0[8]
rlabel metal1 49266 4114 49266 4114 0 chanx_right_out_0[9]
rlabel metal2 21574 24422 21574 24422 0 chany_top_in[0]
rlabel metal1 29256 23698 29256 23698 0 chany_top_in[10]
rlabel metal2 28658 25306 28658 25306 0 chany_top_in[11]
rlabel metal2 32154 23732 32154 23732 0 chany_top_in[12]
rlabel metal1 33442 24174 33442 24174 0 chany_top_in[13]
rlabel metal1 40204 24174 40204 24174 0 chany_top_in[14]
rlabel metal1 33488 23086 33488 23086 0 chany_top_in[15]
rlabel metal1 40204 23698 40204 23698 0 chany_top_in[16]
rlabel metal3 36708 21012 36708 21012 0 chany_top_in[17]
rlabel metal1 42182 22202 42182 22202 0 chany_top_in[18]
rlabel metal2 40710 24327 40710 24327 0 chany_top_in[19]
rlabel metal1 16974 22440 16974 22440 0 chany_top_in[1]
rlabel metal2 41814 23868 41814 23868 0 chany_top_in[20]
rlabel metal2 42182 23868 42182 23868 0 chany_top_in[21]
rlabel metal2 42642 23477 42642 23477 0 chany_top_in[22]
rlabel metal2 43930 23409 43930 23409 0 chany_top_in[23]
rlabel via2 45402 23715 45402 23715 0 chany_top_in[24]
rlabel metal2 41998 23392 41998 23392 0 chany_top_in[25]
rlabel metal1 44114 22644 44114 22644 0 chany_top_in[26]
rlabel metal2 42826 22950 42826 22950 0 chany_top_in[27]
rlabel metal1 44758 22576 44758 22576 0 chany_top_in[28]
rlabel metal1 43470 22576 43470 22576 0 chany_top_in[29]
rlabel metal1 15226 23290 15226 23290 0 chany_top_in[2]
rlabel metal1 22034 23732 22034 23732 0 chany_top_in[3]
rlabel metal1 24472 20910 24472 20910 0 chany_top_in[4]
rlabel metal2 24794 25442 24794 25442 0 chany_top_in[5]
rlabel metal2 25254 24803 25254 24803 0 chany_top_in[6]
rlabel metal1 27094 24174 27094 24174 0 chany_top_in[7]
rlabel metal1 28014 23732 28014 23732 0 chany_top_in[8]
rlabel metal1 28750 24208 28750 24208 0 chany_top_in[9]
rlabel metal2 2254 24252 2254 24252 0 chany_top_out[0]
rlabel metal1 8464 24242 8464 24242 0 chany_top_out[10]
rlabel metal1 9246 23766 9246 23766 0 chany_top_out[11]
rlabel metal2 10258 24429 10258 24429 0 chany_top_out[12]
rlabel metal2 10718 25041 10718 25041 0 chany_top_out[13]
rlabel metal2 11270 24728 11270 24728 0 chany_top_out[14]
rlabel metal1 10994 24276 10994 24276 0 chany_top_out[15]
rlabel metal1 12834 22542 12834 22542 0 chany_top_out[16]
rlabel metal2 13386 24735 13386 24735 0 chany_top_out[17]
rlabel metal1 13708 24242 13708 24242 0 chany_top_out[18]
rlabel metal1 14398 23766 14398 23766 0 chany_top_out[19]
rlabel metal1 3634 23290 3634 23290 0 chany_top_out[1]
rlabel metal1 15272 22542 15272 22542 0 chany_top_out[20]
rlabel metal2 15778 24728 15778 24728 0 chany_top_out[21]
rlabel metal2 16146 25041 16146 25041 0 chany_top_out[22]
rlabel metal1 17618 22134 17618 22134 0 chany_top_out[23]
rlabel metal1 16928 24242 16928 24242 0 chany_top_out[24]
rlabel metal1 18262 23766 18262 23766 0 chany_top_out[25]
rlabel metal1 19458 22134 19458 22134 0 chany_top_out[26]
rlabel metal1 18722 24276 18722 24276 0 chany_top_out[27]
rlabel metal1 21114 24208 21114 24208 0 chany_top_out[28]
rlabel metal2 20930 25272 20930 25272 0 chany_top_out[29]
rlabel metal1 3404 24242 3404 24242 0 chany_top_out[2]
rlabel metal1 4094 23766 4094 23766 0 chany_top_out[3]
rlabel metal1 5060 22542 5060 22542 0 chany_top_out[4]
rlabel metal2 5474 24966 5474 24966 0 chany_top_out[5]
rlabel metal2 6118 24728 6118 24728 0 chany_top_out[6]
rlabel metal1 5842 24276 5842 24276 0 chany_top_out[7]
rlabel metal1 7820 22542 7820 22542 0 chany_top_out[8]
rlabel metal2 7866 24735 7866 24735 0 chany_top_out[9]
rlabel metal1 18492 17646 18492 17646 0 clknet_0_prog_clk
rlabel metal1 13662 8500 13662 8500 0 clknet_4_0_0_prog_clk
rlabel metal2 34086 11730 34086 11730 0 clknet_4_10_0_prog_clk
rlabel metal1 36478 13226 36478 13226 0 clknet_4_11_0_prog_clk
rlabel metal1 32338 17204 32338 17204 0 clknet_4_12_0_prog_clk
rlabel metal2 32614 19040 32614 19040 0 clknet_4_13_0_prog_clk
rlabel metal1 38962 17068 38962 17068 0 clknet_4_14_0_prog_clk
rlabel metal1 35328 20978 35328 20978 0 clknet_4_15_0_prog_clk
rlabel metal1 10626 12274 10626 12274 0 clknet_4_1_0_prog_clk
rlabel metal2 21022 3230 21022 3230 0 clknet_4_2_0_prog_clk
rlabel metal2 21482 11424 21482 11424 0 clknet_4_3_0_prog_clk
rlabel metal2 18630 16592 18630 16592 0 clknet_4_4_0_prog_clk
rlabel metal1 19366 17714 19366 17714 0 clknet_4_5_0_prog_clk
rlabel metal1 19734 20502 19734 20502 0 clknet_4_6_0_prog_clk
rlabel metal2 21206 20400 21206 20400 0 clknet_4_7_0_prog_clk
rlabel metal2 28842 5712 28842 5712 0 clknet_4_8_0_prog_clk
rlabel metal1 29394 13974 29394 13974 0 clknet_4_9_0_prog_clk
rlabel metal2 11730 1622 11730 1622 0 gfpga_pad_io_soc_dir[0]
rlabel metal2 13846 1622 13846 1622 0 gfpga_pad_io_soc_dir[1]
rlabel metal1 17342 2414 17342 2414 0 gfpga_pad_io_soc_dir[2]
rlabel metal2 18078 823 18078 823 0 gfpga_pad_io_soc_dir[3]
rlabel metal1 29118 2414 29118 2414 0 gfpga_pad_io_soc_in[0]
rlabel metal1 30912 2414 30912 2414 0 gfpga_pad_io_soc_in[1]
rlabel metal2 33166 1989 33166 1989 0 gfpga_pad_io_soc_in[2]
rlabel metal1 35144 2414 35144 2414 0 gfpga_pad_io_soc_in[3]
rlabel metal2 20194 1622 20194 1622 0 gfpga_pad_io_soc_out[0]
rlabel metal2 22310 1622 22310 1622 0 gfpga_pad_io_soc_out[1]
rlabel metal2 24426 1622 24426 1622 0 gfpga_pad_io_soc_out[2]
rlabel metal2 26542 1622 26542 1622 0 gfpga_pad_io_soc_out[3]
rlabel metal2 37122 1520 37122 1520 0 isol_n
rlabel metal1 10396 2618 10396 2618 0 net1
rlabel metal1 4393 8466 4393 8466 0 net10
rlabel metal1 35144 16150 35144 16150 0 net100
rlabel metal1 36616 16422 36616 16422 0 net101
rlabel metal1 33672 13294 33672 13294 0 net102
rlabel metal1 35236 19278 35236 19278 0 net103
rlabel metal1 46552 24038 46552 24038 0 net104
rlabel metal1 42090 24106 42090 24106 0 net105
rlabel metal1 47472 24038 47472 24038 0 net106
rlabel metal2 42458 22848 42458 22848 0 net107
rlabel metal2 42182 22678 42182 22678 0 net108
rlabel metal1 44206 22950 44206 22950 0 net109
rlabel metal1 2530 8840 2530 8840 0 net11
rlabel metal1 40526 20570 40526 20570 0 net110
rlabel metal1 39514 2414 39514 2414 0 net111
rlabel metal2 10902 19108 10902 19108 0 net112
rlabel metal1 1794 13328 1794 13328 0 net113
rlabel metal1 3910 18700 3910 18700 0 net114
rlabel metal1 3542 19414 3542 19414 0 net115
rlabel metal2 1794 20026 1794 20026 0 net116
rlabel metal1 1886 20434 1886 20434 0 net117
rlabel metal1 1794 20944 1794 20944 0 net118
rlabel metal1 3542 21454 3542 21454 0 net119
rlabel metal2 14214 9316 14214 9316 0 net12
rlabel metal1 3864 20434 3864 20434 0 net120
rlabel metal1 2277 21998 2277 21998 0 net121
rlabel metal1 15456 19278 15456 19278 0 net122
rlabel metal1 7406 22202 7406 22202 0 net123
rlabel metal1 1794 13940 1794 13940 0 net124
rlabel metal2 4094 21828 4094 21828 0 net125
rlabel metal1 4278 20910 4278 20910 0 net126
rlabel metal1 6256 21998 6256 21998 0 net127
rlabel metal1 5934 20842 5934 20842 0 net128
rlabel metal2 5290 21012 5290 21012 0 net129
rlabel via2 1794 9435 1794 9435 0 net13
rlabel metal1 4554 18734 4554 18734 0 net130
rlabel metal1 6026 19754 6026 19754 0 net131
rlabel metal1 5382 20366 5382 20366 0 net132
rlabel metal1 7176 21386 7176 21386 0 net133
rlabel metal1 7912 22474 7912 22474 0 net134
rlabel metal1 5796 14382 5796 14382 0 net135
rlabel metal2 6578 15164 6578 15164 0 net136
rlabel metal2 10442 15028 10442 15028 0 net137
rlabel metal1 1794 16116 1794 16116 0 net138
rlabel metal2 11086 16796 11086 16796 0 net139
rlabel metal1 19435 2618 19435 2618 0 net14
rlabel metal2 8326 17884 8326 17884 0 net140
rlabel metal2 8602 17136 8602 17136 0 net141
rlabel metal1 3542 18190 3542 18190 0 net142
rlabel metal2 45862 3842 45862 3842 0 net143
rlabel metal1 47472 4590 47472 4590 0 net144
rlabel metal1 47886 5202 47886 5202 0 net145
rlabel metal2 40066 7276 40066 7276 0 net146
rlabel metal1 47840 5678 47840 5678 0 net147
rlabel metal1 47748 6290 47748 6290 0 net148
rlabel metal1 47932 6766 47932 6766 0 net149
rlabel metal2 1886 10438 1886 10438 0 net15
rlabel metal1 42918 9928 42918 9928 0 net150
rlabel metal2 47058 8534 47058 8534 0 net151
rlabel metal2 46966 9180 46966 9180 0 net152
rlabel metal2 46046 9214 46046 9214 0 net153
rlabel metal2 39790 3774 39790 3774 0 net154
rlabel metal2 45770 10540 45770 10540 0 net155
rlabel metal2 43746 10268 43746 10268 0 net156
rlabel metal2 43378 10846 43378 10846 0 net157
rlabel metal2 46322 10812 46322 10812 0 net158
rlabel metal1 47472 10642 47472 10642 0 net159
rlabel metal1 4715 10506 4715 10506 0 net16
rlabel metal1 47518 11118 47518 11118 0 net160
rlabel metal1 46966 11730 46966 11730 0 net161
rlabel metal1 46966 12614 46966 12614 0 net162
rlabel metal1 47518 12818 47518 12818 0 net163
rlabel metal1 47242 13294 47242 13294 0 net164
rlabel metal2 45678 3332 45678 3332 0 net165
rlabel metal2 45770 4318 45770 4318 0 net166
rlabel metal1 46138 3570 46138 3570 0 net167
rlabel metal2 47242 3570 47242 3570 0 net168
rlabel metal2 47334 4454 47334 4454 0 net169
rlabel metal2 1794 10880 1794 10880 0 net17
rlabel metal2 47150 4828 47150 4828 0 net170
rlabel metal1 42090 7208 42090 7208 0 net171
rlabel metal1 47518 4114 47518 4114 0 net172
rlabel metal1 4094 19924 4094 19924 0 net173
rlabel metal2 7406 24225 7406 24225 0 net174
rlabel metal1 8142 23766 8142 23766 0 net175
rlabel metal1 10856 22610 10856 22610 0 net176
rlabel metal1 12696 21114 12696 21114 0 net177
rlabel metal2 12374 22644 12374 22644 0 net178
rlabel metal1 12972 21658 12972 21658 0 net179
rlabel metal2 1794 11169 1794 11169 0 net18
rlabel metal1 13754 22610 13754 22610 0 net180
rlabel metal1 13248 23086 13248 23086 0 net181
rlabel metal1 14260 22066 14260 22066 0 net182
rlabel metal1 13110 23630 13110 23630 0 net183
rlabel metal1 3864 22950 3864 22950 0 net184
rlabel metal1 15870 22610 15870 22610 0 net185
rlabel metal1 18676 19686 18676 19686 0 net186
rlabel metal1 15134 23664 15134 23664 0 net187
rlabel metal1 17618 21964 17618 21964 0 net188
rlabel metal1 19320 21318 19320 21318 0 net189
rlabel metal1 3266 11866 3266 11866 0 net19
rlabel metal1 17158 23766 17158 23766 0 net190
rlabel metal2 19458 23018 19458 23018 0 net191
rlabel metal1 18492 24174 18492 24174 0 net192
rlabel metal2 21298 24004 21298 24004 0 net193
rlabel metal1 20286 24106 20286 24106 0 net194
rlabel metal1 2300 24174 2300 24174 0 net195
rlabel metal1 4094 18258 4094 18258 0 net196
rlabel metal2 4830 23052 4830 23052 0 net197
rlabel metal2 4738 23494 4738 23494 0 net198
rlabel metal1 4278 18394 4278 18394 0 net199
rlabel metal1 43677 23154 43677 23154 0 net2
rlabel metal1 3680 12274 3680 12274 0 net20
rlabel metal2 2162 23970 2162 23970 0 net200
rlabel metal2 7498 23324 7498 23324 0 net201
rlabel metal1 6394 23086 6394 23086 0 net202
rlabel metal1 12420 2414 12420 2414 0 net203
rlabel metal1 15180 2414 15180 2414 0 net204
rlabel metal1 17158 2414 17158 2414 0 net205
rlabel metal1 18354 2958 18354 2958 0 net206
rlabel metal1 20102 2482 20102 2482 0 net207
rlabel metal1 21528 2890 21528 2890 0 net208
rlabel metal2 23230 3026 23230 3026 0 net209
rlabel metal1 4347 11594 4347 11594 0 net21
rlabel metal1 26818 2822 26818 2822 0 net210
rlabel metal1 16698 17646 16698 17646 0 net211
rlabel metal2 23690 13770 23690 13770 0 net212
rlabel metal1 28244 20978 28244 20978 0 net213
rlabel metal1 18860 14042 18860 14042 0 net214
rlabel metal1 24288 19890 24288 19890 0 net215
rlabel metal1 19412 13226 19412 13226 0 net216
rlabel metal1 31234 14246 31234 14246 0 net217
rlabel metal2 30958 7990 30958 7990 0 net218
rlabel metal2 32706 10370 32706 10370 0 net219
rlabel metal1 6854 16626 6854 16626 0 net22
rlabel metal2 33902 15232 33902 15232 0 net220
rlabel metal1 28934 13158 28934 13158 0 net221
rlabel metal2 29762 9282 29762 9282 0 net222
rlabel metal2 31418 7616 31418 7616 0 net223
rlabel metal1 33856 14042 33856 14042 0 net224
rlabel metal1 29164 8874 29164 8874 0 net225
rlabel metal1 26910 11866 26910 11866 0 net226
rlabel metal1 32798 7786 32798 7786 0 net227
rlabel metal1 29394 19482 29394 19482 0 net228
rlabel metal1 31372 15130 31372 15130 0 net229
rlabel metal2 9890 14858 9890 14858 0 net23
rlabel metal1 36386 17306 36386 17306 0 net230
rlabel metal1 36202 15130 36202 15130 0 net231
rlabel metal1 35742 13294 35742 13294 0 net232
rlabel metal1 31280 10778 31280 10778 0 net233
rlabel metal1 33028 21658 33028 21658 0 net234
rlabel metal1 25116 13294 25116 13294 0 net235
rlabel metal1 23966 11050 23966 11050 0 net236
rlabel metal1 20332 11050 20332 11050 0 net237
rlabel metal1 25024 10642 25024 10642 0 net238
rlabel metal2 22678 10880 22678 10880 0 net239
rlabel metal1 19458 18666 19458 18666 0 net24
rlabel metal1 18400 12750 18400 12750 0 net240
rlabel metal1 18446 8398 18446 8398 0 net241
rlabel metal1 19596 10098 19596 10098 0 net242
rlabel metal2 22402 8330 22402 8330 0 net243
rlabel metal1 30912 18258 30912 18258 0 net244
rlabel metal1 12926 13158 12926 13158 0 net245
rlabel metal1 13984 18394 13984 18394 0 net246
rlabel metal1 12788 18734 12788 18734 0 net247
rlabel metal1 10258 18394 10258 18394 0 net248
rlabel metal1 13892 20570 13892 20570 0 net249
rlabel metal2 4370 2448 4370 2448 0 net25
rlabel metal2 9890 21386 9890 21386 0 net250
rlabel metal1 15916 20570 15916 20570 0 net251
rlabel metal1 35512 18802 35512 18802 0 net252
rlabel metal1 40204 20434 40204 20434 0 net253
rlabel metal2 18722 9826 18722 9826 0 net254
rlabel metal1 16698 10710 16698 10710 0 net255
rlabel metal1 11316 13906 11316 13906 0 net256
rlabel metal1 16284 14314 16284 14314 0 net257
rlabel metal1 22402 12240 22402 12240 0 net258
rlabel metal1 21712 12750 21712 12750 0 net259
rlabel metal1 2116 2890 2116 2890 0 net26
rlabel metal1 17158 20774 17158 20774 0 net260
rlabel metal1 17710 24038 17710 24038 0 net261
rlabel metal1 23184 17578 23184 17578 0 net262
rlabel metal2 1886 4284 1886 4284 0 net27
rlabel metal1 2530 4012 2530 4012 0 net28
rlabel metal1 4370 3944 4370 3944 0 net29
rlabel metal1 4991 2618 4991 2618 0 net3
rlabel metal1 1794 4488 1794 4488 0 net30
rlabel metal1 6854 5134 6854 5134 0 net31
rlabel metal1 4738 5882 4738 5882 0 net32
rlabel metal2 48438 14552 48438 14552 0 net33
rlabel metal1 14306 13736 14306 13736 0 net34
rlabel metal4 14444 14892 14444 14892 0 net35
rlabel metal2 48438 18428 48438 18428 0 net36
rlabel metal2 15088 19754 15088 19754 0 net37
rlabel via2 16790 20349 16790 20349 0 net38
rlabel metal1 19412 15674 19412 15674 0 net39
rlabel metal1 1794 5576 1794 5576 0 net4
rlabel metal2 48438 19822 48438 19822 0 net40
rlabel metal1 12742 20774 12742 20774 0 net41
rlabel metal1 12788 20570 12788 20570 0 net42
rlabel via2 15410 19363 15410 19363 0 net43
rlabel metal1 14950 13226 14950 13226 0 net44
rlabel metal1 45034 20910 45034 20910 0 net45
rlabel metal1 48944 22406 48944 22406 0 net46
rlabel metal1 18768 15674 18768 15674 0 net47
rlabel metal2 13754 20808 13754 20808 0 net48
rlabel metal1 44666 21862 44666 21862 0 net49
rlabel metal1 16146 12818 16146 12818 0 net5
rlabel metal1 45770 23494 45770 23494 0 net50
rlabel metal1 48484 22746 48484 22746 0 net51
rlabel metal2 40434 22304 40434 22304 0 net52
rlabel metal2 44206 23154 44206 23154 0 net53
rlabel via2 48806 24157 48806 24157 0 net54
rlabel metal1 17388 14450 17388 14450 0 net55
rlabel metal2 38502 15725 38502 15725 0 net56
rlabel metal1 48944 15674 48944 15674 0 net57
rlabel metal1 21620 13158 21620 13158 0 net58
rlabel metal1 12926 15096 12926 15096 0 net59
rlabel metal2 2346 7854 2346 7854 0 net6
rlabel metal1 15318 18122 15318 18122 0 net60
rlabel metal2 48438 17442 48438 17442 0 net61
rlabel metal1 34454 16728 34454 16728 0 net62
rlabel metal1 32568 14450 32568 14450 0 net63
rlabel metal2 29302 20468 29302 20468 0 net64
rlabel metal1 29670 19720 29670 19720 0 net65
rlabel metal2 32338 24480 32338 24480 0 net66
rlabel metal2 32982 23936 32982 23936 0 net67
rlabel metal2 34362 21182 34362 21182 0 net68
rlabel metal1 33166 19754 33166 19754 0 net69
rlabel metal1 38778 7752 38778 7752 0 net7
rlabel metal1 35144 19822 35144 19822 0 net70
rlabel metal2 34822 21471 34822 21471 0 net71
rlabel metal2 33626 21403 33626 21403 0 net72
rlabel via2 40986 24259 40986 24259 0 net73
rlabel metal2 11362 21709 11362 21709 0 net74
rlabel metal3 35420 19516 35420 19516 0 net75
rlabel metal2 40434 24344 40434 24344 0 net76
rlabel metal2 42826 24344 42826 24344 0 net77
rlabel metal2 44298 24310 44298 24310 0 net78
rlabel via2 45218 23579 45218 23579 0 net79
rlabel metal1 19044 14994 19044 14994 0 net8
rlabel metal2 32430 21267 32430 21267 0 net80
rlabel metal1 34408 19822 34408 19822 0 net81
rlabel via2 42642 22491 42642 22491 0 net82
rlabel metal2 44574 23715 44574 23715 0 net83
rlabel metal1 43056 22406 43056 22406 0 net84
rlabel metal2 17066 24208 17066 24208 0 net85
rlabel metal1 27094 19686 27094 19686 0 net86
rlabel metal1 32706 15538 32706 15538 0 net87
rlabel metal2 33304 17714 33304 17714 0 net88
rlabel metal2 36754 16847 36754 16847 0 net89
rlabel metal1 1794 7752 1794 7752 0 net9
rlabel metal1 32269 18190 32269 18190 0 net90
rlabel metal1 28796 21590 28796 21590 0 net91
rlabel metal2 27830 17204 27830 17204 0 net92
rlabel metal1 28290 2618 28290 2618 0 net93
rlabel metal1 27554 2550 27554 2550 0 net94
rlabel metal1 32936 2618 32936 2618 0 net95
rlabel metal1 34776 2618 34776 2618 0 net96
rlabel metal2 37766 2822 37766 2822 0 net97
rlabel metal1 44528 23018 44528 23018 0 net98
rlabel metal1 39882 2550 39882 2550 0 net99
rlabel metal2 37306 5134 37306 5134 0 prog_clk
rlabel metal1 42412 24174 42412 24174 0 prog_reset_top_in
rlabel metal1 43378 2278 43378 2278 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 45310 3434 45310 3434 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 47702 2336 47702 2336 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 46598 4488 46598 4488 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 32890 12716 32890 12716 0 sb_1__0_.mem_left_track_1.ccff_head
rlabel metal1 24196 17306 24196 17306 0 sb_1__0_.mem_left_track_1.ccff_tail
rlabel metal1 31510 21454 31510 21454 0 sb_1__0_.mem_left_track_1.mem_out\[0\]
rlabel metal1 26404 16218 26404 16218 0 sb_1__0_.mem_left_track_1.mem_out\[1\]
rlabel metal2 21390 14994 21390 14994 0 sb_1__0_.mem_left_track_11.ccff_head
rlabel metal1 20424 18190 20424 18190 0 sb_1__0_.mem_left_track_11.ccff_tail
rlabel via1 26450 19299 26450 19299 0 sb_1__0_.mem_left_track_11.mem_out\[0\]
rlabel metal2 22770 17442 22770 17442 0 sb_1__0_.mem_left_track_11.mem_out\[1\]
rlabel metal1 18860 20774 18860 20774 0 sb_1__0_.mem_left_track_13.ccff_tail
rlabel metal1 21666 18054 21666 18054 0 sb_1__0_.mem_left_track_13.mem_out\[0\]
rlabel metal1 18209 21114 18209 21114 0 sb_1__0_.mem_left_track_13.mem_out\[1\]
rlabel metal1 18262 21454 18262 21454 0 sb_1__0_.mem_left_track_21.ccff_tail
rlabel metal1 25806 22066 25806 22066 0 sb_1__0_.mem_left_track_21.mem_out\[0\]
rlabel metal1 18952 19890 18952 19890 0 sb_1__0_.mem_left_track_21.mem_out\[1\]
rlabel metal1 21390 19244 21390 19244 0 sb_1__0_.mem_left_track_29.ccff_tail
rlabel metal1 24334 20366 24334 20366 0 sb_1__0_.mem_left_track_29.mem_out\[0\]
rlabel metal1 25714 20366 25714 20366 0 sb_1__0_.mem_left_track_29.mem_out\[1\]
rlabel metal1 18860 20570 18860 20570 0 sb_1__0_.mem_left_track_3.ccff_tail
rlabel metal1 25254 18836 25254 18836 0 sb_1__0_.mem_left_track_3.mem_out\[0\]
rlabel metal1 20976 18802 20976 18802 0 sb_1__0_.mem_left_track_3.mem_out\[1\]
rlabel metal2 27370 16966 27370 16966 0 sb_1__0_.mem_left_track_37.ccff_tail
rlabel metal1 32223 19890 32223 19890 0 sb_1__0_.mem_left_track_37.mem_out\[0\]
rlabel metal2 25898 16575 25898 16575 0 sb_1__0_.mem_left_track_37.mem_out\[1\]
rlabel metal1 26312 23154 26312 23154 0 sb_1__0_.mem_left_track_45.ccff_tail
rlabel metal1 32890 22508 32890 22508 0 sb_1__0_.mem_left_track_45.mem_out\[0\]
rlabel metal2 28934 21760 28934 21760 0 sb_1__0_.mem_left_track_45.mem_out\[1\]
rlabel metal2 18906 16286 18906 16286 0 sb_1__0_.mem_left_track_5.ccff_tail
rlabel via1 20562 17595 20562 17595 0 sb_1__0_.mem_left_track_5.mem_out\[0\]
rlabel metal1 18906 13804 18906 13804 0 sb_1__0_.mem_left_track_5.mem_out\[1\]
rlabel metal1 27462 22984 27462 22984 0 sb_1__0_.mem_left_track_53.mem_out\[0\]
rlabel metal2 23230 21947 23230 21947 0 sb_1__0_.mem_left_track_53.mem_out\[1\]
rlabel metal1 25806 15538 25806 15538 0 sb_1__0_.mem_left_track_7.mem_out\[0\]
rlabel metal1 23828 14042 23828 14042 0 sb_1__0_.mem_left_track_7.mem_out\[1\]
rlabel metal3 17572 21964 17572 21964 0 sb_1__0_.mem_right_track_0.ccff_head
rlabel metal2 32614 16456 32614 16456 0 sb_1__0_.mem_right_track_0.ccff_tail
rlabel metal2 32890 13668 32890 13668 0 sb_1__0_.mem_right_track_0.mem_out\[0\]
rlabel metal2 30774 16286 30774 16286 0 sb_1__0_.mem_right_track_0.mem_out\[1\]
rlabel metal1 37352 11866 37352 11866 0 sb_1__0_.mem_right_track_10.ccff_head
rlabel metal2 36662 10948 36662 10948 0 sb_1__0_.mem_right_track_10.ccff_tail
rlabel metal1 33442 15538 33442 15538 0 sb_1__0_.mem_right_track_10.mem_out\[0\]
rlabel metal1 35236 13362 35236 13362 0 sb_1__0_.mem_right_track_10.mem_out\[1\]
rlabel metal1 32798 13192 32798 13192 0 sb_1__0_.mem_right_track_12.ccff_tail
rlabel metal1 32384 16014 32384 16014 0 sb_1__0_.mem_right_track_12.mem_out\[0\]
rlabel metal2 31786 13668 31786 13668 0 sb_1__0_.mem_right_track_12.mem_out\[1\]
rlabel metal1 36754 15674 36754 15674 0 sb_1__0_.mem_right_track_2.ccff_tail
rlabel metal1 33626 21454 33626 21454 0 sb_1__0_.mem_right_track_2.mem_out\[0\]
rlabel metal1 35788 15538 35788 15538 0 sb_1__0_.mem_right_track_2.mem_out\[1\]
rlabel metal1 34086 11730 34086 11730 0 sb_1__0_.mem_right_track_20.ccff_tail
rlabel metal2 32798 14144 32798 14144 0 sb_1__0_.mem_right_track_20.mem_out\[0\]
rlabel metal2 29762 15504 29762 15504 0 sb_1__0_.mem_right_track_20.mem_out\[1\]
rlabel metal1 33166 9520 33166 9520 0 sb_1__0_.mem_right_track_28.ccff_tail
rlabel metal1 30636 14926 30636 14926 0 sb_1__0_.mem_right_track_28.mem_out\[0\]
rlabel metal1 30774 10642 30774 10642 0 sb_1__0_.mem_right_track_28.mem_out\[1\]
rlabel metal2 34086 8806 34086 8806 0 sb_1__0_.mem_right_track_36.ccff_tail
rlabel metal1 32706 14484 32706 14484 0 sb_1__0_.mem_right_track_36.mem_out\[0\]
rlabel metal1 32430 8398 32430 8398 0 sb_1__0_.mem_right_track_36.mem_out\[1\]
rlabel metal1 37996 13158 37996 13158 0 sb_1__0_.mem_right_track_4.ccff_tail
rlabel metal1 36846 16592 36846 16592 0 sb_1__0_.mem_right_track_4.mem_out\[0\]
rlabel metal2 36662 15844 36662 15844 0 sb_1__0_.mem_right_track_4.mem_out\[1\]
rlabel metal1 29762 9622 29762 9622 0 sb_1__0_.mem_right_track_44.ccff_tail
rlabel metal1 29900 16626 29900 16626 0 sb_1__0_.mem_right_track_44.mem_out\[0\]
rlabel metal1 29256 9418 29256 9418 0 sb_1__0_.mem_right_track_52.mem_out\[0\]
rlabel metal1 36156 12750 36156 12750 0 sb_1__0_.mem_right_track_6.mem_out\[0\]
rlabel metal1 36754 12070 36754 12070 0 sb_1__0_.mem_right_track_6.mem_out\[1\]
rlabel metal2 31786 23324 31786 23324 0 sb_1__0_.mem_top_track_0.ccff_tail
rlabel via2 43562 23035 43562 23035 0 sb_1__0_.mem_top_track_0.mem_out\[0\]
rlabel metal2 32614 22559 32614 22559 0 sb_1__0_.mem_top_track_0.mem_out\[1\]
rlabel metal1 37720 20502 37720 20502 0 sb_1__0_.mem_top_track_10.ccff_head
rlabel metal1 34040 18666 34040 18666 0 sb_1__0_.mem_top_track_10.ccff_tail
rlabel metal1 35650 19278 35650 19278 0 sb_1__0_.mem_top_track_10.mem_out\[0\]
rlabel metal2 33902 17646 33902 17646 0 sb_1__0_.mem_top_track_10.mem_out\[1\]
rlabel metal1 39330 18666 39330 18666 0 sb_1__0_.mem_top_track_12.ccff_tail
rlabel via2 38226 19261 38226 19261 0 sb_1__0_.mem_top_track_12.mem_out\[0\]
rlabel metal2 38318 17646 38318 17646 0 sb_1__0_.mem_top_track_12.mem_out\[1\]
rlabel metal1 38548 16150 38548 16150 0 sb_1__0_.mem_top_track_14.ccff_tail
rlabel metal2 40618 17850 40618 17850 0 sb_1__0_.mem_top_track_14.mem_out\[0\]
rlabel metal1 38180 16490 38180 16490 0 sb_1__0_.mem_top_track_14.mem_out\[1\]
rlabel metal2 37858 16932 37858 16932 0 sb_1__0_.mem_top_track_16.ccff_tail
rlabel metal1 40296 16014 40296 16014 0 sb_1__0_.mem_top_track_16.mem_out\[0\]
rlabel metal1 37720 15402 37720 15402 0 sb_1__0_.mem_top_track_16.mem_out\[1\]
rlabel metal1 33442 14926 33442 14926 0 sb_1__0_.mem_top_track_18.ccff_tail
rlabel metal1 38410 14790 38410 14790 0 sb_1__0_.mem_top_track_18.mem_out\[0\]
rlabel metal1 38916 14586 38916 14586 0 sb_1__0_.mem_top_track_18.mem_out\[1\]
rlabel metal1 34178 23494 34178 23494 0 sb_1__0_.mem_top_track_2.ccff_tail
rlabel metal2 35558 23851 35558 23851 0 sb_1__0_.mem_top_track_2.mem_out\[0\]
rlabel metal1 36478 22474 36478 22474 0 sb_1__0_.mem_top_track_2.mem_out\[1\]
rlabel metal2 25162 15538 25162 15538 0 sb_1__0_.mem_top_track_20.ccff_tail
rlabel metal1 25760 13362 25760 13362 0 sb_1__0_.mem_top_track_20.mem_out\[0\]
rlabel metal1 25346 12954 25346 12954 0 sb_1__0_.mem_top_track_22.ccff_tail
rlabel metal1 26588 14042 26588 14042 0 sb_1__0_.mem_top_track_22.mem_out\[0\]
rlabel metal1 24702 11186 24702 11186 0 sb_1__0_.mem_top_track_24.ccff_tail
rlabel metal1 27094 15946 27094 15946 0 sb_1__0_.mem_top_track_24.mem_out\[0\]
rlabel metal1 23276 13362 23276 13362 0 sb_1__0_.mem_top_track_26.ccff_tail
rlabel metal1 27324 15538 27324 15538 0 sb_1__0_.mem_top_track_26.mem_out\[0\]
rlabel metal1 21390 10506 21390 10506 0 sb_1__0_.mem_top_track_28.ccff_tail
rlabel metal1 23276 9486 23276 9486 0 sb_1__0_.mem_top_track_28.mem_out\[0\]
rlabel metal1 19872 7786 19872 7786 0 sb_1__0_.mem_top_track_30.ccff_tail
rlabel metal1 21045 8398 21045 8398 0 sb_1__0_.mem_top_track_30.mem_out\[0\]
rlabel metal1 19596 9622 19596 9622 0 sb_1__0_.mem_top_track_32.ccff_tail
rlabel metal1 19780 8874 19780 8874 0 sb_1__0_.mem_top_track_32.mem_out\[0\]
rlabel metal1 20424 12750 20424 12750 0 sb_1__0_.mem_top_track_34.ccff_tail
rlabel metal1 20700 9962 20700 9962 0 sb_1__0_.mem_top_track_34.mem_out\[0\]
rlabel metal1 21252 12750 21252 12750 0 sb_1__0_.mem_top_track_36.ccff_tail
rlabel metal1 21942 11560 21942 11560 0 sb_1__0_.mem_top_track_36.mem_out\[0\]
rlabel metal1 33442 20978 33442 20978 0 sb_1__0_.mem_top_track_4.ccff_tail
rlabel metal1 35236 20842 35236 20842 0 sb_1__0_.mem_top_track_4.mem_out\[0\]
rlabel metal1 31096 18190 31096 18190 0 sb_1__0_.mem_top_track_4.mem_out\[1\]
rlabel metal1 13340 13838 13340 13838 0 sb_1__0_.mem_top_track_40.ccff_tail
rlabel metal1 14122 10574 14122 10574 0 sb_1__0_.mem_top_track_40.mem_out\[0\]
rlabel metal1 14950 18190 14950 18190 0 sb_1__0_.mem_top_track_42.ccff_tail
rlabel metal1 14720 14042 14720 14042 0 sb_1__0_.mem_top_track_42.mem_out\[0\]
rlabel metal1 13294 18802 13294 18802 0 sb_1__0_.mem_top_track_44.ccff_tail
rlabel metal2 16054 19074 16054 19074 0 sb_1__0_.mem_top_track_44.mem_out\[0\]
rlabel metal1 12328 17850 12328 17850 0 sb_1__0_.mem_top_track_46.ccff_tail
rlabel metal1 12466 14960 12466 14960 0 sb_1__0_.mem_top_track_46.mem_out\[0\]
rlabel metal2 14858 20978 14858 20978 0 sb_1__0_.mem_top_track_48.ccff_tail
rlabel metal1 13846 19958 13846 19958 0 sb_1__0_.mem_top_track_48.mem_out\[0\]
rlabel metal1 15318 22202 15318 22202 0 sb_1__0_.mem_top_track_50.ccff_tail
rlabel metal2 16330 20060 16330 20060 0 sb_1__0_.mem_top_track_50.mem_out\[0\]
rlabel metal1 19550 22746 19550 22746 0 sb_1__0_.mem_top_track_58.mem_out\[0\]
rlabel via1 37575 22202 37575 22202 0 sb_1__0_.mem_top_track_6.ccff_tail
rlabel metal2 34224 20774 34224 20774 0 sb_1__0_.mem_top_track_6.mem_out\[0\]
rlabel metal1 39238 22508 39238 22508 0 sb_1__0_.mem_top_track_6.mem_out\[1\]
rlabel metal1 38226 21454 38226 21454 0 sb_1__0_.mem_top_track_8.mem_out\[0\]
rlabel metal1 37628 20978 37628 20978 0 sb_1__0_.mem_top_track_8.mem_out\[1\]
rlabel metal1 14536 16558 14536 16558 0 sb_1__0_.mux_left_track_1.out
rlabel metal1 26910 18258 26910 18258 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 26772 18394 26772 18394 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 22724 12954 22724 12954 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 23552 16150 23552 16150 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 25070 17884 25070 17884 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 24012 16218 24012 16218 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 21574 17816 21574 17816 0 sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 8372 16218 8372 16218 0 sb_1__0_.mux_left_track_11.out
rlabel metal1 22908 18258 22908 18258 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24150 18394 24150 18394 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 20930 14076 20930 14076 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20378 15062 20378 15062 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 20286 18394 20286 18394 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 19550 16694 19550 16694 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 16606 18394 16606 18394 0 sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 10580 19686 10580 19686 0 sb_1__0_.mux_left_track_13.out
rlabel metal2 21942 21760 21942 21760 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 24794 21658 24794 21658 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20608 15674 20608 15674 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 21482 21896 21482 21896 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 17618 18938 17618 18938 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 14858 19958 14858 19958 0 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 9706 21216 9706 21216 0 sb_1__0_.mux_left_track_21.out
rlabel metal1 26680 23290 26680 23290 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24242 21862 24242 21862 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 21114 19312 21114 19312 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 17894 23154 17894 23154 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 18262 20026 18262 20026 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 12650 21352 12650 21352 0 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 13616 17510 13616 17510 0 sb_1__0_.mux_left_track_29.out
rlabel metal1 26174 21012 26174 21012 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 26818 20434 26818 20434 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23966 15130 23966 15130 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 23874 20264 23874 20264 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 21758 18632 21758 18632 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 13754 17578 13754 17578 0 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 9982 20672 9982 20672 0 sb_1__0_.mux_left_track_3.out
rlabel metal1 26864 21862 26864 21862 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22218 18836 22218 18836 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19780 18938 19780 18938 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17020 17850 17020 17850 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 15916 20026 15916 20026 0 sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 16974 15334 16974 15334 0 sb_1__0_.mux_left_track_37.out
rlabel metal2 32154 19006 32154 19006 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 29256 18258 29256 18258 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23828 16626 23828 16626 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 23368 13498 23368 13498 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 19826 15793 19826 15793 0 sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 8602 18734 8602 18734 0 sb_1__0_.mux_left_track_45.out
rlabel metal1 32108 22406 32108 22406 0 sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 28014 21862 28014 21862 0 sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 28106 21658 28106 21658 0 sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20286 23154 20286 23154 0 sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 10534 19482 10534 19482 0 sb_1__0_.mux_left_track_5.out
rlabel metal1 24058 20026 24058 20026 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24242 18122 24242 18122 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17894 15980 17894 15980 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 18400 14042 18400 14042 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 16192 16218 16192 16218 0 sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 12742 20876 12742 20876 0 sb_1__0_.mux_left_track_53.out
rlabel metal1 28152 21930 28152 21930 0 sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 25990 21352 25990 21352 0 sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20746 20910 20746 20910 0 sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 13754 20944 13754 20944 0 sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 8878 19822 8878 19822 0 sb_1__0_.mux_left_track_7.out
rlabel metal1 25392 15470 25392 15470 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24104 15402 24104 15402 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19826 11594 19826 11594 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 23138 15368 23138 15368 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 20010 13498 20010 13498 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 19918 16320 19918 16320 0 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 39330 14110 39330 14110 0 sb_1__0_.mux_right_track_0.out
rlabel metal1 31050 17102 31050 17102 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 33350 13600 33350 13600 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 30866 14382 30866 14382 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 33994 16592 33994 16592 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 32246 14280 32246 14280 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 39514 14416 39514 14416 0 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 45540 11186 45540 11186 0 sb_1__0_.mux_right_track_10.out
rlabel metal2 35006 14518 35006 14518 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 34684 13906 34684 13906 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 34638 9146 34638 9146 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 32338 8704 32338 8704 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 37720 12716 37720 12716 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 36524 10778 36524 10778 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 40618 11118 40618 11118 0 sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 40802 11934 40802 11934 0 sb_1__0_.mux_right_track_12.out
rlabel metal1 33902 14382 33902 14382 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 33580 14382 33580 14382 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 32269 10574 32269 10574 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 37536 14076 37536 14076 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 32660 10778 32660 10778 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 40986 12274 40986 12274 0 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 45862 14348 45862 14348 0 sb_1__0_.mux_right_track_2.out
rlabel metal2 36386 20366 36386 20366 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 34316 18054 34316 18054 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 33994 14756 33994 14756 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel via2 35926 19499 35926 19499 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 35144 14790 35144 14790 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 40480 14994 40480 14994 0 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 43010 10030 43010 10030 0 sb_1__0_.mux_right_track_20.out
rlabel metal2 31050 18224 31050 18224 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 30958 16592 30958 16592 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 28888 13294 28888 13294 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 33994 11628 33994 11628 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 32430 13464 32430 13464 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 38410 11084 38410 11084 0 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 39606 8670 39606 8670 0 sb_1__0_.mux_right_track_28.out
rlabel metal1 30084 13158 30084 13158 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 29992 13294 29992 13294 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 25714 9214 25714 9214 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 30314 13430 30314 13430 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 31326 10030 31326 10030 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 37858 8976 37858 8976 0 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 40158 7888 40158 7888 0 sb_1__0_.mux_right_track_36.out
rlabel metal2 31464 14892 31464 14892 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 32430 11866 32430 11866 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 35190 8874 35190 8874 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 33534 8024 33534 8024 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 39146 8500 39146 8500 0 sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 46138 12988 46138 12988 0 sb_1__0_.mux_right_track_4.out
rlabel metal2 36478 19414 36478 19414 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 36294 16932 36294 16932 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 33350 11288 33350 11288 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 37812 13974 37812 13974 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 35742 13838 35742 13838 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 41538 13668 41538 13668 0 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 40250 7480 40250 7480 0 sb_1__0_.mux_right_track_44.out
rlabel metal2 32430 15147 32430 15147 0 sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 28612 9146 28612 9146 0 sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 36064 8466 36064 8466 0 sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 43746 6289 43746 6289 0 sb_1__0_.mux_right_track_52.out
rlabel metal2 32798 13158 32798 13158 0 sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 32154 12818 32154 12818 0 sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 33902 12682 33902 12682 0 sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 43493 12070 43493 12070 0 sb_1__0_.mux_right_track_6.out
rlabel metal1 36156 14926 36156 14926 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 36248 14994 36248 14994 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 36432 12682 36432 12682 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 32430 7718 32430 7718 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 36616 14858 36616 14858 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 38686 11968 38686 11968 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 41630 12274 41630 12274 0 sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 25070 24650 25070 24650 0 sb_1__0_.mux_top_track_0.out
rlabel metal1 34914 21896 34914 21896 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 37582 23834 37582 23834 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23368 19958 23368 19958 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 28474 20111 28474 20111 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 35926 23341 35926 23341 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 29256 21114 29256 21114 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 29762 23426 29762 23426 0 sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 21689 21522 21689 21522 0 sb_1__0_.mux_top_track_10.out
rlabel metal1 35190 19482 35190 19482 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 40158 19618 40158 19618 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 31970 19380 31970 19380 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 31878 17544 31878 17544 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 28934 19095 28934 19095 0 sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 29348 22066 29348 22066 0 sb_1__0_.mux_top_track_12.out
rlabel metal1 40480 18394 40480 18394 0 sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 39882 18122 39882 18122 0 sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 37352 17034 37352 17034 0 sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 35604 20298 35604 20298 0 sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 19734 21947 19734 21947 0 sb_1__0_.mux_top_track_14.out
rlabel metal1 40480 17714 40480 17714 0 sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 40526 18190 40526 18190 0 sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 34730 16864 34730 16864 0 sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 38042 18649 38042 18649 0 sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 21482 19312 21482 19312 0 sb_1__0_.mux_top_track_16.out
rlabel metal1 40526 16218 40526 16218 0 sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 38962 15878 38962 15878 0 sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 35466 13498 35466 13498 0 sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 29210 18564 29210 18564 0 sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 25714 17782 25714 17782 0 sb_1__0_.mux_top_track_18.out
rlabel metal2 40158 16218 40158 16218 0 sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 39146 15130 39146 15130 0 sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 32154 15130 32154 15130 0 sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 30406 14960 30406 14960 0 sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 21482 23766 21482 23766 0 sb_1__0_.mux_top_track_2.out
rlabel metal1 37858 23766 37858 23766 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 40066 23494 40066 23494 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 33534 20944 33534 20944 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 36340 23562 36340 23562 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 32890 21862 32890 21862 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 31602 23698 31602 23698 0 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 20746 23970 20746 23970 0 sb_1__0_.mux_top_track_20.out
rlabel metal1 26358 17306 26358 17306 0 sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 25070 13498 25070 13498 0 sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24932 17306 24932 17306 0 sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20102 16456 20102 16456 0 sb_1__0_.mux_top_track_22.out
rlabel metal1 23460 15130 23460 15130 0 sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23368 11254 23368 11254 0 sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21206 16456 21206 16456 0 sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 16146 19788 16146 19788 0 sb_1__0_.mux_top_track_24.out
rlabel metal1 26956 15878 26956 15878 0 sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22908 12138 22908 12138 0 sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21942 13396 21942 13396 0 sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 18400 17850 18400 17850 0 sb_1__0_.mux_top_track_26.out
rlabel metal1 22586 13396 22586 13396 0 sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23690 13192 23690 13192 0 sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 20378 14467 20378 14467 0 sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14490 17306 14490 17306 0 sb_1__0_.mux_top_track_28.out
rlabel metal2 22310 10200 22310 10200 0 sb_1__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 15226 14790 15226 14790 0 sb_1__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12742 17850 12742 17850 0 sb_1__0_.mux_top_track_30.out
rlabel metal1 21298 7514 21298 7514 0 sb_1__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18400 14790 18400 14790 0 sb_1__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 12558 17034 12558 17034 0 sb_1__0_.mux_top_track_32.out
rlabel metal1 18262 10234 18262 10234 0 sb_1__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 13478 14484 13478 14484 0 sb_1__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14950 22440 14950 22440 0 sb_1__0_.mux_top_track_34.out
rlabel metal1 19642 10778 19642 10778 0 sb_1__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18998 12614 18998 12614 0 sb_1__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14352 20026 14352 20026 0 sb_1__0_.mux_top_track_36.out
rlabel metal1 23966 12920 23966 12920 0 sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21528 12818 21528 12818 0 sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20746 12920 20746 12920 0 sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 27186 23290 27186 23290 0 sb_1__0_.mux_top_track_4.out
rlabel metal1 34638 20570 34638 20570 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 40066 21760 40066 21760 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 34546 21216 34546 21216 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 30130 19482 30130 19482 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 30866 21097 30866 21097 0 sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 10028 18122 10028 18122 0 sb_1__0_.mux_top_track_40.out
rlabel metal2 12650 13617 12650 13617 0 sb_1__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11730 14586 11730 14586 0 sb_1__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 10166 21658 10166 21658 0 sb_1__0_.mux_top_track_42.out
rlabel metal1 16698 15674 16698 15674 0 sb_1__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13616 18122 13616 18122 0 sb_1__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 2346 23766 2346 23766 0 sb_1__0_.mux_top_track_44.out
rlabel metal2 15594 17952 15594 17952 0 sb_1__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 11454 19686 11454 19686 0 sb_1__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 3634 18292 3634 18292 0 sb_1__0_.mux_top_track_46.out
rlabel metal1 11684 14858 11684 14858 0 sb_1__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 10442 19244 10442 19244 0 sb_1__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 8510 21114 8510 21114 0 sb_1__0_.mux_top_track_48.out
rlabel metal2 16882 19890 16882 19890 0 sb_1__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13754 20332 13754 20332 0 sb_1__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 8418 22916 8418 22916 0 sb_1__0_.mux_top_track_50.out
rlabel metal1 16744 18938 16744 18938 0 sb_1__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 8602 21964 8602 21964 0 sb_1__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 9200 23086 9200 23086 0 sb_1__0_.mux_top_track_58.out
rlabel metal2 16054 22644 16054 22644 0 sb_1__0_.mux_top_track_58.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 15502 20570 15502 20570 0 sb_1__0_.mux_top_track_58.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20838 24310 20838 24310 0 sb_1__0_.mux_top_track_6.out
rlabel metal1 40204 21658 40204 21658 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 40664 22202 40664 22202 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 33672 18870 33672 18870 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 39698 23494 39698 23494 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 36110 23460 36110 23460 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 30038 24174 30038 24174 0 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 31510 22899 31510 22899 0 sb_1__0_.mux_top_track_8.out
rlabel metal1 40112 20978 40112 20978 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 40848 20842 40848 20842 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 33534 19448 33534 19448 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 40158 21114 40158 21114 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 36156 21862 36156 21862 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 36018 23392 36018 23392 0 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 45402 25289 45402 25289 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
rlabel metal1 46414 24106 46414 24106 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
rlabel metal2 46874 25041 46874 25041 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
rlabel metal1 47564 24174 47564 24174 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
rlabel metal1 47978 23698 47978 23698 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
rlabel metal1 48714 23698 48714 23698 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
rlabel metal1 44206 23086 44206 23086 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
rlabel metal1 45034 24174 45034 24174 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
rlabel metal2 1150 2115 1150 2115 0 top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 3266 1299 3266 1299 0 top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 5382 2387 5382 2387 0 top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal2 7498 2166 7498 2166 0 top_width_0_height_0_subtile_3__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 51000 27000
<< end >>
