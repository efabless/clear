* NGSPICE file created from tile.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__sdfrtp_1 abstract view
.subckt sky130_fd_sc_hd__sdfrtp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__sdfrtp_2 abstract view
.subckt sky130_fd_sc_hd__sdfrtp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

.subckt tile VGND VPWR bottom_width_0_height_0_subtile_0__pin_cout_0_ bottom_width_0_height_0_subtile_0__pin_reg_out_0_
+ ccff_head_1 ccff_head_2 ccff_tail ccff_tail_0 chanx_left_in[0] chanx_left_in[10]
+ chanx_left_in[11] chanx_left_in[12] chanx_left_in[13] chanx_left_in[14] chanx_left_in[15]
+ chanx_left_in[16] chanx_left_in[17] chanx_left_in[18] chanx_left_in[19] chanx_left_in[1]
+ chanx_left_in[20] chanx_left_in[21] chanx_left_in[22] chanx_left_in[23] chanx_left_in[24]
+ chanx_left_in[25] chanx_left_in[26] chanx_left_in[27] chanx_left_in[28] chanx_left_in[29]
+ chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6]
+ chanx_left_in[7] chanx_left_in[8] chanx_left_in[9] chanx_left_out[0] chanx_left_out[10]
+ chanx_left_out[11] chanx_left_out[12] chanx_left_out[13] chanx_left_out[14] chanx_left_out[15]
+ chanx_left_out[16] chanx_left_out[17] chanx_left_out[18] chanx_left_out[19] chanx_left_out[1]
+ chanx_left_out[20] chanx_left_out[21] chanx_left_out[22] chanx_left_out[23] chanx_left_out[24]
+ chanx_left_out[25] chanx_left_out[26] chanx_left_out[27] chanx_left_out[28] chanx_left_out[29]
+ chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6]
+ chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chanx_right_in_0[0] chanx_right_in_0[10]
+ chanx_right_in_0[11] chanx_right_in_0[12] chanx_right_in_0[13] chanx_right_in_0[14]
+ chanx_right_in_0[15] chanx_right_in_0[16] chanx_right_in_0[17] chanx_right_in_0[18]
+ chanx_right_in_0[19] chanx_right_in_0[1] chanx_right_in_0[20] chanx_right_in_0[21]
+ chanx_right_in_0[22] chanx_right_in_0[23] chanx_right_in_0[24] chanx_right_in_0[25]
+ chanx_right_in_0[26] chanx_right_in_0[27] chanx_right_in_0[28] chanx_right_in_0[29]
+ chanx_right_in_0[2] chanx_right_in_0[3] chanx_right_in_0[4] chanx_right_in_0[5]
+ chanx_right_in_0[6] chanx_right_in_0[7] chanx_right_in_0[8] chanx_right_in_0[9]
+ chanx_right_out_0[0] chanx_right_out_0[10] chanx_right_out_0[11] chanx_right_out_0[12]
+ chanx_right_out_0[13] chanx_right_out_0[14] chanx_right_out_0[15] chanx_right_out_0[16]
+ chanx_right_out_0[17] chanx_right_out_0[18] chanx_right_out_0[19] chanx_right_out_0[1]
+ chanx_right_out_0[20] chanx_right_out_0[21] chanx_right_out_0[22] chanx_right_out_0[23]
+ chanx_right_out_0[24] chanx_right_out_0[25] chanx_right_out_0[26] chanx_right_out_0[27]
+ chanx_right_out_0[28] chanx_right_out_0[29] chanx_right_out_0[2] chanx_right_out_0[3]
+ chanx_right_out_0[4] chanx_right_out_0[5] chanx_right_out_0[6] chanx_right_out_0[7]
+ chanx_right_out_0[8] chanx_right_out_0[9] chany_bottom_in[0] chany_bottom_in[10]
+ chany_bottom_in[11] chany_bottom_in[12] chany_bottom_in[13] chany_bottom_in[14]
+ chany_bottom_in[15] chany_bottom_in[16] chany_bottom_in[17] chany_bottom_in[18]
+ chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[20] chany_bottom_in[21] chany_bottom_in[22]
+ chany_bottom_in[23] chany_bottom_in[24] chany_bottom_in[25] chany_bottom_in[26]
+ chany_bottom_in[27] chany_bottom_in[28] chany_bottom_in[29] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[20] chany_bottom_out[21] chany_bottom_out[22]
+ chany_bottom_out[23] chany_bottom_out[24] chany_bottom_out[25] chany_bottom_out[26]
+ chany_bottom_out[27] chany_bottom_out[28] chany_bottom_out[29] chany_bottom_out[2]
+ chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6]
+ chany_bottom_out[7] chany_bottom_out[8] chany_bottom_out[9] chany_top_in_0[0] chany_top_in_0[10]
+ chany_top_in_0[11] chany_top_in_0[12] chany_top_in_0[13] chany_top_in_0[14] chany_top_in_0[15]
+ chany_top_in_0[16] chany_top_in_0[17] chany_top_in_0[18] chany_top_in_0[19] chany_top_in_0[1]
+ chany_top_in_0[20] chany_top_in_0[21] chany_top_in_0[22] chany_top_in_0[23] chany_top_in_0[24]
+ chany_top_in_0[25] chany_top_in_0[26] chany_top_in_0[27] chany_top_in_0[28] chany_top_in_0[29]
+ chany_top_in_0[2] chany_top_in_0[3] chany_top_in_0[4] chany_top_in_0[5] chany_top_in_0[6]
+ chany_top_in_0[7] chany_top_in_0[8] chany_top_in_0[9] chany_top_out_0[0] chany_top_out_0[10]
+ chany_top_out_0[11] chany_top_out_0[12] chany_top_out_0[13] chany_top_out_0[14]
+ chany_top_out_0[15] chany_top_out_0[16] chany_top_out_0[17] chany_top_out_0[18]
+ chany_top_out_0[19] chany_top_out_0[1] chany_top_out_0[20] chany_top_out_0[21] chany_top_out_0[22]
+ chany_top_out_0[23] chany_top_out_0[24] chany_top_out_0[25] chany_top_out_0[26]
+ chany_top_out_0[27] chany_top_out_0[28] chany_top_out_0[29] chany_top_out_0[2] chany_top_out_0[3]
+ chany_top_out_0[4] chany_top_out_0[5] chany_top_out_0[6] chany_top_out_0[7] chany_top_out_0[8]
+ chany_top_out_0[9] clk0 prog_clk prog_reset_bottom_in prog_reset_bottom_out prog_reset_left_in
+ prog_reset_right_out prog_reset_top_in prog_reset_top_out reset_bottom_in reset_bottom_out
+ reset_left_out reset_right_in reset_top_in reset_top_out right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
+ right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_ right_width_0_height_0_subtile_0__pin_O_10_
+ right_width_0_height_0_subtile_0__pin_O_11_ right_width_0_height_0_subtile_0__pin_O_12_
+ right_width_0_height_0_subtile_0__pin_O_13_ right_width_0_height_0_subtile_0__pin_O_14_
+ right_width_0_height_0_subtile_0__pin_O_15_ right_width_0_height_0_subtile_0__pin_O_8_
+ right_width_0_height_0_subtile_0__pin_O_9_ sc_in sc_out test_enable_bottom_in test_enable_bottom_out
+ test_enable_left_out test_enable_right_in test_enable_top_in test_enable_top_out
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_ top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_ top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_ top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_ top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
+ top_width_0_height_0_subtile_0__pin_O_0_ top_width_0_height_0_subtile_0__pin_O_1_
+ top_width_0_height_0_subtile_0__pin_O_2_ top_width_0_height_0_subtile_0__pin_O_3_
+ top_width_0_height_0_subtile_0__pin_O_4_ top_width_0_height_0_subtile_0__pin_O_5_
+ top_width_0_height_0_subtile_0__pin_O_6_ top_width_0_height_0_subtile_0__pin_O_7_
+ top_width_0_height_0_subtile_0__pin_cin_0_ top_width_0_height_0_subtile_0__pin_reg_in_0_
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_left_track_37.mux_l1_in_1_ net68 net38 sb_1__1_.mem_left_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_2.mux_l1_in_0_ sb_1__1_.mux_left_track_5.out net22 cbx_1__1_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_16_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net296 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_53_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_53_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_89_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mux_right_ipin_3.mux_l2_in_3_ net315 net116 cby_1__1_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_45_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_363_ net81 VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_294_ net11 VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__clkbuf_2
XFILLER_95_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_right_track_10.mux_l4_in_0_ sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_10_X
+ sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_9_X sb_1__1_.mem_right_track_10.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_right_track_52.mux_l2_in_0_ sb_1__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_right_track_52.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_83_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__1_.mux_right_ipin_14.mux_l1_in_3_ sb_1__1_.mux_bottom_track_29.out net69 cby_1__1_.mem_right_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_13.mux_l2_in_2_ net14 net35 cbx_1__1_.mem_top_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mux_bottom_track_3.mux_l1_in_0_ net122 net108 sb_1__1_.mem_bottom_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_3.mux_l2_in_0_ sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_left_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_86_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_42_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_39_prog_clk
+ sb_1__1_.mem_bottom_track_13.ccff_tail net298 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_21.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
Xsb_1__1_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_19_prog_clk sb_1__1_.mem_left_track_3.mem_out\[0\]
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_3.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_77_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_73 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_346_ net92 VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__clkbuf_2
X_277_ sb_1__1_.mux_left_track_1.out VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ net144 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_37.mux_l2_in_1__387 VGND VGND VPWR VPWR sb_1__1_.mux_left_track_37.mux_l2_in_1__387/HI
+ net387 sky130_fd_sc_hd__conb_1
XFILLER_68_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_top_track_0.mux_l2_in_3_ net403 net4 sb_1__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_91_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_24_prog_clk sb_1__1_.mem_top_track_28.mem_out\[2\]
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_28.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xoutput242 net242 VGND VGND VPWR VPWR chany_top_out_0[12] sky130_fd_sc_hd__buf_12
Xoutput253 net253 VGND VGND VPWR VPWR chany_top_out_0[22] sky130_fd_sc_hd__buf_12
Xoutput231 net231 VGND VGND VPWR VPWR chany_bottom_out[2] sky130_fd_sc_hd__buf_12
Xoutput220 net220 VGND VGND VPWR VPWR chany_bottom_out[1] sky130_fd_sc_hd__buf_12
Xoutput286 net286 VGND VGND VPWR VPWR test_enable_top_out sky130_fd_sc_hd__buf_12
Xoutput264 net264 VGND VGND VPWR VPWR chany_top_out_0[5] sky130_fd_sc_hd__buf_12
Xoutput275 net275 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_10_
+ sky130_fd_sc_hd__buf_12
XFILLER_87_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_11_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_10.mux_l3_in_1_ sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_right_track_10.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_right_track_52.mux_l1_in_1_ net65 net130 sb_1__1_.mem_right_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_left_track_3.mux_l1_in_1_ net48 net93 sb_1__1_.mem_left_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net124 grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_68_.in net134 VGND
+ VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_64_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_329_ net107 VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_41_prog_clk sb_1__1_.mem_bottom_track_5.mem_out\[2\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_5.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_3.mux_l4_in_0_ cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_3.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_56_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_64_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_75_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__1_.mux_right_ipin_14.mux_l3_in_0_ cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_14.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_55_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_8_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_8_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_3_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_4_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_93_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__341
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__341/HI
+ net341 sky130_fd_sc_hd__conb_1
Xcbx_1__1_.mux_top_ipin_7.mux_l1_in_0_ sb_1__1_.mux_left_track_3.out net23 cbx_1__1_.mem_top_ipin_7.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_57_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_ net143 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_72_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_10.mux_l2_in_2_ net13 sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mem_right_track_10.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_8.mux_l2_in_3_ net320 sb_1__1_.mux_bottom_track_53.out cby_1__1_.mem_right_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_25_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_top_track_0.mux_l4_in_0_ sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_9_X
+ sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_8_X sb_1__1_.mem_top_track_0.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_3.mux_l3_in_1_ cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XANTENNA_5 grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_34_.in VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_11_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net295 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_36_prog_clk sb_1__1_.mem_right_track_28.mem_out\[0\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_28.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
Xcby_1__1_.mux_right_ipin_14.mux_l2_in_1_ cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_2_X cby_1__1_.mem_right_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_13.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_3_X cbx_1__1_.mem_top_ipin_13.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_28_prog_clk sb_1__1_.mem_top_track_2.ccff_tail
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_4.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_5_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_28.mux_l2_in_0_ sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_top_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xinput120 chany_top_in_0[7] VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__buf_2
Xinput142 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_ VGND VGND VPWR
+ VPWR net142 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput131 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_ VGND VGND VPWR
+ VPWR net131 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_15_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net296 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_10.mux_l1_in_3_ net75 net132 sb_1__1_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_8.mux_l1_in_4_ net94 net92 cby_1__1_.mem_right_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_39_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_left_track_37.mux_l1_in_0_ net98 net110 sb_1__1_.mem_left_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_top_track_0.mux_l3_in_1_ sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X sb_1__1_.mem_top_track_0.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_16_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net296 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_22_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_22_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_73_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_3.mux_l2_in_2_ net85 sb_1__1_.mux_bottom_track_37.out cby_1__1_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_45_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_362_ sb_1__1_.mux_top_track_10.out VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_293_ sb_1__1_.mux_right_track_28.out VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_91_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_8.mux_l4_in_0_ cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_9_X cby_1__1_.mem_right_ipin_8.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_64_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_14.mux_l1_in_2_ net107 net76 cby_1__1_.mem_right_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_13.mux_l2_in_1_ net4 cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__1_.mem_top_ipin_13.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_8.mux_l2_in_3__304 VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_8.mux_l2_in_3__304/HI
+ net304 sky130_fd_sc_hd__conb_1
XFILLER_55_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_left_track_21.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_21.out sky130_fd_sc_hd__clkbuf_2
XFILLER_23_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_42_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_top_track_28.mux_l1_in_1_ net44 net61 sb_1__1_.mem_top_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_10_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_19_prog_clk sb_1__1_.mem_left_track_1.ccff_tail
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_3.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_12_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net362 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_58_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_345_ sb_1__1_.mux_top_track_44.out VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__clkbuf_2
X_276_ sb_1__1_.mux_left_track_3.out VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_27_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net298 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_top_track_0.mux_l2_in_2_ net21 net24 sb_1__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_91_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_23_prog_clk sb_1__1_.mem_top_track_28.mem_out\[1\]
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_28.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_32_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput210 net210 VGND VGND VPWR VPWR chany_bottom_out[10] sky130_fd_sc_hd__buf_12
Xoutput243 net243 VGND VGND VPWR VPWR chany_top_out_0[13] sky130_fd_sc_hd__buf_12
Xoutput221 net221 VGND VGND VPWR VPWR chany_bottom_out[20] sky130_fd_sc_hd__buf_12
Xoutput232 net232 VGND VGND VPWR VPWR chany_bottom_out[3] sky130_fd_sc_hd__buf_12
Xoutput254 net254 VGND VGND VPWR VPWR chany_top_out_0[23] sky130_fd_sc_hd__buf_12
Xoutput265 net265 VGND VGND VPWR VPWR chany_top_out_0[6] sky130_fd_sc_hd__buf_12
Xoutput276 net276 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_11_
+ sky130_fd_sc_hd__buf_12
XFILLER_58_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput287 net287 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_0_ sky130_fd_sc_hd__buf_12
XFILLER_59_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_11_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_right_track_10.mux_l3_in_0_ sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_right_track_10.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_8.mux_l3_in_1_ cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_8.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net341 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_right_track_52.mux_l1_in_0_ net117 net95 sb_1__1_.mem_right_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_78_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_13.mux_l1_in_2_ net41 net10 cbx_1__1_.mem_top_ipin_13.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_78_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_53.out sky130_fd_sc_hd__buf_4
XFILLER_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__353
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__353/HI
+ net353 sky130_fd_sc_hd__conb_1
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_left_track_3.mux_l1_in_0_ net122 net108 sb_1__1_.mem_left_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_12.out sky130_fd_sc_hd__clkbuf_1
XFILLER_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_328_ net106 VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__clkbuf_2
X_259_ sb_1__1_.mux_left_track_37.out VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_41_prog_clk sb_1__1_.mem_bottom_track_5.mem_out\[1\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_5.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_2.out sky130_fd_sc_hd__clkbuf_1
XFILLER_49_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_0.mux_l1_in_3_ net64 net81 sb_1__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_50_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_4_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_right_track_10.mux_l2_in_1_ sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_right_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_52_110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mux_right_ipin_8.mux_l2_in_2_ net86 cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mem_right_ipin_8.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_47_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_47_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_4_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_3.mux_l3_in_0_ cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X cby_1__1_.mem_right_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XANTENNA_6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net355 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__mux2_4
Xsb_1__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_37_prog_clk sb_1__1_.mem_right_track_20.ccff_tail
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_28.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mux_right_ipin_14.mux_l2_in_0_ cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_1_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput110 chany_top_in_0[25] VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput143 top_width_0_height_0_subtile_0__pin_cin_0_ VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_1
Xinput121 chany_top_in_0[8] VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput132 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_ VGND VGND VPWR
+ VPWR net132 sky130_fd_sc_hd__clkbuf_2
XFILLER_91_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_15_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net296 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_right_track_10.mux_l1_in_2_ net130 net128 sb_1__1_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_8.mux_l1_in_3_ sb_1__1_.mux_bottom_track_29.out net69 cby_1__1_.mem_right_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_top_track_0.mux_l3_in_0_ sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X sb_1__1_.mem_top_track_0.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_89_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mux_right_ipin_3.mux_l2_in_1_ net65 cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__1_.mem_right_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_12_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net295 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_26_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_361_ sb_1__1_.mux_top_track_12.out VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_left_track_21.mux_l2_in_3_ net384 net294 sb_1__1_.mem_left_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
X_292_ net9 VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_17_prog_clk sb_1__1_.mem_left_track_11.mem_out\[2\]
+ net296 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_11.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_40_prog_clk
+ sb_1__1_.mem_bottom_track_13.mem_out\[2\] net298 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_13.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_67_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__1_.mux_right_ipin_14.mux_l1_in_1_ sb_1__1_.mux_bottom_track_11.out net79 cby_1__1_.mem_right_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_13.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__342
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__342/HI
+ net342 sky130_fd_sc_hd__conb_1
XFILLER_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_42_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_42_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_50_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_top_track_28.mux_l1_in_0_ net39 net135 sb_1__1_.mem_top_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_10_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__365
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__365/HI
+ net365 sky130_fd_sc_hd__conb_1
XFILLER_77_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_344_ net90 VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_275_ sb_1__1_.mux_left_track_5.out VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_27_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net298 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_39_prog_clk
+ sb_1__1_.mem_bottom_track_45.mem_out\[1\] net298 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_45.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_78_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_top_track_0.mux_l2_in_1_ sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_49_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_38_prog_clk sb_1__1_.mem_top_track_28.mem_out\[0\]
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_28.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_32_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_right_track_4.mux_l2_in_3__399 VGND VGND VPWR VPWR sb_1__1_.mux_right_track_4.mux_l2_in_3__399/HI
+ net399 sky130_fd_sc_hd__conb_1
Xcby_1__1_.mux_right_ipin_3.mux_l1_in_2_ net106 net75 cby_1__1_.mem_right_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xoutput200 net200 VGND VGND VPWR VPWR chanx_right_out_0[29] sky130_fd_sc_hd__buf_12
Xoutput244 net244 VGND VGND VPWR VPWR chany_top_out_0[14] sky130_fd_sc_hd__buf_12
Xoutput233 net233 VGND VGND VPWR VPWR chany_bottom_out[4] sky130_fd_sc_hd__buf_12
Xoutput211 net211 VGND VGND VPWR VPWR chany_bottom_out[11] sky130_fd_sc_hd__buf_12
Xoutput222 net222 VGND VGND VPWR VPWR chany_bottom_out[21] sky130_fd_sc_hd__buf_12
Xoutput266 net266 VGND VGND VPWR VPWR chany_top_out_0[7] sky130_fd_sc_hd__buf_12
Xoutput255 net255 VGND VGND VPWR VPWR chany_top_out_0[24] sky130_fd_sc_hd__buf_12
Xoutput277 net277 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_12_
+ sky130_fd_sc_hd__buf_12
Xoutput288 net288 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_1_ sky130_fd_sc_hd__buf_12
XFILLER_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net124 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net134 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_68_.in
+ sky130_fd_sc_hd__sdfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mux_right_ipin_8.mux_l3_in_0_ cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_8.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_right_track_12.mux_l2_in_3__394 VGND VGND VPWR VPWR sb_1__1_.mux_right_track_12.mux_l2_in_3__394/HI
+ net394 sky130_fd_sc_hd__conb_1
Xsb_1__1_.mux_right_track_2.mux_l2_in_3_ net395 net32 sb_1__1_.mem_right_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mux_top_ipin_13.mux_l1_in_1_ net51 net20 cbx_1__1_.mem_top_ipin_13.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_48_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_327_ sb_1__1_.mux_bottom_track_21.out VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_258_ net35 VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_2
Xsb_1__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_41_prog_clk sb_1__1_.mem_bottom_track_5.mem_out\[0\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_5.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_6_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_left_track_21.mux_l4_in_0_ sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_left_track_21.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_77_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_75_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_top_track_0.mux_l1_in_2_ net34 net51 sb_1__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_3_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_left_track_11.mux_l2_in_3__382 VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.mux_l2_in_3__382/HI
+ net382 sky130_fd_sc_hd__conb_1
Xsb_1__1_.mux_left_track_37.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_37.out sky130_fd_sc_hd__buf_4
Xsb_1__1_.mux_right_track_10.mux_l2_in_0_ sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_right_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_8.mux_l2_in_1_ cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_2_X cby_1__1_.mem_right_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_14.mux_l2_in_3__312 VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_14.mux_l2_in_3__312/HI
+ net312 sky130_fd_sc_hd__conb_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_52_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_52_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_16_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_16_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_7 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_left_track_21.mux_l3_in_1_ sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_left_track_21.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_94_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_57_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_right_track_2.mux_l4_in_0_ sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_9_X
+ sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_8_X sb_1__1_.mem_right_track_2.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_30_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_17_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net296 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput111 chany_top_in_0[26] VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__clkbuf_4
Xinput100 chany_top_in_0[16] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput133 sc_in VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_1
Xinput144 top_width_0_height_0_subtile_0__pin_reg_in_0_ VGND VGND VPWR VPWR net144
+ sky130_fd_sc_hd__clkbuf_1
Xinput122 chany_top_in_0[9] VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__buf_2
XFILLER_0_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_28.out sky130_fd_sc_hd__clkbuf_1
XFILLER_48_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_15_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net296 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_10.mux_l1_in_1_ net126 net118 sb_1__1_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_8.mux_l1_in_2_ net107 net76 cby_1__1_.mem_right_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net351 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_54_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_29.mux_l2_in_3__374 VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_29.mux_l2_in_3__374/HI
+ net374 sky130_fd_sc_hd__conb_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mux_right_ipin_3.mux_l2_in_0_ cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_12_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net295 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_26_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_360_ net78 VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__clkbuf_2
XFILLER_53_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_291_ net8 VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__clkbuf_2
Xsb_1__1_.mux_left_track_21.mux_l2_in_2_ net288 net85 sb_1__1_.mem_left_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_31_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_31_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_42_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mux_top_ipin_3.mux_l2_in_3_ net299 net56 cbx_1__1_.mem_top_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_30_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_3_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_17_prog_clk sb_1__1_.mem_left_track_11.mem_out\[1\]
+ net296 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_11.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_76_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_39_prog_clk
+ sb_1__1_.mem_bottom_track_13.mem_out\[1\] net298 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_13.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_77_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_36_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_right_track_2.mux_l3_in_1_ sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_6_X sb_1__1_.mem_right_track_2.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_91_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_14.mux_l1_in_0_ sb_1__1_.mux_bottom_track_5.out net82 cby_1__1_.mem_right_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_51_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_11.mux_l2_in_3__309 VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_11.mux_l2_in_3__309/HI
+ net309 sky130_fd_sc_hd__conb_1
XFILLER_23_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_1.out sky130_fd_sc_hd__buf_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_42_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_50_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_343_ net89 VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__clkbuf_2
X_274_ sb_1__1_.mux_left_track_7.out VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__clkbuf_1
XFILLER_5_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_12.mux_l2_in_3_ net405 net26 sb_1__1_.mem_top_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_5_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_38_prog_clk
+ sb_1__1_.mem_bottom_track_45.mem_out\[0\] net298 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_45.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_78_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_top_track_0.mux_l2_in_0_ sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_64_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_24_prog_clk sb_1__1_.mem_top_track_20.ccff_tail
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_28.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput201 net201 VGND VGND VPWR VPWR chanx_right_out_0[2] sky130_fd_sc_hd__buf_12
Xcby_1__1_.mux_right_ipin_3.mux_l1_in_1_ sb_1__1_.mux_bottom_track_7.out net81 cby_1__1_.mem_right_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xoutput223 net223 VGND VGND VPWR VPWR chany_bottom_out[22] sky130_fd_sc_hd__buf_12
Xoutput212 net212 VGND VGND VPWR VPWR chany_bottom_out[12] sky130_fd_sc_hd__buf_12
Xoutput234 net234 VGND VGND VPWR VPWR chany_bottom_out[5] sky130_fd_sc_hd__buf_12
Xoutput245 net245 VGND VGND VPWR VPWR chany_top_out_0[15] sky130_fd_sc_hd__buf_12
Xoutput267 net267 VGND VGND VPWR VPWR chany_top_out_0[8] sky130_fd_sc_hd__buf_12
Xoutput256 net256 VGND VGND VPWR VPWR chany_top_out_0[25] sky130_fd_sc_hd__buf_12
Xoutput289 net289 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_2_ sky130_fd_sc_hd__buf_12
Xoutput278 net278 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_13_
+ sky130_fd_sc_hd__buf_12
XFILLER_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mux_right_track_2.mux_l2_in_2_ net18 net91 sb_1__1_.mem_right_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_13.mux_l1_in_0_ sb_1__1_.mux_left_track_3.out net23 cbx_1__1_.mem_top_ipin_13.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_78_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net359 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_31_prog_clk sb_1__1_.mem_right_track_2.mem_out\[2\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_48_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_326_ net103 VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_257_ net34 VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_41_prog_clk sb_1__1_.mem_bottom_track_3.ccff_tail
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_5.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_6_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_3.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_3.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_87_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_0.mux_l1_in_1_ net53 net139 sb_1__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_50_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_45_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_93_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_309_ net115 VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__clkbuf_2
XFILLER_69_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_8.mux_l2_in_0_ cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_80_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_right_track_2.mux_l1_in_3_ net92 net78 sb_1__1_.mem_right_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_12.mux_l4_in_0_ sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_top_track_12.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_8.mux_l2_in_3_ net304 sb_1__1_.mux_left_track_53.out cbx_1__1_.mem_top_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_88_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_56_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_56_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_29_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_8 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_left_track_21.mux_l3_in_0_ sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_left_track_21.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_94_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mux_top_ipin_3.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_19_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_58_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_15_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net296 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_29.mux_l2_in_3_ net374 net14 sb_1__1_.mem_bottom_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_53_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_
+ sky130_fd_sc_hd__clkbuf_1
Xinput101 chany_top_in_0[17] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__buf_2
Xinput112 chany_top_in_0[27] VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput123 prog_reset_bottom_in VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_16
Xinput134 test_enable_bottom_in VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__buf_12
XFILLER_91_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_16_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail
+ net296 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net337 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__mux2_2
XFILLER_8_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_10.mux_l1_in_0_ net103 net110 sb_1__1_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_8.mux_l1_in_1_ sb_1__1_.mux_bottom_track_11.out net79 cby_1__1_.mem_right_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_79_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_top_track_12.mux_l3_in_1_ sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_top_track_12.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_94_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_1_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_1_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mux_top_ipin_8.mux_l1_in_4_ net34 net32 cbx_1__1_.mem_top_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_50_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_290_ net7 VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_2
Xsb_1__1_.mux_left_track_21.mux_l2_in_1_ net71 sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_left_track_21.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__338
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__338/HI
+ net338 sky130_fd_sc_hd__conb_1
XFILLER_5_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_3.mux_l2_in_2_ net25 sb_1__1_.mux_left_track_37.out cbx_1__1_.mem_top_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_2.mux_l2_in_3__314 VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_2.mux_l2_in_3__314/HI
+ net314 sky130_fd_sc_hd__conb_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_30_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_17_prog_clk sb_1__1_.mem_left_track_11.mem_out\[0\]
+ net296 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_11.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_67_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_40_prog_clk
+ sb_1__1_.mem_bottom_track_13.mem_out\[0\] net298 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_13.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_76_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_2.mux_l3_in_0_ sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X sb_1__1_.mem_right_track_2.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_64_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mux_top_ipin_8.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_9_X cbx_1__1_.mem_top_ipin_8.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_59_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__331
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__331/HI
+ net331 sky130_fd_sc_hd__conb_1
XFILLER_55_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_342_ net88 VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__clkbuf_2
X_273_ net51 VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_22_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_top_track_12.mux_l2_in_2_ net10 net12 sb_1__1_.mem_top_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_39_prog_clk
+ sb_1__1_.mem_bottom_track_37.ccff_tail net296 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_45.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_78_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_29.mux_l4_in_0_ sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_6_X sb_1__1_.mem_bottom_track_29.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_top_track_52.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_52.out sky130_fd_sc_hd__clkbuf_1
XFILLER_20_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mux_right_ipin_3.mux_l1_in_0_ sb_1__1_.mux_bottom_track_1.out net84 cby_1__1_.mem_right_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_6_prog_clk cby_1__1_.mem_right_ipin_1.mem_out\[2\]
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xoutput202 net202 VGND VGND VPWR VPWR chanx_right_out_0[3] sky130_fd_sc_hd__buf_12
Xoutput235 net235 VGND VGND VPWR VPWR chany_bottom_out[6] sky130_fd_sc_hd__buf_12
Xoutput213 net213 VGND VGND VPWR VPWR chany_bottom_out[13] sky130_fd_sc_hd__buf_12
Xoutput224 net224 VGND VGND VPWR VPWR chany_bottom_out[23] sky130_fd_sc_hd__buf_12
Xoutput257 net257 VGND VGND VPWR VPWR chany_top_out_0[26] sky130_fd_sc_hd__buf_12
Xoutput268 net268 VGND VGND VPWR VPWR chany_top_out_0[9] sky130_fd_sc_hd__buf_12
Xoutput246 net246 VGND VGND VPWR VPWR chany_top_out_0[16] sky130_fd_sc_hd__buf_12
Xoutput279 net279 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_14_
+ sky130_fd_sc_hd__buf_12
XFILLER_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_left_track_21.mux_l1_in_2_ net75 net55 sb_1__1_.mem_left_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_67_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_11_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_right_track_2.mux_l2_in_1_ sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_right_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_2_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_19_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_31_prog_clk sb_1__1_.mem_right_track_2.mem_out\[1\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_2.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_73_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__1_.mux_top_ipin_8.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_8.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_73_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_325_ net102 VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_80_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_256_ net62 VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_top_track_0.mux_l1_in_0_ net136 net141 sb_1__1_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_bottom_track_29.mux_l3_in_1_ sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_4_X sb_1__1_.mem_bottom_track_29.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_47_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_78_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_49_prog_clk cby_1__1_.mem_right_ipin_11.mem_out\[2\]
+ net298 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_11.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_59_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_308_ net104 VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_29_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_84_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_2.mux_l1_in_2_ net132 net129 sb_1__1_.mem_right_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_25_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__350
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__350/HI
+ net350 sky130_fd_sc_hd__conb_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_79_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mux_top_ipin_8.mux_l2_in_2_ net26 cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mem_top_ipin_8.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_25_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_25_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_71_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_bottom_track_5.mux_l2_in_3__378 VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_5.mux_l2_in_3__378/HI
+ net378 sky130_fd_sc_hd__conb_1
XANTENNA_9 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_3.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X cbx_1__1_.mem_top_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_66_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_bottom_track_29.mux_l2_in_2_ net31 net9 sb_1__1_.mem_bottom_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_40_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput102 chany_top_in_0[18] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_4
Xinput135 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_ VGND VGND VPWR
+ VPWR net135 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput113 chany_top_in_0[28] VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput124 reset_bottom_in VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__buf_12
XFILLER_91_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__323
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__323/HI
+ net323 sky130_fd_sc_hd__conb_1
Xcby_1__1_.mux_right_ipin_8.mux_l1_in_0_ sb_1__1_.mux_bottom_track_5.out net82 cby_1__1_.mem_right_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_39_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_top_track_12.mux_l3_in_0_ sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_top_track_12.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_39_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_3_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mux_top_ipin_8.mux_l1_in_3_ sb_1__1_.mux_left_track_29.out net9 cbx_1__1_.mem_top_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_35_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_2_prog_clk cby_1__1_.mem_right_ipin_4.mem_out\[2\]
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_4.ccff_tail sky130_fd_sc_hd__dfrtp_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_left_track_21.mux_l2_in_0_ sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_left_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_3.mux_l2_in_1_ net5 cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__1_.mem_top_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_30_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_17_prog_clk sb_1__1_.mem_left_track_11.ccff_head
+ net296 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_11.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net366 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__mux2_2
Xclkbuf_leaf_40_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_40_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_1__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_41_prog_clk
+ sb_1__1_.mem_bottom_track_11.ccff_tail net297 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_13.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_83_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_2_prog_clk cbx_1__1_.mem_top_ipin_12.mem_out\[2\]
+ net295 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_12.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_50_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_341_ sb_1__1_.mux_top_track_52.out VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_272_ sb_1__1_.mux_left_track_11.out VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__clkbuf_2
Xsb_1__1_.mux_top_track_12.mux_l2_in_1_ net86 sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_top_track_12.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_47_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_48_prog_clk cby_1__1_.mem_right_ipin_14.mem_out\[2\]
+ net298 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_14.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_72_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_55_prog_clk cby_1__1_.mem_right_ipin_1.mem_out\[1\]
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_1.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xoutput203 net203 VGND VGND VPWR VPWR chanx_right_out_0[4] sky130_fd_sc_hd__buf_12
Xoutput214 net214 VGND VGND VPWR VPWR chany_bottom_out[14] sky130_fd_sc_hd__buf_12
Xoutput225 net225 VGND VGND VPWR VPWR chany_bottom_out[24] sky130_fd_sc_hd__buf_12
Xoutput258 net258 VGND VGND VPWR VPWR chany_top_out_0[27] sky130_fd_sc_hd__buf_12
Xoutput247 net247 VGND VGND VPWR VPWR chany_top_out_0[17] sky130_fd_sc_hd__buf_12
Xoutput236 net236 VGND VGND VPWR VPWR chany_bottom_out[7] sky130_fd_sc_hd__buf_12
XFILLER_87_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput269 net269 VGND VGND VPWR VPWR prog_reset_bottom_out sky130_fd_sc_hd__buf_12
XFILLER_87_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_left_track_21.mux_l1_in_1_ net41 net115 sb_1__1_.mem_left_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_right_track_2.mux_l2_in_3__395 VGND VGND VPWR VPWR sb_1__1_.mux_right_track_2.mux_l2_in_3__395/HI
+ net395 sky130_fd_sc_hd__conb_1
XFILLER_28_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mux_top_ipin_3.mux_l1_in_2_ net46 net15 cbx_1__1_.mem_top_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_70_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net332 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_82_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_right_track_2.mux_l2_in_0_ sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_right_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_2_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_31_prog_clk sb_1__1_.mem_right_track_2.mem_out\[0\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_2.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mux_top_ipin_8.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_8.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__345
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__345/HI
+ net345 sky130_fd_sc_hd__conb_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__324
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__324/HI
+ net324 sky130_fd_sc_hd__conb_1
X_324_ net101 VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__clkbuf_2
X_255_ sb_1__1_.mux_left_track_45.out VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_80_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_19_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net298 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__1_.mux_right_ipin_10.mux_l2_in_3_ net308 net115 cby_1__1_.mem_right_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_55_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_12.mux_l1_in_2_ net72 net56 sb_1__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_34_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_29.mux_l3_in_0_ sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_bottom_track_29.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_51_prog_clk cby_1__1_.mem_right_ipin_11.mem_out\[1\]
+ net298 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_11.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_75_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_307_ sb_1__1_.mux_right_track_0.out VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__clkbuf_2
Xsb_1__1_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_4.out sky130_fd_sc_hd__clkbuf_1
XFILLER_6_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_30_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_84_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_2.mux_l1_in_1_ net126 net122 sb_1__1_.mem_right_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_92_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_8.mux_l2_in_1_ cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_2_X cbx_1__1_.mem_top_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_20_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_57_prog_clk cby_1__1_.mem_right_ipin_7.mem_out\[2\]
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_7.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_29_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__335
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__335/HI
+ net335 sky130_fd_sc_hd__conb_1
XFILLER_16_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_10.mux_l1_in_4_ sb_1__1_.mux_bottom_track_45.out net90 cby_1__1_.mem_right_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_13_prog_clk cbx_1__1_.mem_top_ipin_15.mem_out\[2\]
+ net298 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__dfrtp_2
Xsb_1__1_.mux_bottom_track_29.mux_l2_in_1_ net275 net44 sb_1__1_.mem_bottom_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_80_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xinput136 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_ VGND VGND VPWR
+ VPWR net136 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput114 chany_top_in_0[29] VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_1
Xinput103 chany_top_in_0[19] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__buf_2
Xinput125 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_ VGND VGND VPWR
+ VPWR net125 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_55 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__1_.mux_right_ipin_10.mux_l4_in_0_ cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_9_X cby_1__1_.mem_right_ipin_10.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_79_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_3_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net295 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mux_top_ipin_8.mux_l1_in_2_ net47 net16 cbx_1__1_.mem_top_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_62_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_55_prog_clk cby_1__1_.mem_right_ipin_4.mem_out\[1\]
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_4.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_85_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mux_top_ipin_3.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net124 grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_77_.in net134 VGND
+ VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_5_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_right_track_36.mux_l2_in_1__398 VGND VGND VPWR VPWR sb_1__1_.mux_right_track_36.mux_l2_in_1__398/HI
+ net398 sky130_fd_sc_hd__conb_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_30_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_5_prog_clk cbx_1__1_.mem_top_ipin_12.mem_out\[1\]
+ net295 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_12.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_15.mux_l2_in_3_ net313 net122 cby_1__1_.mem_right_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_35_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_6.mux_l2_in_3__302 VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_6.mux_l2_in_3__302/HI
+ net302 sky130_fd_sc_hd__conb_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_340_ net86 VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__clkbuf_2
XFILLER_53_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mux_right_ipin_10.mux_l3_in_1_ cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_10.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_41_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_271_ sb_1__1_.mux_left_track_13.out VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__1_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_23_prog_clk cbx_1__1_.mem_top_ipin_1.mem_out\[2\]
+ net296 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_top_track_12.mux_l2_in_0_ sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_top_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_47_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_78_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_58_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_48_prog_clk cby_1__1_.mem_right_ipin_14.mem_out\[1\]
+ net298 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_14.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_54_prog_clk cby_1__1_.mem_right_ipin_1.mem_out\[0\]
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_1.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_64_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput204 net204 VGND VGND VPWR VPWR chanx_right_out_0[5] sky130_fd_sc_hd__buf_12
Xoutput226 net226 VGND VGND VPWR VPWR chany_bottom_out[25] sky130_fd_sc_hd__buf_12
Xoutput215 net215 VGND VGND VPWR VPWR chany_bottom_out[15] sky130_fd_sc_hd__buf_12
Xoutput259 net259 VGND VGND VPWR VPWR chany_top_out_0[28] sky130_fd_sc_hd__buf_12
Xoutput248 net248 VGND VGND VPWR VPWR chany_top_out_0[18] sky130_fd_sc_hd__buf_12
Xoutput237 net237 VGND VGND VPWR VPWR chany_bottom_out[8] sky130_fd_sc_hd__buf_12
XFILLER_87_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_left_track_21.mux_l1_in_0_ net101 net105 sb_1__1_.mem_left_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_95_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_3.mux_l1_in_1_ sb_1__1_.mux_left_track_7.out net21 cbx_1__1_.mem_top_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_19_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_19_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_1__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_31_prog_clk sb_1__1_.mem_right_track_0.ccff_tail
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_2.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_46_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_323_ sb_1__1_.mux_bottom_track_29.out VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__clkbuf_2
X_254_ net60 VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mux_top_ipin_14.mux_l2_in_3_ net420 sb_1__1_.mux_left_track_53.out cbx_1__1_.mem_top_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_50_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_left_track_45.mux_l3_in_0_ sb_1__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_left_track_45.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_19_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net298 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__347
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__347/HI
+ net347 sky130_fd_sc_hd__conb_1
XFILLER_18_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_10.mux_l2_in_2_ net74 cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mem_right_ipin_10.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_top_track_12.mux_l1_in_1_ net40 net42 sb_1__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_36_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__1_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_51_prog_clk cby_1__1_.mem_right_ipin_11.mem_out\[0\]
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_11.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_19_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_15.mux_l4_in_0_ cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.ccff_tail VGND
+ VGND VPWR VPWR cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_86_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_306_ sb_1__1_.mux_right_track_2.out VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_32_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_right_track_2.mux_l1_in_0_ net108 net114 sb_1__1_.mem_right_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_65_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_8.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_8.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_56_prog_clk cby_1__1_.mem_right_ipin_7.mem_out\[1\]
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_7.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_56_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_14.mux_l1_in_4_ net34 net32 cbx_1__1_.mem_top_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_45_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_34_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_34_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_1__1_.mux_left_track_45.mux_l2_in_1_ net388 sb_1__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_left_track_45.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_10.mux_l1_in_3_ net98 net67 cby_1__1_.mem_right_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_29.mux_l2_in_0_ sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_bottom_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_12_prog_clk cbx_1__1_.mem_top_ipin_15.mem_out\[1\]
+ net298 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_15.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_80_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mux_top_ipin_14.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_9_X cbx_1__1_.mem_top_ipin_14.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_15.mux_l3_in_1_ cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_15.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput115 chany_top_in_0[2] VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_4
Xinput104 chany_top_in_0[1] VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__buf_2
Xinput126 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_ VGND VGND VPWR
+ VPWR net126 sky130_fd_sc_hd__clkbuf_1
Xinput137 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_ VGND VGND VPWR
+ VPWR net137 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_6_prog_clk cbx_1__1_.mem_top_ipin_4.mem_out\[2\]
+ net295 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_4.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_67_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_21.out sky130_fd_sc_hd__clkbuf_2
XFILLER_47_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_8.mux_l1_in_1_ sb_1__1_.mux_left_track_11.out net19 cbx_1__1_.mem_top_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
Xcby_1__1_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_55_prog_clk cby_1__1_.mem_right_ipin_4.mem_out\[0\]
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_4.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_89_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_left_track_45.mux_l1_in_2_ net291 net91 sb_1__1_.mem_left_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_41_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_30_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_29.mux_l1_in_1_ net39 net52 sb_1__1_.mem_bottom_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_79_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__1_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_5_prog_clk cbx_1__1_.mem_top_ipin_12.mem_out\[0\]
+ net295 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_12.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_14.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_14.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_15.mux_l2_in_2_ net91 net99 cby_1__1_.mem_right_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_53_prog_clk
+ sb_1__1_.mem_bottom_track_37.mem_out\[1\] net296 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_37.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ net143 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_34_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net348 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__mux2_4
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__1_.mux_right_ipin_10.mux_l3_in_0_ cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_10.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
X_270_ net48 VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__clkbuf_2
XFILLER_22_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_7_prog_clk cbx_1__1_.mem_top_ipin_1.mem_out\[1\]
+ net296 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_1.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_58_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_94_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_48_prog_clk cby_1__1_.mem_right_ipin_14.mem_out\[0\]
+ net298 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_14.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__359
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__359/HI
+ net359 sky130_fd_sc_hd__conb_1
Xsb_1__1_.mux_left_track_7.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.out sky130_fd_sc_hd__buf_4
Xcby_1__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_55_prog_clk cby_1__1_.mem_right_ipin_0.ccff_tail
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_1.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xoutput216 net216 VGND VGND VPWR VPWR chany_bottom_out[16] sky130_fd_sc_hd__buf_12
Xoutput205 net205 VGND VGND VPWR VPWR chanx_right_out_0[6] sky130_fd_sc_hd__buf_12
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput249 net249 VGND VGND VPWR VPWR chany_top_out_0[19] sky130_fd_sc_hd__buf_12
Xoutput227 net227 VGND VGND VPWR VPWR chany_bottom_out[26] sky130_fd_sc_hd__buf_12
Xoutput238 net238 VGND VGND VPWR VPWR chany_bottom_out[9] sky130_fd_sc_hd__buf_12
XFILLER_95_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mux_top_ipin_3.mux_l1_in_0_ sb_1__1_.mux_left_track_1.out net24 cbx_1__1_.mem_top_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_82_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_top_track_28.mux_l2_in_3__408 VGND VGND VPWR VPWR sb_1__1_.mux_top_track_28.mux_l2_in_3__408/HI
+ net408 sky130_fd_sc_hd__conb_1
Xcby_1__1_.mux_right_ipin_4.mux_l2_in_3_ net316 net115 cby_1__1_.mem_right_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_18_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net296 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_59_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_59_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_322_ net99 VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__clkbuf_2
X_253_ net59 VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
Xcbx_1__1_.mux_top_ipin_14.mux_l2_in_2_ net26 cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mem_top_ipin_14.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_26_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net298 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mux_right_ipin_10.mux_l2_in_1_ cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_2_X cby_1__1_.mem_right_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_95_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_top_track_12.mux_l1_in_0_ net139 net141 sb_1__1_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mem_right_ipin_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_50_prog_clk cby_1__1_.mem_right_ipin_10.ccff_tail
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_11.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_86_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net368 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_305_ sb_1__1_.mux_right_track_4.out VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_12_prog_clk cbx_1__1_.mem_top_ipin_7.mem_out\[2\]
+ net298 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_7.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_69_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mux_right_ipin_4.mux_l1_in_4_ sb_1__1_.mux_bottom_track_45.out net90 cby_1__1_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_80_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_4_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_4_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_65_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_top_track_36.mux_l3_in_0_ sb_1__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_top_track_36.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_45_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mux_right_ipin_12.mux_l2_in_3__310 VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_12.mux_l2_in_3__310/HI
+ net310 sky130_fd_sc_hd__conb_1
Xcby_1__1_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_56_prog_clk cby_1__1_.mem_right_ipin_7.mem_out\[0\]
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_7.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_28_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_14.mux_l1_in_3_ sb_1__1_.mux_left_track_29.out net9 cbx_1__1_.mem_top_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_43_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_left_track_45.mux_l2_in_0_ sb_1__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_left_track_45.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_79_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_1__1_.mux_right_ipin_4.mux_l4_in_0_ cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_9_X cby_1__1_.mem_right_ipin_4.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_10.mux_l1_in_2_ sb_1__1_.mux_bottom_track_21.out net73 cby_1__1_.mem_right_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net322 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_9_prog_clk cbx_1__1_.mem_top_ipin_15.mem_out\[0\]
+ net298 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_15.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_80_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mux_right_ipin_15.mux_l3_in_0_ cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_3_X cby_1__1_.mem_right_ipin_15.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput105 chany_top_in_0[20] VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput116 chany_top_in_0[3] VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_4
Xinput127 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_ VGND VGND VPWR
+ VPWR net127 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput138 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_ VGND VGND VPWR
+ VPWR net138 sky130_fd_sc_hd__clkbuf_1
XFILLER_29_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_6_prog_clk cbx_1__1_.mem_top_ipin_4.mem_out\[1\]
+ net295 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_4.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_top_track_36.mux_l2_in_1_ net409 sb_1__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_top_track_36.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_11.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.out sky130_fd_sc_hd__buf_4
XFILLER_67_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mux_top_ipin_8.mux_l1_in_0_ sb_1__1_.mux_left_track_5.out net22 cbx_1__1_.mem_top_ipin_8.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net124 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net134 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_77_.in
+ sky130_fd_sc_hd__sdfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
Xcby_1__1_.mux_right_ipin_9.mux_l2_in_3_ net321 net119 cby_1__1_.mem_right_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mem_right_ipin_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_6_prog_clk cby_1__1_.mem_right_ipin_3.ccff_tail
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_4.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_11_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net295 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_
+ sky130_fd_sc_hd__clkbuf_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xload_slew295 net123 VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__buf_12
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_45.mux_l1_in_1_ net67 net37 sb_1__1_.mem_left_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_13_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_30_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_4.mux_l3_in_1_ cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_4.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_67_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_29.mux_l1_in_0_ net104 net99 sb_1__1_.mem_bottom_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_4_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mem_top_ipin_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_10_prog_clk cbx_1__1_.mem_top_ipin_11.ccff_tail
+ net295 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_12.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xcbx_1__1_.mux_top_ipin_14.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_14.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_15.mux_l2_in_1_ net68 cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__1_.mem_right_ipin_15.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_53_prog_clk
+ sb_1__1_.mem_bottom_track_37.mem_out\[0\] net296 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_37.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_43_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_52_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_right_track_44.mux_l2_in_1__400 VGND VGND VPWR VPWR sb_1__1_.mux_right_track_44.mux_l2_in_1__400/HI
+ net400 sky130_fd_sc_hd__conb_1
XFILLER_58_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_8_prog_clk cbx_1__1_.mem_top_ipin_1.mem_out\[0\]
+ net296 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_1.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xsb_1__1_.mux_top_track_36.mux_l1_in_2_ net8 net20 sb_1__1_.mem_top_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_top_track_6.mux_l2_in_3_ net413 net29 sb_1__1_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_78_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ net424 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net124 net133 net134 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_94_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_58_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f_clk0 clknet_0_clk0 VGND VGND VPWR VPWR clknet_1_0__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
Xcby_1__1_.mem_right_ipin_14.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_52_prog_clk cby_1__1_.mem_right_ipin_13.ccff_tail
+ net298 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_14.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_60_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput217 net217 VGND VGND VPWR VPWR chany_bottom_out[17] sky130_fd_sc_hd__buf_12
Xoutput206 net206 VGND VGND VPWR VPWR chanx_right_out_0[7] sky130_fd_sc_hd__buf_12
Xsb_1__1_.mux_bottom_track_13.mux_l2_in_3__372 VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_13.mux_l2_in_3__372/HI
+ net372 sky130_fd_sc_hd__conb_1
Xoutput239 net239 VGND VGND VPWR VPWR chany_top_out_0[0] sky130_fd_sc_hd__buf_12
Xoutput228 net228 VGND VGND VPWR VPWR chany_bottom_out[27] sky130_fd_sc_hd__buf_12
XFILLER_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__1_.mux_right_ipin_4.mux_l2_in_2_ net74 cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mem_right_ipin_4.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_18_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net298 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_right_track_10.mux_l2_in_3__393 VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.mux_l2_in_3__393/HI
+ net393 sky130_fd_sc_hd__conb_1
XFILLER_73_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_28_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_28_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_321_ net98 VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__clkbuf_2
XFILLER_80_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_252_ net58 VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
Xcby_1__1_.mux_right_ipin_9.mux_l4_in_0_ cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_10.ccff_head
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_89_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__1_.mux_right_ipin_15.mux_l1_in_2_ sb_1__1_.mux_bottom_track_13.out net78 cby_1__1_.mem_right_ipin_15.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_14.mux_l2_in_1_ cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_2_X cbx_1__1_.mem_top_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_89_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_37.out sky130_fd_sc_hd__buf_4
XFILLER_49_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_26_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net298 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__367
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__367/HI
+ net367 sky130_fd_sc_hd__conb_1
Xcby_1__1_.mux_right_ipin_10.mux_l2_in_0_ cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_28_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_top_track_6.mux_l1_in_4_ net16 net89 sb_1__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_11_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_46_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mux_top_ipin_0.mux_l2_in_3__414 VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_0.mux_l2_in_3__414/HI
+ net414 sky130_fd_sc_hd__conb_1
X_304_ sb_1__1_.mux_right_track_6.out VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_9_prog_clk cbx_1__1_.mem_top_ipin_7.mem_out\[1\]
+ net296 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_7.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_37_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__1_.mux_right_ipin_4.mux_l1_in_3_ net98 net67 cby_1__1_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_top_track_6.mux_l4_in_0_ sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_10_X
+ sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_9_X sb_1__1_.mem_top_track_10.ccff_head
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mem_right_ipin_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_56_prog_clk cby_1__1_.mem_right_ipin_6.ccff_tail
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_7.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xcby_1__1_.mux_right_ipin_9.mux_l3_in_1_ cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_9.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__1_.mux_top_ipin_14.mux_l1_in_2_ net47 net16 cbx_1__1_.mem_top_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_43_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_3.mux_l2_in_3__375 VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_3.mux_l2_in_3__375/HI
+ net375 sky130_fd_sc_hd__conb_1
XFILLER_86_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_43_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_43_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_1__1_.mux_right_ipin_10.mux_l1_in_1_ net111 net80 cby_1__1_.mem_right_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__1_.mem_top_ipin_15.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_4_prog_clk cbx_1__1_.mem_top_ipin_14.ccff_tail
+ net295 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_15.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_53_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_86_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput117 chany_top_in_0[4] VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput106 chany_top_in_0[21] VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput139 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_ VGND VGND VPWR
+ VPWR net139 sky130_fd_sc_hd__clkbuf_1
Xinput128 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_ VGND VGND VPWR
+ VPWR net128 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_7_prog_clk cbx_1__1_.mem_top_ipin_4.mem_out\[0\]
+ net295 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_4.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_90 net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_top_track_36.mux_l2_in_0_ sb_1__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_top_track_36.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_79_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_6.mux_l3_in_1_ sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_top_track_6.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_28_prog_clk sb_1__1_.mem_top_track_0.mem_out\[2\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_62_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_right_track_28.mux_l2_in_3_ net397 net14 sb_1__1_.mem_right_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
Xcby_1__1_.mux_right_ipin_9.mux_l2_in_2_ net88 net99 cby_1__1_.mem_right_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_12_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net295 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xload_slew296 net298 VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__buf_12
XFILLER_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_left_track_45.mux_l1_in_0_ net97 net112 sb_1__1_.mem_left_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_38_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_30_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_4.mux_l3_in_0_ cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_4.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_61_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_70_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mux_right_ipin_15.mux_l2_in_0_ cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_67_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_54_prog_clk
+ sb_1__1_.mem_bottom_track_29.ccff_tail net298 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_37.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_90_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_bottom_track_13.mux_l2_in_3_ net372 net26 sb_1__1_.mem_bottom_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_top_track_36.mux_l1_in_1_ net68 net57 sb_1__1_.mem_top_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_21_prog_clk cbx_1__1_.mem_top_ipin_0.ccff_tail
+ net296 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_1.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xsb_1__1_.mux_top_track_6.mux_l2_in_2_ net31 sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mem_top_track_6.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net330 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__mux2_2
Xoutput207 net207 VGND VGND VPWR VPWR chanx_right_out_0[8] sky130_fd_sc_hd__buf_12
Xoutput218 net218 VGND VGND VPWR VPWR chany_bottom_out[18] sky130_fd_sc_hd__buf_12
Xoutput229 net229 VGND VGND VPWR VPWR chany_bottom_out[28] sky130_fd_sc_hd__buf_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_3_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net357 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_right_track_0.mux_l2_in_3__392 VGND VGND VPWR VPWR sb_1__1_.mux_right_track_0.mux_l2_in_3__392/HI
+ net392 sky130_fd_sc_hd__conb_1
XFILLER_90_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__1_.mux_right_ipin_4.mux_l2_in_1_ cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_2_X cby_1__1_.mem_right_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_18_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net298 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_86_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_28.mux_l4_in_0_ sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_6_X sb_1__1_.mem_right_track_28.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_64_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_320_ net97 VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__clkbuf_2
X_251_ sb_1__1_.mux_left_track_53.out VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mux_right_ipin_15.mux_l1_in_1_ sb_1__1_.mux_bottom_track_7.out net81 cby_1__1_.mem_right_ipin_15.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_14.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_14.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_89_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_26_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net298 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_top_track_6.mux_l1_in_3_ net76 net59 sb_1__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_24_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__368
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__368/HI
+ net368 sky130_fd_sc_hd__conb_1
Xcby_1__1_.mux_right_ipin_7.mux_l2_in_3__319 VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_7.mux_l2_in_3__319/HI
+ net319 sky130_fd_sc_hd__conb_1
XFILLER_51_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_75_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_303_ net21 VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_13.mux_l4_in_0_ sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_bottom_track_13.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_9_prog_clk cbx_1__1_.mem_top_ipin_7.mem_out\[0\]
+ net296 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_7.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_77_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mux_right_ipin_4.mux_l1_in_2_ sb_1__1_.mux_bottom_track_21.out net73 cby_1__1_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_65_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_20_prog_clk sb_1__1_.mem_left_track_21.mem_out\[2\]
+ net296 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_21.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_28.mux_l3_in_1_ sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_4_X sb_1__1_.mem_right_track_28.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_9.mux_l3_in_0_ cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_3_X cby_1__1_.mem_right_ipin_9.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_56_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__1_.mux_top_ipin_14.mux_l1_in_1_ sb_1__1_.mux_left_track_11.out net19 cbx_1__1_.mem_top_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_12_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_12_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mux_right_ipin_10.mux_l1_in_0_ sb_1__1_.mux_bottom_track_3.out net83 cby_1__1_.mem_right_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_51_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_21_prog_clk sb_1__1_.mem_left_track_53.mem_out\[1\]
+ net296 VGND VGND VPWR VPWR cbx_1__1_.ccff_head sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net340 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_20.out sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xinput118 chany_top_in_0[5] VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_4
Xinput107 chany_top_in_0[22] VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_4
Xinput129 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_ VGND VGND VPWR
+ VPWR net129 sky130_fd_sc_hd__dlymetal6s2s_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_57_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_13.mux_l3_in_1_ sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_bottom_track_13.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_52_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_80 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__1_.mem_top_ipin_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_54_prog_clk cbx_1__1_.mem_top_ipin_3.ccff_tail
+ net298 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_4.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_91 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_6.mux_l3_in_0_ sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_top_track_6.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_28_prog_clk sb_1__1_.mem_top_track_0.mem_out\[1\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_0.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_47_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_right_track_28.mux_l2_in_2_ net9 net74 sb_1__1_.mem_right_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_62_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_7.mux_l2_in_3__391 VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.mux_l2_in_3__391/HI
+ net391 sky130_fd_sc_hd__conb_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
Xcby_1__1_.mux_right_ipin_9.mux_l2_in_1_ net68 cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__1_.mem_right_ipin_9.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xload_slew297 net298 VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__clkbuf_16
XFILLER_38_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_79_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_88_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_58_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_bottom_track_13.mux_l2_in_2_ net10 net12 sb_1__1_.mem_bottom_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_top_track_36.mux_l1_in_0_ net38 net136 sb_1__1_.mem_top_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_22_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_6.mux_l2_in_1_ sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_89_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_9.mux_l1_in_2_ net106 net75 cby_1__1_.mem_right_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput208 net208 VGND VGND VPWR VPWR chanx_right_out_0[9] sky130_fd_sc_hd__buf_12
Xoutput219 net219 VGND VGND VPWR VPWR chany_bottom_out[19] sky130_fd_sc_hd__buf_12
XFILLER_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_3_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_right_track_52.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_52.out sky130_fd_sc_hd__clkbuf_1
XFILLER_51_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_28_prog_clk sb_1__1_.mem_top_track_6.mem_out\[2\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_10.ccff_head sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mux_right_ipin_4.mux_l2_in_0_ cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_18_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net298 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_2_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_
+ sky130_fd_sc_hd__clkbuf_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__1_.mux_top_ipin_4.mux_l2_in_3_ net300 net55 cbx_1__1_.mem_top_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_86_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_250_ net56 VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_15.mux_l1_in_0_ sb_1__1_.mux_bottom_track_1.out net84 cby_1__1_.mem_right_ipin_15.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_15.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_37_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_37_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_27_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net298 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_5.mux_l2_in_3_ net378 net30 sb_1__1_.mem_bottom_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_68_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_top_track_6.mux_l1_in_2_ net46 net49 sb_1__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_34_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_302_ sb_1__1_.mux_right_track_10.out VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mem_top_ipin_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_13_prog_clk cbx_1__1_.mem_top_ipin_6.ccff_tail
+ net296 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_7.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_77_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__1_.mux_right_ipin_4.mux_l1_in_1_ net111 net80 cby_1__1_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_65_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_20_prog_clk sb_1__1_.mem_left_track_21.mem_out\[1\]
+ net296 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_21.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_45_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_13_prog_clk sb_1__1_.mem_left_track_5.mem_out\[2\]
+ net296 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_5.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mux_top_ipin_4.mux_l1_in_4_ sb_1__1_.mux_left_track_45.out net30 cbx_1__1_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_right_track_28.mux_l3_in_0_ sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_right_track_28.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_68_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_14.mux_l1_in_0_ sb_1__1_.mux_left_track_5.out net22 cbx_1__1_.mem_top_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_14.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_24_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_1.mux_l2_in_3__370 VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_1.mux_l2_in_3__370/HI
+ net370 sky130_fd_sc_hd__conb_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__332
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__332/HI
+ net332 sky130_fd_sc_hd__conb_1
XFILLER_74_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_52_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_52_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcbx_1__1_.mux_top_ipin_4.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_9_X cbx_1__1_.mem_top_ipin_4.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__329
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0__329/HI
+ net329 sky130_fd_sc_hd__conb_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_20_prog_clk sb_1__1_.mem_left_track_53.mem_out\[0\]
+ net296 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_53.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_38_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xinput108 chany_top_in_0[23] VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_4
Xinput119 chany_top_in_0[6] VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__buf_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_57_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_bottom_track_13.mux_l3_in_0_ sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_bottom_track_13.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_81 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_70 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_92 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_5.mux_l4_in_0_ sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_bottom_track_5.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_29_prog_clk sb_1__1_.mem_top_track_0.mem_out\[0\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_0.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_90_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_right_track_28.mux_l2_in_1_ net69 net82 sb_1__1_.mem_right_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_50_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mux_right_ipin_9.mux_l2_in_0_ cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_7_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xload_slew298 net123 VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__clkbuf_16
XFILLER_93_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mux_top_ipin_9.mux_l2_in_3_ net305 net59 cbx_1__1_.mem_top_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_38_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput90 chany_bottom_in[7] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__buf_4
Xsb_1__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_54_prog_clk
+ sb_1__1_.mem_bottom_track_29.mem_out\[2\] net298 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_29.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mux_top_ipin_4.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_4.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_58_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_90_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__340
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__340/HI
+ net340 sky130_fd_sc_hd__conb_1
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_4.mux_l2_in_3__300 VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_4.mux_l2_in_3__300/HI
+ net300 sky130_fd_sc_hd__conb_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_bottom_track_13.mux_l2_in_1_ net279 sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_bottom_track_13.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_58_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_bottom_track_5.mux_l3_in_1_ sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_bottom_track_5.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_top_track_6.mux_l2_in_0_ sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_9.mux_l1_in_1_ sb_1__1_.mux_bottom_track_7.out net81 cby_1__1_.mem_right_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_43_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_top_track_20.mux_l2_in_3_ net407 net25 sb_1__1_.mem_top_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xoutput209 net209 VGND VGND VPWR VPWR chany_bottom_out[0] sky130_fd_sc_hd__buf_12
XFILLER_95_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_36.out sky130_fd_sc_hd__clkbuf_1
XFILLER_63_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_7_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_7_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_1__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_28_prog_clk sb_1__1_.mem_top_track_6.mem_out\[1\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_6.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_19_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net298 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__1_.mux_top_ipin_4.mux_l2_in_2_ net14 cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mem_top_ipin_4.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.out sky130_fd_sc_hd__buf_4
XFILLER_89_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_9.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_10.ccff_head
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_38_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_27_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net298 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_bottom_track_13.mux_l1_in_2_ net281 net56 sb_1__1_.mem_bottom_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_9_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_bottom_track_5.mux_l2_in_2_ net17 net20 sb_1__1_.mem_bottom_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_95_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__327
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__327/HI
+ net327 sky130_fd_sc_hd__conb_1
XFILLER_36_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_6.mux_l1_in_1_ net139 net137 sb_1__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_40_prog_clk sb_1__1_.mem_bottom_track_1.mem_out\[2\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_51_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_301_ sb_1__1_.mux_right_track_12.out VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__clkbuf_2
XFILLER_24_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__1_.mux_right_ipin_4.mux_l1_in_0_ sb_1__1_.mux_bottom_track_3.out net83 cby_1__1_.mem_right_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_top_track_12.mux_l2_in_3__405 VGND VGND VPWR VPWR sb_1__1_.mux_top_track_12.mux_l2_in_3__405/HI
+ net405 sky130_fd_sc_hd__conb_1
XFILLER_92_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_20_prog_clk sb_1__1_.mem_left_track_21.mem_out\[0\]
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_21.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_33_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_21_prog_clk sb_1__1_.mem_left_track_5.mem_out\[1\]
+ net296 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_5.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mux_top_ipin_4.mux_l1_in_3_ net38 net7 cbx_1__1_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_14_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net295 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net124 grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_86_.in net134 VGND
+ VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_56_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net338 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_top_track_20.mux_l4_in_0_ sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_top_track_20.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_9.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_9.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_10_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_5.mux_l2_in_3_ net389 net292 sb_1__1_.mem_left_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_21_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_21_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__349
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__349/HI
+ net349 sky130_fd_sc_hd__conb_1
XFILLER_65_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_20_prog_clk sb_1__1_.mem_left_track_45.ccff_tail
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_53.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_65_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net358 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput109 chany_top_in_0[24] VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__clkbuf_1
XFILLER_84_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_60 net291 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_71 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_82 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_93 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__352
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__352/HI
+ net352 sky130_fd_sc_hd__conb_1
Xsb_1__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_30_prog_clk net2
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_0.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_46_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_right_track_28.mux_l2_in_0_ sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_right_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_15_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mux_bottom_track_37.mux_l2_in_1__376 VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_37.mux_l2_in_1__376/HI
+ net376 sky130_fd_sc_hd__conb_1
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_top_track_20.mux_l3_in_1_ sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_top_track_20.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_9.mux_l2_in_2_ net28 net39 cbx_1__1_.mem_top_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_81_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net329 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
Xinput91 chany_bottom_in[8] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__buf_2
Xinput80 chany_bottom_in[25] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_4
Xsb_1__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_54_prog_clk
+ sb_1__1_.mem_bottom_track_29.mem_out\[1\] net298 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_29.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_44_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__1_.mux_top_ipin_4.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_4.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_0.out sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mux_top_track_6.mux_l2_in_3__413 VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.mux_l2_in_3__413/HI
+ net413 sky130_fd_sc_hd__conb_1
XFILLER_67_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_bottom_track_13.mux_l2_in_0_ sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_bottom_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_bottom_track_5.mux_l3_in_0_ sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_bottom_track_5.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_left_track_5.mux_l4_in_0_ sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_left_track_5.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_78_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_28.mux_l1_in_1_ net127 net104 sb_1__1_.mem_right_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_89_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__1_.mux_right_ipin_9.mux_l1_in_0_ sb_1__1_.mux_bottom_track_1.out net84 cby_1__1_.mem_right_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_9.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_20.mux_l2_in_2_ net11 net15 sb_1__1_.mem_top_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_28_prog_clk sb_1__1_.mem_top_track_6.mem_out\[0\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_6.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_19_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net298 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__1_.mux_top_ipin_4.mux_l2_in_1_ cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_2_X cbx_1__1_.mem_top_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_58_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net367 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__mux2_2
XFILLER_22_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_46_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_46_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_27_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net298 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_377_ net134 VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__clkbuf_2
Xsb_1__1_.mux_bottom_track_13.mux_l1_in_1_ net42 net49 sb_1__1_.mem_bottom_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_9_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_5.mux_l2_in_1_ net278 sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_bottom_track_5.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_68_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_left_track_5.mux_l3_in_1_ sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_left_track_5.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_95_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_top_track_6.mux_l1_in_0_ net135 net141 sb_1__1_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_40_prog_clk sb_1__1_.mem_bottom_track_1.mem_out\[1\]
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_1.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_48_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_300_ net18 VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__clkbuf_2
XFILLER_24_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_19_prog_clk sb_1__1_.mem_left_track_13.ccff_tail
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_21.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_20_prog_clk sb_1__1_.mem_left_track_5.mem_out\[0\]
+ net296 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_5.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
Xcbx_1__1_.mux_top_ipin_4.mux_l1_in_2_ sb_1__1_.mux_left_track_21.out net13 cbx_1__1_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_14_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net295 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_56_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput1 ccff_head_1 VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_9.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_3_X cbx_1__1_.mem_top_ipin_9.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__364
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__364/HI
+ net364 sky130_fd_sc_hd__conb_1
Xclkbuf_0_prog_clk prog_clk VGND VGND VPWR VPWR clknet_0_prog_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_10_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_bottom_track_5.mux_l1_in_2_ net275 net60 sb_1__1_.mem_bottom_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_5.mux_l2_in_2_ net289 net90 sb_1__1_.mem_left_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_top_track_52.mux_l2_in_1__412 VGND VGND VPWR VPWR sb_1__1_.mux_top_track_52.mux_l2_in_1__412/HI
+ net412 sky130_fd_sc_hd__conb_1
XFILLER_80_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_0_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mux_right_ipin_11.mux_l2_in_3_ net309 sb_1__1_.mux_bottom_track_53.out
+ cby_1__1_.mem_right_ipin_11.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_44_prog_clk sb_1__1_.mem_bottom_track_7.mem_out\[2\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_11.ccff_head sky130_fd_sc_hd__dfrtp_1
XANTENNA_50 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_61 net294 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_83 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_72 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_94 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xoutput190 net190 VGND VGND VPWR VPWR chanx_right_out_0[1] sky130_fd_sc_hd__buf_12
XFILLER_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_top_track_20.mux_l3_in_0_ sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_top_track_20.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_41_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__1_.mux_top_ipin_9.mux_l2_in_1_ net8 cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__1_.mem_top_ipin_9.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_27_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
Xinput70 chany_bottom_in[16] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_2
Xinput81 chany_bottom_in[26] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__buf_4
Xsb_1__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_38_prog_clk
+ sb_1__1_.mem_bottom_track_29.mem_out\[0\] net296 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_29.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xinput92 chany_bottom_in[9] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__buf_4
XFILLER_88_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_94_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_10.mux_l2_in_3_ net416 net55 cbx_1__1_.mem_top_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_57_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_3_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net295 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_89_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_right_track_28.mux_l1_in_0_ net99 net100 sb_1__1_.mem_right_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_94_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_11.mux_l4_in_0_ cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_11.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_13_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_20.mux_l2_in_1_ net85 sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_top_track_20.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_9.mux_l1_in_2_ net46 net15 cbx_1__1_.mem_top_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_4_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_34_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_90_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_25_prog_clk sb_1__1_.mem_top_track_4.ccff_tail
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_6.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_19_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net298 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_29_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__1_.mux_top_ipin_4.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_4.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_31_prog_clk sb_1__1_.mem_right_track_10.mem_out\[2\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_10.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_10.mux_l1_in_4_ sb_1__1_.mux_left_track_45.out net30 cbx_1__1_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_89_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_27_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net298 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_72_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_15_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_15_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_60_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net327 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
X_376_ net134 VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__clkbuf_2
Xsb_1__1_.mux_bottom_track_13.mux_l1_in_0_ net116 net102 sb_1__1_.mem_bottom_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_5.mux_l2_in_0_ sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_bottom_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_5.mux_l3_in_0_ sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_left_track_5.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_68_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_40_prog_clk sb_1__1_.mem_bottom_track_1.mem_out\[0\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_1.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_63_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mux_top_ipin_15.mux_l2_in_3__421 VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_15.mux_l2_in_3__421/HI
+ net421 sky130_fd_sc_hd__conb_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
Xcby_1__1_.mux_right_ipin_11.mux_l3_in_1_ cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_11.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_10.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_9_X cbx_1__1_.mem_top_ipin_10.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_86_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_20.mux_l1_in_2_ net71 net55 sb_1__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_39_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_37.mux_l3_in_0_ sb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_bottom_track_37.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net124 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net134 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_86_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_2_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_20_prog_clk sb_1__1_.mem_left_track_3.ccff_tail
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_5.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xcbx_1__1_.mux_top_ipin_4.mux_l1_in_1_ net51 net20 cbx_1__1_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
X_359_ net77 VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_14_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net295 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ net146 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xinput2 ccff_head_2 VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_right_track_6.mux_l2_in_3__402 VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.mux_l2_in_3__402/HI
+ net402 sky130_fd_sc_hd__conb_1
XFILLER_83_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.out sky130_fd_sc_hd__buf_4
XFILLER_10_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mux_top_ipin_15.mux_l2_in_3_ net421 net62 cbx_1__1_.mem_top_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_bottom_track_5.mux_l1_in_1_ net36 net47 sb_1__1_.mem_bottom_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_7_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_left_track_5.mux_l2_in_1_ net77 sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_left_track_5.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_3.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_3.out sky130_fd_sc_hd__buf_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_12_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net295 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_30_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_30_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_0_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_61_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_11.mux_l2_in_2_ net86 net97 cby_1__1_.mem_right_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_10.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_10.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_29_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_bottom_track_37.mux_l2_in_1_ net376 sb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_bottom_track_37.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_64_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ net424 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net124 grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_32_.in net134 VGND
+ VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_43_prog_clk sb_1__1_.mem_bottom_track_7.mem_out\[1\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_7.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_40 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_62 chanx_right_in_0[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_84 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_73 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_51 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_95 net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput180 net180 VGND VGND VPWR VPWR chanx_right_out_0[10] sky130_fd_sc_hd__buf_12
Xoutput191 net191 VGND VGND VPWR VPWR chanx_right_out_0[20] sky130_fd_sc_hd__buf_12
XFILLER_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_13_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net298 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_75_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_494 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_9.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_9.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_29_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
Xcbx_1__1_.mux_top_ipin_12.mux_l2_in_3__418 VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_12.mux_l2_in_3__418/HI
+ net418 sky130_fd_sc_hd__conb_1
Xinput71 chany_bottom_in[17] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__buf_4
Xinput82 chany_bottom_in[27] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_4
Xsb_1__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_39_prog_clk
+ sb_1__1_.mem_bottom_track_21.ccff_tail net296 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_29.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput60 chanx_right_in_0[7] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_2
Xinput93 chany_top_in_0[0] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net347 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_8.mux_l2_in_3__320 VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_8.mux_l2_in_3__320/HI
+ net320 sky130_fd_sc_hd__conb_1
XFILLER_88_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mux_right_ipin_0.mux_l2_in_3_ net306 net119 cby_1__1_.mem_right_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_0.mux_l2_in_3__306 VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_0.mux_l2_in_3__306/HI
+ net306 sky130_fd_sc_hd__conb_1
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_left_track_5.mux_l1_in_2_ net83 net60 sb_1__1_.mem_left_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_83_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_10.mux_l2_in_2_ net14 cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mem_top_ipin_10.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_37.mux_l1_in_2_ net27 net8 sb_1__1_.mem_bottom_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_4_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__1_.mux_top_ipin_15.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_7_X net148 VGND VGND VPWR VPWR
+ cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_54_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_42_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_22_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_1_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_top_track_20.mux_l2_in_0_ sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_top_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_9.mux_l1_in_1_ sb_1__1_.mux_left_track_7.out net21 cbx_1__1_.mem_top_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__361
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__361/HI
+ net361 sky130_fd_sc_hd__conb_1
XFILLER_4_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_11.mux_l2_in_3__371 VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.mux_l2_in_3__371/HI
+ net371 sky130_fd_sc_hd__conb_1
Xsb_1__1_.mux_right_track_12.mux_l2_in_3_ net394 net26 sb_1__1_.mem_right_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_36_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_0.mux_l1_in_4_ sb_1__1_.mux_bottom_track_37.out net65 cby_1__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_31_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_29_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_32_prog_clk sb_1__1_.mem_right_track_10.mem_out\[1\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_10.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_81_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_10.mux_l1_in_3_ net38 net7 cbx_1__1_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_27_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail
+ net298 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_375_ net134 VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_55_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_55_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcbx_1__1_.mux_top_ipin_15.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_15.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_0.mux_l4_in_0_ cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X cby_1__1_.mem_right_ipin_0.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_68_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_41_prog_clk sb_1__1_.mem_bottom_track_1.ccff_head
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_1.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xsb_1__1_.mux_left_track_53.mux_l3_in_0_ sb_1__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_3_X cbx_1__1_.ccff_head VGND
+ VGND VPWR VPWR sb_1__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_48_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net349 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__mux2_4
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_5.mux_l2_in_3__317 VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_5.mux_l2_in_3__317/HI
+ net317 sky130_fd_sc_hd__conb_1
Xsb_1__1_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_19_prog_clk sb_1__1_.mem_left_track_13.mem_out\[2\]
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_13.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
Xcby_1__1_.mux_right_ipin_11.mux_l3_in_0_ cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_3_X cby_1__1_.mem_right_ipin_11.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_86_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_58_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_top_track_20.mux_l1_in_1_ net36 net41 sb_1__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_27_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_358_ net76 VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__1_.mux_top_ipin_4.mux_l1_in_0_ sb_1__1_.mux_left_track_3.out net23 cbx_1__1_.mem_top_ipin_4.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_4.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_15_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net295 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_289_ sb_1__1_.mux_right_track_36.out VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_2
XFILLER_46_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mux_right_ipin_5.mux_l2_in_3_ net317 net104 cby_1__1_.mem_right_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_56_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput3 chanx_left_in[0] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_2
XFILLER_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_20_prog_clk sb_1__1_.mem_left_track_45.mem_out\[1\]
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_45.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_3_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_0_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_1__1_.mux_right_track_12.mux_l4_in_0_ sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_right_track_12.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_15.mux_l2_in_2_ net31 net39 cbx_1__1_.mem_top_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_19_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_0.mux_l3_in_1_ cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_bottom_track_5.mux_l1_in_0_ net120 net107 sb_1__1_.mem_bottom_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_left_track_5.mux_l2_in_0_ sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_left_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_53.mux_l2_in_1_ net390 sb_1__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_left_track_53.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_13_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net298 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_0_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_92_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mux_right_ipin_11.mux_l2_in_1_ net66 cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__1_.mem_right_ipin_11.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_10.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_10.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_29_prog_clk sb_1__1_.mem_top_track_10.mem_out\[2\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_10.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_29_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_37.mux_l2_in_0_ sb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_bottom_track_37.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_43_prog_clk sb_1__1_.mem_bottom_track_7.mem_out\[0\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_7.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_30 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_41 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_63 sb_1__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_74 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_52 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_85 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_96 net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xoutput170 net170 VGND VGND VPWR VPWR chanx_left_out[29] sky130_fd_sc_hd__buf_12
Xoutput181 net181 VGND VGND VPWR VPWR chanx_right_out_0[11] sky130_fd_sc_hd__buf_12
Xoutput192 net192 VGND VGND VPWR VPWR chanx_right_out_0[21] sky130_fd_sc_hd__buf_12
XFILLER_75_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_2.mux_l2_in_3_ net406 net3 sb_1__1_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_14_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net298 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_right_track_12.mux_l3_in_1_ sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_right_track_12.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
Xinput72 chany_bottom_in[18] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_4
Xinput61 chanx_right_in_0[8] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_1
Xinput50 chanx_right_in_0[25] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_1
Xinput94 chany_top_in_0[10] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_4
Xinput83 chany_bottom_in[28] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_4
XFILLER_88_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__1_.mux_right_ipin_0.mux_l2_in_2_ net88 cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mem_right_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_5.mux_l1_in_1_ net47 net117 sb_1__1_.mem_left_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_29_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_53.mux_l1_in_2_ net292 net87 sb_1__1_.mem_left_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mux_right_ipin_5.mux_l4_in_0_ cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_5.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_94_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_11.mux_l1_in_2_ net103 net72 cby_1__1_.mem_right_ipin_11.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_10.mux_l2_in_1_ cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_2_X cbx_1__1_.mem_top_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_48_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_37.mux_l1_in_1_ net276 net38 sb_1__1_.mem_bottom_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_42_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mux_top_ipin_9.mux_l1_in_0_ sb_1__1_.mux_left_track_1.out net24 cbx_1__1_.mem_top_ipin_9.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_top_track_36.mux_l2_in_1__409 VGND VGND VPWR VPWR sb_1__1_.mux_top_track_36.mux_l2_in_1__409/HI
+ net409 sky130_fd_sc_hd__conb_1
XFILLER_48_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_12.mux_l2_in_2_ net12 net86 sb_1__1_.mem_right_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_75_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_49_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_61_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_47_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mux_right_ipin_0.mux_l1_in_3_ net102 net71 cby_1__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_11.mux_l2_in_3_ net382 net294 sb_1__1_.mem_left_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_top_track_2.mux_l4_in_0_ sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_9_X
+ sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_8_X sb_1__1_.mem_top_track_2.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_32_prog_clk sb_1__1_.mem_right_track_10.mem_out\[0\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_10.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_54_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_5.mux_l3_in_1_ cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_5.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_13_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_10.mux_l1_in_2_ sb_1__1_.mux_left_track_21.out net13 cbx_1__1_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_89_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__322
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__322/HI
+ net322 sky130_fd_sc_hd__conb_1
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_374_ net146 VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__clkbuf_1
Xcbx_1__1_.mux_top_ipin_15.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_3_X cbx_1__1_.mem_top_ipin_15.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_24_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_24_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_83_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_19_prog_clk sb_1__1_.mem_left_track_13.mem_out\[1\]
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_13.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__354
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__354/HI
+ net354 sky130_fd_sc_hd__conb_1
XFILLER_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_top_track_20.mux_l1_in_0_ net140 net142 sb_1__1_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_58_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_67_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_11.mux_l1_in_4_ net290 net288 sb_1__1_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_45_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_120 net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_top_track_2.mux_l3_in_1_ sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_6_X sb_1__1_.mem_top_track_2.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_41_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_357_ sb_1__1_.mux_top_track_20.out VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_15_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net295 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_288_ net5 VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_2
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__1_.mux_right_ipin_5.mux_l2_in_2_ net63 net94 cby_1__1_.mem_right_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xinput4 chanx_left_in[10] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_2
Xsb_1__1_.mux_top_track_44.mux_l3_in_0_ sb_1__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_top_track_44.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_36_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net363 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_26_prog_clk sb_1__1_.mem_left_track_45.mem_out\[0\]
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_45.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__1_.mux_top_ipin_15.mux_l2_in_1_ net8 cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__1_.mem_top_ipin_15.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_1__1_.mux_right_ipin_0.mux_l3_in_0_ cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_11.mux_l4_in_0_ sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_10_X
+ sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_9_X sb_1__1_.mem_left_track_11.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_53.mux_l2_in_0_ sb_1__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_left_track_53.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_68_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_0_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ net424 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net124 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net134 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_32_.in
+ sky130_fd_sc_hd__sdfrtp_1
Xcby_1__1_.mux_right_ipin_11.mux_l2_in_0_ cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_33_prog_clk sb_1__1_.mem_right_track_4.mem_out\[2\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_4.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_31_prog_clk sb_1__1_.mem_top_track_10.mem_out\[1\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_10.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_37_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_right_track_20.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_20.out sky130_fd_sc_hd__clkbuf_1
XFILLER_52_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_31 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_42_prog_clk sb_1__1_.mem_bottom_track_5.ccff_tail
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_7.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_20 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_75 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_42 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_64 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_53 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_86 net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_97 net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput160 net160 VGND VGND VPWR VPWR chanx_left_out[1] sky130_fd_sc_hd__buf_12
Xoutput182 net182 VGND VGND VPWR VPWR chanx_right_out_0[12] sky130_fd_sc_hd__buf_12
Xoutput193 net193 VGND VGND VPWR VPWR chanx_right_out_0[22] sky130_fd_sc_hd__buf_12
Xoutput171 net171 VGND VGND VPWR VPWR chanx_left_out[2] sky130_fd_sc_hd__buf_12
Xsb_1__1_.mux_top_track_2.mux_l2_in_2_ net32 net18 sb_1__1_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_47_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_3_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_top_track_44.mux_l2_in_1_ net411 sb_1__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_top_track_44.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_12.mux_l3_in_0_ sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_right_track_12.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_30_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput40 chanx_right_in_0[16] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_1
Xinput51 chanx_right_in_0[26] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__buf_4
Xinput73 chany_bottom_in[19] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_4
Xcbx_1__1_.mux_top_ipin_15.mux_l1_in_2_ sb_1__1_.mux_left_track_13.out net18 cbx_1__1_.mem_top_ipin_15.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xinput62 chanx_right_in_0[9] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_2
Xinput95 chany_top_in_0[11] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__buf_2
Xinput84 chany_bottom_in[29] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_4
XFILLER_88_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net365 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_0.mux_l2_in_1_ cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X cby_1__1_.mem_right_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_left_track_5.mux_l1_in_0_ net120 net107 sb_1__1_.mem_left_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_11.mux_l3_in_1_ sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_left_track_11.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_44_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_left_track_53.mux_l1_in_1_ net65 net35 sb_1__1_.mem_left_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_58_prog_clk cby_1__1_.mem_right_ipin_0.mem_out\[2\]
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_11.mux_l1_in_1_ sb_1__1_.mux_bottom_track_11.out net79 cby_1__1_.mem_right_ipin_11.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_10.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_10.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_57_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_top_track_4.mux_l2_in_3__410 VGND VGND VPWR VPWR sb_1__1_.mux_top_track_4.mux_l2_in_3__410/HI
+ net410 sky130_fd_sc_hd__conb_1
XFILLER_63_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_49_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_49_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_28_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_37.mux_l1_in_0_ net53 net98 sb_1__1_.mem_bottom_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_34_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_4.out sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mux_top_track_2.mux_l1_in_3_ net92 net78 sb_1__1_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_30_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__334
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__334/HI
+ net334 sky130_fd_sc_hd__conb_1
XFILLER_94_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__362
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__362/HI
+ net362 sky130_fd_sc_hd__conb_1
XFILLER_84_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mux_top_track_44.mux_l1_in_2_ net7 net22 sb_1__1_.mem_top_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_3.mux_l2_in_3__299 VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_3.mux_l2_in_3__299/HI
+ net299 sky130_fd_sc_hd__conb_1
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_right_track_12.mux_l2_in_1_ net72 sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_right_track_12.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_50_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_84_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_49_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mux_right_ipin_0.mux_l1_in_2_ sb_1__1_.mux_bottom_track_13.out net78 cby_1__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_31_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_11.mux_l2_in_2_ net292 sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mem_left_track_11.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_51_prog_clk cby_1__1_.mem_right_ipin_10.mem_out\[2\]
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_10.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_33_prog_clk sb_1__1_.mem_right_track_10.ccff_head
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_10.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mux_right_ipin_5.mux_l3_in_0_ cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_3_X cby_1__1_.mem_right_ipin_5.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_22_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mux_top_ipin_10.mux_l1_in_1_ net51 net20 cbx_1__1_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_13_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_373_ net124 VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__clkbuf_1
XFILLER_70_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_26_prog_clk sb_1__1_.mem_left_track_13.mem_out\[0\]
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_13.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_right_track_12.mux_l1_in_2_ net79 net131 sb_1__1_.mem_right_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_49_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.out sky130_fd_sc_hd__clkbuf_1
XFILLER_92_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net331 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__mux2_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_110 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_121 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_11.mux_l1_in_3_ net88 net73 sb_1__1_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_81_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_top_track_2.mux_l3_in_0_ sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X sb_1__1_.mem_top_track_2.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_9.mux_l2_in_3__305 VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_9.mux_l2_in_3__305/HI
+ net305 sky130_fd_sc_hd__conb_1
XFILLER_60_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_356_ net73 VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_15_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net295 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_287_ net4 VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__clkbuf_2
Xcby_1__1_.mux_right_ipin_5.mux_l2_in_1_ net92 cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__1_.mem_right_ipin_5.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_68_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput5 chanx_left_in[11] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_4
XFILLER_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_20_prog_clk sb_1__1_.mem_left_track_37.ccff_tail
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_45.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_10_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mux_top_ipin_15.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_15.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_2_prog_clk cby_1__1_.mem_right_ipin_3.mem_out\[2\]
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_3.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_51_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_0_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_339_ net85 VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__clkbuf_2
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_32_prog_clk sb_1__1_.mem_right_track_4.mem_out\[1\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_4.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_29_prog_clk sb_1__1_.mem_top_track_10.mem_out\[0\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_10.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_10 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_32 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_21 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_65 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_54 net116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_43 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_87 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_98 net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_76 net66 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_10_prog_clk cbx_1__1_.mem_top_ipin_11.mem_out\[2\]
+ net295 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_11.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xoutput150 net150 VGND VGND VPWR VPWR chanx_left_out[10] sky130_fd_sc_hd__buf_12
Xoutput161 net161 VGND VGND VPWR VPWR chanx_left_out[20] sky130_fd_sc_hd__buf_12
Xoutput183 net183 VGND VGND VPWR VPWR chanx_right_out_0[13] sky130_fd_sc_hd__buf_12
Xoutput194 net194 VGND VGND VPWR VPWR chanx_right_out_0[23] sky130_fd_sc_hd__buf_12
Xoutput172 net172 VGND VGND VPWR VPWR chanx_left_out[3] sky130_fd_sc_hd__buf_12
Xsb_1__1_.mux_top_track_2.mux_l2_in_1_ sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mux_right_ipin_5.mux_l1_in_2_ net103 net72 cby_1__1_.mem_right_ipin_5.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_3_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_top_track_44.mux_l2_in_0_ sb_1__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_top_track_44.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__357
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__357/HI
+ net357 sky130_fd_sc_hd__conb_1
XFILLER_34_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_right_track_4.mux_l2_in_3_ net399 net30 sb_1__1_.mem_right_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_30_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__346
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__346/HI
+ net346 sky130_fd_sc_hd__conb_1
Xinput30 chanx_left_in[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__buf_4
Xinput52 chanx_right_in_0[27] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput63 chany_bottom_in[0] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__1_.mux_top_ipin_15.mux_l1_in_1_ sb_1__1_.mux_left_track_7.out net21 cbx_1__1_.mem_top_ipin_15.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xinput41 chanx_right_in_0[17] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__buf_2
Xinput96 chany_top_in_0[12] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput85 chany_bottom_in[2] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_4
Xinput74 chany_bottom_in[1] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__buf_4
Xcby_1__1_.mux_right_ipin_0.mux_l2_in_0_ cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_52_prog_clk cby_1__1_.mem_right_ipin_13.mem_out\[2\]
+ net298 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_13.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_left_track_11.mux_l3_in_0_ sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_left_track_11.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_53.mux_l1_in_0_ net95 net113 sb_1__1_.mem_left_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_16_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_55_prog_clk cby_1__1_.mem_right_ipin_0.mem_out\[1\]
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_0.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_0.mux_l2_in_3_ net414 net59 cbx_1__1_.mem_top_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_32_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_11.mux_l1_in_0_ sb_1__1_.mux_bottom_track_5.out net82 cby_1__1_.mem_right_ipin_11.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_11.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_75_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_45.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_45.out sky130_fd_sc_hd__clkbuf_2
XFILLER_16_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_18_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_18_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_34_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_bottom_track_1.mux_l2_in_3_ net370 net4 sb_1__1_.mem_bottom_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_34_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_top_track_2.mux_l1_in_2_ net62 net48 sb_1__1_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_89_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_bottom_track_21.mux_l2_in_3_ net373 net25 sb_1__1_.mem_bottom_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_44.mux_l1_in_1_ net67 net33 sb_1__1_.mem_top_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_13_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_12.mux_l2_in_0_ sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_right_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_68_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_0.mux_l1_in_1_ sb_1__1_.mux_bottom_track_7.out net81 cby_1__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_88_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__1_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_51_prog_clk cby_1__1_.mem_right_ipin_10.mem_out\[1\]
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_10.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_left_track_11.mux_l2_in_1_ sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_left_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__1_.mux_top_ipin_0.mux_l1_in_4_ sb_1__1_.mux_left_track_37.out net5 cbx_1__1_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_86_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_right_track_36.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_36.out sky130_fd_sc_hd__clkbuf_1
XFILLER_54_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_10.mux_l1_in_0_ sb_1__1_.mux_left_track_3.out net23 cbx_1__1_.mem_top_ipin_10.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_10.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_85_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_372_ net124 VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__clkbuf_1
XFILLER_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_right_track_4.mux_l4_in_0_ sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_right_track_4.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_13_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__1_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_56_prog_clk cby_1__1_.mem_right_ipin_6.mem_out\[2\]
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_6.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_5_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_0.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X cbx_1__1_.mem_top_ipin_0.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_33_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_33_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_20_prog_clk sb_1__1_.mem_left_track_11.ccff_tail
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_13.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_39_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_12.mux_l1_in_1_ net125 net116 sb_1__1_.mem_right_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__343
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__343/HI
+ net343 sky130_fd_sc_hd__conb_1
XFILLER_2_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_4_prog_clk cbx_1__1_.mem_top_ipin_14.mem_out\[2\]
+ net295 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_14.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_85_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_1.mux_l4_in_0_ sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_9_X
+ sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_8_X sb_1__1_.mem_bottom_track_1.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_100 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_11.mux_l1_in_2_ net80 net58 sb_1__1_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_122 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_111 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_top_track_10.mux_l2_in_3__404 VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.mux_l2_in_3__404/HI
+ net404 sky130_fd_sc_hd__conb_1
X_355_ net72 VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_286_ net32 VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_15_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net295 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_21.mux_l4_in_0_ sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_bottom_track_21.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_5.mux_l2_in_0_ cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xinput6 chanx_left_in[12] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_2
XFILLER_64_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__1_.mux_top_ipin_5.mux_l2_in_3_ net301 net44 cbx_1__1_.mem_top_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_87_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_right_track_4.mux_l3_in_1_ sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_right_track_4.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_19_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_55_prog_clk cby_1__1_.mem_right_ipin_3.mem_out\[1\]
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_3.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net360 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__mux2_2
XFILLER_51_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__1_.mux_top_ipin_0.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_93_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_1_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__358
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__358/HI
+ net358 sky130_fd_sc_hd__conb_1
XFILLER_92_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_338_ net74 VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__clkbuf_2
X_269_ net47 VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__clkbuf_2
Xsb_1__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_28_prog_clk sb_1__1_.mem_top_track_10.ccff_head
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_10.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_44_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_32_prog_clk sb_1__1_.mem_right_track_4.mem_out\[0\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_4.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_69_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_11 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_22 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_44 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_33 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_66 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_55 net116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_77 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_99 net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_88 net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_41_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_bottom_track_1.mux_l3_in_1_ sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_6_X sb_1__1_.mem_bottom_track_1.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_10_prog_clk cbx_1__1_.mem_top_ipin_11.mem_out\[1\]
+ net295 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_11.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xoutput151 net151 VGND VGND VPWR VPWR chanx_left_out[11] sky130_fd_sc_hd__buf_12
Xsb_1__1_.mux_top_track_2.mux_l2_in_0_ sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xoutput184 net184 VGND VGND VPWR VPWR chanx_right_out_0[14] sky130_fd_sc_hd__buf_12
Xsb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_3.out sky130_fd_sc_hd__buf_4
Xoutput195 net195 VGND VGND VPWR VPWR chanx_right_out_0[24] sky130_fd_sc_hd__buf_12
Xoutput173 net173 VGND VGND VPWR VPWR chanx_left_out[4] sky130_fd_sc_hd__buf_12
Xoutput162 net162 VGND VGND VPWR VPWR chanx_left_out[21] sky130_fd_sc_hd__buf_12
XFILLER_75_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_21.mux_l3_in_1_ sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_bottom_track_21.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_70_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_5.mux_l1_in_1_ sb_1__1_.mux_bottom_track_11.out net79 cby_1__1_.mem_right_ipin_5.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_2_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_21_prog_clk cbx_1__1_.mem_top_ipin_0.mem_out\[2\]
+ net296 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_46_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_30_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_right_track_4.mux_l2_in_2_ net17 net90 sb_1__1_.mem_right_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xinput31 chanx_left_in[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_2
Xinput20 chanx_left_in[25] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_4
Xinput53 chanx_right_in_0[28] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput64 chany_bottom_in[10] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__buf_4
Xcbx_1__1_.mux_top_ipin_15.mux_l1_in_0_ sb_1__1_.mux_left_track_1.out net24 cbx_1__1_.mem_top_ipin_15.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xinput42 chanx_right_in_0[18] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_4
Xinput97 chany_top_in_0[13] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__buf_2
Xinput75 chany_bottom_in[20] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__buf_2
Xinput86 chany_bottom_in[3] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__buf_4
Xcby_1__1_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_53_prog_clk cby_1__1_.mem_right_ipin_13.mem_out\[1\]
+ net298 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_13.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_69_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_55_prog_clk cby_1__1_.mem_right_ipin_0.mem_out\[0\]
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_0.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_25_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mux_top_ipin_0.mux_l2_in_2_ net28 cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mem_top_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net344 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_5.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_5.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_31_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_58_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_58_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcby_1__1_.mux_right_ipin_15.mux_l2_in_3__313 VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_15.mux_l2_in_3__313/HI
+ net313 sky130_fd_sc_hd__conb_1
XFILLER_7_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_1__1_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_48_prog_clk cby_1__1_.mem_right_ipin_9.mem_out\[2\]
+ net298 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_10.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_3_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_42_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_81_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_bottom_track_1.mux_l2_in_2_ net21 net23 sb_1__1_.mem_bottom_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_34_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_top_track_2.mux_l1_in_1_ net52 net140 sb_1__1_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_30_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_21.mux_l2_in_2_ net6 net11 sb_1__1_.mem_bottom_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_44.mux_l1_in_0_ net37 net137 sb_1__1_.mem_top_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_13_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mux_right_ipin_0.mux_l1_in_0_ sb_1__1_.mux_bottom_track_1.out net84 cby_1__1_.mem_right_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_83_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_left_track_21.mux_l2_in_3__384 VGND VGND VPWR VPWR sb_1__1_.mux_left_track_21.mux_l2_in_3__384/HI
+ net384 sky130_fd_sc_hd__conb_1
XFILLER_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_51_prog_clk cby_1__1_.mem_right_ipin_10.mem_out\[0\]
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_10.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xsb_1__1_.mux_left_track_11.mux_l2_in_0_ sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_left_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_58_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mux_top_ipin_0.mux_l1_in_3_ net42 net11 cbx_1__1_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_3_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_3_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcbx_1__1_.mux_top_ipin_5.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_5.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_38_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_371_ net124 VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__clkbuf_1
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_56_prog_clk cby_1__1_.mem_right_ipin_6.mem_out\[1\]
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_6.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_bottom_track_1.mux_l1_in_3_ net279 net276 sb_1__1_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_1.mux_l2_in_3_ net381 net293 sb_1__1_.mem_left_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_right_track_12.mux_l1_in_0_ net102 net109 sb_1__1_.mem_right_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_40_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_4_prog_clk cbx_1__1_.mem_top_ipin_14.mem_out\[1\]
+ net295 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_14.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_57_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_49_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_123 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_101 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_112 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_left_track_11.mux_l1_in_1_ net43 net118 sb_1__1_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_8.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_60_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_354_ net71 VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__clkbuf_2
X_285_ sb_1__1_.mux_right_track_44.out VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput7 chanx_left_in[13] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_4
XFILLER_49_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_7_prog_clk cbx_1__1_.mem_top_ipin_3.mem_out\[2\]
+ net298 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_3.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_5.mux_l2_in_2_ net3 net34 cbx_1__1_.mem_top_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_right_track_36.mux_l3_in_0_ sb_1__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_right_track_36.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_87_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_4.mux_l3_in_0_ sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_right_track_4.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_59_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_54_prog_clk cby_1__1_.mem_right_ipin_3.mem_out\[0\]
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_3.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_0.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_1_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_337_ sb_1__1_.mux_bottom_track_1.out VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__clkbuf_2
X_268_ net46 VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__clkbuf_2
Xsb_1__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_31_prog_clk sb_1__1_.mem_right_track_2.ccff_tail
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_4.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__336
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__336/HI
+ net336 sky130_fd_sc_hd__conb_1
XFILLER_56_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_12 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_23 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_45 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_34 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_56 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_78 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_67 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_89 net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__1_.mux_bottom_track_1.mux_l3_in_0_ sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X sb_1__1_.mem_bottom_track_1.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_5_prog_clk cbx_1__1_.mem_top_ipin_11.mem_out\[0\]
+ net295 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_11.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xsb_1__1_.mux_left_track_1.mux_l4_in_0_ sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_9_X
+ sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_8_X sb_1__1_.mem_left_track_1.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
Xoutput152 net152 VGND VGND VPWR VPWR chanx_left_out[12] sky130_fd_sc_hd__buf_12
Xoutput185 net185 VGND VGND VPWR VPWR chanx_right_out_0[15] sky130_fd_sc_hd__buf_12
Xoutput174 net174 VGND VGND VPWR VPWR chanx_left_out[5] sky130_fd_sc_hd__buf_12
Xoutput163 net163 VGND VGND VPWR VPWR chanx_left_out[22] sky130_fd_sc_hd__buf_12
Xoutput196 net196 VGND VGND VPWR VPWR chanx_right_out_0[25] sky130_fd_sc_hd__buf_12
XFILLER_87_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
Xsb_1__1_.mux_bottom_track_21.mux_l3_in_0_ sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_bottom_track_21.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_5.mux_l1_in_0_ sb_1__1_.mux_bottom_track_5.out net82 cby_1__1_.mem_right_ipin_5.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_5.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_1_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_9.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_78_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_21_prog_clk cbx_1__1_.mem_top_ipin_0.mem_out\[1\]
+ net296 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_0.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_46_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_right_track_36.mux_l2_in_1_ net398 sb_1__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_right_track_36.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_30_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_right_track_4.mux_l2_in_1_ net66 sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_right_track_4.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xinput10 chanx_left_in[16] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_2
Xinput21 chanx_left_in[26] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_4
Xinput54 chanx_right_in_0[29] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput32 chanx_left_in[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_4
Xinput43 chanx_right_in_0[19] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__buf_2
Xinput98 chany_top_in_0[14] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_4
Xinput76 chany_bottom_in[21] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_4
Xinput65 chany_bottom_in[11] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_4
Xinput87 chany_bottom_in[4] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_2
Xcby_1__1_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_52_prog_clk cby_1__1_.mem_right_ipin_13.mem_out\[0\]
+ net298 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_13.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xcbx_1__1_.mux_top_ipin_10.mux_l2_in_3__416 VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_10.mux_l2_in_3__416/HI
+ net416 sky130_fd_sc_hd__conb_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_59_prog_clk net1
+ net123 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_0.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_37_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__1_.mux_top_ipin_0.mux_l2_in_1_ cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X cbx_1__1_.mem_top_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_87_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_77 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__1_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_44_prog_clk cby_1__1_.mem_right_ipin_9.mem_out\[1\]
+ net298 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_9.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_27_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_27_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_44_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_42_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_1.mux_l2_in_1_ sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_bottom_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_1.mux_l3_in_1_ sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_6_X sb_1__1_.mem_left_track_1.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_22_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_top_track_2.mux_l1_in_0_ net137 net142 sb_1__1_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_8_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_bottom_track_21.mux_l2_in_1_ net280 sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_bottom_track_21.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net124 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net134 VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__sdfrtp_2
XFILLER_25_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_right_track_36.mux_l1_in_2_ net8 net68 sb_1__1_.mem_right_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_68_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_4.mux_l1_in_2_ net77 net130 sb_1__1_.mem_right_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_75_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mem_right_ipin_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_48_prog_clk cby_1__1_.mem_right_ipin_10.ccff_head
+ net298 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_10.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_58_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__1_.mux_top_ipin_0.mux_l1_in_2_ sb_1__1_.mux_left_track_13.out net18 cbx_1__1_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_50_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_54_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_13_prog_clk cbx_1__1_.mem_top_ipin_6.mem_out\[2\]
+ net298 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_6.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_30_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mux_top_ipin_5.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_3_X cbx_1__1_.mem_top_ipin_5.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_370_ net297 VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__clkbuf_1
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_51_prog_clk cby_1__1_.mem_right_ipin_6.mem_out\[0\]
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_6.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_79_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_1.mux_l1_in_2_ net281 net57 sb_1__1_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_1.mux_l2_in_2_ net290 net287 sb_1__1_.mem_left_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_95_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_21.mux_l1_in_2_ net282 net55 sb_1__1_.mem_bottom_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ net424 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net124 grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_41_.in net134 VGND
+ VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
Xclkbuf_leaf_42_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_42_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_67_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_3.mux_l2_in_3__315 VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_3.mux_l2_in_3__315/HI
+ net315 sky130_fd_sc_hd__conb_1
XFILLER_67_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_57_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_5_prog_clk cbx_1__1_.mem_top_ipin_14.mem_out\[0\]
+ net295 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_14.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_26_prog_clk sb_1__1_.mem_left_track_37.mem_out\[1\]
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_37.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_18_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_left_track_11.mux_l1_in_0_ net96 net103 sb_1__1_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_113 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_124 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_102 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_353_ sb_1__1_.mux_top_track_28.out VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_15_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net296 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
X_284_ net30 VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput8 chanx_left_in[14] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_4
XFILLER_39_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_7_prog_clk cbx_1__1_.mem_top_ipin_3.mem_out\[1\]
+ net298 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_3.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_20_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_5.mux_l2_in_1_ net32 cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__1_.mem_top_ipin_5.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
Xcby_1__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_55_prog_clk cby_1__1_.mem_right_ipin_2.ccff_tail
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_3.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xsb_1__1_.mux_left_track_1.mux_l1_in_3_ net63 net64 sb_1__1_.mem_left_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_23_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_336_ sb_1__1_.mux_bottom_track_3.out VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__clkbuf_2
X_267_ sb_1__1_.mux_left_track_21.out VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net333 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_13 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net342 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net294 sky130_fd_sc_hd__mux2_4
XFILLER_32_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_35 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_24 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_57 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_46 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_68 net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_79 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mem_top_ipin_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_4_prog_clk cbx_1__1_.mem_top_ipin_10.ccff_tail
+ net295 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_11.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
Xoutput186 net186 VGND VGND VPWR VPWR chanx_right_out_0[16] sky130_fd_sc_hd__buf_12
Xoutput175 net175 VGND VGND VPWR VPWR chanx_left_out[6] sky130_fd_sc_hd__buf_12
Xoutput153 net153 VGND VGND VPWR VPWR chanx_left_out[13] sky130_fd_sc_hd__buf_12
Xoutput164 net164 VGND VGND VPWR VPWR chanx_left_out[23] sky130_fd_sc_hd__buf_12
Xoutput197 net197 VGND VGND VPWR VPWR chanx_right_out_0[26] sky130_fd_sc_hd__buf_12
XFILLER_28_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_1_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_5.mux_l1_in_2_ net43 net12 cbx_1__1_.mem_top_ipin_5.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_9_prog_clk cbx_1__1_.mem_top_ipin_0.mem_out\[0\]
+ net296 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_0.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_93_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_right_track_36.mux_l2_in_0_ sb_1__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_right_track_36.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_61_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_31_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_4.mux_l2_in_0_ sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_right_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
X_319_ sb_1__1_.mux_bottom_track_37.out VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__clkbuf_2
Xinput11 chanx_left_in[17] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_4
Xinput22 chanx_left_in[27] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_2
Xinput55 chanx_right_in_0[2] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_4
Xinput44 chanx_right_in_0[1] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__buf_2
Xinput33 chanx_right_in_0[0] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput66 chany_bottom_in[12] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_2
Xinput77 chany_bottom_in[22] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_4
Xinput88 chany_bottom_in[5] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__buf_4
Xinput99 chany_top_in_0[15] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__buf_2
Xcby_1__1_.mem_right_ipin_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_52_prog_clk cby_1__1_.mem_right_ipin_12.ccff_tail
+ net298 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_13.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_69_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__1_.mux_top_ipin_0.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_33_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_11_prog_clk cbx_1__1_.mem_top_ipin_9.mem_out\[2\]
+ net298 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_10.ccff_head sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_52_prog_clk cby_1__1_.mem_right_ipin_9.mem_out\[0\]
+ net298 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_9.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_1__1_.mux_right_ipin_12.mux_l2_in_3_ net310 net119 cby_1__1_.mem_right_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_45_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_42_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_1.mux_l2_in_0_ sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_bottom_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_62_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_left_track_1.mux_l3_in_0_ sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_4_X sb_1__1_.mem_left_track_1.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_30_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_bottom_track_21.mux_l2_in_0_ sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_bottom_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_1_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_right_track_36.mux_l1_in_1_ net83 net128 sb_1__1_.mem_right_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_88_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_4.mux_l1_in_1_ net127 net120 sb_1__1_.mem_right_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_90_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__1_.mux_top_ipin_0.mux_l1_in_1_ sb_1__1_.mux_left_track_7.out net21 cbx_1__1_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.out sky130_fd_sc_hd__clkbuf_1
XFILLER_94_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_
+ sky130_fd_sc_hd__clkbuf_1
Xcbx_1__1_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_13_prog_clk cbx_1__1_.mem_top_ipin_6.mem_out\[1\]
+ net298 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_6.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_0_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_4_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_12.mux_l1_in_4_ sb_1__1_.mux_bottom_track_37.out net65 cby_1__1_.mem_right_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_11.mux_l2_in_3_ net417 sb_1__1_.mux_left_track_53.out cbx_1__1_.mem_top_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__1_.mem_right_ipin_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_55_prog_clk cby_1__1_.mem_right_ipin_5.ccff_tail
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_6.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_79_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_1.mux_l1_in_1_ net34 net51 sb_1__1_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_bottom_track_53.mux_l2_in_1__379 VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_53.mux_l2_in_1__379/HI
+ net379 sky130_fd_sc_hd__conb_1
XFILLER_79_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_left_track_1.mux_l2_in_1_ sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_left_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_88_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net328 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_44_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_bottom_track_21.mux_l1_in_1_ net41 net50 sb_1__1_.mem_bottom_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_12_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_11_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_11_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_79_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mux_right_ipin_12.mux_l4_in_0_ cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_9_X cby_1__1_.mem_right_ipin_12.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mem_top_ipin_14.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_6_prog_clk cbx_1__1_.mem_top_ipin_13.ccff_tail
+ net295 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_14.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_25_prog_clk sb_1__1_.mem_left_track_37.mem_out\[0\]
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_37.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_103 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_125 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_114 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_352_ net69 VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_15_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net296 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_283_ net29 VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput9 chanx_left_in[15] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_4
XFILLER_17_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_8_prog_clk cbx_1__1_.mem_top_ipin_3.mem_out\[0\]
+ net298 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_3.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_44_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_5.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_5.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_87_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_left_track_1.mux_l1_in_2_ net81 net34 sb_1__1_.mem_left_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_335_ sb_1__1_.mux_bottom_track_5.out VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__clkbuf_2
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_266_ net43 VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__1_.mux_right_ipin_12.mux_l3_in_1_ cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_12.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_11.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_11.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XANTENNA_14 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_47 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_36 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_25 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_69 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_58 net121 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__325
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__325/HI
+ net325 sky130_fd_sc_hd__conb_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
Xoutput176 net176 VGND VGND VPWR VPWR chanx_left_out[7] sky130_fd_sc_hd__buf_12
Xoutput154 net154 VGND VGND VPWR VPWR chanx_left_out[14] sky130_fd_sc_hd__buf_12
Xoutput165 net165 VGND VGND VPWR VPWR chanx_left_out[24] sky130_fd_sc_hd__buf_12
XFILLER_87_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput187 net187 VGND VGND VPWR VPWR chanx_right_out_0[17] sky130_fd_sc_hd__buf_12
Xoutput198 net198 VGND VGND VPWR VPWR chanx_right_out_0[27] sky130_fd_sc_hd__buf_12
XFILLER_87_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_35_prog_clk sb_1__1_.mem_right_track_20.mem_out\[2\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_20.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_0_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_78_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_5.mux_l1_in_1_ sb_1__1_.mux_left_track_11.out net19 cbx_1__1_.mem_top_ipin_5.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_21_prog_clk cbx_1__1_.ccff_head
+ net296 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_0.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_46_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_61_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_30_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_318_ net95 VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__clkbuf_2
Xinput12 chanx_left_in[18] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_4
Xinput23 chanx_left_in[28] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_4
X_249_ net55 VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__clkbuf_2
Xinput34 chanx_right_in_0[10] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_4
Xinput45 chanx_right_in_0[20] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_1
Xinput67 chany_bottom_in[13] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__buf_4
Xinput78 chany_bottom_in[23] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__buf_4
Xinput89 chany_bottom_in[6] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_2
Xinput56 chanx_right_in_0[3] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__buf_2
XFILLER_6_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_10_prog_clk cbx_1__1_.mem_top_ipin_9.mem_out\[1\]
+ net298 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_9.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_35_prog_clk sb_1__1_.mem_right_track_52.mem_out\[1\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_1.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mem_right_ipin_9.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_49_prog_clk cby_1__1_.mem_right_ipin_8.ccff_tail
+ net298 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_9.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_78_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_1__1_.mux_right_ipin_12.mux_l2_in_2_ net88 cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mem_right_ipin_12.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_11.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_11.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_93_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_42_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_66_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_49_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_74_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_36_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_36_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_30_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_right_track_36.mux_l1_in_0_ net96 net98 sb_1__1_.mem_right_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_right_track_4.mux_l1_in_0_ net107 net113 sb_1__1_.mem_right_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__328
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__328/HI
+ net328 sky130_fd_sc_hd__conb_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__1_.mux_top_ipin_0.mux_l1_in_0_ sb_1__1_.mux_left_track_1.out net24 cbx_1__1_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_
+ sky130_fd_sc_hd__clkbuf_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1 cby_1__1_.mem_right_ipin_4.ccff_tail VGND VGND VPWR VPWR net423 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_94_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__1_.mux_right_ipin_1.mux_l2_in_3_ net307 net118 cby_1__1_.mem_right_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_50_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_0_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_13_prog_clk cbx_1__1_.mem_top_ipin_6.mem_out\[0\]
+ net296 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_6.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_11_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_27_prog_clk sb_1__1_.mem_top_track_2.mem_out\[2\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_57_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_12.mux_l1_in_3_ net102 net71 cby_1__1_.mem_right_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_11.mux_l2_in_2_ net26 net37 cbx_1__1_.mem_top_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_70_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ net424 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net124 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net134 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_41_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_5_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_1.mux_l1_in_0_ net94 net111 sb_1__1_.mem_bottom_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_1.mux_l2_in_0_ sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_left_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_0_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_48_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net298 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_48_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_21.mux_l1_in_0_ net115 net101 sb_1__1_.mem_bottom_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_44_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_51_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_51_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_82_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_22_prog_clk sb_1__1_.mem_left_track_29.ccff_tail
+ net296 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_37.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_104 net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_115 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_126 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_351_ net68 VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__clkbuf_2
XFILLER_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_282_ net28 VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_45.mux_l3_in_0_ sb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_bottom_track_45.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_7.mux_l2_in_3__303 VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_7.mux_l2_in_3__303/HI
+ net303 sky130_fd_sc_hd__conb_1
XFILLER_5_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_8_prog_clk cbx_1__1_.mem_top_ipin_2.ccff_tail
+ net296 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_3.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_17_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_19_prog_clk sb_1__1_.mem_left_track_1.mem_out\[2\]
+ net296 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_55_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_left_track_1.mux_l1_in_1_ net51 net94 sb_1__1_.mem_left_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_11_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__1_.mux_right_ipin_1.mux_l4_in_0_ cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_1.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_58_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_334_ sb_1__1_.mux_bottom_track_7.out VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__clkbuf_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_265_ net42 VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mux_right_ipin_12.mux_l3_in_0_ cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_12.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_15 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_26 net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_37 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_48 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_59 net125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
Xoutput177 net177 VGND VGND VPWR VPWR chanx_left_out[8] sky130_fd_sc_hd__buf_12
Xoutput155 net155 VGND VGND VPWR VPWR chanx_left_out[15] sky130_fd_sc_hd__buf_12
Xoutput166 net166 VGND VGND VPWR VPWR chanx_left_out[25] sky130_fd_sc_hd__buf_12
Xoutput188 net188 VGND VGND VPWR VPWR chanx_right_out_0[18] sky130_fd_sc_hd__buf_12
Xoutput199 net199 VGND VGND VPWR VPWR chanx_right_out_0[28] sky130_fd_sc_hd__buf_12
XFILLER_87_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_45.mux_l2_in_1_ net377 sb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_bottom_track_45.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_55_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_44_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_36_prog_clk sb_1__1_.mem_right_track_20.mem_out\[1\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_20.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_1_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_3_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_5.mux_l1_in_0_ sb_1__1_.mux_left_track_5.out net22 cbx_1__1_.mem_top_ipin_5.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net324 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__mux2_4
XFILLER_27_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_31_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_left_track_45.mux_l2_in_1__388 VGND VGND VPWR VPWR sb_1__1_.mux_left_track_45.mux_l2_in_1__388/HI
+ net388 sky130_fd_sc_hd__conb_1
X_317_ net94 VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_6.mux_l2_in_3_ net318 net119 cby_1__1_.mem_right_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xinput13 chanx_left_in[19] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_4
X_248_ net44 VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_2
Xinput24 chanx_left_in[29] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_4
Xinput35 chanx_right_in_0[11] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_2
Xinput46 chanx_right_in_0[21] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_2
Xinput68 chany_bottom_in[14] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__buf_4
Xinput79 chany_bottom_in[24] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_4
Xinput57 chanx_right_in_0[4] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net369 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ net147 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_10_prog_clk cbx_1__1_.mem_top_ipin_9.mem_out\[0\]
+ net298 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_9.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xcby_1__1_.mux_right_ipin_1.mux_l3_in_1_ cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_6_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_6_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_87_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_35_prog_clk sb_1__1_.mem_right_track_52.mem_out\[0\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_52.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcby_1__1_.mux_right_ipin_12.mux_l2_in_1_ cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_2_X cby_1__1_.mem_right_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_11.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_3_X cbx_1__1_.mem_top_ipin_11.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_3_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_43_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_49_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_bottom_track_45.mux_l1_in_2_ net3 net7 sb_1__1_.mem_bottom_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_6_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mux_right_ipin_6.mux_l1_in_4_ sb_1__1_.mux_bottom_track_37.out net65 cby_1__1_.mem_right_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__344
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__344/HI
+ net344 sky130_fd_sc_hd__conb_1
Xsb_1__1_.mux_right_track_20.mux_l2_in_3_ net396 net25 sb_1__1_.mem_right_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_66_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_1.mux_l2_in_2_ net87 net98 cby_1__1_.mem_right_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_0_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mem_top_ipin_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_9_prog_clk cbx_1__1_.mem_top_ipin_5.ccff_tail
+ net298 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_6.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_62_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_28_prog_clk sb_1__1_.mem_top_track_2.mem_out\[1\]
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_2.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mux_right_ipin_6.mux_l4_in_0_ cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_9_X cby_1__1_.mem_right_ipin_6.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_24_prog_clk sb_1__1_.mem_top_track_20.mem_out\[2\]
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_20.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_80_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__1_.mux_right_ipin_12.mux_l1_in_2_ sb_1__1_.mux_bottom_track_13.out net78 cby_1__1_.mem_right_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_11.mux_l2_in_1_ net6 cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__1_.mem_top_ipin_11.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net346 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_20_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_20_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_62_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_27_prog_clk sb_1__1_.mem_top_track_52.mem_out\[1\]
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_0.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_85_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_105 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_116 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_127 net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_350_ net67 VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__clkbuf_2
X_281_ sb_1__1_.mux_right_track_52.out VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_14_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net295 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.out sky130_fd_sc_hd__clkbuf_1
XFILLER_1_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_left_track_13.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_13.out sky130_fd_sc_hd__buf_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_0.out sky130_fd_sc_hd__clkbuf_1
XFILLER_65_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_6.mux_l3_in_1_ cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_6.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_59_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_20_prog_clk sb_1__1_.mem_left_track_1.mem_out\[1\]
+ net296 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_1.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mux_top_ipin_11.mux_l1_in_2_ net43 net12 cbx_1__1_.mem_top_ipin_11.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_55_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_1.mux_l1_in_0_ net111 net114 sb_1__1_.mem_left_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_50_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_right_track_20.mux_l4_in_0_ sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_right_track_20.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_46_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_333_ net111 VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_264_ net41 VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__clkbuf_2
XFILLER_1_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_27 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_16 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_38 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_49 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput145 net145 VGND VGND VPWR VPWR bottom_width_0_height_0_subtile_0__pin_cout_0_
+ sky130_fd_sc_hd__buf_12
Xoutput156 net156 VGND VGND VPWR VPWR chanx_left_out[16] sky130_fd_sc_hd__buf_12
Xoutput167 net167 VGND VGND VPWR VPWR chanx_left_out[26] sky130_fd_sc_hd__buf_12
Xoutput189 net189 VGND VGND VPWR VPWR chanx_right_out_0[19] sky130_fd_sc_hd__buf_12
Xoutput178 net178 VGND VGND VPWR VPWR chanx_left_out[9] sky130_fd_sc_hd__buf_12
XFILLER_87_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_45.out sky130_fd_sc_hd__clkbuf_2
Xsb_1__1_.mux_bottom_track_45.mux_l2_in_0_ sb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_bottom_track_45.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_55_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_44_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_32_prog_clk sb_1__1_.mem_right_track_20.mem_out\[0\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_20.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_7_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_6.mux_l2_in_2_ net88 cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mem_right_ipin_6.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_42_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_31_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_316_ net122 VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput14 chanx_left_in[1] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_4
Xinput25 chanx_left_in[2] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__buf_2
Xinput36 chanx_right_in_0[12] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_1
Xinput47 chanx_right_in_0[22] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_4
Xinput69 chany_bottom_in[15] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__clkbuf_4
Xinput58 chanx_right_in_0[5] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_2
XFILLER_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_right_track_20.mux_l3_in_1_ sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_right_track_20.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_60_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__1_.mem_top_ipin_9.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_11_prog_clk cbx_1__1_.mem_top_ipin_8.ccff_tail
+ net298 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_9.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xcby_1__1_.mux_right_ipin_1.mux_l3_in_0_ cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X cby_1__1_.mem_right_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_0_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__339
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__339/HI
+ net339 sky130_fd_sc_hd__conb_1
XFILLER_28_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_34_prog_clk sb_1__1_.mem_right_track_44.ccff_tail
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_52.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xsb_1__1_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_16_prog_clk sb_1__1_.mem_left_track_7.mem_out\[2\]
+ net296 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_11.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mux_right_ipin_12.mux_l2_in_0_ cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_13.mux_l2_in_3__311 VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_13.mux_l2_in_3__311/HI
+ net311 sky130_fd_sc_hd__conb_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_43_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ccff_tail
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_45.mux_l1_in_1_ net277 net37 sb_1__1_.mem_bottom_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_45_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_45_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_1_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_6.mux_l1_in_3_ net102 net71 cby_1__1_.mem_right_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_right_track_20.mux_l2_in_2_ net11 net85 sb_1__1_.mem_right_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_39_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_81_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_1.mux_l2_in_1_ net67 cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__1_.mem_right_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_0_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_22_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_28_prog_clk sb_1__1_.mem_top_track_2.mem_out\[0\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_2.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_24_prog_clk sb_1__1_.mem_top_track_20.mem_out\[1\]
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_20.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_12.mux_l1_in_1_ sb_1__1_.mux_bottom_track_7.out net81 cby_1__1_.mem_right_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_11.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_11.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_22_prog_clk sb_1__1_.mem_left_track_29.mem_out\[2\]
+ net296 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_29.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_8_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_50_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_27_prog_clk sb_1__1_.mem_top_track_52.mem_out\[0\]
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_52.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_106 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_128 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_117 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_280_ net26 VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_14_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net295 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_1_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mux_right_ipin_10.mux_l2_in_3__308 VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_10.mux_l2_in_3__308/HI
+ net308 sky130_fd_sc_hd__conb_1
Xcby_1__1_.mux_right_ipin_1.mux_l1_in_2_ net108 net77 cby_1__1_.mem_right_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_49_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_55_82 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__351
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__351/HI
+ net351 sky130_fd_sc_hd__conb_1
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__1_.mux_right_ipin_6.mux_l3_in_0_ cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_6.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_right_track_0.mux_l2_in_3_ net392 net4 sb_1__1_.mem_right_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_11.mux_l1_in_1_ sb_1__1_.mux_left_track_11.out net19 cbx_1__1_.mem_top_ipin_11.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_22_prog_clk sb_1__1_.mem_left_track_1.mem_out\[0\]
+ net296 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_1.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_82_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_52.mux_l3_in_0_ sb_1__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_right_track_0.ccff_head
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xwire1 clknet_1_1__leaf_clk0 VGND VGND VPWR VPWR net424 sky130_fd_sc_hd__buf_4
XFILLER_58_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_332_ sb_1__1_.mux_bottom_track_11.out VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__clkbuf_1
XFILLER_25_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_263_ sb_1__1_.mux_left_track_29.out VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_2
XFILLER_41_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_28 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_17 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_39 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput146 net146 VGND VGND VPWR VPWR bottom_width_0_height_0_subtile_0__pin_reg_out_0_
+ sky130_fd_sc_hd__buf_12
Xoutput157 net157 VGND VGND VPWR VPWR chanx_left_out[17] sky130_fd_sc_hd__buf_12
Xoutput168 net168 VGND VGND VPWR VPWR chanx_left_out[27] sky130_fd_sc_hd__buf_12
XFILLER_87_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput179 net179 VGND VGND VPWR VPWR chanx_right_out_0[0] sky130_fd_sc_hd__buf_12
XFILLER_87_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_33_prog_clk sb_1__1_.mem_right_track_12.ccff_tail
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_20.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_11_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_35_prog_clk sb_1__1_.mem_bottom_track_3.mem_out\[2\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_3.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_93_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_31_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mux_right_ipin_6.mux_l2_in_1_ cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_2_X cby_1__1_.mem_right_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
X_315_ sb_1__1_.mux_bottom_track_45.out VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__clkbuf_2
Xinput26 chanx_left_in[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__buf_4
Xinput15 chanx_left_in[20] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_2
Xinput37 chanx_right_in_0[13] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_4
Xinput48 chanx_right_in_0[23] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_4
Xinput59 chanx_right_in_0[6] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_4
Xsb_1__1_.mux_top_track_52.mux_l2_in_1_ net412 sb_1__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_top_track_52.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_20.mux_l3_in_0_ sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_right_track_20.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_20_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_1.mux_l2_in_3__415 VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_1.mux_l2_in_3__415/HI
+ net415 sky130_fd_sc_hd__conb_1
XFILLER_87_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_16_prog_clk sb_1__1_.mem_left_track_7.mem_out\[1\]
+ net296 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_7.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_right_track_0.mux_l4_in_0_ sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_9_X
+ sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_8_X sb_1__1_.mem_right_track_0.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_78_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mux_left_track_29.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_29.out sky130_fd_sc_hd__clkbuf_2
XFILLER_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_45.mux_l1_in_0_ net54 net97 sb_1__1_.mem_bottom_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xclkbuf_3_7__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_7__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_14_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_14_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_1_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_88_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_6.mux_l1_in_2_ sb_1__1_.mux_bottom_track_13.out net78 cby_1__1_.mem_right_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_88_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_top_track_52.mux_l1_in_2_ net5 net23 sb_1__1_.mem_top_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_71_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_right_track_20.mux_l2_in_1_ net71 sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_right_track_20.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_1.mux_l2_in_0_ cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_50_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_0_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mux_top_ipin_1.mux_l2_in_3_ net415 net58 cbx_1__1_.mem_top_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_28_prog_clk sb_1__1_.mem_top_track_0.ccff_tail
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_2.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_37_prog_clk sb_1__1_.mem_top_track_20.mem_out\[0\]
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_20.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_80_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_right_track_0.mux_l3_in_1_ sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_6_X sb_1__1_.mem_right_track_0.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_80_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_12.mux_l1_in_0_ sb_1__1_.mux_bottom_track_1.out net84 cby_1__1_.mem_right_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_12.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_5_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net350 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net364 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_22_prog_clk sb_1__1_.mem_left_track_29.mem_out\[1\]
+ net296 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_29.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_60_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_49_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_94_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_57_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_top_track_10.mux_l2_in_3_ net404 net28 sb_1__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_26_prog_clk sb_1__1_.mem_top_track_44.ccff_tail
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_52.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_107 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_118 net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_20.mux_l1_in_2_ net80 net132 sb_1__1_.mem_right_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__330
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__330/HI
+ net330 sky130_fd_sc_hd__conb_1
Xcby_1__1_.mux_right_ipin_1.mux_l1_in_1_ net111 net80 cby_1__1_.mem_right_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_1_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_left_track_29.mux_l2_in_3_ net385 net289 sb_1__1_.mem_left_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_39_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net335 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_right_track_0.mux_l2_in_2_ net21 net87 sb_1__1_.mem_right_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_11.mux_l1_in_0_ sb_1__1_.mux_left_track_5.out net22 cbx_1__1_.mem_top_ipin_11.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_38_prog_clk sb_1__1_.mem_bottom_track_53.ccff_tail
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_1.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_82_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mux_bottom_track_7.mux_l2_in_3__380 VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.mux_l2_in_3__380/HI
+ net380 sky130_fd_sc_hd__conb_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_46_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_331_ sb_1__1_.mux_bottom_track_13.out VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__clkbuf_2
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_262_ net39 VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__1_.mux_top_ipin_1.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_1.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_1_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_39_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_39_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_1__1_.mux_top_track_10.mux_l1_in_4_ net13 net88 sb_1__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_20_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_18 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_29 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput147 net147 VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__buf_12
Xoutput158 net158 VGND VGND VPWR VPWR chanx_left_out[18] sky130_fd_sc_hd__buf_12
XFILLER_87_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput169 net169 VGND VGND VPWR VPWR chanx_left_out[28] sky130_fd_sc_hd__buf_12
XFILLER_28_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_36_prog_clk sb_1__1_.mem_bottom_track_3.mem_out\[1\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_3.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_74_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_6.mux_l2_in_0_ cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_42_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_33_prog_clk cby_1__1_.ccff_tail net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_right_track_0.mux_l1_in_3_ net64 net81 sb_1__1_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_14_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_314_ net120 VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput27 chanx_left_in[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_2
Xinput16 chanx_left_in[21] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_4
XFILLER_6_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_6__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_6__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xinput38 chanx_right_in_0[14] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_4
Xinput49 chanx_right_in_0[24] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mux_top_track_52.mux_l2_in_0_ sb_1__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_top_track_52.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_top_track_10.mux_l4_in_0_ sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_10_X
+ sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_9_X sb_1__1_.mem_top_track_10.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_6_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_6.mux_l2_in_3_ net302 net59 cbx_1__1_.mem_top_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_left_track_29.mux_l4_in_0_ sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_6_X sb_1__1_.mem_left_track_29.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_87_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net361 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__mux2_2
XFILLER_83_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mux_top_ipin_1.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_17_prog_clk sb_1__1_.mem_left_track_7.mem_out\[0\]
+ net296 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_7.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
Xsb_1__1_.mux_right_track_20.mux_l2_in_3__396 VGND VGND VPWR VPWR sb_1__1_.mux_right_track_20.mux_l2_in_3__396/HI
+ net396 sky130_fd_sc_hd__conb_1
XFILLER_11_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_4.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_11_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_bottom_track_7.mux_l2_in_3_ net380 net29 sb_1__1_.mem_bottom_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ net424 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net124 grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_50_.in net134 VGND
+ VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_66_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_54_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_54_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_92_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mux_right_ipin_6.mux_l1_in_1_ sb_1__1_.mux_bottom_track_7.out net81 cby_1__1_.mem_right_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_10.mux_l3_in_1_ sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_top_track_10.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_71_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_top_track_52.mux_l1_in_1_ net65 net35 sb_1__1_.mem_top_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_71_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mux_top_ipin_6.mux_l1_in_4_ sb_1__1_.mux_left_track_37.out net5 cbx_1__1_.mem_top_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_8_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_right_track_20.mux_l2_in_0_ sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_right_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_47_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_29.mux_l3_in_1_ sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_4_X sb_1__1_.mem_left_track_29.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_0_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_1.mux_l2_in_2_ net27 net38 cbx_1__1_.mem_top_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_25_prog_clk sb_1__1_.mem_top_track_12.ccff_tail
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_20.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xsb_1__1_.mux_right_track_0.mux_l3_in_0_ sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X sb_1__1_.mem_right_track_0.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_27_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_80_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_bottom_track_7.mux_l1_in_4_ net19 net279 sb_1__1_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_6.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_9_X cbx_1__1_.mem_top_ipin_6.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_5.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_22_prog_clk sb_1__1_.mem_left_track_29.mem_out\[0\]
+ net296 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_29.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_5_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_57_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_bottom_track_7.mux_l4_in_0_ sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_10_X
+ sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_9_X sb_1__1_.mem_bottom_track_11.ccff_head
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_top_track_10.mux_l2_in_2_ net6 sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mem_top_track_10.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_108 net66 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_119 net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_41_prog_clk
+ sb_1__1_.mem_bottom_track_11.mem_out\[2\] net297 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_11.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_right_track_20.mux_l1_in_1_ net126 net115 sb_1__1_.mem_right_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_5_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_34_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_43_.in
+ sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_1.mux_l1_in_0_ sb_1__1_.mux_bottom_track_3.out net83 cby_1__1_.mem_right_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_1_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_left_track_29.mux_l2_in_2_ net74 net69 sb_1__1_.mem_left_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_45_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__dfrtp_1
XFILLER_76_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_right_track_0.mux_l2_in_1_ sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_right_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_82_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_59_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_46_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mux_top_ipin_6.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_6.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_23_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_76_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_9_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_9_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_44.out sky130_fd_sc_hd__clkbuf_1
XFILLER_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_330_ net108 VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__clkbuf_2
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_261_ net38 VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_41_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_5__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_5__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_1__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_33_prog_clk sb_1__1_.mem_right_track_12.mem_out\[2\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_12.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_2_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_7.mux_l3_in_1_ sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_bottom_track_7.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_10.mux_l1_in_3_ net73 net58 sb_1__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_19 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput148 net148 VGND VGND VPWR VPWR ccff_tail_0 sky130_fd_sc_hd__buf_12
Xoutput159 net159 VGND VGND VPWR VPWR chanx_left_out[19] sky130_fd_sc_hd__buf_12
XFILLER_55_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_left_track_5.mux_l2_in_3__389 VGND VGND VPWR VPWR sb_1__1_.mux_left_track_5.mux_l2_in_3__389/HI
+ net389 sky130_fd_sc_hd__conb_1
Xsb_1__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_41_prog_clk sb_1__1_.mem_bottom_track_3.mem_out\[0\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_3.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_46_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_43_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_0.mux_l1_in_2_ net131 net128 sb_1__1_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
X_313_ net119 VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput28 chanx_left_in[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_4
Xinput17 chanx_left_in[22] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_2
XFILLER_6_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput39 chanx_right_in_0[15] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_2
Xsb_1__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_33_prog_clk sb_1__1_.mem_right_track_44.mem_out\[1\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_44.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mux_top_ipin_6.mux_l2_in_2_ net28 cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mem_top_ipin_6.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mux_top_ipin_1.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X cbx_1__1_.mem_top_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_83_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_13_prog_clk sb_1__1_.mem_left_track_5.ccff_tail
+ net296 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_7.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_24_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_7.mux_l2_in_2_ net16 sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mem_bottom_track_7.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_93_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net339 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_23_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_23_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__1_.mux_right_ipin_6.mux_l1_in_0_ sb_1__1_.mux_bottom_track_1.out net84 cby_1__1_.mem_right_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_6.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_29_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_top_track_10.mux_l3_in_0_ sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_top_track_10.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_71_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_top_track_52.mux_l1_in_0_ net54 net138 sb_1__1_.mem_top_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_6.mux_l1_in_3_ net42 net11 cbx_1__1_.mem_top_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_left_track_29.mux_l3_in_0_ sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_left_track_29.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_3_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_86_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mux_top_ipin_1.mux_l2_in_1_ net7 cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__1_.mem_top_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_29_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_bottom_track_7.mux_l1_in_3_ net277 net275 sb_1__1_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_7.mux_l2_in_3_ net391 net293 sb_1__1_.mem_left_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_88_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_21_prog_clk sb_1__1_.mem_left_track_21.ccff_tail
+ net296 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_29.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_60_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_58_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_top_track_10.mux_l2_in_1_ sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_109 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_41_prog_clk
+ sb_1__1_.mem_bottom_track_11.mem_out\[1\] net297 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_11.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_4__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_4__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_1__1_.mux_right_track_20.mux_l1_in_0_ net101 net105 sb_1__1_.mem_right_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_52_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_61_.in
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_left_track_29.mux_l2_in_1_ net70 net44 sb_1__1_.mem_left_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_5.mux_l2_in_3__301 VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_5.mux_l2_in_3__301/HI
+ net301 sky130_fd_sc_hd__conb_1
XFILLER_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_45_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mux_top_ipin_1.mux_l1_in_2_ net48 net17 cbx_1__1_.mem_top_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_44_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_0.mux_l2_in_0_ sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_right_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net353 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_7.mux_l1_in_4_ net289 net287 sb_1__1_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_46_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mux_top_ipin_6.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_6.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_50_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_44.mux_l3_in_0_ sb_1__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_right_track_44.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_58_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_260_ net37 VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_2
XFILLER_2_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_32_prog_clk sb_1__1_.mem_right_track_12.mem_out\[1\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_12.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_2.out sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mux_bottom_track_7.mux_l3_in_0_ sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_bottom_track_7.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_7.mux_l4_in_0_ sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_10_X
+ sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_9_X sb_1__1_.mem_left_track_11.ccff_head
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_17_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_top_track_10.mux_l1_in_2_ net43 net45 sb_1__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_10.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput149 net149 VGND VGND VPWR VPWR chanx_left_out[0] sky130_fd_sc_hd__buf_12
Xclkbuf_leaf_48_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_48_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_83_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_32_prog_clk sb_1__1_.mem_right_track_0.mem_out\[2\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_70_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_40_prog_clk sb_1__1_.mem_bottom_track_1.ccff_tail
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_3.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_19_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_right_track_0.mux_l1_in_1_ net125 net93 sb_1__1_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
X_312_ net118 VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput18 chanx_left_in[23] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_4
Xinput29 chanx_left_in[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__buf_2
Xsb_1__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_33_prog_clk sb_1__1_.mem_right_track_44.mem_out\[0\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_44.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mux_top_ipin_6.mux_l2_in_1_ cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_2_X cbx_1__1_.mem_top_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_44.mux_l2_in_1_ net400 sb_1__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_right_track_44.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_44.mux_l2_in_1__411 VGND VGND VPWR VPWR sb_1__1_.mux_top_track_44.mux_l2_in_1__411/HI
+ net411 sky130_fd_sc_hd__conb_1
XFILLER_87_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ net424 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net124 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net134 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_50_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_bottom_track_7.mux_l2_in_1_ sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_bottom_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_7.mux_l3_in_1_ sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_left_track_7.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_3_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net343 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__mux2_4
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_18_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net296 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_left_track_29.mux_l2_in_3__385 VGND VGND VPWR VPWR sb_1__1_.mux_left_track_29.mux_l2_in_3__385/HI
+ net385 sky130_fd_sc_hd__conb_1
XFILLER_24_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_6.mux_l1_in_2_ sb_1__1_.mux_left_track_13.out net18 cbx_1__1_.mem_top_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_8_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_28_prog_clk sb_1__1_.mem_top_track_12.mem_out\[2\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_12.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_right_track_44.mux_l1_in_2_ net7 net67 sb_1__1_.mem_right_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_94_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_3_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mux_top_ipin_1.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_7_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_bottom_track_7.mux_l1_in_2_ net281 net59 sb_1__1_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_7.mux_l2_in_2_ net291 sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mem_left_track_7.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_3__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_3__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mux_right_ipin_13.mux_l2_in_3_ net311 net115 cby_1__1_.mem_right_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_0_clk0 clk0 VGND VGND VPWR VPWR clknet_0_clk0 sky130_fd_sc_hd__clkbuf_16
XFILLER_52_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_26_prog_clk sb_1__1_.mem_top_track_44.mem_out\[1\]
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_44.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_8_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_57_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_10.mux_l2_in_0_ sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_41_prog_clk
+ sb_1__1_.mem_bottom_track_11.mem_out\[0\] net297 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_11.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_53_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_70_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_79_.in
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_29.mux_l2_in_0_ sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_left_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_39_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_1.mux_l1_in_1_ net51 net20 cbx_1__1_.mem_top_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_71_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_left_track_7.mux_l1_in_3_ net89 net76 sb_1__1_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_90_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_46_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_50_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_12.mux_l2_in_3_ net418 net59 cbx_1__1_.mem_top_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_86_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_58_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_32_prog_clk sb_1__1_.mem_right_track_12.mem_out\[0\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_12.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_top_track_10.mux_l1_in_1_ net140 net138 sb_1__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_72_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_45_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_17_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_17_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_48_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mux_right_ipin_13.mux_l4_in_0_ cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_13.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_32_prog_clk sb_1__1_.mem_right_track_0.mem_out\[1\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_0.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_51_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_left_track_29.mux_l1_in_1_ net39 net104 sb_1__1_.mem_left_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_15.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l1_in_0_
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_70_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_right_track_0.mux_l1_in_0_ net94 net111 sb_1__1_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_14_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_311_ sb_1__1_.mux_bottom_track_53.out VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__clkbuf_2
Xinput19 chanx_left_in[24] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_2
XFILLER_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_33_prog_clk sb_1__1_.mem_right_track_36.ccff_tail
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_44.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xcbx_1__1_.mux_top_ipin_6.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_6.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_right_track_44.mux_l2_in_0_ sb_1__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_right_track_44.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__1_.mux_top_ipin_12.mux_l1_in_4_ sb_1__1_.mux_left_track_37.out net5 cbx_1__1_.mem_top_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_60_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_bottom_track_7.mux_l2_in_0_ sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_bottom_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_7.mux_l3_in_0_ sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_left_track_7.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_3_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_13.mux_l3_in_1_ cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_13.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_12.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_9_X cbx_1__1_.mem_top_ipin_12.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_2__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_2__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_21_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_32_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_32_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_16_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net296 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_68_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mux_top_ipin_6.mux_l1_in_1_ sb_1__1_.mux_left_track_7.out net21 cbx_1__1_.mem_top_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_8_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_25_prog_clk sb_1__1_.mem_top_track_12.mem_out\[1\]
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_12.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_3_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_32_prog_clk sb_1__1_.mem_right_track_6.mem_out\[2\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_10.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_right_track_44.mux_l1_in_1_ net84 net129 sb_1__1_.mem_right_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_94_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_3_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_70_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_7.mux_l1_in_1_ net40 net46 sb_1__1_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_80_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_left_track_7.mux_l2_in_1_ sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_left_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_21_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__326
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__326/HI
+ net326 sky130_fd_sc_hd__conb_1
XFILLER_95_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_13.out sky130_fd_sc_hd__clkbuf_2
XFILLER_44_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_12.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_12.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_13.mux_l2_in_2_ net74 net95 cby_1__1_.mem_right_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_44_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_59_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_26_prog_clk sb_1__1_.mem_top_track_44.mem_out\[0\]
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_44.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_4_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_55_prog_clk cby_1__1_.mem_right_ipin_2.mem_out\[2\]
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_left_track_5.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_5.out sky130_fd_sc_hd__buf_4
XFILLER_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_58_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__369
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__369/HI
+ net369 sky130_fd_sc_hd__conb_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_43_prog_clk
+ sb_1__1_.mem_bottom_track_11.ccff_head net297 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_11.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__carry_follower_0.sky130_fd_sc_hd__mux2_1_wrapper_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_88_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__mux2_1
XFILLER_41_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_1.mux_l1_in_0_ sb_1__1_.mux_left_track_3.out net23 cbx_1__1_.mem_top_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_55_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_4_prog_clk cbx_1__1_.mem_top_ipin_10.mem_out\[2\]
+ net295 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_10.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_71_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_2.mux_l2_in_3_ net314 sb_1__1_.mux_bottom_track_53.out cby_1__1_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_47_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_left_track_7.mux_l1_in_2_ net82 net59 sb_1__1_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_48_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_46_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_12.mux_l2_in_2_ net28 cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mem_top_ipin_12.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_48_prog_clk cby_1__1_.mem_right_ipin_12.mem_out\[2\]
+ net298 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_12.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_33_prog_clk sb_1__1_.mem_right_track_10.ccff_tail
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_12.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_89_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_10.mux_l1_in_0_ net136 net142 sb_1__1_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_17_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_46_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_43_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_32_prog_clk sb_1__1_.mem_right_track_0.mem_out\[0\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_0.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_57_prog_clk clknet_3_0__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_57_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_23_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_29.mux_l1_in_0_ net99 net109 sb_1__1_.mem_left_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_310_ net116 VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__clkbuf_2
Xcby_1__1_.mux_right_ipin_2.mux_l1_in_4_ net94 net92 cby_1__1_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_54_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__366
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__366/HI
+ net366 sky130_fd_sc_hd__conb_1
XFILLER_77_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_1__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_1__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_20_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__1_.mux_top_ipin_12.mux_l1_in_3_ net42 net11 cbx_1__1_.mem_top_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_60_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__1_.mux_right_ipin_2.mux_l4_in_0_ cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X cby_1__1_.mem_right_ipin_2.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_2_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_2_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcby_1__1_.mux_right_ipin_13.mux_l3_in_0_ cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_3_X cby_1__1_.mem_right_ipin_13.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_88_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__1_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_55_prog_clk cby_1__1_.mem_right_ipin_5.mem_out\[2\]
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_5.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_73_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_6.mux_l1_in_0_ sb_1__1_.mux_left_track_1.out net24 cbx_1__1_.mem_top_ipin_6.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_6.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_64_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_32_prog_clk sb_1__1_.mem_top_track_12.mem_out\[0\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_12.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
Xsb_1__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_33_prog_clk sb_1__1_.mem_right_track_6.mem_out\[1\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_6.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0_
+ net325 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__mux2_4
Xsb_1__1_.mux_right_track_44.mux_l1_in_0_ net121 net97 sb_1__1_.mem_right_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__1_.mux_right_ipin_7.mux_l2_in_3_ net319 sb_1__1_.mux_bottom_track_45.out cby_1__1_.mem_right_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xoutput290 net290 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_3_ sky130_fd_sc_hd__buf_12
XFILLER_58_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_4_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_62_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_2_prog_clk cbx_1__1_.mem_top_ipin_13.mem_out\[2\]
+ net295 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_13.ccff_tail sky130_fd_sc_hd__dfrtp_1
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_2.mux_l3_in_1_ cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_80_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_7.mux_l1_in_0_ net119 net106 sb_1__1_.mem_bottom_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_7.mux_l2_in_0_ sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_left_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_13.mux_l2_in_1_ net64 cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__1_.mem_right_ipin_13.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_12.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_12.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_52_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_25_prog_clk sb_1__1_.mem_top_track_36.ccff_tail
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_44.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_8_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_34_prog_clk cby_1__1_.mem_right_ipin_15.mem_out\[2\]
+ net297 VGND VGND VPWR VPWR cby_1__1_.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_69_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_13.mux_l2_in_3__419 VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_13.mux_l2_in_3__419/HI
+ net419 sky130_fd_sc_hd__conb_1
XFILLER_75_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_56_prog_clk cby_1__1_.mem_right_ipin_2.mem_out\[1\]
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_2.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_47_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_9.mux_l2_in_3__321 VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_9.mux_l2_in_3__321/HI
+ net321 sky130_fd_sc_hd__conb_1
XFILLER_75_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_1.mux_l2_in_3__307 VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_1.mux_l2_in_3__307/HI
+ net307 sky130_fd_sc_hd__conb_1
XFILLER_43_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_top_track_4.mux_l2_in_3_ net410 net27 sb_1__1_.mem_top_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_8.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_5_prog_clk cbx_1__1_.mem_top_ipin_10.mem_out\[1\]
+ net295 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_10.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_44_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_53.mux_l3_in_0_ sb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_bottom_track_53.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_47_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net298 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__1_.mux_right_ipin_2.mux_l2_in_2_ net86 cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mem_right_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_left_track_7.mux_l1_in_1_ net46 net119 sb_1__1_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_67_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_46_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_63_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_7.mux_l4_in_0_ cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_7.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_13.mux_l1_in_2_ net101 net70 cby_1__1_.mem_right_ipin_13.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_12.mux_l2_in_1_ cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_2_X cbx_1__1_.mem_top_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
Xcby_1__1_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_48_prog_clk cby_1__1_.mem_right_ipin_12.mem_out\[1\]
+ net298 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_12.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__333
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__333/HI
+ net333 sky130_fd_sc_hd__conb_1
XFILLER_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_0__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_0__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_32_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_46_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_27_prog_clk sb_1__1_.mem_right_track_0.ccff_head
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_0.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_49_prog_clk cby_1__1_.mem_right_ipin_8.mem_out\[2\]
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_8.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_26_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_26_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_1__1_.mux_right_track_52.mux_l2_in_1__401 VGND VGND VPWR VPWR sb_1__1_.mux_right_track_52.mux_l2_in_1__401/HI
+ net401 sky130_fd_sc_hd__conb_1
Xsb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_29.out sky130_fd_sc_hd__clkbuf_2
XFILLER_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_bottom_track_53.mux_l2_in_1_ net379 sb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_bottom_track_53.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_3.mux_l2_in_3__386 VGND VGND VPWR VPWR sb_1__1_.mux_left_track_3.mux_l2_in_3__386/HI
+ net386 sky130_fd_sc_hd__conb_1
Xcby_1__1_.mux_right_ipin_2.mux_l1_in_3_ sb_1__1_.mux_bottom_track_29.out net69 cby_1__1_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_14_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_left_track_13.mux_l2_in_3_ net383 net293 sb_1__1_.mem_left_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_top_track_4.mux_l4_in_0_ sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_top_track_4.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_6.mux_l2_in_3__318 VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_6.mux_l2_in_3__318/HI
+ net318 sky130_fd_sc_hd__conb_1
XFILLER_65_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__1_.mux_right_ipin_7.mux_l3_in_1_ cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_7.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_33_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_21.mux_l2_in_3__373 VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_21.mux_l2_in_3__373/HI
+ net373 sky130_fd_sc_hd__conb_1
XFILLER_26_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mux_top_ipin_12.mux_l1_in_2_ sb_1__1_.mux_left_track_13.out net18 cbx_1__1_.mem_top_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
X_369_ net297 VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__clkbuf_1
XFILLER_9_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_2.mux_l2_in_3__406 VGND VGND VPWR VPWR sb_1__1_.mux_top_track_2.mux_l2_in_3__406/HI
+ net406 sky130_fd_sc_hd__conb_1
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__1_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_55_prog_clk cby_1__1_.mem_right_ipin_5.mem_out\[1\]
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_5.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_33_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_53.mux_l1_in_2_ net5 net24 sb_1__1_.mem_bottom_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_56_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_4.mux_l3_in_1_ sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_top_track_4.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_41_prog_clk clknet_3_3__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_41_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_12_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_32_prog_clk sb_1__1_.mem_right_track_6.mem_out\[0\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_6.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
Xsb_1__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_31_prog_clk sb_1__1_.mem_top_track_10.ccff_tail
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_12.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xoutput280 net280 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_15_
+ sky130_fd_sc_hd__buf_12
Xcby_1__1_.mux_right_ipin_7.mux_l2_in_2_ net90 net101 cby_1__1_.mem_right_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xoutput291 net291 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_4_ sky130_fd_sc_hd__buf_12
XFILLER_59_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_6_prog_clk cbx_1__1_.mem_top_ipin_13.mem_out\[1\]
+ net295 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_13.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_11_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mux_right_ipin_2.mux_l3_in_0_ cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X cby_1__1_.mem_right_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_80_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_left_track_13.mux_l4_in_0_ sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_left_track_13.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_8_prog_clk cbx_1__1_.mem_top_ipin_2.mem_out\[2\]
+ net296 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_29_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net354 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__mux2_4
XFILLER_44_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__1_.mux_right_ipin_13.mux_l2_in_0_ cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_37_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_41_prog_clk cby_1__1_.mem_right_ipin_15.mem_out\[1\]
+ net297 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_15.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_69_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcby_1__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_56_prog_clk cby_1__1_.mem_right_ipin_2.mem_out\[0\]
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_2.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_75_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_bottom_track_11.mux_l2_in_3_ net371 net28 sb_1__1_.mem_bottom_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_47_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_58_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_top_track_4.mux_l2_in_2_ net30 net17 sb_1__1_.mem_top_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_32_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_16_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net296 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_6_prog_clk cbx_1__1_.mem_top_ipin_10.mem_out\[0\]
+ net295 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_10.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_40_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_2.mux_l2_in_1_ cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X cby_1__1_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_4_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_left_track_7.mux_l1_in_0_ net121 net106 sb_1__1_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_13.mux_l3_in_1_ sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_left_track_13.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_3_
+ clknet_leaf_47_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mux_right_ipin_13.mux_l1_in_1_ net111 net80 cby_1__1_.mem_right_ipin_13.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_12.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_12.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ net124 grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_59_.in net134 VGND
+ VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ sky130_fd_sc_hd__sdfrtp_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_51_prog_clk cby_1__1_.mem_right_ipin_12.mem_out\[0\]
+ net298 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_12.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_22_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_bottom_track_11.mux_l1_in_4_ net15 net280 sb_1__1_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_89_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net356 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_46_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_40_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_33_prog_clk sb_1__1_.mem_right_track_36.mem_out\[1\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_36.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_51_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_50_prog_clk cby_1__1_.mem_right_ipin_8.mem_out\[1\]
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_8.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_15_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net295 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_6.out sky130_fd_sc_hd__clkbuf_1
XFILLER_86_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_bottom_track_11.mux_l4_in_0_ sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_10_X
+ sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_9_X sb_1__1_.mem_bottom_track_11.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_bottom_track_53.mux_l2_in_0_ sb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_bottom_track_53.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__1_.mux_right_ipin_2.mux_l1_in_2_ net107 net76 cby_1__1_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_42_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_left_track_13.mux_l2_in_2_ net287 net86 sb_1__1_.mem_left_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_77_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_7.mux_l3_in_0_ cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_3_X cby_1__1_.mem_right_ipin_7.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__355
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__355/HI
+ net355 sky130_fd_sc_hd__conb_1
Xcbx_1__1_.mux_top_ipin_12.mux_l1_in_1_ sb_1__1_.mux_left_track_7.out net21 cbx_1__1_.mem_top_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_9_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_368_ net123 VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__clkbuf_1
XFILLER_41_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_299_ net17 VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_2
XFILLER_5_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_10_prog_clk cbx_1__1_.mem_top_ipin_5.mem_out\[2\]
+ net298 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_5.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_15_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__1_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_55_prog_clk cby_1__1_.mem_right_ipin_5.mem_out\[0\]
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_5.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_18_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_11.mux_l3_in_1_ sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_bottom_track_11.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_bottom_track_53.mux_l1_in_1_ net278 net33 sb_1__1_.mem_bottom_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_88_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_4.mux_l3_in_0_ sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_top_track_4.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_24_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_10_prog_clk clknet_3_4__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_10_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xsb_1__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_33_prog_clk sb_1__1_.mem_right_track_4.ccff_tail
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_6.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xcby_1__1_.mux_right_ipin_7.mux_l2_in_1_ net70 cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_2_X
+ cby_1__1_.mem_right_ipin_7.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xoutput270 net270 VGND VGND VPWR VPWR prog_reset_right_out sky130_fd_sc_hd__buf_12
XFILLER_79_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput292 net292 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_5_ sky130_fd_sc_hd__buf_12
Xoutput281 net281 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_8_ sky130_fd_sc_hd__buf_12
XFILLER_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_12.out sky130_fd_sc_hd__clkbuf_1
Xcbx_1__1_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_5_prog_clk cbx_1__1_.mem_top_ipin_13.mem_out\[0\]
+ net295 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_13.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_90_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_16_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net296 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_93_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_8_prog_clk cbx_1__1_.mem_top_ipin_2.mem_out\[1\]
+ net298 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_2.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_84_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_40_prog_clk cby_1__1_.mem_right_ipin_15.mem_out\[0\]
+ net298 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_15.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_4_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_55_prog_clk cby_1__1_.mem_right_ipin_1.ccff_tail
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_2.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_85_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_11.mux_l2_in_2_ net13 sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mem_bottom_track_11.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_top_track_4.mux_l2_in_1_ net90 sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_top_track_4.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_left_track_53.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_53.out sky130_fd_sc_hd__clkbuf_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_16_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ net296 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mux_right_ipin_7.mux_l1_in_2_ net108 net77 cby_1__1_.mem_right_ipin_7.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_39_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_410 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mem_top_ipin_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_10_prog_clk cbx_1__1_.mem_top_ipin_10.ccff_head
+ net298 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_10.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_13_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_6.mux_l2_in_3_ net402 net29 sb_1__1_.mem_right_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_2.mux_l2_in_0_ cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_20_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_left_track_13.mux_l3_in_0_ sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_left_track_13.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_0_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_2_
+ clknet_leaf_47_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mux_top_ipin_2.mux_l2_in_3_ net422 sb_1__1_.mux_left_track_53.out cbx_1__1_.mem_top_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_90_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcby_1__1_.mux_right_ipin_13.mux_l1_in_0_ sb_1__1_.mux_bottom_track_3.out net83 cby_1__1_.mem_right_ipin_13.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_13.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mem_right_ipin_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_49_prog_clk cby_1__1_.mem_right_ipin_11.ccff_tail
+ net298 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_12.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_11.mux_l1_in_3_ net278 net276 sb_1__1_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_3.mux_l2_in_3_ net375 net32 sb_1__1_.mem_bottom_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_44.out sky130_fd_sc_hd__clkbuf_1
Xcbx_1__1_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_11_prog_clk cbx_1__1_.mem_top_ipin_8.mem_out\[2\]
+ net295 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_8.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_72_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_4.mux_l1_in_2_ net77 net60 sb_1__1_.mem_top_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_9_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_13_
+ clknet_leaf_46_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_48_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_35_prog_clk sb_1__1_.mem_right_track_36.mem_out\[0\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_36.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_63_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcby_1__1_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_50_prog_clk cby_1__1_.mem_right_ipin_8.mem_out\[0\]
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_8.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_8_
+ clknet_leaf_15_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ net295 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_1_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_right_track_6.mux_l1_in_4_ net89 net70 sb_1__1_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_59_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_35_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_35_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_2.mux_l1_in_1_ sb_1__1_.mux_bottom_track_11.out net79 cby_1__1_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_left_track_1.mux_l2_in_3__381 VGND VGND VPWR VPWR sb_1__1_.mux_left_track_1.mux_l2_in_3__381/HI
+ net381 sky130_fd_sc_hd__conb_1
XFILLER_10_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_left_track_13.mux_l2_in_1_ net72 sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_left_track_13.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_2.mux_l1_in_4_ net34 net32 cbx_1__1_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_12.mux_l1_in_0_ sb_1__1_.mux_left_track_1.out net24 cbx_1__1_.mem_top_ipin_12.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_12.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_9_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_367_ sb_1__1_.mux_top_track_0.out VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_298_ net16 VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__clkbuf_2
XFILLER_68_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_right_track_6.mux_l4_in_0_ sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_10_X
+ sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_9_X sb_1__1_.mem_right_track_10.ccff_head
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_68_.in grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_6_prog_clk cbx_1__1_.mem_top_ipin_5.mem_out\[1\]
+ net295 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_5.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mux_top_ipin_2.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X cbx_1__1_.mem_top_ipin_2.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_67_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_10_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mem_right_ipin_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_55_prog_clk net423
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_5.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_58_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_11.mux_l3_in_0_ sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_bottom_track_11.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_bottom_track_53.mux_l1_in_0_ net35 net95 sb_1__1_.mem_bottom_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_88_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_3.mux_l4_in_0_ sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_9_X
+ sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_8_X sb_1__1_.mem_bottom_track_3.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_83_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_left_track_13.mux_l1_in_2_ net79 net56 sb_1__1_.mem_left_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_49_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__348
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__348/HI
+ net348 sky130_fd_sc_hd__conb_1
Xclkbuf_leaf_50_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_50_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcby_1__1_.mux_right_ipin_7.mux_l2_in_0_ cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_1_X
+ cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_0_X cby_1__1_.mem_right_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xoutput271 net271 VGND VGND VPWR VPWR prog_reset_top_out sky130_fd_sc_hd__buf_12
Xoutput260 net260 VGND VGND VPWR VPWR chany_top_out_0[29] sky130_fd_sc_hd__buf_12
Xoutput293 net293 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_6_ sky130_fd_sc_hd__buf_12
Xoutput282 net282 VGND VGND VPWR VPWR right_width_0_height_0_subtile_0__pin_O_9_ sky130_fd_sc_hd__buf_12
XFILLER_59_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_7.mux_l2_in_3_ net303 sb_1__1_.mux_left_track_45.out cbx_1__1_.mem_top_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mem_top_ipin_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_5_prog_clk cbx_1__1_.mem_top_ipin_12.ccff_tail
+ net295 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_13.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_30_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_right_track_6.mux_l3_in_1_ sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_8_X
+ sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_7_X sb_1__1_.mem_right_track_6.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_25_prog_clk sb_1__1_.mem_top_track_36.mem_out\[1\]
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_36.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_93_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_16_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net296 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__1_.mux_top_ipin_2.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__1_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_8_prog_clk cbx_1__1_.mem_top_ipin_2.mem_out\[0\]
+ net298 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_2.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_69_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mem_right_ipin_15.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_48_prog_clk cby_1__1_.mem_right_ipin_14.ccff_tail
+ net298 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_15.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_79_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_49_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_bottom_track_11.mux_l2_in_1_ sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_bottom_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_43_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_bottom_track_3.mux_l3_in_1_ sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_6_X sb_1__1_.mem_bottom_track_3.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_top_track_4.mux_l2_in_0_ sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_top_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0_
+ net345 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ sky130_fd_sc_hd__mux2_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_left_track_13.mux_l2_in_3__383 VGND VGND VPWR VPWR sb_1__1_.mux_left_track_13.mux_l2_in_3__383/HI
+ net383 sky130_fd_sc_hd__conb_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0_
+ net336 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__mux2_2
XFILLER_38_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_7.mux_l1_in_1_ net111 net80 cby_1__1_.mem_right_ipin_7.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_5.out sky130_fd_sc_hd__buf_4
XFILLER_13_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_6.mux_l2_in_2_ net16 sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mem_right_track_6.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_47_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.sky130_fd_sc_hd__sdfrtp_1_0_
+ clknet_1_0__leaf_clk0 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_1.ff_D
+ net124 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ net134 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.direct_interc_59_.in
+ sky130_fd_sc_hd__sdfrtp_1
XFILLER_29_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mux_top_ipin_2.mux_l2_in_2_ net26 cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mem_top_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1 chanx_right_in_0[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mux_top_ipin_7.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_7.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_66_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_22_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_bottom_track_11.mux_l1_in_2_ net282 net58 sb_1__1_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_89_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_bottom_track_3.mux_l2_in_2_ net18 net22 sb_1__1_.mem_bottom_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_57_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_28.out sky130_fd_sc_hd__clkbuf_1
XFILLER_17_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_11_prog_clk cbx_1__1_.mem_top_ipin_8.mem_out\[1\]
+ net295 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_8.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_72_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_top_track_4.mux_l1_in_1_ net47 net50 sb_1__1_.mem_top_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_9_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_12_
+ clknet_leaf_46_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_5_prog_clk clknet_3_1__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_5_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_35_prog_clk sb_1__1_.mem_right_track_28.ccff_tail
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_36.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_63_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mem_right_ipin_8.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_56_prog_clk cby_1__1_.mem_right_ipin_7.ccff_tail
+ net295 VGND VGND VPWR VPWR cby_1__1_.mem_right_ipin_8.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_7_
+ clknet_leaf_15_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ net296 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_50_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_1_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mux_right_track_6.mux_l1_in_3_ net76 net131 sb_1__1_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcby_1__1_.mux_right_ipin_2.mux_l1_in_0_ sb_1__1_.mux_bottom_track_5.out net82 cby_1__1_.mem_right_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_13.mux_l2_in_0_ sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_left_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_10_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_2.mux_l1_in_3_ sb_1__1_.mux_left_track_29.out net9 cbx_1__1_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_77_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_366_ sb_1__1_.mux_top_track_2.out VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__clkbuf_1
XFILLER_41_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_297_ sb_1__1_.mux_right_track_20.out VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__1_.mux_top_ipin_7.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_7.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[12\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_36_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_bottom_track_3.mux_l1_in_3_ net280 net277 sb_1__1_.mem_bottom_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_3.mux_l2_in_3_ net386 net294 sb_1__1_.mem_left_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_6_prog_clk cbx_1__1_.mem_top_ipin_5.mem_out\[0\]
+ net295 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_5.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_47_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net334 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_63_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_4_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_16_
+ clknet_leaf_43_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_53_prog_clk
+ sb_1__1_.mem_bottom_track_21.mem_out\[2\] net298 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_21.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_349_ sb_1__1_.mux_top_track_36.out VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__clkbuf_2
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_left_track_13.mux_l1_in_1_ net42 net116 sb_1__1_.mem_left_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_83_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput261 net261 VGND VGND VPWR VPWR chany_top_out_0[2] sky130_fd_sc_hd__buf_12
Xoutput250 net250 VGND VGND VPWR VPWR chany_top_out_0[1] sky130_fd_sc_hd__buf_12
Xoutput294 net294 VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_O_7_ sky130_fd_sc_hd__buf_12
Xoutput272 net272 VGND VGND VPWR VPWR reset_bottom_out sky130_fd_sc_hd__buf_12
Xoutput283 net283 VGND VGND VPWR VPWR sc_out sky130_fd_sc_hd__buf_12
XFILLER_58_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_7.mux_l2_in_2_ net30 net41 cbx_1__1_.mem_top_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_15_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_38_prog_clk
+ sb_1__1_.mem_bottom_track_53.mem_out\[1\] net298 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_53.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_X
+ sky130_fd_sc_hd__clkbuf_1
Xsb_1__1_.mux_right_track_6.mux_l3_in_0_ sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_6_X
+ sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_5_X sb_1__1_.mem_right_track_6.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_25_prog_clk sb_1__1_.mem_top_track_36.mem_out\[0\]
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_36.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_2.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_3_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_23_prog_clk cbx_1__1_.mem_top_ipin_1.ccff_tail
+ net296 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_2.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_88_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_71_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.ccff_tail
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_ VGND VGND VPWR
+ VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_X
+ sky130_fd_sc_hd__or2_1
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_49_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mux_bottom_track_11.mux_l2_in_0_ sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_bottom_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_3.mux_l3_in_0_ sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X sb_1__1_.mem_bottom_track_3.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_3.mux_l4_in_0_ sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_9_X
+ sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_8_X sb_1__1_.mem_left_track_3.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_3_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_7.mux_l1_in_0_ sb_1__1_.mux_bottom_track_3.out net83 cby_1__1_.mem_right_ipin_7.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_7.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_61_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_29_prog_clk clknet_3_7__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_29_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_30_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_29_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_right_track_6.mux_l2_in_1_ sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_right_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_80_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_44_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_75_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_49_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_48_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__1_.mux_top_ipin_2.mux_l2_in_1_ cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X cbx_1__1_.mem_top_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_bottom_track_45.mux_l2_in_1__377 VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_45.mux_l2_in_1__377/HI
+ net377 sky130_fd_sc_hd__conb_1
XFILLER_50_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_2 chanx_right_in_0[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_left_track_53.mux_l2_in_1__390 VGND VGND VPWR VPWR sb_1__1_.mux_left_track_53.mux_l2_in_1__390/HI
+ net390 sky130_fd_sc_hd__conb_1
XFILLER_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_11.mux_l1_in_1_ net43 net45 sb_1__1_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_1_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_bottom_track_3.mux_l2_in_1_ sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_bottom_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_3.mux_l3_in_1_ sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_6_X sb_1__1_.mem_left_track_3.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_17_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__1_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_10_prog_clk cbx_1__1_.mem_top_ipin_8.mem_out\[0\]
+ net295 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_8.mem_out\[1\] sky130_fd_sc_hd__dfrtp_2
Xsb_1__1_.mux_top_track_4.mux_l1_in_0_ net138 net135 sb_1__1_.mem_top_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_72_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_11_
+ clknet_leaf_46_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_0_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.direct_interc_11_.in
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_45_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_25_prog_clk sb_1__1_.mem_top_track_4.mem_out\[2\]
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_4.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_95_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_top_track_28.mux_l2_in_3_ net408 net14 sb_1__1_.mem_top_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_0_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_6_
+ clknet_leaf_15_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ net296 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_57_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__356
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0__356/HI
+ net356 sky130_fd_sc_hd__conb_1
Xsb_1__1_.mux_right_track_6.mux_l1_in_2_ net129 net127 sb_1__1_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_44_prog_clk clknet_3_2__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_44_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_2.mux_l1_in_2_ net47 net16 cbx_1__1_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_89_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_14.mux_l2_in_3__420 VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_14.mux_l2_in_3__420/HI
+ net420 sky130_fd_sc_hd__conb_1
XFILLER_60_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_365_ sb_1__1_.mux_top_track_4.out VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_296_ net13 VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__1_.mux_top_ipin_7.mux_l3_in_0_ cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_3_X cbx_1__1_.mem_top_ipin_7.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_right_track_28.mux_l2_in_3__397 VGND VGND VPWR VPWR sb_1__1_.mux_right_track_28.mux_l2_in_3__397/HI
+ net397 sky130_fd_sc_hd__conb_1
XFILLER_68_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[11\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_bottom_track_3.mux_l1_in_2_ net282 net61 sb_1__1_.mem_bottom_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_top_track_0.mux_l2_in_3__403 VGND VGND VPWR VPWR sb_1__1_.mux_top_track_0.mux_l2_in_3__403/HI
+ net403 sky130_fd_sc_hd__conb_1
Xsb_1__1_.mux_left_track_3.mux_l2_in_2_ net291 net288 sb_1__1_.mem_left_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mem_top_ipin_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_6_prog_clk cbx_1__1_.mem_top_ipin_4.ccff_tail
+ net295 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_5.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_59_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_15_
+ clknet_leaf_43_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_53_prog_clk
+ sb_1__1_.mem_bottom_track_21.mem_out\[1\] net298 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_21.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_18_prog_clk sb_1__1_.mem_left_track_3.mem_out\[2\]
+ net296 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_3.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_77_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_348_ net65 VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_495 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_279_ net25 VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__clkbuf_2
XFILLER_45_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_left_track_13.mux_l1_in_0_ net100 net102 sb_1__1_.mem_left_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput251 net251 VGND VGND VPWR VPWR chany_top_out_0[20] sky130_fd_sc_hd__buf_12
Xoutput262 net262 VGND VGND VPWR VPWR chany_top_out_0[3] sky130_fd_sc_hd__buf_12
Xoutput240 net240 VGND VGND VPWR VPWR chany_top_out_0[10] sky130_fd_sc_hd__buf_12
Xsb_1__1_.mux_top_track_28.mux_l4_in_0_ sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_7_X
+ sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_6_X sb_1__1_.mem_top_track_28.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_87_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput273 net273 VGND VGND VPWR VPWR reset_left_out sky130_fd_sc_hd__buf_12
Xoutput284 net284 VGND VGND VPWR VPWR test_enable_bottom_out sky130_fd_sc_hd__buf_12
XFILLER_59_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_7.mux_l2_in_1_ net10 cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_2_X
+ cbx_1__1_.mem_top_ipin_7.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_38_prog_clk
+ sb_1__1_.mem_bottom_track_53.mem_out\[0\] net298 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_53.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__337
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_1.mux_l2_in_0__337/HI
+ net337 sky130_fd_sc_hd__conb_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_top_track_20.mux_l2_in_3__407 VGND VGND VPWR VPWR sb_1__1_.mux_top_track_20.mux_l2_in_3__407/HI
+ net407 sky130_fd_sc_hd__conb_1
XFILLER_2_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_24_prog_clk sb_1__1_.mem_top_track_28.ccff_tail
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_36.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_37.mux_l3_in_0_ sb_1__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_left_track_37.ccff_tail
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_3.mux_l1_in_3_ net92 net78 sb_1__1_.mem_left_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_9_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut3_out\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out\[0\]
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_88_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0_ cbx_1__1_.mux_top_ipin_11.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_71_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mux_top_ipin_11.mux_l2_in_3__417 VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_11.mux_l2_in_3__417/HI
+ net417 sky130_fd_sc_hd__conb_1
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_2.mux_l2_in_3__422 VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_2.mux_l2_in_3__422/HI
+ net422 sky130_fd_sc_hd__conb_1
XFILLER_66_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_28.mux_l3_in_1_ sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_4_X sb_1__1_.mem_top_track_28.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_7_X sky130_fd_sc_hd__mux2_1
XFILLER_89_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mux_top_ipin_7.mux_l1_in_2_ net48 net17 cbx_1__1_.mem_top_ipin_7.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_27_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_57_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_right_track_6.mux_l2_in_0_ sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_right_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_37.mux_l2_in_1_ net387 sb_1__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_left_track_37.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_44_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ net297 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__1_.mux_top_ipin_2.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_90_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[2\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_3 chanx_right_in_0[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_5_.in
+ sky130_fd_sc_hd__clkbuf_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__360
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_fabric_out_0.mux_l2_in_0__360/HI
+ net360 sky130_fd_sc_hd__conb_1
XFILLER_62_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_6_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_right_track_52.mux_l3_in_0_ sb_1__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_3_X sb_1__1_.mem_bottom_track_1.ccff_head
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_bottom_track_11.mux_l1_in_0_ net118 net103 sb_1__1_.mem_bottom_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_3_ clknet_leaf_35_prog_clk sb_1__1_.mem_right_track_28.mem_out\[2\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_28.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xcby_1__1_.mux_right_ipin_14.mux_l2_in_3_ net312 sb_1__1_.mux_bottom_track_53.out
+ cby_1__1_.mem_right_ipin_14.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__1_.mux_bottom_track_3.mux_l2_in_0_ sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_bottom_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_66_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_left_track_3.mux_l3_in_0_ sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_4_X sb_1__1_.mem_left_track_3.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_57_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__1_.mem_top_ipin_8.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_12_prog_clk cbx_1__1_.mem_top_ipin_7.ccff_tail
+ net298 VGND VGND VPWR VPWR cbx_1__1_.mem_top_ipin_8.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_53_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_10_
+ clknet_leaf_46_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_25_prog_clk sb_1__1_.mem_top_track_4.mem_out\[1\]
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_4.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_leaf_45_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.ccff_tail
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__1_.mux_top_track_28.mux_l2_in_2_ net9 net19 sb_1__1_.mem_top_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_95_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput140 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_ VGND VGND VPWR
+ VPWR net140 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_5_
+ clknet_leaf_15_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ net296 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_right_track_6.mux_l1_in_1_ net125 net119 sb_1__1_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_86_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.mux_l2_in_0_
+ net326 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_0_D_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__ff_0.ff_D
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_left_track_37.mux_l1_in_2_ net290 net66 sb_1__1_.mem_left_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_22_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_13_prog_clk clknet_3_5__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_13_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xcbx_1__1_.mux_top_ipin_2.mux_l1_in_1_ sb_1__1_.mux_left_track_11.out net19 cbx_1__1_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_77_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_left_track_1.sky130_fd_sc_hd__buf_4_0_ sb_1__1_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_1.out sky130_fd_sc_hd__buf_4
XFILLER_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcby_1__1_.mux_right_ipin_4.mux_l2_in_3__316 VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_4.mux_l2_in_3__316/HI
+ net316 sky130_fd_sc_hd__conb_1
X_364_ sb_1__1_.mux_top_track_6.out VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__clkbuf_2
X_295_ net12 VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f_clk0 clknet_0_clk0 VGND VGND VPWR VPWR clknet_1_1__leaf_clk0 sky130_fd_sc_hd__clkbuf_16
XFILLER_5_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_76_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mux_right_track_52.mux_l2_in_1_ net401 sb_1__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__1_.mem_right_track_52.mem_out\[1\] VGND VGND VPWR VPWR sb_1__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcby_1__1_.mux_right_ipin_14.mux_l1_in_4_ net94 net92 cby_1__1_.mem_right_ipin_14.mem_out\[0\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xcbx_1__1_.mux_top_ipin_13.mux_l2_in_3_ net419 net55 cbx_1__1_.mem_top_ipin_13.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_32_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mux_bottom_track_3.mux_l1_in_1_ net62 net48 sb_1__1_.mem_bottom_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_left_track_3.mux_l2_in_1_ sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_left_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_67_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ net352 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_logic_out_0.out
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_14_
+ clknet_leaf_43_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[13\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_39_prog_clk
+ sb_1__1_.mem_bottom_track_21.mem_out\[0\] net298 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_21.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_12_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_19_prog_clk sb_1__1_.mem_left_track_3.mem_out\[1\]
+ net296 VGND VGND VPWR VPWR sb_1__1_.mem_left_track_3.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_12_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ sky130_fd_sc_hd__mux2_1
X_347_ net64 VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__clkbuf_2
Xcby_1__1_.mux_right_ipin_14.mux_l4_in_0_ cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_10_X
+ cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_9_X cby_1__1_.mem_right_ipin_14.ccff_tail
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
X_278_ net14 VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__clkbuf_2
XFILLER_38_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_9_
+ clknet_leaf_59_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[8\]
+ net123 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__363
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mux_ff_1_D_0.mux_l2_in_0__363/HI
+ net363 sky130_fd_sc_hd__conb_1
XFILLER_20_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput241 net241 VGND VGND VPWR VPWR chany_top_out_0[11] sky130_fd_sc_hd__buf_12
Xoutput252 net252 VGND VGND VPWR VPWR chany_top_out_0[21] sky130_fd_sc_hd__buf_12
Xoutput230 net230 VGND VGND VPWR VPWR chany_bottom_out[29] sky130_fd_sc_hd__buf_12
Xoutput274 net274 VGND VGND VPWR VPWR reset_top_out sky130_fd_sc_hd__buf_12
Xoutput285 net285 VGND VGND VPWR VPWR test_enable_left_out sky130_fd_sc_hd__buf_12
Xoutput263 net263 VGND VGND VPWR VPWR chany_top_out_0[4] sky130_fd_sc_hd__buf_12
XFILLER_87_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__1_.mux_top_ipin_7.mux_l2_in_0_ cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_0_X cbx_1__1_.mem_top_ipin_7.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_0_ clknet_leaf_38_prog_clk
+ sb_1__1_.mem_bottom_track_45.ccff_tail net298 VGND VGND VPWR VPWR sb_1__1_.mem_bottom_track_53.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_11_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_14_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.lut4_out
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.mux_l2_in_0_
+ net323 grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.sky130_fd_sc_hd__mux2_1_0_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.ccff_tail
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mux_frac_lut4_0_in_2.out
+ sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_right_track_52.mux_l1_in_2_ net5 net63 sb_1__1_.mem_right_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_left_track_3.mux_l1_in_2_ net84 net62 sb_1__1_.mem_left_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_9_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[15\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[14\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ cbx_1__1_.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_71_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_11_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_13_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcby_1__1_.mux_right_ipin_14.mux_l3_in_1_ cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_8_X
+ cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_7_X cby_1__1_.mem_right_ipin_14.mem_out\[2\]
+ VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_10_X sky130_fd_sc_hd__mux2_1
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__1_.mux_top_ipin_13.mux_l4_in_0_ cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_7_X cbx_1__1_.mem_top_ipin_13.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_9_X sky130_fd_sc_hd__mux2_1
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__1_.mux_top_track_28.mux_l3_in_0_ sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_2_X sb_1__1_.mem_top_track_28.mem_out\[2\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_89_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_1__1_.mux_top_ipin_7.mux_l1_in_1_ net51 net20 cbx_1__1_.mem_top_ipin_7.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_7.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_84_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_38_prog_clk clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR clknet_leaf_38_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_ VGND VGND VPWR VPWR
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_84_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__1_.mux_right_track_10.mux_l2_in_3_ net393 net28 sb_1__1_.mem_right_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
XFILLER_13_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_left_track_37.mux_l2_in_0_ sb_1__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_0_X sb_1__1_.mem_left_track_37.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_0_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[1\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[0\]
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_4 chanx_right_in_0[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_ cby_1__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ VGND VGND VPWR VPWR cby_1__1_.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_
+ sky130_fd_sc_hd__clkbuf_1
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.direct_interc_7_.in
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.sky130_fd_sc_hd__dfrtp_1_1_
+ clknet_leaf_11_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out\[0\]
+ net295 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_5_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_4_X
+ grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_X
+ VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_2_ clknet_leaf_36_prog_clk sb_1__1_.mem_right_track_28.mem_out\[1\]
+ net297 VGND VGND VPWR VPWR sb_1__1_.mem_right_track_28.mem_out\[2\] sky130_fd_sc_hd__dfrtp_1
Xcbx_1__1_.mux_top_ipin_13.mux_l3_in_1_ cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_5_X cbx_1__1_.mem_top_ipin_13.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__1_.mux_top_ipin_13.sky130_fd_sc_hd__mux2_1_8_X sky130_fd_sc_hd__mux2_1
Xcby_1__1_.mux_right_ipin_14.mux_l2_in_2_ net86 cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_4_X
+ cby_1__1_.mem_right_ipin_14.mem_out\[1\] VGND VGND VPWR VPWR cby_1__1_.mux_right_ipin_14.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_leaf_25_prog_clk sb_1__1_.mem_top_track_4.mem_out\[0\]
+ net298 VGND VGND VPWR VPWR sb_1__1_.mem_top_track_4.mem_out\[1\] sky130_fd_sc_hd__dfrtp_4
Xsb_1__1_.mux_top_track_28.mux_l2_in_1_ net74 net69 sb_1__1_.mem_top_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xinput141 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_ VGND VGND VPWR
+ VPWR net141 sky130_fd_sc_hd__clkbuf_1
Xinput130 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_ VGND VGND VPWR
+ VPWR net130 sky130_fd_sc_hd__clkbuf_2
XFILLER_29_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xgrid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_4_
+ clknet_leaf_15_prog_clk grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[3\]
+ net296 VGND VGND VPWR VPWR grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__1_.mux_right_track_10.mux_l1_in_4_ net88 net73 sb_1__1_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xsb_1__1_.mux_right_track_6.mux_l1_in_0_ net106 net112 sb_1__1_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_86_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
.ends

