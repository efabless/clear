magic
tech sky130A
magscale 1 2
timestamp 1656943399
<< viali >>
rect 4537 20009 4571 20043
rect 5641 20009 5675 20043
rect 7389 19873 7423 19907
rect 4721 19805 4755 19839
rect 5825 19805 5859 19839
rect 7665 19805 7699 19839
rect 4537 19465 4571 19499
rect 8585 19397 8619 19431
rect 4721 19329 4755 19363
rect 8861 19329 8895 19363
rect 4629 18921 4663 18955
rect 4813 18717 4847 18751
rect 4813 18377 4847 18411
rect 4997 18241 5031 18275
rect 1961 17833 1995 17867
rect 3985 17833 4019 17867
rect 4721 17833 4755 17867
rect 7113 17697 7147 17731
rect 2145 17629 2179 17663
rect 4169 17629 4203 17663
rect 4905 17629 4939 17663
rect 7389 17629 7423 17663
rect 1593 17289 1627 17323
rect 3709 17289 3743 17323
rect 2237 17221 2271 17255
rect 7481 17221 7515 17255
rect 1777 17153 1811 17187
rect 2513 17153 2547 17187
rect 3893 17153 3927 17187
rect 5181 17153 5215 17187
rect 5457 17153 5491 17187
rect 7757 17153 7791 17187
rect 9413 16609 9447 16643
rect 9597 16609 9631 16643
rect 10517 16609 10551 16643
rect 4445 16541 4479 16575
rect 4721 16541 4755 16575
rect 6193 16541 6227 16575
rect 6469 16541 6503 16575
rect 7205 16541 7239 16575
rect 7665 16541 7699 16575
rect 7941 16541 7975 16575
rect 6929 16473 6963 16507
rect 8953 16405 8987 16439
rect 9321 16405 9355 16439
rect 9965 16405 9999 16439
rect 1961 16201 1995 16235
rect 2145 16065 2179 16099
rect 5181 15861 5215 15895
rect 1685 15657 1719 15691
rect 2789 15657 2823 15691
rect 5917 15657 5951 15691
rect 7297 15657 7331 15691
rect 2237 15589 2271 15623
rect 4537 15521 4571 15555
rect 5365 15521 5399 15555
rect 7941 15521 7975 15555
rect 1869 15453 1903 15487
rect 2421 15453 2455 15487
rect 2973 15453 3007 15487
rect 4813 15453 4847 15487
rect 5641 15453 5675 15487
rect 7665 15385 7699 15419
rect 8309 15385 8343 15419
rect 7757 15317 7791 15351
rect 4261 15113 4295 15147
rect 4721 15113 4755 15147
rect 5273 15113 5307 15147
rect 6929 15113 6963 15147
rect 2973 15045 3007 15079
rect 3709 15045 3743 15079
rect 2145 14977 2179 15011
rect 3249 14977 3283 15011
rect 3985 14977 4019 15011
rect 4629 14977 4663 15011
rect 5641 14977 5675 15011
rect 7297 14977 7331 15011
rect 7941 14977 7975 15011
rect 4813 14909 4847 14943
rect 5733 14909 5767 14943
rect 5825 14909 5859 14943
rect 7389 14909 7423 14943
rect 7573 14909 7607 14943
rect 1961 14773 1995 14807
rect 6377 14773 6411 14807
rect 1501 14569 1535 14603
rect 9321 14569 9355 14603
rect 3801 14501 3835 14535
rect 2145 14433 2179 14467
rect 4445 14433 4479 14467
rect 9965 14433 9999 14467
rect 1685 14365 1719 14399
rect 2421 14365 2455 14399
rect 3433 14365 3467 14399
rect 8953 14365 8987 14399
rect 9781 14365 9815 14399
rect 12449 14365 12483 14399
rect 3157 14297 3191 14331
rect 4169 14229 4203 14263
rect 4261 14229 4295 14263
rect 4813 14229 4847 14263
rect 5457 14229 5491 14263
rect 6193 14229 6227 14263
rect 8493 14229 8527 14263
rect 9689 14229 9723 14263
rect 11161 14229 11195 14263
rect 11713 14229 11747 14263
rect 12817 14229 12851 14263
rect 1961 14025 1995 14059
rect 2605 14025 2639 14059
rect 4077 14025 4111 14059
rect 4905 14025 4939 14059
rect 7941 14025 7975 14059
rect 8309 14025 8343 14059
rect 9413 14025 9447 14059
rect 10425 14025 10459 14059
rect 10793 14025 10827 14059
rect 11529 14025 11563 14059
rect 12541 14025 12575 14059
rect 12909 14025 12943 14059
rect 5365 13957 5399 13991
rect 7665 13957 7699 13991
rect 9873 13957 9907 13991
rect 11897 13957 11931 13991
rect 13001 13957 13035 13991
rect 2145 13889 2179 13923
rect 2421 13889 2455 13923
rect 3617 13889 3651 13923
rect 3709 13889 3743 13923
rect 4353 13889 4387 13923
rect 5273 13889 5307 13923
rect 8401 13889 8435 13923
rect 9781 13889 9815 13923
rect 10885 13889 10919 13923
rect 3525 13821 3559 13855
rect 5549 13821 5583 13855
rect 5917 13821 5951 13855
rect 6653 13821 6687 13855
rect 8585 13821 8619 13855
rect 9045 13821 9079 13855
rect 10057 13821 10091 13855
rect 11069 13821 11103 13855
rect 11989 13821 12023 13855
rect 12173 13821 12207 13855
rect 13185 13821 13219 13855
rect 2973 13685 3007 13719
rect 4169 13481 4203 13515
rect 7757 13481 7791 13515
rect 12081 13481 12115 13515
rect 6837 13413 6871 13447
rect 10241 13413 10275 13447
rect 1961 13345 1995 13379
rect 3157 13345 3191 13379
rect 4813 13345 4847 13379
rect 5365 13345 5399 13379
rect 6285 13345 6319 13379
rect 6469 13345 6503 13379
rect 8217 13345 8251 13379
rect 8309 13345 8343 13379
rect 9781 13345 9815 13379
rect 10885 13345 10919 13379
rect 12725 13345 12759 13379
rect 3433 13277 3467 13311
rect 6193 13277 6227 13311
rect 9505 13277 9539 13311
rect 12449 13277 12483 13311
rect 2145 13209 2179 13243
rect 3893 13209 3927 13243
rect 8125 13209 8159 13243
rect 8953 13209 8987 13243
rect 11345 13209 11379 13243
rect 12541 13209 12575 13243
rect 1409 13141 1443 13175
rect 2053 13141 2087 13175
rect 2513 13141 2547 13175
rect 4537 13141 4571 13175
rect 4629 13141 4663 13175
rect 5825 13141 5859 13175
rect 7297 13141 7331 13175
rect 10609 13141 10643 13175
rect 10701 13141 10735 13175
rect 11805 13141 11839 13175
rect 2697 12937 2731 12971
rect 5641 12937 5675 12971
rect 7389 12937 7423 12971
rect 7757 12937 7791 12971
rect 11713 12937 11747 12971
rect 12173 12937 12207 12971
rect 2053 12869 2087 12903
rect 1777 12801 1811 12835
rect 2513 12801 2547 12835
rect 3525 12801 3559 12835
rect 7849 12801 7883 12835
rect 10149 12801 10183 12835
rect 10793 12801 10827 12835
rect 12541 12801 12575 12835
rect 13185 12801 13219 12835
rect 3249 12733 3283 12767
rect 5733 12733 5767 12767
rect 5825 12733 5859 12767
rect 7113 12733 7147 12767
rect 8033 12733 8067 12767
rect 9413 12733 9447 12767
rect 9965 12733 9999 12767
rect 10057 12733 10091 12767
rect 12633 12733 12667 12767
rect 12817 12733 12851 12767
rect 10517 12665 10551 12699
rect 1501 12597 1535 12631
rect 4997 12597 5031 12631
rect 5273 12597 5307 12631
rect 6561 12597 6595 12631
rect 8401 12597 8435 12631
rect 9137 12597 9171 12631
rect 1685 12393 1719 12427
rect 4353 12393 4387 12427
rect 5825 12393 5859 12427
rect 6837 12393 6871 12427
rect 9321 12393 9355 12427
rect 2329 12257 2363 12291
rect 4997 12257 5031 12291
rect 6469 12257 6503 12291
rect 7297 12257 7331 12291
rect 7481 12257 7515 12291
rect 8493 12257 8527 12291
rect 9873 12257 9907 12291
rect 10885 12257 10919 12291
rect 1869 12189 1903 12223
rect 4813 12189 4847 12223
rect 6193 12189 6227 12223
rect 7205 12189 7239 12223
rect 8309 12189 8343 12223
rect 9045 12189 9079 12223
rect 10793 12189 10827 12223
rect 11805 12189 11839 12223
rect 17049 12189 17083 12223
rect 2421 12121 2455 12155
rect 9689 12121 9723 12155
rect 11345 12121 11379 12155
rect 12050 12121 12084 12155
rect 16804 12121 16838 12155
rect 2513 12053 2547 12087
rect 2881 12053 2915 12087
rect 3157 12053 3191 12087
rect 3985 12053 4019 12087
rect 4721 12053 4755 12087
rect 5365 12053 5399 12087
rect 6285 12053 6319 12087
rect 7849 12053 7883 12087
rect 8217 12053 8251 12087
rect 9781 12053 9815 12087
rect 10333 12053 10367 12087
rect 10701 12053 10735 12087
rect 13185 12053 13219 12087
rect 13553 12053 13587 12087
rect 15669 12053 15703 12087
rect 17417 12053 17451 12087
rect 19901 12053 19935 12087
rect 21373 12053 21407 12087
rect 2513 11849 2547 11883
rect 3341 11849 3375 11883
rect 4353 11849 4387 11883
rect 4997 11849 5031 11883
rect 5365 11849 5399 11883
rect 5457 11849 5491 11883
rect 6377 11849 6411 11883
rect 6837 11849 6871 11883
rect 7757 11849 7791 11883
rect 8217 11849 8251 11883
rect 8769 11849 8803 11883
rect 9781 11849 9815 11883
rect 15577 11849 15611 11883
rect 19993 11849 20027 11883
rect 1593 11781 1627 11815
rect 16926 11781 16960 11815
rect 18604 11781 18638 11815
rect 1869 11713 1903 11747
rect 6745 11713 6779 11747
rect 8125 11713 8159 11747
rect 9137 11713 9171 11747
rect 10905 11713 10939 11747
rect 12348 11713 12382 11747
rect 14197 11713 14231 11747
rect 14453 11713 14487 11747
rect 15945 11713 15979 11747
rect 16313 11713 16347 11747
rect 16681 11713 16715 11747
rect 21106 11713 21140 11747
rect 21373 11713 21407 11747
rect 2605 11645 2639 11679
rect 2697 11645 2731 11679
rect 3709 11645 3743 11679
rect 4445 11645 4479 11679
rect 4629 11645 4663 11679
rect 5641 11645 5675 11679
rect 7021 11645 7055 11679
rect 8401 11645 8435 11679
rect 9229 11645 9263 11679
rect 9413 11645 9447 11679
rect 11161 11645 11195 11679
rect 11529 11645 11563 11679
rect 12081 11645 12115 11679
rect 18337 11645 18371 11679
rect 3985 11577 4019 11611
rect 2145 11509 2179 11543
rect 7389 11509 7423 11543
rect 13461 11509 13495 11543
rect 13737 11509 13771 11543
rect 18061 11509 18095 11543
rect 19717 11509 19751 11543
rect 1777 11305 1811 11339
rect 3341 11305 3375 11339
rect 4537 11305 4571 11339
rect 7573 11305 7607 11339
rect 12081 11305 12115 11339
rect 17509 11305 17543 11339
rect 19349 11305 19383 11339
rect 21097 11305 21131 11339
rect 5549 11237 5583 11271
rect 7849 11237 7883 11271
rect 14473 11237 14507 11271
rect 2237 11169 2271 11203
rect 2421 11169 2455 11203
rect 4997 11169 5031 11203
rect 5181 11169 5215 11203
rect 6193 11169 6227 11203
rect 6745 11169 6779 11203
rect 8401 11169 8435 11203
rect 8953 11169 8987 11203
rect 20729 11169 20763 11203
rect 5917 11101 5951 11135
rect 8217 11101 8251 11135
rect 8309 11101 8343 11135
rect 9781 11101 9815 11135
rect 10701 11101 10735 11135
rect 13470 11101 13504 11135
rect 13737 11101 13771 11135
rect 15853 11101 15887 11135
rect 16129 11101 16163 11135
rect 16385 11101 16419 11135
rect 20462 11101 20496 11135
rect 1409 11033 1443 11067
rect 9413 11033 9447 11067
rect 10149 11033 10183 11067
rect 10946 11033 10980 11067
rect 15586 11033 15620 11067
rect 17877 11033 17911 11067
rect 2145 10965 2179 10999
rect 2789 10965 2823 10999
rect 3893 10965 3927 10999
rect 4905 10965 4939 10999
rect 6009 10965 6043 10999
rect 12357 10965 12391 10999
rect 14197 10965 14231 10999
rect 18153 10965 18187 10999
rect 18521 10965 18555 10999
rect 1961 10761 1995 10795
rect 2329 10761 2363 10795
rect 3893 10761 3927 10795
rect 4261 10761 4295 10795
rect 5457 10761 5491 10795
rect 7205 10761 7239 10795
rect 8953 10761 8987 10795
rect 10057 10761 10091 10795
rect 16681 10761 16715 10795
rect 18337 10761 18371 10795
rect 2421 10693 2455 10727
rect 3801 10693 3835 10727
rect 14228 10693 14262 10727
rect 5089 10625 5123 10659
rect 7297 10625 7331 10659
rect 7941 10625 7975 10659
rect 9597 10625 9631 10659
rect 15862 10625 15896 10659
rect 17794 10625 17828 10659
rect 18061 10625 18095 10659
rect 19450 10625 19484 10659
rect 19717 10625 19751 10659
rect 21106 10625 21140 10659
rect 21373 10625 21407 10659
rect 2605 10557 2639 10591
rect 3709 10557 3743 10591
rect 4905 10557 4939 10591
rect 4997 10557 5031 10591
rect 7113 10557 7147 10591
rect 8769 10557 8803 10591
rect 8861 10557 8895 10591
rect 14473 10557 14507 10591
rect 16129 10557 16163 10591
rect 3249 10489 3283 10523
rect 9321 10489 9355 10523
rect 19993 10489 20027 10523
rect 5733 10421 5767 10455
rect 6561 10421 6595 10455
rect 7665 10421 7699 10455
rect 12265 10421 12299 10455
rect 13093 10421 13127 10455
rect 14749 10421 14783 10455
rect 2697 10217 2731 10251
rect 3433 10217 3467 10251
rect 6193 10217 6227 10251
rect 7481 10217 7515 10251
rect 8953 10217 8987 10251
rect 12449 10217 12483 10251
rect 14657 10217 14691 10251
rect 16221 10217 16255 10251
rect 17325 10217 17359 10251
rect 21005 10217 21039 10251
rect 21373 10217 21407 10251
rect 5089 10081 5123 10115
rect 5549 10081 5583 10115
rect 8401 10081 8435 10115
rect 9505 10081 9539 10115
rect 10333 10081 10367 10115
rect 10793 10081 10827 10115
rect 3801 10013 3835 10047
rect 4813 10013 4847 10047
rect 5733 10013 5767 10047
rect 8217 10013 8251 10047
rect 18705 10013 18739 10047
rect 19257 10013 19291 10047
rect 6745 9945 6779 9979
rect 8309 9945 8343 9979
rect 11060 9945 11094 9979
rect 18438 9945 18472 9979
rect 19502 9945 19536 9979
rect 2973 9877 3007 9911
rect 3985 9877 4019 9911
rect 4445 9877 4479 9911
rect 4905 9877 4939 9911
rect 5825 9877 5859 9911
rect 7113 9877 7147 9911
rect 7849 9877 7883 9911
rect 9321 9877 9355 9911
rect 9413 9877 9447 9911
rect 9965 9877 9999 9911
rect 12173 9877 12207 9911
rect 20637 9877 20671 9911
rect 6377 9673 6411 9707
rect 10885 9673 10919 9707
rect 11529 9673 11563 9707
rect 19349 9673 19383 9707
rect 21373 9673 21407 9707
rect 6837 9605 6871 9639
rect 9873 9605 9907 9639
rect 12642 9605 12676 9639
rect 20462 9605 20496 9639
rect 3893 9537 3927 9571
rect 4997 9537 5031 9571
rect 6745 9537 6779 9571
rect 7757 9537 7791 9571
rect 8401 9537 8435 9571
rect 9137 9537 9171 9571
rect 9781 9537 9815 9571
rect 10793 9537 10827 9571
rect 18162 9537 18196 9571
rect 18429 9537 18463 9571
rect 18797 9537 18831 9571
rect 20729 9537 20763 9571
rect 3985 9469 4019 9503
rect 4077 9469 4111 9503
rect 5089 9469 5123 9503
rect 5273 9469 5307 9503
rect 6929 9469 6963 9503
rect 7849 9469 7883 9503
rect 8033 9469 8067 9503
rect 10057 9469 10091 9503
rect 11069 9469 11103 9503
rect 12909 9469 12943 9503
rect 3525 9401 3559 9435
rect 7389 9401 7423 9435
rect 17049 9401 17083 9435
rect 3157 9333 3191 9367
rect 4629 9333 4663 9367
rect 5917 9333 5951 9367
rect 9413 9333 9447 9367
rect 10425 9333 10459 9367
rect 13277 9333 13311 9367
rect 3249 9129 3283 9163
rect 4261 9129 4295 9163
rect 15945 9129 15979 9163
rect 19717 9129 19751 9163
rect 2237 9061 2271 9095
rect 6101 9061 6135 9095
rect 2697 8993 2731 9027
rect 4721 8993 4755 9027
rect 4905 8993 4939 9027
rect 6929 8993 6963 9027
rect 8033 8993 8067 9027
rect 21097 8993 21131 9027
rect 2789 8925 2823 8959
rect 4629 8925 4663 8959
rect 7757 8925 7791 8959
rect 8953 8925 8987 8959
rect 10894 8925 10928 8959
rect 11161 8925 11195 8959
rect 12817 8925 12851 8959
rect 15310 8925 15344 8959
rect 15577 8925 15611 8959
rect 17325 8925 17359 8959
rect 17693 8925 17727 8959
rect 18245 8925 18279 8959
rect 18613 8925 18647 8959
rect 19441 8925 19475 8959
rect 3893 8857 3927 8891
rect 7849 8857 7883 8891
rect 12550 8857 12584 8891
rect 17080 8857 17114 8891
rect 20830 8857 20864 8891
rect 2881 8789 2915 8823
rect 5365 8789 5399 8823
rect 6653 8789 6687 8823
rect 7389 8789 7423 8823
rect 8401 8789 8435 8823
rect 9505 8789 9539 8823
rect 9781 8789 9815 8823
rect 11437 8789 11471 8823
rect 13185 8789 13219 8823
rect 14197 8789 14231 8823
rect 2789 8585 2823 8619
rect 3525 8585 3559 8619
rect 5273 8585 5307 8619
rect 7481 8585 7515 8619
rect 9781 8585 9815 8619
rect 11161 8585 11195 8619
rect 13369 8585 13403 8619
rect 15761 8585 15795 8619
rect 18061 8585 18095 8619
rect 21373 8585 21407 8619
rect 5365 8517 5399 8551
rect 20238 8517 20272 8551
rect 4261 8449 4295 8483
rect 6837 8449 6871 8483
rect 8493 8449 8527 8483
rect 12826 8449 12860 8483
rect 14482 8449 14516 8483
rect 14749 8449 14783 8483
rect 15117 8449 15151 8483
rect 16681 8449 16715 8483
rect 16937 8449 16971 8483
rect 18337 8449 18371 8483
rect 18593 8449 18627 8483
rect 19993 8449 20027 8483
rect 4353 8381 4387 8415
rect 4445 8381 4479 8415
rect 5457 8381 5491 8415
rect 7573 8381 7607 8415
rect 7665 8381 7699 8415
rect 8585 8381 8619 8415
rect 8769 8381 8803 8415
rect 9873 8381 9907 8415
rect 10057 8381 10091 8415
rect 13093 8381 13127 8415
rect 3893 8313 3927 8347
rect 5917 8313 5951 8347
rect 7113 8313 7147 8347
rect 8125 8313 8159 8347
rect 11713 8313 11747 8347
rect 19717 8313 19751 8347
rect 4905 8245 4939 8279
rect 9413 8245 9447 8279
rect 4169 8041 4203 8075
rect 6837 8041 6871 8075
rect 7205 8041 7239 8075
rect 8493 8041 8527 8075
rect 10057 8041 10091 8075
rect 11345 8041 11379 8075
rect 15669 8041 15703 8075
rect 17325 8041 17359 8075
rect 17693 8041 17727 8075
rect 20913 8041 20947 8075
rect 21281 8041 21315 8075
rect 18153 7973 18187 8007
rect 4629 7905 4663 7939
rect 4813 7905 4847 7939
rect 5365 7905 5399 7939
rect 7665 7905 7699 7939
rect 7849 7905 7883 7939
rect 9505 7905 9539 7939
rect 15945 7905 15979 7939
rect 19257 7905 19291 7939
rect 6469 7837 6503 7871
rect 7573 7837 7607 7871
rect 9689 7837 9723 7871
rect 12725 7837 12759 7871
rect 13277 7837 13311 7871
rect 13645 7837 13679 7871
rect 14289 7837 14323 7871
rect 3433 7769 3467 7803
rect 5549 7769 5583 7803
rect 12480 7769 12514 7803
rect 14534 7769 14568 7803
rect 16212 7769 16246 7803
rect 19524 7769 19558 7803
rect 3065 7701 3099 7735
rect 3893 7701 3927 7735
rect 4537 7701 4571 7735
rect 5457 7701 5491 7735
rect 5917 7701 5951 7735
rect 9045 7701 9079 7735
rect 9597 7701 9631 7735
rect 20637 7701 20671 7735
rect 2421 7497 2455 7531
rect 4445 7497 4479 7531
rect 5089 7497 5123 7531
rect 7113 7497 7147 7531
rect 7573 7497 7607 7531
rect 11529 7497 11563 7531
rect 15301 7497 15335 7531
rect 15761 7497 15795 7531
rect 16129 7497 16163 7531
rect 17417 7497 17451 7531
rect 19073 7497 19107 7531
rect 20729 7497 20763 7531
rect 21097 7497 21131 7531
rect 3433 7429 3467 7463
rect 3985 7429 4019 7463
rect 5733 7429 5767 7463
rect 14166 7429 14200 7463
rect 1869 7361 1903 7395
rect 4077 7361 4111 7395
rect 6837 7361 6871 7395
rect 7481 7361 7515 7395
rect 8585 7361 8619 7395
rect 12642 7361 12676 7395
rect 12909 7361 12943 7395
rect 13277 7361 13311 7395
rect 13921 7361 13955 7395
rect 18530 7361 18564 7395
rect 18797 7361 18831 7395
rect 20186 7361 20220 7395
rect 20453 7361 20487 7395
rect 3893 7293 3927 7327
rect 4813 7293 4847 7327
rect 4997 7293 5031 7327
rect 7757 7293 7791 7327
rect 8309 7293 8343 7327
rect 2053 7225 2087 7259
rect 2973 7157 3007 7191
rect 5457 7157 5491 7191
rect 5181 6953 5215 6987
rect 8493 6953 8527 6987
rect 8953 6953 8987 6987
rect 13369 6953 13403 6987
rect 13737 6953 13771 6987
rect 16313 6953 16347 6987
rect 18429 6953 18463 6987
rect 19257 6953 19291 6987
rect 19625 6953 19659 6987
rect 21281 6953 21315 6987
rect 2237 6817 2271 6851
rect 3893 6817 3927 6851
rect 4077 6817 4111 6851
rect 5825 6817 5859 6851
rect 6837 6817 6871 6851
rect 9597 6817 9631 6851
rect 16037 6817 16071 6851
rect 18153 6817 18187 6851
rect 21005 6817 21039 6851
rect 3433 6749 3467 6783
rect 5549 6749 5583 6783
rect 7757 6749 7791 6783
rect 11989 6749 12023 6783
rect 15781 6749 15815 6783
rect 20738 6749 20772 6783
rect 4169 6681 4203 6715
rect 6653 6681 6687 6715
rect 7481 6681 7515 6715
rect 9321 6681 9355 6715
rect 9965 6681 9999 6715
rect 12234 6681 12268 6715
rect 17886 6681 17920 6715
rect 1685 6613 1719 6647
rect 2329 6613 2363 6647
rect 2421 6613 2455 6647
rect 2789 6613 2823 6647
rect 4537 6613 4571 6647
rect 4905 6613 4939 6647
rect 5641 6613 5675 6647
rect 6285 6613 6319 6647
rect 6745 6613 6779 6647
rect 8033 6613 8067 6647
rect 9413 6613 9447 6647
rect 14657 6613 14691 6647
rect 16773 6613 16807 6647
rect 2513 6409 2547 6443
rect 5641 6409 5675 6443
rect 6745 6409 6779 6443
rect 8677 6409 8711 6443
rect 9045 6409 9079 6443
rect 15485 6409 15519 6443
rect 18061 6409 18095 6443
rect 18337 6409 18371 6443
rect 19073 6409 19107 6443
rect 20821 6409 20855 6443
rect 21097 6409 21131 6443
rect 6377 6341 6411 6375
rect 4537 6273 4571 6307
rect 7113 6273 7147 6307
rect 13010 6273 13044 6307
rect 13277 6273 13311 6307
rect 14850 6273 14884 6307
rect 15117 6273 15151 6307
rect 16681 6273 16715 6307
rect 16937 6273 16971 6307
rect 19441 6273 19475 6307
rect 19708 6273 19742 6307
rect 2973 6205 3007 6239
rect 4721 6205 4755 6239
rect 5733 6205 5767 6239
rect 5917 6205 5951 6239
rect 7205 6205 7239 6239
rect 7389 6205 7423 6239
rect 8493 6205 8527 6239
rect 8585 6205 8619 6239
rect 9321 6205 9355 6239
rect 4261 6137 4295 6171
rect 5273 6069 5307 6103
rect 8033 6069 8067 6103
rect 11897 6069 11931 6103
rect 13737 6069 13771 6103
rect 3801 5865 3835 5899
rect 5273 5865 5307 5899
rect 13461 5865 13495 5899
rect 15761 5865 15795 5899
rect 18705 5865 18739 5899
rect 19349 5865 19383 5899
rect 21097 5865 21131 5899
rect 6929 5797 6963 5831
rect 8033 5797 8067 5831
rect 11437 5797 11471 5831
rect 18429 5797 18463 5831
rect 1593 5729 1627 5763
rect 3065 5729 3099 5763
rect 4169 5729 4203 5763
rect 4721 5729 4755 5763
rect 6101 5729 6135 5763
rect 7481 5729 7515 5763
rect 9413 5729 9447 5763
rect 9597 5729 9631 5763
rect 12817 5729 12851 5763
rect 15485 5729 15519 5763
rect 17049 5729 17083 5763
rect 20729 5729 20763 5763
rect 1685 5661 1719 5695
rect 1777 5661 1811 5695
rect 6285 5661 6319 5695
rect 7665 5661 7699 5695
rect 9321 5661 9355 5695
rect 17305 5661 17339 5695
rect 20462 5661 20496 5695
rect 2789 5593 2823 5627
rect 12572 5593 12606 5627
rect 15240 5593 15274 5627
rect 2145 5525 2179 5559
rect 2421 5525 2455 5559
rect 2881 5525 2915 5559
rect 4813 5525 4847 5559
rect 4905 5525 4939 5559
rect 5549 5525 5583 5559
rect 6193 5525 6227 5559
rect 6653 5525 6687 5559
rect 7573 5525 7607 5559
rect 8585 5525 8619 5559
rect 8953 5525 8987 5559
rect 9965 5525 9999 5559
rect 11161 5525 11195 5559
rect 14105 5525 14139 5559
rect 1501 5321 1535 5355
rect 2605 5321 2639 5355
rect 2973 5321 3007 5355
rect 3249 5321 3283 5355
rect 3709 5321 3743 5355
rect 4721 5321 4755 5355
rect 5089 5321 5123 5355
rect 6745 5321 6779 5355
rect 7481 5321 7515 5355
rect 9137 5321 9171 5355
rect 13277 5321 13311 5355
rect 13553 5321 13587 5355
rect 16221 5321 16255 5355
rect 18337 5321 18371 5355
rect 18981 5321 19015 5355
rect 19349 5321 19383 5355
rect 19717 5321 19751 5355
rect 9229 5253 9263 5287
rect 12642 5253 12676 5287
rect 15678 5253 15712 5287
rect 20830 5253 20864 5287
rect 3617 5185 3651 5219
rect 4445 5185 4479 5219
rect 5181 5185 5215 5219
rect 6009 5185 6043 5219
rect 6837 5185 6871 5219
rect 8217 5185 8251 5219
rect 10894 5185 10928 5219
rect 11161 5185 11195 5219
rect 12909 5185 12943 5219
rect 15945 5185 15979 5219
rect 16681 5185 16715 5219
rect 16948 5185 16982 5219
rect 21097 5185 21131 5219
rect 2421 5117 2455 5151
rect 2513 5117 2547 5151
rect 3893 5117 3927 5151
rect 5365 5117 5399 5151
rect 6929 5117 6963 5151
rect 7941 5117 7975 5151
rect 9413 5117 9447 5151
rect 9781 5049 9815 5083
rect 11529 5049 11563 5083
rect 1869 4981 1903 5015
rect 6377 4981 6411 5015
rect 8769 4981 8803 5015
rect 14565 4981 14599 5015
rect 18061 4981 18095 5015
rect 4629 4777 4663 4811
rect 5181 4777 5215 4811
rect 8585 4777 8619 4811
rect 10885 4777 10919 4811
rect 12633 4777 12667 4811
rect 13001 4777 13035 4811
rect 14105 4777 14139 4811
rect 16497 4777 16531 4811
rect 17141 4777 17175 4811
rect 21005 4777 21039 4811
rect 21281 4777 21315 4811
rect 3341 4709 3375 4743
rect 4261 4709 4295 4743
rect 17509 4709 17543 4743
rect 1869 4641 1903 4675
rect 1961 4641 1995 4675
rect 5641 4641 5675 4675
rect 5733 4641 5767 4675
rect 7297 4641 7331 4675
rect 9597 4641 9631 4675
rect 9781 4641 9815 4675
rect 11253 4641 11287 4675
rect 16129 4641 16163 4675
rect 18889 4641 18923 4675
rect 20637 4641 20671 4675
rect 2053 4573 2087 4607
rect 8125 4573 8159 4607
rect 15862 4573 15896 4607
rect 16773 4573 16807 4607
rect 2881 4505 2915 4539
rect 7113 4505 7147 4539
rect 7849 4505 7883 4539
rect 11498 4505 11532 4539
rect 18622 4505 18656 4539
rect 20370 4505 20404 4539
rect 2421 4437 2455 4471
rect 3893 4437 3927 4471
rect 5825 4437 5859 4471
rect 6193 4437 6227 4471
rect 6653 4437 6687 4471
rect 7021 4437 7055 4471
rect 9137 4437 9171 4471
rect 9505 4437 9539 4471
rect 10149 4437 10183 4471
rect 14749 4437 14783 4471
rect 19257 4437 19291 4471
rect 5549 4233 5583 4267
rect 9413 4233 9447 4267
rect 11161 4233 11195 4267
rect 16037 4233 16071 4267
rect 18061 4233 18095 4267
rect 19993 4233 20027 4267
rect 9321 4165 9355 4199
rect 2697 4097 2731 4131
rect 4813 4097 4847 4131
rect 5641 4097 5675 4131
rect 6837 4097 6871 4131
rect 7389 4097 7423 4131
rect 8677 4097 8711 4131
rect 13746 4097 13780 4131
rect 14013 4097 14047 4131
rect 15402 4097 15436 4131
rect 15669 4097 15703 4131
rect 16681 4097 16715 4131
rect 16937 4097 16971 4131
rect 19450 4097 19484 4131
rect 19717 4097 19751 4131
rect 21106 4097 21140 4131
rect 21373 4097 21407 4131
rect 2973 4029 3007 4063
rect 5825 4029 5859 4063
rect 6653 4029 6687 4063
rect 7665 4029 7699 4063
rect 8401 4029 8435 4063
rect 9597 4029 9631 4063
rect 4169 3961 4203 3995
rect 5181 3961 5215 3995
rect 8953 3961 8987 3995
rect 14289 3961 14323 3995
rect 18337 3961 18371 3995
rect 3801 3893 3835 3927
rect 4537 3893 4571 3927
rect 12633 3893 12667 3927
rect 4353 3689 4387 3723
rect 5825 3689 5859 3723
rect 13001 3689 13035 3723
rect 15853 3689 15887 3723
rect 16957 3689 16991 3723
rect 18705 3689 18739 3723
rect 20913 3689 20947 3723
rect 21281 3689 21315 3723
rect 9229 3621 9263 3655
rect 11253 3621 11287 3655
rect 3985 3553 4019 3587
rect 6285 3553 6319 3587
rect 6469 3553 6503 3587
rect 7757 3553 7791 3587
rect 10977 3553 11011 3587
rect 12633 3553 12667 3587
rect 15485 3553 15519 3587
rect 18337 3553 18371 3587
rect 20637 3553 20671 3587
rect 5089 3485 5123 3519
rect 5365 3485 5399 3519
rect 8585 3485 8619 3519
rect 9045 3485 9079 3519
rect 10710 3485 10744 3519
rect 15218 3485 15252 3519
rect 18070 3485 18104 3519
rect 20370 3485 20404 3519
rect 6193 3417 6227 3451
rect 7481 3417 7515 3451
rect 7573 3417 7607 3451
rect 8309 3417 8343 3451
rect 12366 3417 12400 3451
rect 4813 3349 4847 3383
rect 7113 3349 7147 3383
rect 9597 3349 9631 3383
rect 14105 3349 14139 3383
rect 19257 3349 19291 3383
rect 1501 3145 1535 3179
rect 5273 3145 5307 3179
rect 6929 3145 6963 3179
rect 7389 3145 7423 3179
rect 9781 3145 9815 3179
rect 12909 3145 12943 3179
rect 13369 3145 13403 3179
rect 16681 3145 16715 3179
rect 17141 3145 17175 3179
rect 18245 3145 18279 3179
rect 19901 3145 19935 3179
rect 9321 3077 9355 3111
rect 17877 3077 17911 3111
rect 1869 3009 1903 3043
rect 2421 3009 2455 3043
rect 2973 3009 3007 3043
rect 4629 3009 4663 3043
rect 5457 3009 5491 3043
rect 6009 3009 6043 3043
rect 7021 3009 7055 3043
rect 8033 3009 8067 3043
rect 8769 3009 8803 3043
rect 9045 3009 9079 3043
rect 10894 3009 10928 3043
rect 11161 3009 11195 3043
rect 11529 3009 11563 3043
rect 11785 3009 11819 3043
rect 13185 3009 13219 3043
rect 13737 3009 13771 3043
rect 14749 3009 14783 3043
rect 15025 3009 15059 3043
rect 15577 3009 15611 3043
rect 16313 3009 16347 3043
rect 17049 3009 17083 3043
rect 18521 3009 18555 3043
rect 18788 3009 18822 3043
rect 20361 3009 20395 3043
rect 6837 2941 6871 2975
rect 8585 2941 8619 2975
rect 14565 2941 14599 2975
rect 17233 2941 17267 2975
rect 20637 2941 20671 2975
rect 4813 2873 4847 2907
rect 5825 2873 5859 2907
rect 7849 2873 7883 2907
rect 15209 2873 15243 2907
rect 15761 2873 15795 2907
rect 2053 2805 2087 2839
rect 2605 2805 2639 2839
rect 13921 2805 13955 2839
rect 11161 2601 11195 2635
rect 17601 2601 17635 2635
rect 17969 2601 18003 2635
rect 21097 2601 21131 2635
rect 6745 2533 6779 2567
rect 8493 2533 8527 2567
rect 10057 2533 10091 2567
rect 11529 2533 11563 2567
rect 20821 2533 20855 2567
rect 9413 2465 9447 2499
rect 12909 2465 12943 2499
rect 13185 2465 13219 2499
rect 13553 2465 13587 2499
rect 1961 2397 1995 2431
rect 2513 2397 2547 2431
rect 5181 2397 5215 2431
rect 6009 2397 6043 2431
rect 6929 2397 6963 2431
rect 7205 2397 7239 2431
rect 8309 2397 8343 2431
rect 9597 2397 9631 2431
rect 10339 2397 10373 2431
rect 15117 2397 15151 2431
rect 18337 2397 18371 2431
rect 18613 2397 18647 2431
rect 19441 2397 19475 2431
rect 7481 2329 7515 2363
rect 9045 2329 9079 2363
rect 12642 2329 12676 2363
rect 19686 2329 19720 2363
rect 2145 2261 2179 2295
rect 4813 2261 4847 2295
rect 5365 2261 5399 2295
rect 5825 2261 5859 2295
rect 7941 2261 7975 2295
rect 9689 2261 9723 2295
rect 10517 2261 10551 2295
rect 15301 2261 15335 2295
rect 18797 2261 18831 2295
<< metal1 >>
rect 2958 20952 2964 21004
rect 3016 20992 3022 21004
rect 5902 20992 5908 21004
rect 3016 20964 5908 20992
rect 3016 20952 3022 20964
rect 5902 20952 5908 20964
rect 5960 20952 5966 21004
rect 3878 20748 3884 20800
rect 3936 20788 3942 20800
rect 5626 20788 5632 20800
rect 3936 20760 5632 20788
rect 3936 20748 3942 20760
rect 5626 20748 5632 20760
rect 5684 20748 5690 20800
rect 1104 20698 22056 20720
rect 1104 20646 6148 20698
rect 6200 20646 6212 20698
rect 6264 20646 6276 20698
rect 6328 20646 6340 20698
rect 6392 20646 6404 20698
rect 6456 20646 11346 20698
rect 11398 20646 11410 20698
rect 11462 20646 11474 20698
rect 11526 20646 11538 20698
rect 11590 20646 11602 20698
rect 11654 20646 16544 20698
rect 16596 20646 16608 20698
rect 16660 20646 16672 20698
rect 16724 20646 16736 20698
rect 16788 20646 16800 20698
rect 16852 20646 21742 20698
rect 21794 20646 21806 20698
rect 21858 20646 21870 20698
rect 21922 20646 21934 20698
rect 21986 20646 21998 20698
rect 22050 20646 22056 20698
rect 1104 20624 22056 20646
rect 1104 20154 21896 20176
rect 1104 20102 3549 20154
rect 3601 20102 3613 20154
rect 3665 20102 3677 20154
rect 3729 20102 3741 20154
rect 3793 20102 3805 20154
rect 3857 20102 8747 20154
rect 8799 20102 8811 20154
rect 8863 20102 8875 20154
rect 8927 20102 8939 20154
rect 8991 20102 9003 20154
rect 9055 20102 13945 20154
rect 13997 20102 14009 20154
rect 14061 20102 14073 20154
rect 14125 20102 14137 20154
rect 14189 20102 14201 20154
rect 14253 20102 19143 20154
rect 19195 20102 19207 20154
rect 19259 20102 19271 20154
rect 19323 20102 19335 20154
rect 19387 20102 19399 20154
rect 19451 20102 21896 20154
rect 1104 20080 21896 20102
rect 4062 20000 4068 20052
rect 4120 20040 4126 20052
rect 4525 20043 4583 20049
rect 4525 20040 4537 20043
rect 4120 20012 4537 20040
rect 4120 20000 4126 20012
rect 4525 20009 4537 20012
rect 4571 20009 4583 20043
rect 5626 20040 5632 20052
rect 5587 20012 5632 20040
rect 4525 20003 4583 20009
rect 5626 20000 5632 20012
rect 5684 20000 5690 20052
rect 7377 19907 7435 19913
rect 7377 19904 7389 19907
rect 4724 19876 7389 19904
rect 4724 19845 4752 19876
rect 7377 19873 7389 19876
rect 7423 19873 7435 19907
rect 7377 19867 7435 19873
rect 4709 19839 4767 19845
rect 4709 19805 4721 19839
rect 4755 19805 4767 19839
rect 5810 19836 5816 19848
rect 5771 19808 5816 19836
rect 4709 19799 4767 19805
rect 5810 19796 5816 19808
rect 5868 19796 5874 19848
rect 7653 19839 7711 19845
rect 7653 19805 7665 19839
rect 7699 19836 7711 19839
rect 10410 19836 10416 19848
rect 7699 19808 10416 19836
rect 7699 19805 7711 19808
rect 7653 19799 7711 19805
rect 10410 19796 10416 19808
rect 10468 19796 10474 19848
rect 1104 19610 22056 19632
rect 1104 19558 6148 19610
rect 6200 19558 6212 19610
rect 6264 19558 6276 19610
rect 6328 19558 6340 19610
rect 6392 19558 6404 19610
rect 6456 19558 11346 19610
rect 11398 19558 11410 19610
rect 11462 19558 11474 19610
rect 11526 19558 11538 19610
rect 11590 19558 11602 19610
rect 11654 19558 16544 19610
rect 16596 19558 16608 19610
rect 16660 19558 16672 19610
rect 16724 19558 16736 19610
rect 16788 19558 16800 19610
rect 16852 19558 21742 19610
rect 21794 19558 21806 19610
rect 21858 19558 21870 19610
rect 21922 19558 21934 19610
rect 21986 19558 21998 19610
rect 22050 19558 22056 19610
rect 1104 19536 22056 19558
rect 3234 19456 3240 19508
rect 3292 19496 3298 19508
rect 4525 19499 4583 19505
rect 4525 19496 4537 19499
rect 3292 19468 4537 19496
rect 3292 19456 3298 19468
rect 4525 19465 4537 19468
rect 4571 19465 4583 19499
rect 4525 19459 4583 19465
rect 5810 19388 5816 19440
rect 5868 19428 5874 19440
rect 8573 19431 8631 19437
rect 8573 19428 8585 19431
rect 5868 19400 8585 19428
rect 5868 19388 5874 19400
rect 8573 19397 8585 19400
rect 8619 19397 8631 19431
rect 8573 19391 8631 19397
rect 4706 19360 4712 19372
rect 4667 19332 4712 19360
rect 4706 19320 4712 19332
rect 4764 19320 4770 19372
rect 8849 19363 8907 19369
rect 8849 19329 8861 19363
rect 8895 19360 8907 19363
rect 9122 19360 9128 19372
rect 8895 19332 9128 19360
rect 8895 19329 8907 19332
rect 8849 19323 8907 19329
rect 9122 19320 9128 19332
rect 9180 19320 9186 19372
rect 1104 19066 21896 19088
rect 1104 19014 3549 19066
rect 3601 19014 3613 19066
rect 3665 19014 3677 19066
rect 3729 19014 3741 19066
rect 3793 19014 3805 19066
rect 3857 19014 8747 19066
rect 8799 19014 8811 19066
rect 8863 19014 8875 19066
rect 8927 19014 8939 19066
rect 8991 19014 9003 19066
rect 9055 19014 13945 19066
rect 13997 19014 14009 19066
rect 14061 19014 14073 19066
rect 14125 19014 14137 19066
rect 14189 19014 14201 19066
rect 14253 19014 19143 19066
rect 19195 19014 19207 19066
rect 19259 19014 19271 19066
rect 19323 19014 19335 19066
rect 19387 19014 19399 19066
rect 19451 19014 21896 19066
rect 1104 18992 21896 19014
rect 4154 18912 4160 18964
rect 4212 18952 4218 18964
rect 4617 18955 4675 18961
rect 4617 18952 4629 18955
rect 4212 18924 4629 18952
rect 4212 18912 4218 18924
rect 4617 18921 4629 18924
rect 4663 18921 4675 18955
rect 4617 18915 4675 18921
rect 4801 18751 4859 18757
rect 4801 18717 4813 18751
rect 4847 18748 4859 18751
rect 5810 18748 5816 18760
rect 4847 18720 5816 18748
rect 4847 18717 4859 18720
rect 4801 18711 4859 18717
rect 5810 18708 5816 18720
rect 5868 18708 5874 18760
rect 1104 18522 22056 18544
rect 1104 18470 6148 18522
rect 6200 18470 6212 18522
rect 6264 18470 6276 18522
rect 6328 18470 6340 18522
rect 6392 18470 6404 18522
rect 6456 18470 11346 18522
rect 11398 18470 11410 18522
rect 11462 18470 11474 18522
rect 11526 18470 11538 18522
rect 11590 18470 11602 18522
rect 11654 18470 16544 18522
rect 16596 18470 16608 18522
rect 16660 18470 16672 18522
rect 16724 18470 16736 18522
rect 16788 18470 16800 18522
rect 16852 18470 21742 18522
rect 21794 18470 21806 18522
rect 21858 18470 21870 18522
rect 21922 18470 21934 18522
rect 21986 18470 21998 18522
rect 22050 18470 22056 18522
rect 1104 18448 22056 18470
rect 4062 18368 4068 18420
rect 4120 18408 4126 18420
rect 4801 18411 4859 18417
rect 4801 18408 4813 18411
rect 4120 18380 4813 18408
rect 4120 18368 4126 18380
rect 4801 18377 4813 18380
rect 4847 18377 4859 18411
rect 4801 18371 4859 18377
rect 4985 18275 5043 18281
rect 4985 18241 4997 18275
rect 5031 18272 5043 18275
rect 7650 18272 7656 18284
rect 5031 18244 7656 18272
rect 5031 18241 5043 18244
rect 4985 18235 5043 18241
rect 7650 18232 7656 18244
rect 7708 18232 7714 18284
rect 1104 17978 21896 18000
rect 1104 17926 3549 17978
rect 3601 17926 3613 17978
rect 3665 17926 3677 17978
rect 3729 17926 3741 17978
rect 3793 17926 3805 17978
rect 3857 17926 8747 17978
rect 8799 17926 8811 17978
rect 8863 17926 8875 17978
rect 8927 17926 8939 17978
rect 8991 17926 9003 17978
rect 9055 17926 13945 17978
rect 13997 17926 14009 17978
rect 14061 17926 14073 17978
rect 14125 17926 14137 17978
rect 14189 17926 14201 17978
rect 14253 17926 19143 17978
rect 19195 17926 19207 17978
rect 19259 17926 19271 17978
rect 19323 17926 19335 17978
rect 19387 17926 19399 17978
rect 19451 17926 21896 17978
rect 1104 17904 21896 17926
rect 1946 17864 1952 17876
rect 1907 17836 1952 17864
rect 1946 17824 1952 17836
rect 2004 17824 2010 17876
rect 3970 17864 3976 17876
rect 3931 17836 3976 17864
rect 3970 17824 3976 17836
rect 4028 17824 4034 17876
rect 4154 17824 4160 17876
rect 4212 17864 4218 17876
rect 4709 17867 4767 17873
rect 4709 17864 4721 17867
rect 4212 17836 4721 17864
rect 4212 17824 4218 17836
rect 4709 17833 4721 17836
rect 4755 17833 4767 17867
rect 4709 17827 4767 17833
rect 5810 17688 5816 17740
rect 5868 17728 5874 17740
rect 7101 17731 7159 17737
rect 7101 17728 7113 17731
rect 5868 17700 7113 17728
rect 5868 17688 5874 17700
rect 7101 17697 7113 17700
rect 7147 17697 7159 17731
rect 7101 17691 7159 17697
rect 2133 17663 2191 17669
rect 2133 17629 2145 17663
rect 2179 17660 2191 17663
rect 2222 17660 2228 17672
rect 2179 17632 2228 17660
rect 2179 17629 2191 17632
rect 2133 17623 2191 17629
rect 2222 17620 2228 17632
rect 2280 17620 2286 17672
rect 4157 17663 4215 17669
rect 4157 17629 4169 17663
rect 4203 17629 4215 17663
rect 4157 17623 4215 17629
rect 4893 17663 4951 17669
rect 4893 17629 4905 17663
rect 4939 17660 4951 17663
rect 6730 17660 6736 17672
rect 4939 17632 6736 17660
rect 4939 17629 4951 17632
rect 4893 17623 4951 17629
rect 4172 17592 4200 17623
rect 6730 17620 6736 17632
rect 6788 17620 6794 17672
rect 7377 17663 7435 17669
rect 7377 17629 7389 17663
rect 7423 17660 7435 17663
rect 9398 17660 9404 17672
rect 7423 17632 9404 17660
rect 7423 17629 7435 17632
rect 7377 17623 7435 17629
rect 9398 17620 9404 17632
rect 9456 17620 9462 17672
rect 5994 17592 6000 17604
rect 4172 17564 6000 17592
rect 5994 17552 6000 17564
rect 6052 17552 6058 17604
rect 1104 17434 22056 17456
rect 1104 17382 6148 17434
rect 6200 17382 6212 17434
rect 6264 17382 6276 17434
rect 6328 17382 6340 17434
rect 6392 17382 6404 17434
rect 6456 17382 11346 17434
rect 11398 17382 11410 17434
rect 11462 17382 11474 17434
rect 11526 17382 11538 17434
rect 11590 17382 11602 17434
rect 11654 17382 16544 17434
rect 16596 17382 16608 17434
rect 16660 17382 16672 17434
rect 16724 17382 16736 17434
rect 16788 17382 16800 17434
rect 16852 17382 21742 17434
rect 21794 17382 21806 17434
rect 21858 17382 21870 17434
rect 21922 17382 21934 17434
rect 21986 17382 21998 17434
rect 22050 17382 22056 17434
rect 1104 17360 22056 17382
rect 1578 17320 1584 17332
rect 1539 17292 1584 17320
rect 1578 17280 1584 17292
rect 1636 17280 1642 17332
rect 3694 17320 3700 17332
rect 3655 17292 3700 17320
rect 3694 17280 3700 17292
rect 3752 17280 3758 17332
rect 2222 17252 2228 17264
rect 2183 17224 2228 17252
rect 2222 17212 2228 17224
rect 2280 17212 2286 17264
rect 4706 17212 4712 17264
rect 4764 17252 4770 17264
rect 7469 17255 7527 17261
rect 7469 17252 7481 17255
rect 4764 17224 7481 17252
rect 4764 17212 4770 17224
rect 7469 17221 7481 17224
rect 7515 17221 7527 17255
rect 7469 17215 7527 17221
rect 1765 17187 1823 17193
rect 1765 17153 1777 17187
rect 1811 17153 1823 17187
rect 1765 17147 1823 17153
rect 2501 17187 2559 17193
rect 2501 17153 2513 17187
rect 2547 17153 2559 17187
rect 2501 17147 2559 17153
rect 3881 17187 3939 17193
rect 3881 17153 3893 17187
rect 3927 17184 3939 17187
rect 5169 17187 5227 17193
rect 5169 17184 5181 17187
rect 3927 17156 5181 17184
rect 3927 17153 3939 17156
rect 3881 17147 3939 17153
rect 5169 17153 5181 17156
rect 5215 17153 5227 17187
rect 5169 17147 5227 17153
rect 5445 17187 5503 17193
rect 5445 17153 5457 17187
rect 5491 17184 5503 17187
rect 6638 17184 6644 17196
rect 5491 17156 6644 17184
rect 5491 17153 5503 17156
rect 5445 17147 5503 17153
rect 1780 17048 1808 17147
rect 2516 17116 2544 17147
rect 6638 17144 6644 17156
rect 6696 17144 6702 17196
rect 7745 17187 7803 17193
rect 7745 17153 7757 17187
rect 7791 17184 7803 17187
rect 12158 17184 12164 17196
rect 7791 17156 12164 17184
rect 7791 17153 7803 17156
rect 7745 17147 7803 17153
rect 12158 17144 12164 17156
rect 12216 17144 12222 17196
rect 4246 17116 4252 17128
rect 2516 17088 4252 17116
rect 4246 17076 4252 17088
rect 4304 17076 4310 17128
rect 4430 17048 4436 17060
rect 1780 17020 4436 17048
rect 4430 17008 4436 17020
rect 4488 17008 4494 17060
rect 1104 16890 21896 16912
rect 1104 16838 3549 16890
rect 3601 16838 3613 16890
rect 3665 16838 3677 16890
rect 3729 16838 3741 16890
rect 3793 16838 3805 16890
rect 3857 16838 8747 16890
rect 8799 16838 8811 16890
rect 8863 16838 8875 16890
rect 8927 16838 8939 16890
rect 8991 16838 9003 16890
rect 9055 16838 13945 16890
rect 13997 16838 14009 16890
rect 14061 16838 14073 16890
rect 14125 16838 14137 16890
rect 14189 16838 14201 16890
rect 14253 16838 19143 16890
rect 19195 16838 19207 16890
rect 19259 16838 19271 16890
rect 19323 16838 19335 16890
rect 19387 16838 19399 16890
rect 19451 16838 21896 16890
rect 1104 16816 21896 16838
rect 10870 16708 10876 16720
rect 9416 16680 10876 16708
rect 9416 16649 9444 16680
rect 10870 16668 10876 16680
rect 10928 16668 10934 16720
rect 9401 16643 9459 16649
rect 9401 16609 9413 16643
rect 9447 16609 9459 16643
rect 9401 16603 9459 16609
rect 9585 16643 9643 16649
rect 9585 16609 9597 16643
rect 9631 16640 9643 16643
rect 10505 16643 10563 16649
rect 10505 16640 10517 16643
rect 9631 16612 10517 16640
rect 9631 16609 9643 16612
rect 9585 16603 9643 16609
rect 10505 16609 10517 16612
rect 10551 16640 10563 16643
rect 21450 16640 21456 16652
rect 10551 16612 21456 16640
rect 10551 16609 10563 16612
rect 10505 16603 10563 16609
rect 21450 16600 21456 16612
rect 21508 16600 21514 16652
rect 4430 16572 4436 16584
rect 4391 16544 4436 16572
rect 4430 16532 4436 16544
rect 4488 16532 4494 16584
rect 4709 16575 4767 16581
rect 4709 16541 4721 16575
rect 4755 16572 4767 16575
rect 5810 16572 5816 16584
rect 4755 16544 5816 16572
rect 4755 16541 4767 16544
rect 4709 16535 4767 16541
rect 5810 16532 5816 16544
rect 5868 16532 5874 16584
rect 5994 16532 6000 16584
rect 6052 16572 6058 16584
rect 6181 16575 6239 16581
rect 6181 16572 6193 16575
rect 6052 16544 6193 16572
rect 6052 16532 6058 16544
rect 6181 16541 6193 16544
rect 6227 16541 6239 16575
rect 6181 16535 6239 16541
rect 6457 16575 6515 16581
rect 6457 16541 6469 16575
rect 6503 16572 6515 16575
rect 6822 16572 6828 16584
rect 6503 16544 6828 16572
rect 6503 16541 6515 16544
rect 6457 16535 6515 16541
rect 6822 16532 6828 16544
rect 6880 16532 6886 16584
rect 7190 16572 7196 16584
rect 7151 16544 7196 16572
rect 7190 16532 7196 16544
rect 7248 16532 7254 16584
rect 7650 16572 7656 16584
rect 7611 16544 7656 16572
rect 7650 16532 7656 16544
rect 7708 16532 7714 16584
rect 7929 16575 7987 16581
rect 7929 16541 7941 16575
rect 7975 16572 7987 16575
rect 8570 16572 8576 16584
rect 7975 16544 8576 16572
rect 7975 16541 7987 16544
rect 7929 16535 7987 16541
rect 8570 16532 8576 16544
rect 8628 16532 8634 16584
rect 6730 16464 6736 16516
rect 6788 16504 6794 16516
rect 6917 16507 6975 16513
rect 6917 16504 6929 16507
rect 6788 16476 6929 16504
rect 6788 16464 6794 16476
rect 6917 16473 6929 16476
rect 6963 16473 6975 16507
rect 6917 16467 6975 16473
rect 8941 16439 8999 16445
rect 8941 16405 8953 16439
rect 8987 16436 8999 16439
rect 9122 16436 9128 16448
rect 8987 16408 9128 16436
rect 8987 16405 8999 16408
rect 8941 16399 8999 16405
rect 9122 16396 9128 16408
rect 9180 16396 9186 16448
rect 9309 16439 9367 16445
rect 9309 16405 9321 16439
rect 9355 16436 9367 16439
rect 9953 16439 10011 16445
rect 9953 16436 9965 16439
rect 9355 16408 9965 16436
rect 9355 16405 9367 16408
rect 9309 16399 9367 16405
rect 9953 16405 9965 16408
rect 9999 16405 10011 16439
rect 9953 16399 10011 16405
rect 1104 16346 22056 16368
rect 1104 16294 6148 16346
rect 6200 16294 6212 16346
rect 6264 16294 6276 16346
rect 6328 16294 6340 16346
rect 6392 16294 6404 16346
rect 6456 16294 11346 16346
rect 11398 16294 11410 16346
rect 11462 16294 11474 16346
rect 11526 16294 11538 16346
rect 11590 16294 11602 16346
rect 11654 16294 16544 16346
rect 16596 16294 16608 16346
rect 16660 16294 16672 16346
rect 16724 16294 16736 16346
rect 16788 16294 16800 16346
rect 16852 16294 21742 16346
rect 21794 16294 21806 16346
rect 21858 16294 21870 16346
rect 21922 16294 21934 16346
rect 21986 16294 21998 16346
rect 22050 16294 22056 16346
rect 1104 16272 22056 16294
rect 1946 16232 1952 16244
rect 1907 16204 1952 16232
rect 1946 16192 1952 16204
rect 2004 16192 2010 16244
rect 2133 16099 2191 16105
rect 2133 16065 2145 16099
rect 2179 16096 2191 16099
rect 5350 16096 5356 16108
rect 2179 16068 5356 16096
rect 2179 16065 2191 16068
rect 2133 16059 2191 16065
rect 5350 16056 5356 16068
rect 5408 16056 5414 16108
rect 5166 15892 5172 15904
rect 5127 15864 5172 15892
rect 5166 15852 5172 15864
rect 5224 15852 5230 15904
rect 1104 15802 21896 15824
rect 1104 15750 3549 15802
rect 3601 15750 3613 15802
rect 3665 15750 3677 15802
rect 3729 15750 3741 15802
rect 3793 15750 3805 15802
rect 3857 15750 8747 15802
rect 8799 15750 8811 15802
rect 8863 15750 8875 15802
rect 8927 15750 8939 15802
rect 8991 15750 9003 15802
rect 9055 15750 13945 15802
rect 13997 15750 14009 15802
rect 14061 15750 14073 15802
rect 14125 15750 14137 15802
rect 14189 15750 14201 15802
rect 14253 15750 19143 15802
rect 19195 15750 19207 15802
rect 19259 15750 19271 15802
rect 19323 15750 19335 15802
rect 19387 15750 19399 15802
rect 19451 15750 21896 15802
rect 1104 15728 21896 15750
rect 1670 15688 1676 15700
rect 1631 15660 1676 15688
rect 1670 15648 1676 15660
rect 1728 15648 1734 15700
rect 2774 15688 2780 15700
rect 2735 15660 2780 15688
rect 2774 15648 2780 15660
rect 2832 15648 2838 15700
rect 5902 15688 5908 15700
rect 5863 15660 5908 15688
rect 5902 15648 5908 15660
rect 5960 15648 5966 15700
rect 6638 15648 6644 15700
rect 6696 15688 6702 15700
rect 7285 15691 7343 15697
rect 7285 15688 7297 15691
rect 6696 15660 7297 15688
rect 6696 15648 6702 15660
rect 7285 15657 7297 15660
rect 7331 15657 7343 15691
rect 7285 15651 7343 15657
rect 2222 15620 2228 15632
rect 2183 15592 2228 15620
rect 2222 15580 2228 15592
rect 2280 15580 2286 15632
rect 4525 15555 4583 15561
rect 4525 15552 4537 15555
rect 1872 15524 4537 15552
rect 1872 15493 1900 15524
rect 4525 15521 4537 15524
rect 4571 15521 4583 15555
rect 5350 15552 5356 15564
rect 5311 15524 5356 15552
rect 4525 15515 4583 15521
rect 5350 15512 5356 15524
rect 5408 15512 5414 15564
rect 7929 15555 7987 15561
rect 7929 15521 7941 15555
rect 7975 15552 7987 15555
rect 11790 15552 11796 15564
rect 7975 15524 11796 15552
rect 7975 15521 7987 15524
rect 7929 15515 7987 15521
rect 11790 15512 11796 15524
rect 11848 15512 11854 15564
rect 1857 15487 1915 15493
rect 1857 15453 1869 15487
rect 1903 15453 1915 15487
rect 1857 15447 1915 15453
rect 2409 15487 2467 15493
rect 2409 15453 2421 15487
rect 2455 15484 2467 15487
rect 2866 15484 2872 15496
rect 2455 15456 2872 15484
rect 2455 15453 2467 15456
rect 2409 15447 2467 15453
rect 2866 15444 2872 15456
rect 2924 15444 2930 15496
rect 2961 15487 3019 15493
rect 2961 15453 2973 15487
rect 3007 15484 3019 15487
rect 3694 15484 3700 15496
rect 3007 15456 3700 15484
rect 3007 15453 3019 15456
rect 2961 15447 3019 15453
rect 3694 15444 3700 15456
rect 3752 15444 3758 15496
rect 4801 15487 4859 15493
rect 4801 15453 4813 15487
rect 4847 15453 4859 15487
rect 4801 15447 4859 15453
rect 5629 15487 5687 15493
rect 5629 15453 5641 15487
rect 5675 15484 5687 15487
rect 7742 15484 7748 15496
rect 5675 15456 7748 15484
rect 5675 15453 5687 15456
rect 5629 15447 5687 15453
rect 4816 15416 4844 15447
rect 7742 15444 7748 15456
rect 7800 15444 7806 15496
rect 5994 15416 6000 15428
rect 4816 15388 6000 15416
rect 5994 15376 6000 15388
rect 6052 15376 6058 15428
rect 7653 15419 7711 15425
rect 7653 15385 7665 15419
rect 7699 15416 7711 15419
rect 8297 15419 8355 15425
rect 8297 15416 8309 15419
rect 7699 15388 8309 15416
rect 7699 15385 7711 15388
rect 7653 15379 7711 15385
rect 8297 15385 8309 15388
rect 8343 15385 8355 15419
rect 8297 15379 8355 15385
rect 7745 15351 7803 15357
rect 7745 15317 7757 15351
rect 7791 15348 7803 15351
rect 9306 15348 9312 15360
rect 7791 15320 9312 15348
rect 7791 15317 7803 15320
rect 7745 15311 7803 15317
rect 9306 15308 9312 15320
rect 9364 15308 9370 15360
rect 1104 15258 22056 15280
rect 1104 15206 6148 15258
rect 6200 15206 6212 15258
rect 6264 15206 6276 15258
rect 6328 15206 6340 15258
rect 6392 15206 6404 15258
rect 6456 15206 11346 15258
rect 11398 15206 11410 15258
rect 11462 15206 11474 15258
rect 11526 15206 11538 15258
rect 11590 15206 11602 15258
rect 11654 15206 16544 15258
rect 16596 15206 16608 15258
rect 16660 15206 16672 15258
rect 16724 15206 16736 15258
rect 16788 15206 16800 15258
rect 16852 15206 21742 15258
rect 21794 15206 21806 15258
rect 21858 15206 21870 15258
rect 21922 15206 21934 15258
rect 21986 15206 21998 15258
rect 22050 15206 22056 15258
rect 1104 15184 22056 15206
rect 4246 15144 4252 15156
rect 4207 15116 4252 15144
rect 4246 15104 4252 15116
rect 4304 15104 4310 15156
rect 4709 15147 4767 15153
rect 4709 15113 4721 15147
rect 4755 15144 4767 15147
rect 5261 15147 5319 15153
rect 5261 15144 5273 15147
rect 4755 15116 5273 15144
rect 4755 15113 4767 15116
rect 4709 15107 4767 15113
rect 5261 15113 5273 15116
rect 5307 15113 5319 15147
rect 5261 15107 5319 15113
rect 5810 15104 5816 15156
rect 5868 15144 5874 15156
rect 6917 15147 6975 15153
rect 6917 15144 6929 15147
rect 5868 15116 6929 15144
rect 5868 15104 5874 15116
rect 6917 15113 6929 15116
rect 6963 15113 6975 15147
rect 6917 15107 6975 15113
rect 2866 15036 2872 15088
rect 2924 15076 2930 15088
rect 2961 15079 3019 15085
rect 2961 15076 2973 15079
rect 2924 15048 2973 15076
rect 2924 15036 2930 15048
rect 2961 15045 2973 15048
rect 3007 15045 3019 15079
rect 3694 15076 3700 15088
rect 3655 15048 3700 15076
rect 2961 15039 3019 15045
rect 3694 15036 3700 15048
rect 3752 15036 3758 15088
rect 7098 15076 7104 15088
rect 3988 15048 7104 15076
rect 2130 15008 2136 15020
rect 2091 14980 2136 15008
rect 2130 14968 2136 14980
rect 2188 14968 2194 15020
rect 3237 15011 3295 15017
rect 3237 14977 3249 15011
rect 3283 15008 3295 15011
rect 3878 15008 3884 15020
rect 3283 14980 3884 15008
rect 3283 14977 3295 14980
rect 3237 14971 3295 14977
rect 3878 14968 3884 14980
rect 3936 14968 3942 15020
rect 3988 15017 4016 15048
rect 7098 15036 7104 15048
rect 7156 15036 7162 15088
rect 3973 15011 4031 15017
rect 3973 14977 3985 15011
rect 4019 14977 4031 15011
rect 3973 14971 4031 14977
rect 4617 15011 4675 15017
rect 4617 14977 4629 15011
rect 4663 15008 4675 15011
rect 4890 15008 4896 15020
rect 4663 14980 4896 15008
rect 4663 14977 4675 14980
rect 4617 14971 4675 14977
rect 4890 14968 4896 14980
rect 4948 14968 4954 15020
rect 5629 15011 5687 15017
rect 5629 14977 5641 15011
rect 5675 15008 5687 15011
rect 5902 15008 5908 15020
rect 5675 14980 5908 15008
rect 5675 14977 5687 14980
rect 5629 14971 5687 14977
rect 5902 14968 5908 14980
rect 5960 14968 5966 15020
rect 7285 15011 7343 15017
rect 7285 14977 7297 15011
rect 7331 15008 7343 15011
rect 7929 15011 7987 15017
rect 7929 15008 7941 15011
rect 7331 14980 7941 15008
rect 7331 14977 7343 14980
rect 7285 14971 7343 14977
rect 7929 14977 7941 14980
rect 7975 14977 7987 15011
rect 7929 14971 7987 14977
rect 4801 14943 4859 14949
rect 4801 14909 4813 14943
rect 4847 14940 4859 14943
rect 5166 14940 5172 14952
rect 4847 14912 5172 14940
rect 4847 14909 4859 14912
rect 4801 14903 4859 14909
rect 5166 14900 5172 14912
rect 5224 14900 5230 14952
rect 5718 14940 5724 14952
rect 5679 14912 5724 14940
rect 5718 14900 5724 14912
rect 5776 14900 5782 14952
rect 5813 14943 5871 14949
rect 5813 14909 5825 14943
rect 5859 14909 5871 14943
rect 7374 14940 7380 14952
rect 7335 14912 7380 14940
rect 5813 14903 5871 14909
rect 1946 14804 1952 14816
rect 1907 14776 1952 14804
rect 1946 14764 1952 14776
rect 2004 14764 2010 14816
rect 5534 14764 5540 14816
rect 5592 14804 5598 14816
rect 5828 14804 5856 14903
rect 7374 14900 7380 14912
rect 7432 14900 7438 14952
rect 7561 14943 7619 14949
rect 7561 14909 7573 14943
rect 7607 14940 7619 14943
rect 15562 14940 15568 14952
rect 7607 14912 15568 14940
rect 7607 14909 7619 14912
rect 7561 14903 7619 14909
rect 15562 14900 15568 14912
rect 15620 14900 15626 14952
rect 6365 14807 6423 14813
rect 6365 14804 6377 14807
rect 5592 14776 6377 14804
rect 5592 14764 5598 14776
rect 6365 14773 6377 14776
rect 6411 14773 6423 14807
rect 6365 14767 6423 14773
rect 1104 14714 21896 14736
rect 1104 14662 3549 14714
rect 3601 14662 3613 14714
rect 3665 14662 3677 14714
rect 3729 14662 3741 14714
rect 3793 14662 3805 14714
rect 3857 14662 8747 14714
rect 8799 14662 8811 14714
rect 8863 14662 8875 14714
rect 8927 14662 8939 14714
rect 8991 14662 9003 14714
rect 9055 14662 13945 14714
rect 13997 14662 14009 14714
rect 14061 14662 14073 14714
rect 14125 14662 14137 14714
rect 14189 14662 14201 14714
rect 14253 14662 19143 14714
rect 19195 14662 19207 14714
rect 19259 14662 19271 14714
rect 19323 14662 19335 14714
rect 19387 14662 19399 14714
rect 19451 14662 21896 14714
rect 1104 14640 21896 14662
rect 1486 14600 1492 14612
rect 1447 14572 1492 14600
rect 1486 14560 1492 14572
rect 1544 14560 1550 14612
rect 9306 14600 9312 14612
rect 9267 14572 9312 14600
rect 9306 14560 9312 14572
rect 9364 14560 9370 14612
rect 3789 14535 3847 14541
rect 3789 14501 3801 14535
rect 3835 14501 3847 14535
rect 3789 14495 3847 14501
rect 2130 14464 2136 14476
rect 2091 14436 2136 14464
rect 2130 14424 2136 14436
rect 2188 14424 2194 14476
rect 3804 14464 3832 14495
rect 7834 14492 7840 14544
rect 7892 14532 7898 14544
rect 11882 14532 11888 14544
rect 7892 14504 11888 14532
rect 7892 14492 7898 14504
rect 11882 14492 11888 14504
rect 11940 14492 11946 14544
rect 2424 14436 3832 14464
rect 4433 14467 4491 14473
rect 2424 14405 2452 14436
rect 4433 14433 4445 14467
rect 4479 14464 4491 14467
rect 9953 14467 10011 14473
rect 4479 14436 9904 14464
rect 4479 14433 4491 14436
rect 4433 14427 4491 14433
rect 1673 14399 1731 14405
rect 1673 14365 1685 14399
rect 1719 14365 1731 14399
rect 1673 14359 1731 14365
rect 2409 14399 2467 14405
rect 2409 14365 2421 14399
rect 2455 14365 2467 14399
rect 2409 14359 2467 14365
rect 1688 14328 1716 14359
rect 3326 14356 3332 14408
rect 3384 14396 3390 14408
rect 3421 14399 3479 14405
rect 3421 14396 3433 14399
rect 3384 14368 3433 14396
rect 3384 14356 3390 14368
rect 3421 14365 3433 14368
rect 3467 14365 3479 14399
rect 3421 14359 3479 14365
rect 8386 14356 8392 14408
rect 8444 14396 8450 14408
rect 8941 14399 8999 14405
rect 8941 14396 8953 14399
rect 8444 14368 8953 14396
rect 8444 14356 8450 14368
rect 8941 14365 8953 14368
rect 8987 14396 8999 14399
rect 9769 14399 9827 14405
rect 9769 14396 9781 14399
rect 8987 14368 9781 14396
rect 8987 14365 8999 14368
rect 8941 14359 8999 14365
rect 9769 14365 9781 14368
rect 9815 14365 9827 14399
rect 9876 14396 9904 14436
rect 9953 14433 9965 14467
rect 9999 14464 10011 14467
rect 10594 14464 10600 14476
rect 9999 14436 10600 14464
rect 9999 14433 10011 14436
rect 9953 14427 10011 14433
rect 10594 14424 10600 14436
rect 10652 14424 10658 14476
rect 10318 14396 10324 14408
rect 9876 14368 10324 14396
rect 9769 14359 9827 14365
rect 10318 14356 10324 14368
rect 10376 14356 10382 14408
rect 11146 14356 11152 14408
rect 11204 14396 11210 14408
rect 12342 14396 12348 14408
rect 11204 14368 12348 14396
rect 11204 14356 11210 14368
rect 12342 14356 12348 14368
rect 12400 14396 12406 14408
rect 12437 14399 12495 14405
rect 12437 14396 12449 14399
rect 12400 14368 12449 14396
rect 12400 14356 12406 14368
rect 12437 14365 12449 14368
rect 12483 14365 12495 14399
rect 12437 14359 12495 14365
rect 3145 14331 3203 14337
rect 3145 14328 3157 14331
rect 1688 14300 3157 14328
rect 3145 14297 3157 14300
rect 3191 14297 3203 14331
rect 3145 14291 3203 14297
rect 8202 14288 8208 14340
rect 8260 14328 8266 14340
rect 8260 14300 12848 14328
rect 8260 14288 8266 14300
rect 4062 14220 4068 14272
rect 4120 14260 4126 14272
rect 4157 14263 4215 14269
rect 4157 14260 4169 14263
rect 4120 14232 4169 14260
rect 4120 14220 4126 14232
rect 4157 14229 4169 14232
rect 4203 14229 4215 14263
rect 4157 14223 4215 14229
rect 4246 14220 4252 14272
rect 4304 14260 4310 14272
rect 4798 14260 4804 14272
rect 4304 14232 4349 14260
rect 4759 14232 4804 14260
rect 4304 14220 4310 14232
rect 4798 14220 4804 14232
rect 4856 14260 4862 14272
rect 5445 14263 5503 14269
rect 5445 14260 5457 14263
rect 4856 14232 5457 14260
rect 4856 14220 4862 14232
rect 5445 14229 5457 14232
rect 5491 14229 5503 14263
rect 5445 14223 5503 14229
rect 5718 14220 5724 14272
rect 5776 14260 5782 14272
rect 6181 14263 6239 14269
rect 6181 14260 6193 14263
rect 5776 14232 6193 14260
rect 5776 14220 5782 14232
rect 6181 14229 6193 14232
rect 6227 14260 6239 14263
rect 6546 14260 6552 14272
rect 6227 14232 6552 14260
rect 6227 14229 6239 14232
rect 6181 14223 6239 14229
rect 6546 14220 6552 14232
rect 6604 14220 6610 14272
rect 8478 14260 8484 14272
rect 8439 14232 8484 14260
rect 8478 14220 8484 14232
rect 8536 14260 8542 14272
rect 9674 14260 9680 14272
rect 8536 14232 9680 14260
rect 8536 14220 8542 14232
rect 9674 14220 9680 14232
rect 9732 14220 9738 14272
rect 10778 14220 10784 14272
rect 10836 14260 10842 14272
rect 11149 14263 11207 14269
rect 11149 14260 11161 14263
rect 10836 14232 11161 14260
rect 10836 14220 10842 14232
rect 11149 14229 11161 14232
rect 11195 14229 11207 14263
rect 11149 14223 11207 14229
rect 11701 14263 11759 14269
rect 11701 14229 11713 14263
rect 11747 14260 11759 14263
rect 11882 14260 11888 14272
rect 11747 14232 11888 14260
rect 11747 14229 11759 14232
rect 11701 14223 11759 14229
rect 11882 14220 11888 14232
rect 11940 14220 11946 14272
rect 12820 14269 12848 14300
rect 12805 14263 12863 14269
rect 12805 14229 12817 14263
rect 12851 14260 12863 14263
rect 12894 14260 12900 14272
rect 12851 14232 12900 14260
rect 12851 14229 12863 14232
rect 12805 14223 12863 14229
rect 12894 14220 12900 14232
rect 12952 14220 12958 14272
rect 1104 14170 22056 14192
rect 1104 14118 6148 14170
rect 6200 14118 6212 14170
rect 6264 14118 6276 14170
rect 6328 14118 6340 14170
rect 6392 14118 6404 14170
rect 6456 14118 11346 14170
rect 11398 14118 11410 14170
rect 11462 14118 11474 14170
rect 11526 14118 11538 14170
rect 11590 14118 11602 14170
rect 11654 14118 16544 14170
rect 16596 14118 16608 14170
rect 16660 14118 16672 14170
rect 16724 14118 16736 14170
rect 16788 14118 16800 14170
rect 16852 14118 21742 14170
rect 21794 14118 21806 14170
rect 21858 14118 21870 14170
rect 21922 14118 21934 14170
rect 21986 14118 21998 14170
rect 22050 14118 22056 14170
rect 1104 14096 22056 14118
rect 1946 14056 1952 14068
rect 1907 14028 1952 14056
rect 1946 14016 1952 14028
rect 2004 14016 2010 14068
rect 2593 14059 2651 14065
rect 2593 14025 2605 14059
rect 2639 14056 2651 14059
rect 2774 14056 2780 14068
rect 2639 14028 2780 14056
rect 2639 14025 2651 14028
rect 2593 14019 2651 14025
rect 2774 14016 2780 14028
rect 2832 14016 2838 14068
rect 4062 14056 4068 14068
rect 4023 14028 4068 14056
rect 4062 14016 4068 14028
rect 4120 14016 4126 14068
rect 4890 14056 4896 14068
rect 4851 14028 4896 14056
rect 4890 14016 4896 14028
rect 4948 14016 4954 14068
rect 7374 14016 7380 14068
rect 7432 14056 7438 14068
rect 7929 14059 7987 14065
rect 7929 14056 7941 14059
rect 7432 14028 7941 14056
rect 7432 14016 7438 14028
rect 7929 14025 7941 14028
rect 7975 14025 7987 14059
rect 7929 14019 7987 14025
rect 8202 14016 8208 14068
rect 8260 14056 8266 14068
rect 8297 14059 8355 14065
rect 8297 14056 8309 14059
rect 8260 14028 8309 14056
rect 8260 14016 8266 14028
rect 8297 14025 8309 14028
rect 8343 14025 8355 14059
rect 9398 14056 9404 14068
rect 9359 14028 9404 14056
rect 8297 14019 8355 14025
rect 9398 14016 9404 14028
rect 9456 14016 9462 14068
rect 10410 14056 10416 14068
rect 10371 14028 10416 14056
rect 10410 14016 10416 14028
rect 10468 14016 10474 14068
rect 10778 14056 10784 14068
rect 10739 14028 10784 14056
rect 10778 14016 10784 14028
rect 10836 14016 10842 14068
rect 11517 14059 11575 14065
rect 11517 14025 11529 14059
rect 11563 14025 11575 14059
rect 12529 14059 12587 14065
rect 12529 14056 12541 14059
rect 11517 14019 11575 14025
rect 11716 14028 12541 14056
rect 4798 13988 4804 14000
rect 3620 13960 4804 13988
rect 2133 13923 2191 13929
rect 2133 13889 2145 13923
rect 2179 13889 2191 13923
rect 2406 13920 2412 13932
rect 2367 13892 2412 13920
rect 2133 13883 2191 13889
rect 2148 13852 2176 13883
rect 2406 13880 2412 13892
rect 2464 13880 2470 13932
rect 3620 13929 3648 13960
rect 4798 13948 4804 13960
rect 4856 13988 4862 14000
rect 5353 13991 5411 13997
rect 5353 13988 5365 13991
rect 4856 13960 5365 13988
rect 4856 13948 4862 13960
rect 5353 13957 5365 13960
rect 5399 13988 5411 13991
rect 6178 13988 6184 14000
rect 5399 13960 6184 13988
rect 5399 13957 5411 13960
rect 5353 13951 5411 13957
rect 6178 13948 6184 13960
rect 6236 13948 6242 14000
rect 7650 13988 7656 14000
rect 7563 13960 7656 13988
rect 7650 13948 7656 13960
rect 7708 13988 7714 14000
rect 8220 13988 8248 14016
rect 7708 13960 8248 13988
rect 9861 13991 9919 13997
rect 7708 13948 7714 13960
rect 9861 13957 9873 13991
rect 9907 13988 9919 13991
rect 11532 13988 11560 14019
rect 9907 13960 11560 13988
rect 9907 13957 9919 13960
rect 9861 13951 9919 13957
rect 3605 13923 3663 13929
rect 3605 13920 3617 13923
rect 3436 13892 3617 13920
rect 3142 13852 3148 13864
rect 2148 13824 3148 13852
rect 3142 13812 3148 13824
rect 3200 13812 3206 13864
rect 3436 13784 3464 13892
rect 3605 13889 3617 13892
rect 3651 13889 3663 13923
rect 3605 13883 3663 13889
rect 3697 13923 3755 13929
rect 3697 13889 3709 13923
rect 3743 13920 3755 13923
rect 4341 13923 4399 13929
rect 4341 13920 4353 13923
rect 3743 13892 4353 13920
rect 3743 13889 3755 13892
rect 3697 13883 3755 13889
rect 4341 13889 4353 13892
rect 4387 13889 4399 13923
rect 5258 13920 5264 13932
rect 5219 13892 5264 13920
rect 4341 13883 4399 13889
rect 5258 13880 5264 13892
rect 5316 13880 5322 13932
rect 8389 13923 8447 13929
rect 8389 13889 8401 13923
rect 8435 13920 8447 13923
rect 9766 13920 9772 13932
rect 8435 13892 9076 13920
rect 9727 13892 9772 13920
rect 8435 13889 8447 13892
rect 8389 13883 8447 13889
rect 9048 13864 9076 13892
rect 9766 13880 9772 13892
rect 9824 13880 9830 13932
rect 10873 13923 10931 13929
rect 10873 13889 10885 13923
rect 10919 13920 10931 13923
rect 11716 13920 11744 14028
rect 12529 14025 12541 14028
rect 12575 14025 12587 14059
rect 12894 14056 12900 14068
rect 12855 14028 12900 14056
rect 12529 14019 12587 14025
rect 12894 14016 12900 14028
rect 12952 14016 12958 14068
rect 11882 13988 11888 14000
rect 11843 13960 11888 13988
rect 11882 13948 11888 13960
rect 11940 13948 11946 14000
rect 12342 13948 12348 14000
rect 12400 13988 12406 14000
rect 12989 13991 13047 13997
rect 12989 13988 13001 13991
rect 12400 13960 13001 13988
rect 12400 13948 12406 13960
rect 12989 13957 13001 13960
rect 13035 13957 13047 13991
rect 12989 13951 13047 13957
rect 10919 13892 11744 13920
rect 13096 13892 13400 13920
rect 10919 13889 10931 13892
rect 10873 13883 10931 13889
rect 3513 13855 3571 13861
rect 3513 13821 3525 13855
rect 3559 13821 3571 13855
rect 5534 13852 5540 13864
rect 5495 13824 5540 13852
rect 3513 13815 3571 13821
rect 2976 13756 3464 13784
rect 3528 13784 3556 13815
rect 5534 13812 5540 13824
rect 5592 13852 5598 13864
rect 5905 13855 5963 13861
rect 5905 13852 5917 13855
rect 5592 13824 5917 13852
rect 5592 13812 5598 13824
rect 5905 13821 5917 13824
rect 5951 13821 5963 13855
rect 6638 13852 6644 13864
rect 6599 13824 6644 13852
rect 5905 13815 5963 13821
rect 6638 13812 6644 13824
rect 6696 13812 6702 13864
rect 8573 13855 8631 13861
rect 8573 13821 8585 13855
rect 8619 13821 8631 13855
rect 9030 13852 9036 13864
rect 8991 13824 9036 13852
rect 8573 13815 8631 13821
rect 4798 13784 4804 13796
rect 3528 13756 4804 13784
rect 2130 13676 2136 13728
rect 2188 13716 2194 13728
rect 2976 13725 3004 13756
rect 4798 13744 4804 13756
rect 4856 13744 4862 13796
rect 8588 13784 8616 13815
rect 9030 13812 9036 13824
rect 9088 13812 9094 13864
rect 10045 13855 10103 13861
rect 10045 13821 10057 13855
rect 10091 13852 10103 13855
rect 11057 13855 11115 13861
rect 10091 13824 10180 13852
rect 10091 13821 10103 13824
rect 10045 13815 10103 13821
rect 10152 13796 10180 13824
rect 11057 13821 11069 13855
rect 11103 13821 11115 13855
rect 11974 13852 11980 13864
rect 11935 13824 11980 13852
rect 11057 13815 11115 13821
rect 9950 13784 9956 13796
rect 8588 13756 9956 13784
rect 9950 13744 9956 13756
rect 10008 13744 10014 13796
rect 10134 13744 10140 13796
rect 10192 13744 10198 13796
rect 11072 13784 11100 13815
rect 11974 13812 11980 13824
rect 12032 13812 12038 13864
rect 12161 13855 12219 13861
rect 12161 13821 12173 13855
rect 12207 13821 12219 13855
rect 12161 13815 12219 13821
rect 12176 13784 12204 13815
rect 13096 13784 13124 13892
rect 13173 13855 13231 13861
rect 13173 13821 13185 13855
rect 13219 13821 13231 13855
rect 13173 13815 13231 13821
rect 11072 13756 11192 13784
rect 12176 13756 13124 13784
rect 2961 13719 3019 13725
rect 2961 13716 2973 13719
rect 2188 13688 2973 13716
rect 2188 13676 2194 13688
rect 2961 13685 2973 13688
rect 3007 13685 3019 13719
rect 2961 13679 3019 13685
rect 3234 13676 3240 13728
rect 3292 13716 3298 13728
rect 8478 13716 8484 13728
rect 3292 13688 8484 13716
rect 3292 13676 3298 13688
rect 8478 13676 8484 13688
rect 8536 13676 8542 13728
rect 11164 13716 11192 13756
rect 13078 13716 13084 13728
rect 11164 13688 13084 13716
rect 13078 13676 13084 13688
rect 13136 13676 13142 13728
rect 13188 13716 13216 13815
rect 13372 13784 13400 13892
rect 19978 13784 19984 13796
rect 13372 13756 19984 13784
rect 19978 13744 19984 13756
rect 20036 13744 20042 13796
rect 15654 13716 15660 13728
rect 13188 13688 15660 13716
rect 15654 13676 15660 13688
rect 15712 13676 15718 13728
rect 1104 13626 21896 13648
rect 1104 13574 3549 13626
rect 3601 13574 3613 13626
rect 3665 13574 3677 13626
rect 3729 13574 3741 13626
rect 3793 13574 3805 13626
rect 3857 13574 8747 13626
rect 8799 13574 8811 13626
rect 8863 13574 8875 13626
rect 8927 13574 8939 13626
rect 8991 13574 9003 13626
rect 9055 13574 13945 13626
rect 13997 13574 14009 13626
rect 14061 13574 14073 13626
rect 14125 13574 14137 13626
rect 14189 13574 14201 13626
rect 14253 13574 19143 13626
rect 19195 13574 19207 13626
rect 19259 13574 19271 13626
rect 19323 13574 19335 13626
rect 19387 13574 19399 13626
rect 19451 13574 21896 13626
rect 1104 13552 21896 13574
rect 4157 13515 4215 13521
rect 4157 13481 4169 13515
rect 4203 13512 4215 13515
rect 4246 13512 4252 13524
rect 4203 13484 4252 13512
rect 4203 13481 4215 13484
rect 4157 13475 4215 13481
rect 4246 13472 4252 13484
rect 4304 13472 4310 13524
rect 7190 13472 7196 13524
rect 7248 13512 7254 13524
rect 7745 13515 7803 13521
rect 7745 13512 7757 13515
rect 7248 13484 7757 13512
rect 7248 13472 7254 13484
rect 7745 13481 7757 13484
rect 7791 13481 7803 13515
rect 7745 13475 7803 13481
rect 10870 13472 10876 13524
rect 10928 13512 10934 13524
rect 12069 13515 12127 13521
rect 12069 13512 12081 13515
rect 10928 13484 12081 13512
rect 10928 13472 10934 13484
rect 12069 13481 12081 13484
rect 12115 13481 12127 13515
rect 12069 13475 12127 13481
rect 6825 13447 6883 13453
rect 6825 13444 6837 13447
rect 2332 13416 6837 13444
rect 1946 13376 1952 13388
rect 1907 13348 1952 13376
rect 1946 13336 1952 13348
rect 2004 13336 2010 13388
rect 1486 13200 1492 13252
rect 1544 13240 1550 13252
rect 2130 13240 2136 13252
rect 1544 13212 2136 13240
rect 1544 13200 1550 13212
rect 2130 13200 2136 13212
rect 2188 13200 2194 13252
rect 1397 13175 1455 13181
rect 1397 13141 1409 13175
rect 1443 13172 1455 13175
rect 1578 13172 1584 13184
rect 1443 13144 1584 13172
rect 1443 13141 1455 13144
rect 1397 13135 1455 13141
rect 1578 13132 1584 13144
rect 1636 13172 1642 13184
rect 2041 13175 2099 13181
rect 2041 13172 2053 13175
rect 1636 13144 2053 13172
rect 1636 13132 1642 13144
rect 2041 13141 2053 13144
rect 2087 13172 2099 13175
rect 2332 13172 2360 13416
rect 3142 13376 3148 13388
rect 3103 13348 3148 13376
rect 3142 13336 3148 13348
rect 3200 13336 3206 13388
rect 4798 13376 4804 13388
rect 4759 13348 4804 13376
rect 4798 13336 4804 13348
rect 4856 13336 4862 13388
rect 5258 13336 5264 13388
rect 5316 13376 5322 13388
rect 6288 13385 6316 13416
rect 6825 13413 6837 13416
rect 6871 13444 6883 13447
rect 7650 13444 7656 13456
rect 6871 13416 7656 13444
rect 6871 13413 6883 13416
rect 6825 13407 6883 13413
rect 7650 13404 7656 13416
rect 7708 13404 7714 13456
rect 10229 13447 10287 13453
rect 10229 13444 10241 13447
rect 8220 13416 10241 13444
rect 5353 13379 5411 13385
rect 5353 13376 5365 13379
rect 5316 13348 5365 13376
rect 5316 13336 5322 13348
rect 5353 13345 5365 13348
rect 5399 13345 5411 13379
rect 5353 13339 5411 13345
rect 6273 13379 6331 13385
rect 6273 13345 6285 13379
rect 6319 13345 6331 13379
rect 6273 13339 6331 13345
rect 6457 13379 6515 13385
rect 6457 13345 6469 13379
rect 6503 13376 6515 13379
rect 6546 13376 6552 13388
rect 6503 13348 6552 13376
rect 6503 13345 6515 13348
rect 6457 13339 6515 13345
rect 6546 13336 6552 13348
rect 6604 13336 6610 13388
rect 8220 13385 8248 13416
rect 10229 13413 10241 13416
rect 10275 13413 10287 13447
rect 10229 13407 10287 13413
rect 8205 13379 8263 13385
rect 8205 13345 8217 13379
rect 8251 13345 8263 13379
rect 8205 13339 8263 13345
rect 8294 13336 8300 13388
rect 8352 13376 8358 13388
rect 9766 13376 9772 13388
rect 8352 13348 8397 13376
rect 9727 13348 9772 13376
rect 8352 13336 8358 13348
rect 9766 13336 9772 13348
rect 9824 13336 9830 13388
rect 10870 13376 10876 13388
rect 10831 13348 10876 13376
rect 10870 13336 10876 13348
rect 10928 13336 10934 13388
rect 12713 13379 12771 13385
rect 12713 13345 12725 13379
rect 12759 13376 12771 13379
rect 17954 13376 17960 13388
rect 12759 13348 17960 13376
rect 12759 13345 12771 13348
rect 12713 13339 12771 13345
rect 17954 13336 17960 13348
rect 18012 13336 18018 13388
rect 3421 13311 3479 13317
rect 3421 13277 3433 13311
rect 3467 13308 3479 13311
rect 4522 13308 4528 13320
rect 3467 13280 4528 13308
rect 3467 13277 3479 13280
rect 3421 13271 3479 13277
rect 4522 13268 4528 13280
rect 4580 13268 4586 13320
rect 6178 13308 6184 13320
rect 6139 13280 6184 13308
rect 6178 13268 6184 13280
rect 6236 13268 6242 13320
rect 9493 13311 9551 13317
rect 9493 13277 9505 13311
rect 9539 13308 9551 13311
rect 10686 13308 10692 13320
rect 9539 13280 10692 13308
rect 9539 13277 9551 13280
rect 9493 13271 9551 13277
rect 10686 13268 10692 13280
rect 10744 13268 10750 13320
rect 11698 13268 11704 13320
rect 11756 13308 11762 13320
rect 12437 13311 12495 13317
rect 12437 13308 12449 13311
rect 11756 13280 12449 13308
rect 11756 13268 11762 13280
rect 12437 13277 12449 13280
rect 12483 13277 12495 13311
rect 12437 13271 12495 13277
rect 3881 13243 3939 13249
rect 3881 13209 3893 13243
rect 3927 13240 3939 13243
rect 4062 13240 4068 13252
rect 3927 13212 4068 13240
rect 3927 13209 3939 13212
rect 3881 13203 3939 13209
rect 4062 13200 4068 13212
rect 4120 13240 4126 13252
rect 5902 13240 5908 13252
rect 4120 13212 5908 13240
rect 4120 13200 4126 13212
rect 2498 13172 2504 13184
rect 2087 13144 2360 13172
rect 2459 13144 2504 13172
rect 2087 13141 2099 13144
rect 2041 13135 2099 13141
rect 2498 13132 2504 13144
rect 2556 13132 2562 13184
rect 4540 13181 4568 13212
rect 5902 13200 5908 13212
rect 5960 13200 5966 13252
rect 8113 13243 8171 13249
rect 8113 13209 8125 13243
rect 8159 13240 8171 13243
rect 8941 13243 8999 13249
rect 8941 13240 8953 13243
rect 8159 13212 8953 13240
rect 8159 13209 8171 13212
rect 8113 13203 8171 13209
rect 8941 13209 8953 13212
rect 8987 13209 8999 13243
rect 8941 13203 8999 13209
rect 10502 13200 10508 13252
rect 10560 13240 10566 13252
rect 11333 13243 11391 13249
rect 11333 13240 11345 13243
rect 10560 13212 11345 13240
rect 10560 13200 10566 13212
rect 11333 13209 11345 13212
rect 11379 13240 11391 13243
rect 11974 13240 11980 13252
rect 11379 13212 11980 13240
rect 11379 13209 11391 13212
rect 11333 13203 11391 13209
rect 11974 13200 11980 13212
rect 12032 13200 12038 13252
rect 12529 13243 12587 13249
rect 12529 13240 12541 13243
rect 12084 13212 12541 13240
rect 12084 13184 12112 13212
rect 12529 13209 12541 13212
rect 12575 13209 12587 13243
rect 12529 13203 12587 13209
rect 4525 13175 4583 13181
rect 4525 13141 4537 13175
rect 4571 13141 4583 13175
rect 4525 13135 4583 13141
rect 4617 13175 4675 13181
rect 4617 13141 4629 13175
rect 4663 13172 4675 13175
rect 4982 13172 4988 13184
rect 4663 13144 4988 13172
rect 4663 13141 4675 13144
rect 4617 13135 4675 13141
rect 4982 13132 4988 13144
rect 5040 13132 5046 13184
rect 5810 13172 5816 13184
rect 5771 13144 5816 13172
rect 5810 13132 5816 13144
rect 5868 13132 5874 13184
rect 7285 13175 7343 13181
rect 7285 13141 7297 13175
rect 7331 13172 7343 13175
rect 7926 13172 7932 13184
rect 7331 13144 7932 13172
rect 7331 13141 7343 13144
rect 7285 13135 7343 13141
rect 7926 13132 7932 13144
rect 7984 13172 7990 13184
rect 10597 13175 10655 13181
rect 10597 13172 10609 13175
rect 7984 13144 10609 13172
rect 7984 13132 7990 13144
rect 10597 13141 10609 13144
rect 10643 13141 10655 13175
rect 10597 13135 10655 13141
rect 10686 13132 10692 13184
rect 10744 13172 10750 13184
rect 11793 13175 11851 13181
rect 10744 13144 10789 13172
rect 10744 13132 10750 13144
rect 11793 13141 11805 13175
rect 11839 13172 11851 13175
rect 12066 13172 12072 13184
rect 11839 13144 12072 13172
rect 11839 13141 11851 13144
rect 11793 13135 11851 13141
rect 12066 13132 12072 13144
rect 12124 13132 12130 13184
rect 1104 13082 22056 13104
rect 1104 13030 6148 13082
rect 6200 13030 6212 13082
rect 6264 13030 6276 13082
rect 6328 13030 6340 13082
rect 6392 13030 6404 13082
rect 6456 13030 11346 13082
rect 11398 13030 11410 13082
rect 11462 13030 11474 13082
rect 11526 13030 11538 13082
rect 11590 13030 11602 13082
rect 11654 13030 16544 13082
rect 16596 13030 16608 13082
rect 16660 13030 16672 13082
rect 16724 13030 16736 13082
rect 16788 13030 16800 13082
rect 16852 13030 21742 13082
rect 21794 13030 21806 13082
rect 21858 13030 21870 13082
rect 21922 13030 21934 13082
rect 21986 13030 21998 13082
rect 22050 13030 22056 13082
rect 1104 13008 22056 13030
rect 2685 12971 2743 12977
rect 2685 12937 2697 12971
rect 2731 12968 2743 12971
rect 2774 12968 2780 12980
rect 2731 12940 2780 12968
rect 2731 12937 2743 12940
rect 2685 12931 2743 12937
rect 2774 12928 2780 12940
rect 2832 12928 2838 12980
rect 5629 12971 5687 12977
rect 5629 12937 5641 12971
rect 5675 12968 5687 12971
rect 7377 12971 7435 12977
rect 7377 12968 7389 12971
rect 5675 12940 7389 12968
rect 5675 12937 5687 12940
rect 5629 12931 5687 12937
rect 7377 12937 7389 12940
rect 7423 12937 7435 12971
rect 7377 12931 7435 12937
rect 7650 12928 7656 12980
rect 7708 12968 7714 12980
rect 7745 12971 7803 12977
rect 7745 12968 7757 12971
rect 7708 12940 7757 12968
rect 7708 12928 7714 12940
rect 7745 12937 7757 12940
rect 7791 12968 7803 12971
rect 7834 12968 7840 12980
rect 7791 12940 7840 12968
rect 7791 12937 7803 12940
rect 7745 12931 7803 12937
rect 7834 12928 7840 12940
rect 7892 12928 7898 12980
rect 7944 12940 9628 12968
rect 2041 12903 2099 12909
rect 2041 12869 2053 12903
rect 2087 12900 2099 12903
rect 2406 12900 2412 12912
rect 2087 12872 2412 12900
rect 2087 12869 2099 12872
rect 2041 12863 2099 12869
rect 2406 12860 2412 12872
rect 2464 12860 2470 12912
rect 4798 12860 4804 12912
rect 4856 12900 4862 12912
rect 7944 12900 7972 12940
rect 4856 12872 7972 12900
rect 9600 12900 9628 12940
rect 9674 12928 9680 12980
rect 9732 12968 9738 12980
rect 11698 12968 11704 12980
rect 9732 12940 11704 12968
rect 9732 12928 9738 12940
rect 11698 12928 11704 12940
rect 11756 12928 11762 12980
rect 12158 12968 12164 12980
rect 12119 12940 12164 12968
rect 12158 12928 12164 12940
rect 12216 12928 12222 12980
rect 11974 12900 11980 12912
rect 9600 12872 11980 12900
rect 4856 12860 4862 12872
rect 11974 12860 11980 12872
rect 12032 12860 12038 12912
rect 1762 12832 1768 12844
rect 1723 12804 1768 12832
rect 1762 12792 1768 12804
rect 1820 12792 1826 12844
rect 2314 12792 2320 12844
rect 2372 12832 2378 12844
rect 2501 12835 2559 12841
rect 2501 12832 2513 12835
rect 2372 12804 2513 12832
rect 2372 12792 2378 12804
rect 2501 12801 2513 12804
rect 2547 12801 2559 12835
rect 2501 12795 2559 12801
rect 3513 12835 3571 12841
rect 3513 12801 3525 12835
rect 3559 12832 3571 12835
rect 4338 12832 4344 12844
rect 3559 12804 4344 12832
rect 3559 12801 3571 12804
rect 3513 12795 3571 12801
rect 4338 12792 4344 12804
rect 4396 12792 4402 12844
rect 7837 12835 7895 12841
rect 7837 12801 7849 12835
rect 7883 12832 7895 12835
rect 7926 12832 7932 12844
rect 7883 12804 7932 12832
rect 7883 12801 7895 12804
rect 7837 12795 7895 12801
rect 7926 12792 7932 12804
rect 7984 12832 7990 12844
rect 7984 12804 8524 12832
rect 7984 12792 7990 12804
rect 3234 12764 3240 12776
rect 3195 12736 3240 12764
rect 3234 12724 3240 12736
rect 3292 12724 3298 12776
rect 5718 12764 5724 12776
rect 5679 12736 5724 12764
rect 5718 12724 5724 12736
rect 5776 12724 5782 12776
rect 5813 12767 5871 12773
rect 5813 12733 5825 12767
rect 5859 12733 5871 12767
rect 7098 12764 7104 12776
rect 7059 12736 7104 12764
rect 5813 12727 5871 12733
rect 5626 12656 5632 12708
rect 5684 12696 5690 12708
rect 5828 12696 5856 12727
rect 7098 12724 7104 12736
rect 7156 12724 7162 12776
rect 8018 12764 8024 12776
rect 7979 12736 8024 12764
rect 8018 12724 8024 12736
rect 8076 12724 8082 12776
rect 8496 12764 8524 12804
rect 9122 12792 9128 12844
rect 9180 12832 9186 12844
rect 10137 12835 10195 12841
rect 10137 12832 10149 12835
rect 9180 12804 10149 12832
rect 9180 12792 9186 12804
rect 10137 12801 10149 12804
rect 10183 12801 10195 12835
rect 10781 12835 10839 12841
rect 10781 12832 10793 12835
rect 10137 12795 10195 12801
rect 10244 12804 10793 12832
rect 10244 12776 10272 12804
rect 10781 12801 10793 12804
rect 10827 12801 10839 12835
rect 10781 12795 10839 12801
rect 12529 12835 12587 12841
rect 12529 12801 12541 12835
rect 12575 12832 12587 12835
rect 13173 12835 13231 12841
rect 13173 12832 13185 12835
rect 12575 12804 13185 12832
rect 12575 12801 12587 12804
rect 12529 12795 12587 12801
rect 13173 12801 13185 12804
rect 13219 12801 13231 12835
rect 13173 12795 13231 12801
rect 9401 12767 9459 12773
rect 9401 12764 9413 12767
rect 8496 12736 9413 12764
rect 9401 12733 9413 12736
rect 9447 12733 9459 12767
rect 9401 12727 9459 12733
rect 9953 12767 10011 12773
rect 9953 12733 9965 12767
rect 9999 12733 10011 12767
rect 9953 12727 10011 12733
rect 10045 12767 10103 12773
rect 10045 12733 10057 12767
rect 10091 12764 10103 12767
rect 10226 12764 10232 12776
rect 10091 12736 10232 12764
rect 10091 12733 10103 12736
rect 10045 12727 10103 12733
rect 5684 12668 5856 12696
rect 9968 12696 9996 12727
rect 10226 12724 10232 12736
rect 10284 12724 10290 12776
rect 12621 12767 12679 12773
rect 12621 12764 12633 12767
rect 10520 12736 12633 12764
rect 10520 12705 10548 12736
rect 12621 12733 12633 12736
rect 12667 12733 12679 12767
rect 12621 12727 12679 12733
rect 12805 12767 12863 12773
rect 12805 12733 12817 12767
rect 12851 12733 12863 12767
rect 17126 12764 17132 12776
rect 12805 12727 12863 12733
rect 16546 12736 17132 12764
rect 10505 12699 10563 12705
rect 9968 12668 10088 12696
rect 5684 12656 5690 12668
rect 1486 12628 1492 12640
rect 1447 12600 1492 12628
rect 1486 12588 1492 12600
rect 1544 12588 1550 12640
rect 4982 12628 4988 12640
rect 4943 12600 4988 12628
rect 4982 12588 4988 12600
rect 5040 12588 5046 12640
rect 5258 12628 5264 12640
rect 5219 12600 5264 12628
rect 5258 12588 5264 12600
rect 5316 12588 5322 12640
rect 6362 12588 6368 12640
rect 6420 12628 6426 12640
rect 6549 12631 6607 12637
rect 6549 12628 6561 12631
rect 6420 12600 6561 12628
rect 6420 12588 6426 12600
rect 6549 12597 6561 12600
rect 6595 12628 6607 12631
rect 7650 12628 7656 12640
rect 6595 12600 7656 12628
rect 6595 12597 6607 12600
rect 6549 12591 6607 12597
rect 7650 12588 7656 12600
rect 7708 12588 7714 12640
rect 8110 12588 8116 12640
rect 8168 12628 8174 12640
rect 8389 12631 8447 12637
rect 8389 12628 8401 12631
rect 8168 12600 8401 12628
rect 8168 12588 8174 12600
rect 8389 12597 8401 12600
rect 8435 12597 8447 12631
rect 9122 12628 9128 12640
rect 9083 12600 9128 12628
rect 8389 12591 8447 12597
rect 9122 12588 9128 12600
rect 9180 12588 9186 12640
rect 10060 12628 10088 12668
rect 10505 12665 10517 12699
rect 10551 12665 10563 12699
rect 12820 12696 12848 12727
rect 16546 12696 16574 12736
rect 17126 12724 17132 12736
rect 17184 12724 17190 12776
rect 12820 12668 16574 12696
rect 10505 12659 10563 12665
rect 12710 12628 12716 12640
rect 10060 12600 12716 12628
rect 12710 12588 12716 12600
rect 12768 12588 12774 12640
rect 1104 12538 21896 12560
rect 1104 12486 3549 12538
rect 3601 12486 3613 12538
rect 3665 12486 3677 12538
rect 3729 12486 3741 12538
rect 3793 12486 3805 12538
rect 3857 12486 8747 12538
rect 8799 12486 8811 12538
rect 8863 12486 8875 12538
rect 8927 12486 8939 12538
rect 8991 12486 9003 12538
rect 9055 12486 13945 12538
rect 13997 12486 14009 12538
rect 14061 12486 14073 12538
rect 14125 12486 14137 12538
rect 14189 12486 14201 12538
rect 14253 12486 19143 12538
rect 19195 12486 19207 12538
rect 19259 12486 19271 12538
rect 19323 12486 19335 12538
rect 19387 12486 19399 12538
rect 19451 12486 21896 12538
rect 1104 12464 21896 12486
rect 1670 12424 1676 12436
rect 1631 12396 1676 12424
rect 1670 12384 1676 12396
rect 1728 12384 1734 12436
rect 4338 12424 4344 12436
rect 4299 12396 4344 12424
rect 4338 12384 4344 12396
rect 4396 12384 4402 12436
rect 5166 12384 5172 12436
rect 5224 12424 5230 12436
rect 5442 12424 5448 12436
rect 5224 12396 5448 12424
rect 5224 12384 5230 12396
rect 5442 12384 5448 12396
rect 5500 12384 5506 12436
rect 5718 12384 5724 12436
rect 5776 12424 5782 12436
rect 5813 12427 5871 12433
rect 5813 12424 5825 12427
rect 5776 12396 5825 12424
rect 5776 12384 5782 12396
rect 5813 12393 5825 12396
rect 5859 12393 5871 12427
rect 5813 12387 5871 12393
rect 6362 12384 6368 12436
rect 6420 12384 6426 12436
rect 6822 12424 6828 12436
rect 6783 12396 6828 12424
rect 6822 12384 6828 12396
rect 6880 12384 6886 12436
rect 8018 12424 8024 12436
rect 6932 12396 8024 12424
rect 2682 12316 2688 12368
rect 2740 12356 2746 12368
rect 6380 12356 6408 12384
rect 6546 12356 6552 12368
rect 2740 12328 6408 12356
rect 6472 12328 6552 12356
rect 2740 12316 2746 12328
rect 1946 12248 1952 12300
rect 2004 12288 2010 12300
rect 2317 12291 2375 12297
rect 2317 12288 2329 12291
rect 2004 12260 2329 12288
rect 2004 12248 2010 12260
rect 2317 12257 2329 12260
rect 2363 12288 2375 12291
rect 2406 12288 2412 12300
rect 2363 12260 2412 12288
rect 2363 12257 2375 12260
rect 2317 12251 2375 12257
rect 2406 12248 2412 12260
rect 2464 12248 2470 12300
rect 4985 12291 5043 12297
rect 4985 12257 4997 12291
rect 5031 12288 5043 12291
rect 5166 12288 5172 12300
rect 5031 12260 5172 12288
rect 5031 12257 5043 12260
rect 4985 12251 5043 12257
rect 5166 12248 5172 12260
rect 5224 12248 5230 12300
rect 6472 12297 6500 12328
rect 6546 12316 6552 12328
rect 6604 12356 6610 12368
rect 6932 12356 6960 12396
rect 8018 12384 8024 12396
rect 8076 12424 8082 12436
rect 8076 12396 8432 12424
rect 8076 12384 8082 12396
rect 8294 12356 8300 12368
rect 6604 12328 6960 12356
rect 7300 12328 8300 12356
rect 6604 12316 6610 12328
rect 7300 12297 7328 12328
rect 8294 12316 8300 12328
rect 8352 12316 8358 12368
rect 8404 12356 8432 12396
rect 8570 12384 8576 12436
rect 8628 12424 8634 12436
rect 9309 12427 9367 12433
rect 9309 12424 9321 12427
rect 8628 12396 9321 12424
rect 8628 12384 8634 12396
rect 9309 12393 9321 12396
rect 9355 12393 9367 12427
rect 9309 12387 9367 12393
rect 9950 12384 9956 12436
rect 10008 12424 10014 12436
rect 13170 12424 13176 12436
rect 10008 12396 13176 12424
rect 10008 12384 10014 12396
rect 13170 12384 13176 12396
rect 13228 12384 13234 12436
rect 8404 12328 11008 12356
rect 6457 12291 6515 12297
rect 6457 12257 6469 12291
rect 6503 12257 6515 12291
rect 6457 12251 6515 12257
rect 7285 12291 7343 12297
rect 7285 12257 7297 12291
rect 7331 12257 7343 12291
rect 7466 12288 7472 12300
rect 7427 12260 7472 12288
rect 7285 12251 7343 12257
rect 7466 12248 7472 12260
rect 7524 12248 7530 12300
rect 8018 12248 8024 12300
rect 8076 12288 8082 12300
rect 8202 12288 8208 12300
rect 8076 12260 8208 12288
rect 8076 12248 8082 12260
rect 8202 12248 8208 12260
rect 8260 12248 8266 12300
rect 8481 12291 8539 12297
rect 8481 12257 8493 12291
rect 8527 12288 8539 12291
rect 8570 12288 8576 12300
rect 8527 12260 8576 12288
rect 8527 12257 8539 12260
rect 8481 12251 8539 12257
rect 8570 12248 8576 12260
rect 8628 12248 8634 12300
rect 9582 12248 9588 12300
rect 9640 12288 9646 12300
rect 9861 12291 9919 12297
rect 9861 12288 9873 12291
rect 9640 12260 9873 12288
rect 9640 12248 9646 12260
rect 9861 12257 9873 12260
rect 9907 12257 9919 12291
rect 10410 12288 10416 12300
rect 9861 12251 9919 12257
rect 10060 12260 10416 12288
rect 10060 12232 10088 12260
rect 10410 12248 10416 12260
rect 10468 12248 10474 12300
rect 10870 12288 10876 12300
rect 10831 12260 10876 12288
rect 10870 12248 10876 12260
rect 10928 12248 10934 12300
rect 10980 12288 11008 12328
rect 10980 12260 11928 12288
rect 1857 12223 1915 12229
rect 1857 12189 1869 12223
rect 1903 12220 1915 12223
rect 3234 12220 3240 12232
rect 1903 12192 3240 12220
rect 1903 12189 1915 12192
rect 1857 12183 1915 12189
rect 3234 12180 3240 12192
rect 3292 12180 3298 12232
rect 4801 12223 4859 12229
rect 4801 12189 4813 12223
rect 4847 12220 4859 12223
rect 5258 12220 5264 12232
rect 4847 12192 5264 12220
rect 4847 12189 4859 12192
rect 4801 12183 4859 12189
rect 5258 12180 5264 12192
rect 5316 12180 5322 12232
rect 5902 12180 5908 12232
rect 5960 12220 5966 12232
rect 6181 12223 6239 12229
rect 6181 12220 6193 12223
rect 5960 12192 6193 12220
rect 5960 12180 5966 12192
rect 6181 12189 6193 12192
rect 6227 12189 6239 12223
rect 6181 12183 6239 12189
rect 7098 12180 7104 12232
rect 7156 12220 7162 12232
rect 7193 12223 7251 12229
rect 7193 12220 7205 12223
rect 7156 12192 7205 12220
rect 7156 12180 7162 12192
rect 7193 12189 7205 12192
rect 7239 12189 7251 12223
rect 7193 12183 7251 12189
rect 8110 12180 8116 12232
rect 8168 12220 8174 12232
rect 8297 12223 8355 12229
rect 8297 12220 8309 12223
rect 8168 12192 8309 12220
rect 8168 12180 8174 12192
rect 8297 12189 8309 12192
rect 8343 12189 8355 12223
rect 8297 12183 8355 12189
rect 9033 12223 9091 12229
rect 9033 12189 9045 12223
rect 9079 12220 9091 12223
rect 10042 12220 10048 12232
rect 9079 12192 10048 12220
rect 9079 12189 9091 12192
rect 9033 12183 9091 12189
rect 10042 12180 10048 12192
rect 10100 12180 10106 12232
rect 10134 12180 10140 12232
rect 10192 12220 10198 12232
rect 10781 12223 10839 12229
rect 10781 12220 10793 12223
rect 10192 12192 10793 12220
rect 10192 12180 10198 12192
rect 10781 12189 10793 12192
rect 10827 12189 10839 12223
rect 11790 12220 11796 12232
rect 11751 12192 11796 12220
rect 10781 12183 10839 12189
rect 11790 12180 11796 12192
rect 11848 12180 11854 12232
rect 11900 12220 11928 12260
rect 17037 12223 17095 12229
rect 11900 12192 12388 12220
rect 12360 12164 12388 12192
rect 17037 12189 17049 12223
rect 17083 12220 17095 12223
rect 17083 12192 17448 12220
rect 17083 12189 17095 12192
rect 17037 12183 17095 12189
rect 2409 12155 2467 12161
rect 2409 12121 2421 12155
rect 2455 12152 2467 12155
rect 2455 12124 3096 12152
rect 2455 12121 2467 12124
rect 2409 12115 2467 12121
rect 3068 12096 3096 12124
rect 7650 12112 7656 12164
rect 7708 12152 7714 12164
rect 9677 12155 9735 12161
rect 7708 12124 8248 12152
rect 7708 12112 7714 12124
rect 8220 12096 8248 12124
rect 9677 12121 9689 12155
rect 9723 12152 9735 12155
rect 11333 12155 11391 12161
rect 11333 12152 11345 12155
rect 9723 12124 11345 12152
rect 9723 12121 9735 12124
rect 9677 12115 9735 12121
rect 11333 12121 11345 12124
rect 11379 12121 11391 12155
rect 11333 12115 11391 12121
rect 11698 12112 11704 12164
rect 11756 12152 11762 12164
rect 12038 12155 12096 12161
rect 12038 12152 12050 12155
rect 11756 12124 12050 12152
rect 11756 12112 11762 12124
rect 12038 12121 12050 12124
rect 12084 12121 12096 12155
rect 12038 12115 12096 12121
rect 12342 12112 12348 12164
rect 12400 12152 12406 12164
rect 16792 12155 16850 12161
rect 12400 12124 16712 12152
rect 12400 12112 12406 12124
rect 1394 12044 1400 12096
rect 1452 12084 1458 12096
rect 2501 12087 2559 12093
rect 2501 12084 2513 12087
rect 1452 12056 2513 12084
rect 1452 12044 1458 12056
rect 2501 12053 2513 12056
rect 2547 12084 2559 12087
rect 2682 12084 2688 12096
rect 2547 12056 2688 12084
rect 2547 12053 2559 12056
rect 2501 12047 2559 12053
rect 2682 12044 2688 12056
rect 2740 12044 2746 12096
rect 2866 12084 2872 12096
rect 2827 12056 2872 12084
rect 2866 12044 2872 12056
rect 2924 12044 2930 12096
rect 3050 12044 3056 12096
rect 3108 12084 3114 12096
rect 3145 12087 3203 12093
rect 3145 12084 3157 12087
rect 3108 12056 3157 12084
rect 3108 12044 3114 12056
rect 3145 12053 3157 12056
rect 3191 12053 3203 12087
rect 3970 12084 3976 12096
rect 3931 12056 3976 12084
rect 3145 12047 3203 12053
rect 3970 12044 3976 12056
rect 4028 12044 4034 12096
rect 4706 12084 4712 12096
rect 4667 12056 4712 12084
rect 4706 12044 4712 12056
rect 4764 12044 4770 12096
rect 5350 12084 5356 12096
rect 5311 12056 5356 12084
rect 5350 12044 5356 12056
rect 5408 12044 5414 12096
rect 6273 12087 6331 12093
rect 6273 12053 6285 12087
rect 6319 12084 6331 12087
rect 6638 12084 6644 12096
rect 6319 12056 6644 12084
rect 6319 12053 6331 12056
rect 6273 12047 6331 12053
rect 6638 12044 6644 12056
rect 6696 12044 6702 12096
rect 7374 12044 7380 12096
rect 7432 12084 7438 12096
rect 7837 12087 7895 12093
rect 7837 12084 7849 12087
rect 7432 12056 7849 12084
rect 7432 12044 7438 12056
rect 7837 12053 7849 12056
rect 7883 12053 7895 12087
rect 8202 12084 8208 12096
rect 8163 12056 8208 12084
rect 7837 12047 7895 12053
rect 8202 12044 8208 12056
rect 8260 12044 8266 12096
rect 9769 12087 9827 12093
rect 9769 12053 9781 12087
rect 9815 12084 9827 12087
rect 10321 12087 10379 12093
rect 10321 12084 10333 12087
rect 9815 12056 10333 12084
rect 9815 12053 9827 12056
rect 9769 12047 9827 12053
rect 10321 12053 10333 12056
rect 10367 12053 10379 12087
rect 10321 12047 10379 12053
rect 10410 12044 10416 12096
rect 10468 12084 10474 12096
rect 10689 12087 10747 12093
rect 10689 12084 10701 12087
rect 10468 12056 10701 12084
rect 10468 12044 10474 12056
rect 10689 12053 10701 12056
rect 10735 12053 10747 12087
rect 13170 12084 13176 12096
rect 13131 12056 13176 12084
rect 10689 12047 10747 12053
rect 13170 12044 13176 12056
rect 13228 12044 13234 12096
rect 13541 12087 13599 12093
rect 13541 12053 13553 12087
rect 13587 12084 13599 12087
rect 13722 12084 13728 12096
rect 13587 12056 13728 12084
rect 13587 12053 13599 12056
rect 13541 12047 13599 12053
rect 13722 12044 13728 12056
rect 13780 12044 13786 12096
rect 15654 12084 15660 12096
rect 15615 12056 15660 12084
rect 15654 12044 15660 12056
rect 15712 12044 15718 12096
rect 16684 12084 16712 12124
rect 16792 12121 16804 12155
rect 16838 12152 16850 12155
rect 17126 12152 17132 12164
rect 16838 12124 17132 12152
rect 16838 12121 16850 12124
rect 16792 12115 16850 12121
rect 17126 12112 17132 12124
rect 17184 12112 17190 12164
rect 17034 12084 17040 12096
rect 16684 12056 17040 12084
rect 17034 12044 17040 12056
rect 17092 12044 17098 12096
rect 17420 12093 17448 12192
rect 17405 12087 17463 12093
rect 17405 12053 17417 12087
rect 17451 12084 17463 12087
rect 18322 12084 18328 12096
rect 17451 12056 18328 12084
rect 17451 12053 17463 12056
rect 17405 12047 17463 12053
rect 18322 12044 18328 12056
rect 18380 12044 18386 12096
rect 19889 12087 19947 12093
rect 19889 12053 19901 12087
rect 19935 12084 19947 12087
rect 21358 12084 21364 12096
rect 19935 12056 21364 12084
rect 19935 12053 19947 12056
rect 19889 12047 19947 12053
rect 21358 12044 21364 12056
rect 21416 12044 21422 12096
rect 1104 11994 22056 12016
rect 1104 11942 6148 11994
rect 6200 11942 6212 11994
rect 6264 11942 6276 11994
rect 6328 11942 6340 11994
rect 6392 11942 6404 11994
rect 6456 11942 11346 11994
rect 11398 11942 11410 11994
rect 11462 11942 11474 11994
rect 11526 11942 11538 11994
rect 11590 11942 11602 11994
rect 11654 11942 16544 11994
rect 16596 11942 16608 11994
rect 16660 11942 16672 11994
rect 16724 11942 16736 11994
rect 16788 11942 16800 11994
rect 16852 11942 21742 11994
rect 21794 11942 21806 11994
rect 21858 11942 21870 11994
rect 21922 11942 21934 11994
rect 21986 11942 21998 11994
rect 22050 11942 22056 11994
rect 1104 11920 22056 11942
rect 2501 11883 2559 11889
rect 2501 11849 2513 11883
rect 2547 11880 2559 11883
rect 2866 11880 2872 11892
rect 2547 11852 2872 11880
rect 2547 11849 2559 11852
rect 2501 11843 2559 11849
rect 2866 11840 2872 11852
rect 2924 11840 2930 11892
rect 3329 11883 3387 11889
rect 3329 11849 3341 11883
rect 3375 11880 3387 11883
rect 3970 11880 3976 11892
rect 3375 11852 3976 11880
rect 3375 11849 3387 11852
rect 3329 11843 3387 11849
rect 3970 11840 3976 11852
rect 4028 11880 4034 11892
rect 4341 11883 4399 11889
rect 4341 11880 4353 11883
rect 4028 11852 4353 11880
rect 4028 11840 4034 11852
rect 4341 11849 4353 11852
rect 4387 11849 4399 11883
rect 4341 11843 4399 11849
rect 4706 11840 4712 11892
rect 4764 11880 4770 11892
rect 4985 11883 5043 11889
rect 4985 11880 4997 11883
rect 4764 11852 4997 11880
rect 4764 11840 4770 11852
rect 4985 11849 4997 11852
rect 5031 11849 5043 11883
rect 5350 11880 5356 11892
rect 5311 11852 5356 11880
rect 4985 11843 5043 11849
rect 5350 11840 5356 11852
rect 5408 11840 5414 11892
rect 5445 11883 5503 11889
rect 5445 11849 5457 11883
rect 5491 11880 5503 11883
rect 5810 11880 5816 11892
rect 5491 11852 5816 11880
rect 5491 11849 5503 11852
rect 5445 11843 5503 11849
rect 5810 11840 5816 11852
rect 5868 11840 5874 11892
rect 5994 11840 6000 11892
rect 6052 11880 6058 11892
rect 6365 11883 6423 11889
rect 6365 11880 6377 11883
rect 6052 11852 6377 11880
rect 6052 11840 6058 11852
rect 6365 11849 6377 11852
rect 6411 11849 6423 11883
rect 6365 11843 6423 11849
rect 6825 11883 6883 11889
rect 6825 11849 6837 11883
rect 6871 11880 6883 11883
rect 7374 11880 7380 11892
rect 6871 11852 7380 11880
rect 6871 11849 6883 11852
rect 6825 11843 6883 11849
rect 7374 11840 7380 11852
rect 7432 11840 7438 11892
rect 7742 11880 7748 11892
rect 7703 11852 7748 11880
rect 7742 11840 7748 11852
rect 7800 11840 7806 11892
rect 8205 11883 8263 11889
rect 8205 11849 8217 11883
rect 8251 11880 8263 11883
rect 8757 11883 8815 11889
rect 8757 11880 8769 11883
rect 8251 11852 8769 11880
rect 8251 11849 8263 11852
rect 8205 11843 8263 11849
rect 8757 11849 8769 11852
rect 8803 11849 8815 11883
rect 8757 11843 8815 11849
rect 9769 11883 9827 11889
rect 9769 11849 9781 11883
rect 9815 11880 9827 11883
rect 11698 11880 11704 11892
rect 9815 11852 11704 11880
rect 9815 11849 9827 11852
rect 9769 11843 9827 11849
rect 1581 11815 1639 11821
rect 1581 11781 1593 11815
rect 1627 11812 1639 11815
rect 2314 11812 2320 11824
rect 1627 11784 2320 11812
rect 1627 11781 1639 11784
rect 1581 11775 1639 11781
rect 2314 11772 2320 11784
rect 2372 11772 2378 11824
rect 2406 11772 2412 11824
rect 2464 11812 2470 11824
rect 8386 11812 8392 11824
rect 2464 11784 4660 11812
rect 2464 11772 2470 11784
rect 1854 11744 1860 11756
rect 1815 11716 1860 11744
rect 1854 11704 1860 11716
rect 1912 11704 1918 11756
rect 2593 11679 2651 11685
rect 2593 11645 2605 11679
rect 2639 11645 2651 11679
rect 2593 11639 2651 11645
rect 2608 11608 2636 11639
rect 2682 11636 2688 11688
rect 2740 11676 2746 11688
rect 4632 11685 4660 11784
rect 5460 11784 8392 11812
rect 3697 11679 3755 11685
rect 2740 11648 2785 11676
rect 2740 11636 2746 11648
rect 3697 11645 3709 11679
rect 3743 11676 3755 11679
rect 4433 11679 4491 11685
rect 4433 11676 4445 11679
rect 3743 11648 4445 11676
rect 3743 11645 3755 11648
rect 3697 11639 3755 11645
rect 4433 11645 4445 11648
rect 4479 11645 4491 11679
rect 4433 11639 4491 11645
rect 4617 11679 4675 11685
rect 4617 11645 4629 11679
rect 4663 11676 4675 11679
rect 5460 11676 5488 11784
rect 8386 11772 8392 11784
rect 8444 11772 8450 11824
rect 9784 11812 9812 11843
rect 11698 11840 11704 11852
rect 11756 11840 11762 11892
rect 13170 11840 13176 11892
rect 13228 11880 13234 11892
rect 15562 11880 15568 11892
rect 13228 11852 14320 11880
rect 15523 11852 15568 11880
rect 13228 11840 13234 11852
rect 9048 11784 9812 11812
rect 6730 11744 6736 11756
rect 6691 11716 6736 11744
rect 6730 11704 6736 11716
rect 6788 11704 6794 11756
rect 8113 11747 8171 11753
rect 8113 11713 8125 11747
rect 8159 11744 8171 11747
rect 8662 11744 8668 11756
rect 8159 11716 8668 11744
rect 8159 11713 8171 11716
rect 8113 11707 8171 11713
rect 8662 11704 8668 11716
rect 8720 11704 8726 11756
rect 5626 11676 5632 11688
rect 4663 11648 5488 11676
rect 5587 11648 5632 11676
rect 4663 11645 4675 11648
rect 4617 11639 4675 11645
rect 3973 11611 4031 11617
rect 3973 11608 3985 11611
rect 2608 11580 3985 11608
rect 3973 11577 3985 11580
rect 4019 11577 4031 11611
rect 4448 11608 4476 11639
rect 5626 11636 5632 11648
rect 5684 11636 5690 11688
rect 7009 11679 7067 11685
rect 7009 11645 7021 11679
rect 7055 11645 7067 11679
rect 7009 11639 7067 11645
rect 8389 11679 8447 11685
rect 8389 11645 8401 11679
rect 8435 11676 8447 11679
rect 9048 11676 9076 11784
rect 10778 11772 10784 11824
rect 10836 11812 10842 11824
rect 11330 11812 11336 11824
rect 10836 11784 11336 11812
rect 10836 11772 10842 11784
rect 11330 11772 11336 11784
rect 11388 11772 11394 11824
rect 12084 11784 13768 11812
rect 9122 11704 9128 11756
rect 9180 11744 9186 11756
rect 10893 11747 10951 11753
rect 10893 11744 10905 11747
rect 9180 11716 9225 11744
rect 9416 11716 10905 11744
rect 9180 11704 9186 11716
rect 8435 11648 9076 11676
rect 9217 11679 9275 11685
rect 8435 11645 8447 11648
rect 8389 11639 8447 11645
rect 9217 11645 9229 11679
rect 9263 11676 9275 11679
rect 9306 11676 9312 11688
rect 9263 11648 9312 11676
rect 9263 11645 9275 11648
rect 9217 11639 9275 11645
rect 5350 11608 5356 11620
rect 4448 11580 5356 11608
rect 3973 11571 4031 11577
rect 5350 11568 5356 11580
rect 5408 11568 5414 11620
rect 7024 11608 7052 11639
rect 9306 11636 9312 11648
rect 9364 11636 9370 11688
rect 9416 11685 9444 11716
rect 10893 11713 10905 11716
rect 10939 11744 10951 11747
rect 11698 11744 11704 11756
rect 10939 11716 11704 11744
rect 10939 11713 10951 11716
rect 10893 11707 10951 11713
rect 11698 11704 11704 11716
rect 11756 11704 11762 11756
rect 9401 11679 9459 11685
rect 9401 11645 9413 11679
rect 9447 11645 9459 11679
rect 9401 11639 9459 11645
rect 11149 11679 11207 11685
rect 11149 11645 11161 11679
rect 11195 11676 11207 11679
rect 11517 11679 11575 11685
rect 11517 11676 11529 11679
rect 11195 11648 11529 11676
rect 11195 11645 11207 11648
rect 11149 11639 11207 11645
rect 11517 11645 11529 11648
rect 11563 11676 11575 11679
rect 11790 11676 11796 11688
rect 11563 11648 11796 11676
rect 11563 11645 11575 11648
rect 11517 11639 11575 11645
rect 9950 11608 9956 11620
rect 7024 11580 9956 11608
rect 9950 11568 9956 11580
rect 10008 11568 10014 11620
rect 2133 11543 2191 11549
rect 2133 11509 2145 11543
rect 2179 11540 2191 11543
rect 2222 11540 2228 11552
rect 2179 11512 2228 11540
rect 2179 11509 2191 11512
rect 2133 11503 2191 11509
rect 2222 11500 2228 11512
rect 2280 11500 2286 11552
rect 7374 11540 7380 11552
rect 7335 11512 7380 11540
rect 7374 11500 7380 11512
rect 7432 11540 7438 11552
rect 7926 11540 7932 11552
rect 7432 11512 7932 11540
rect 7432 11500 7438 11512
rect 7926 11500 7932 11512
rect 7984 11540 7990 11552
rect 9122 11540 9128 11552
rect 7984 11512 9128 11540
rect 7984 11500 7990 11512
rect 9122 11500 9128 11512
rect 9180 11500 9186 11552
rect 10778 11500 10784 11552
rect 10836 11540 10842 11552
rect 11164 11540 11192 11639
rect 11790 11636 11796 11648
rect 11848 11676 11854 11688
rect 12084 11685 12112 11784
rect 13740 11756 13768 11784
rect 12342 11753 12348 11756
rect 12336 11744 12348 11753
rect 12303 11716 12348 11744
rect 12336 11707 12348 11716
rect 12342 11704 12348 11707
rect 12400 11704 12406 11756
rect 13722 11704 13728 11756
rect 13780 11744 13786 11756
rect 14185 11747 14243 11753
rect 14185 11744 14197 11747
rect 13780 11716 14197 11744
rect 13780 11704 13786 11716
rect 14185 11713 14197 11716
rect 14231 11713 14243 11747
rect 14292 11744 14320 11852
rect 15562 11840 15568 11852
rect 15620 11840 15626 11892
rect 19978 11880 19984 11892
rect 19939 11852 19984 11880
rect 19978 11840 19984 11852
rect 20036 11840 20042 11892
rect 16482 11772 16488 11824
rect 16540 11812 16546 11824
rect 18598 11821 18604 11824
rect 16914 11815 16972 11821
rect 16914 11812 16926 11815
rect 16540 11784 16926 11812
rect 16540 11772 16546 11784
rect 16914 11781 16926 11784
rect 16960 11781 16972 11815
rect 18592 11812 18604 11821
rect 18559 11784 18604 11812
rect 16914 11775 16972 11781
rect 18592 11775 18604 11784
rect 18598 11772 18604 11775
rect 18656 11772 18662 11824
rect 14441 11747 14499 11753
rect 14441 11744 14453 11747
rect 14292 11716 14453 11744
rect 14185 11707 14243 11713
rect 14441 11713 14453 11716
rect 14487 11713 14499 11747
rect 14441 11707 14499 11713
rect 15933 11747 15991 11753
rect 15933 11713 15945 11747
rect 15979 11744 15991 11747
rect 16114 11744 16120 11756
rect 15979 11716 16120 11744
rect 15979 11713 15991 11716
rect 15933 11707 15991 11713
rect 16114 11704 16120 11716
rect 16172 11744 16178 11756
rect 16301 11747 16359 11753
rect 16301 11744 16313 11747
rect 16172 11716 16313 11744
rect 16172 11704 16178 11716
rect 16301 11713 16313 11716
rect 16347 11744 16359 11747
rect 16669 11747 16727 11753
rect 16669 11744 16681 11747
rect 16347 11716 16681 11744
rect 16347 11713 16359 11716
rect 16301 11707 16359 11713
rect 16669 11713 16681 11716
rect 16715 11744 16727 11747
rect 16715 11716 18368 11744
rect 16715 11713 16727 11716
rect 16669 11707 16727 11713
rect 18340 11688 18368 11716
rect 21082 11704 21088 11756
rect 21140 11753 21146 11756
rect 21140 11744 21152 11753
rect 21358 11744 21364 11756
rect 21140 11716 21185 11744
rect 21319 11716 21364 11744
rect 21140 11707 21152 11716
rect 21140 11704 21146 11707
rect 21358 11704 21364 11716
rect 21416 11704 21422 11756
rect 12069 11679 12127 11685
rect 12069 11676 12081 11679
rect 11848 11648 12081 11676
rect 11848 11636 11854 11648
rect 12069 11645 12081 11648
rect 12115 11645 12127 11679
rect 18322 11676 18328 11688
rect 18283 11648 18328 11676
rect 12069 11639 12127 11645
rect 18322 11636 18328 11648
rect 18380 11636 18386 11688
rect 13372 11580 14228 11608
rect 10836 11512 11192 11540
rect 10836 11500 10842 11512
rect 11330 11500 11336 11552
rect 11388 11540 11394 11552
rect 13372 11540 13400 11580
rect 11388 11512 13400 11540
rect 11388 11500 11394 11512
rect 13446 11500 13452 11552
rect 13504 11540 13510 11552
rect 13722 11540 13728 11552
rect 13504 11512 13549 11540
rect 13683 11512 13728 11540
rect 13504 11500 13510 11512
rect 13722 11500 13728 11512
rect 13780 11500 13786 11552
rect 14200 11540 14228 11580
rect 17788 11580 18184 11608
rect 17788 11540 17816 11580
rect 18046 11540 18052 11552
rect 14200 11512 17816 11540
rect 18007 11512 18052 11540
rect 18046 11500 18052 11512
rect 18104 11500 18110 11552
rect 18156 11540 18184 11580
rect 19705 11543 19763 11549
rect 19705 11540 19717 11543
rect 18156 11512 19717 11540
rect 19705 11509 19717 11512
rect 19751 11540 19763 11543
rect 20622 11540 20628 11552
rect 19751 11512 20628 11540
rect 19751 11509 19763 11512
rect 19705 11503 19763 11509
rect 20622 11500 20628 11512
rect 20680 11500 20686 11552
rect 1104 11450 21896 11472
rect 1104 11398 3549 11450
rect 3601 11398 3613 11450
rect 3665 11398 3677 11450
rect 3729 11398 3741 11450
rect 3793 11398 3805 11450
rect 3857 11398 8747 11450
rect 8799 11398 8811 11450
rect 8863 11398 8875 11450
rect 8927 11398 8939 11450
rect 8991 11398 9003 11450
rect 9055 11398 13945 11450
rect 13997 11398 14009 11450
rect 14061 11398 14073 11450
rect 14125 11398 14137 11450
rect 14189 11398 14201 11450
rect 14253 11398 19143 11450
rect 19195 11398 19207 11450
rect 19259 11398 19271 11450
rect 19323 11398 19335 11450
rect 19387 11398 19399 11450
rect 19451 11398 21896 11450
rect 1104 11376 21896 11398
rect 1762 11336 1768 11348
rect 1723 11308 1768 11336
rect 1762 11296 1768 11308
rect 1820 11296 1826 11348
rect 3142 11296 3148 11348
rect 3200 11336 3206 11348
rect 3329 11339 3387 11345
rect 3329 11336 3341 11339
rect 3200 11308 3341 11336
rect 3200 11296 3206 11308
rect 3329 11305 3341 11308
rect 3375 11305 3387 11339
rect 4522 11336 4528 11348
rect 4483 11308 4528 11336
rect 3329 11299 3387 11305
rect 4522 11296 4528 11308
rect 4580 11296 4586 11348
rect 7561 11339 7619 11345
rect 7561 11305 7573 11339
rect 7607 11336 7619 11339
rect 8202 11336 8208 11348
rect 7607 11308 8208 11336
rect 7607 11305 7619 11308
rect 7561 11299 7619 11305
rect 8202 11296 8208 11308
rect 8260 11296 8266 11348
rect 8386 11296 8392 11348
rect 8444 11336 8450 11348
rect 8444 11308 11836 11336
rect 8444 11296 8450 11308
rect 5537 11271 5595 11277
rect 5537 11268 5549 11271
rect 5000 11240 5549 11268
rect 2222 11200 2228 11212
rect 2183 11172 2228 11200
rect 2222 11160 2228 11172
rect 2280 11160 2286 11212
rect 2406 11200 2412 11212
rect 2367 11172 2412 11200
rect 2406 11160 2412 11172
rect 2464 11160 2470 11212
rect 5000 11209 5028 11240
rect 5537 11237 5549 11240
rect 5583 11237 5595 11271
rect 7837 11271 7895 11277
rect 7837 11268 7849 11271
rect 5537 11231 5595 11237
rect 6840 11240 7849 11268
rect 4985 11203 5043 11209
rect 4985 11169 4997 11203
rect 5031 11169 5043 11203
rect 4985 11163 5043 11169
rect 5169 11203 5227 11209
rect 5169 11169 5181 11203
rect 5215 11200 5227 11203
rect 5626 11200 5632 11212
rect 5215 11172 5632 11200
rect 5215 11169 5227 11172
rect 5169 11163 5227 11169
rect 5626 11160 5632 11172
rect 5684 11160 5690 11212
rect 5718 11160 5724 11212
rect 5776 11200 5782 11212
rect 6178 11200 6184 11212
rect 5776 11172 6184 11200
rect 5776 11160 5782 11172
rect 6178 11160 6184 11172
rect 6236 11160 6242 11212
rect 6730 11200 6736 11212
rect 6691 11172 6736 11200
rect 6730 11160 6736 11172
rect 6788 11160 6794 11212
rect 4062 11092 4068 11144
rect 4120 11132 4126 11144
rect 5905 11135 5963 11141
rect 4120 11104 5856 11132
rect 4120 11092 4126 11104
rect 1394 11064 1400 11076
rect 1355 11036 1400 11064
rect 1394 11024 1400 11036
rect 1452 11024 1458 11076
rect 3418 11024 3424 11076
rect 3476 11064 3482 11076
rect 4338 11064 4344 11076
rect 3476 11036 4344 11064
rect 3476 11024 3482 11036
rect 4338 11024 4344 11036
rect 4396 11024 4402 11076
rect 5828 11064 5856 11104
rect 5905 11101 5917 11135
rect 5951 11132 5963 11135
rect 6840 11132 6868 11240
rect 7837 11237 7849 11240
rect 7883 11237 7895 11271
rect 7837 11231 7895 11237
rect 7926 11228 7932 11280
rect 7984 11268 7990 11280
rect 7984 11240 8248 11268
rect 7984 11228 7990 11240
rect 8220 11141 8248 11240
rect 8386 11200 8392 11212
rect 8347 11172 8392 11200
rect 8386 11160 8392 11172
rect 8444 11160 8450 11212
rect 8662 11160 8668 11212
rect 8720 11200 8726 11212
rect 8941 11203 8999 11209
rect 8941 11200 8953 11203
rect 8720 11172 8953 11200
rect 8720 11160 8726 11172
rect 8941 11169 8953 11172
rect 8987 11169 8999 11203
rect 11808 11200 11836 11308
rect 11882 11296 11888 11348
rect 11940 11336 11946 11348
rect 12069 11339 12127 11345
rect 12069 11336 12081 11339
rect 11940 11308 12081 11336
rect 11940 11296 11946 11308
rect 12069 11305 12081 11308
rect 12115 11336 12127 11339
rect 13814 11336 13820 11348
rect 12115 11308 12434 11336
rect 12115 11305 12127 11308
rect 12069 11299 12127 11305
rect 12406 11268 12434 11308
rect 12820 11308 13820 11336
rect 12820 11268 12848 11308
rect 13814 11296 13820 11308
rect 13872 11296 13878 11348
rect 15470 11296 15476 11348
rect 15528 11336 15534 11348
rect 16482 11336 16488 11348
rect 15528 11308 16488 11336
rect 15528 11296 15534 11308
rect 16482 11296 16488 11308
rect 16540 11336 16546 11348
rect 17497 11339 17555 11345
rect 17497 11336 17509 11339
rect 16540 11308 17509 11336
rect 16540 11296 16546 11308
rect 17497 11305 17509 11308
rect 17543 11305 17555 11339
rect 17497 11299 17555 11305
rect 19337 11339 19395 11345
rect 19337 11305 19349 11339
rect 19383 11336 19395 11339
rect 19518 11336 19524 11348
rect 19383 11308 19524 11336
rect 19383 11305 19395 11308
rect 19337 11299 19395 11305
rect 19518 11296 19524 11308
rect 19576 11336 19582 11348
rect 20714 11336 20720 11348
rect 19576 11308 20720 11336
rect 19576 11296 19582 11308
rect 20714 11296 20720 11308
rect 20772 11296 20778 11348
rect 21085 11339 21143 11345
rect 21085 11305 21097 11339
rect 21131 11336 21143 11339
rect 21358 11336 21364 11348
rect 21131 11308 21364 11336
rect 21131 11305 21143 11308
rect 21085 11299 21143 11305
rect 14458 11268 14464 11280
rect 12406 11240 12848 11268
rect 14419 11240 14464 11268
rect 14458 11228 14464 11240
rect 14516 11228 14522 11280
rect 20717 11203 20775 11209
rect 11808 11172 12572 11200
rect 8941 11163 8999 11169
rect 5951 11104 6868 11132
rect 8205 11135 8263 11141
rect 5951 11101 5963 11104
rect 5905 11095 5963 11101
rect 8205 11101 8217 11135
rect 8251 11101 8263 11135
rect 8205 11095 8263 11101
rect 8297 11135 8355 11141
rect 8297 11101 8309 11135
rect 8343 11132 8355 11135
rect 9769 11135 9827 11141
rect 9769 11132 9781 11135
rect 8343 11104 9781 11132
rect 8343 11101 8355 11104
rect 8297 11095 8355 11101
rect 8404 11076 8432 11104
rect 9769 11101 9781 11104
rect 9815 11132 9827 11135
rect 10042 11132 10048 11144
rect 9815 11104 10048 11132
rect 9815 11101 9827 11104
rect 9769 11095 9827 11101
rect 10042 11092 10048 11104
rect 10100 11092 10106 11144
rect 10689 11135 10747 11141
rect 10689 11101 10701 11135
rect 10735 11132 10747 11135
rect 10778 11132 10784 11144
rect 10735 11104 10784 11132
rect 10735 11101 10747 11104
rect 10689 11095 10747 11101
rect 10778 11092 10784 11104
rect 10836 11092 10842 11144
rect 12544 11132 12572 11172
rect 20717 11169 20729 11203
rect 20763 11200 20775 11203
rect 21100 11200 21128 11299
rect 21358 11296 21364 11308
rect 21416 11296 21422 11348
rect 20763 11172 21128 11200
rect 20763 11169 20775 11172
rect 20717 11163 20775 11169
rect 13458 11135 13516 11141
rect 13458 11132 13470 11135
rect 12544 11104 13470 11132
rect 13372 11076 13400 11104
rect 13458 11101 13470 11104
rect 13504 11101 13516 11135
rect 13458 11095 13516 11101
rect 13722 11092 13728 11144
rect 13780 11132 13786 11144
rect 15841 11135 15899 11141
rect 13780 11104 14228 11132
rect 13780 11092 13786 11104
rect 7466 11064 7472 11076
rect 5828 11036 7472 11064
rect 7466 11024 7472 11036
rect 7524 11024 7530 11076
rect 8386 11024 8392 11076
rect 8444 11024 8450 11076
rect 9306 11024 9312 11076
rect 9364 11064 9370 11076
rect 9401 11067 9459 11073
rect 9401 11064 9413 11067
rect 9364 11036 9413 11064
rect 9364 11024 9370 11036
rect 9401 11033 9413 11036
rect 9447 11033 9459 11067
rect 10134 11064 10140 11076
rect 10095 11036 10140 11064
rect 9401 11027 9459 11033
rect 10134 11024 10140 11036
rect 10192 11024 10198 11076
rect 10594 11024 10600 11076
rect 10652 11064 10658 11076
rect 10934 11067 10992 11073
rect 10934 11064 10946 11067
rect 10652 11036 10946 11064
rect 10652 11024 10658 11036
rect 10934 11033 10946 11036
rect 10980 11033 10992 11067
rect 10934 11027 10992 11033
rect 13354 11024 13360 11076
rect 13412 11024 13418 11076
rect 2130 10996 2136 11008
rect 2091 10968 2136 10996
rect 2130 10956 2136 10968
rect 2188 10956 2194 11008
rect 2774 10956 2780 11008
rect 2832 10996 2838 11008
rect 3878 10996 3884 11008
rect 2832 10968 2877 10996
rect 3839 10968 3884 10996
rect 2832 10956 2838 10968
rect 3878 10956 3884 10968
rect 3936 10956 3942 11008
rect 4890 10996 4896 11008
rect 4851 10968 4896 10996
rect 4890 10956 4896 10968
rect 4948 10956 4954 11008
rect 5994 10956 6000 11008
rect 6052 10996 6058 11008
rect 6052 10968 6097 10996
rect 6052 10956 6058 10968
rect 6178 10956 6184 11008
rect 6236 10996 6242 11008
rect 11054 10996 11060 11008
rect 6236 10968 11060 10996
rect 6236 10956 6242 10968
rect 11054 10956 11060 10968
rect 11112 10956 11118 11008
rect 12250 10956 12256 11008
rect 12308 10996 12314 11008
rect 14200 11005 14228 11104
rect 15841 11101 15853 11135
rect 15887 11132 15899 11135
rect 16114 11132 16120 11144
rect 15887 11104 16120 11132
rect 15887 11101 15899 11104
rect 15841 11095 15899 11101
rect 16114 11092 16120 11104
rect 16172 11092 16178 11144
rect 16373 11135 16431 11141
rect 16373 11132 16385 11135
rect 16316 11104 16385 11132
rect 15562 11024 15568 11076
rect 15620 11073 15626 11076
rect 15620 11064 15632 11073
rect 15620 11036 15665 11064
rect 15620 11027 15632 11036
rect 15620 11024 15626 11027
rect 16316 11008 16344 11104
rect 16373 11101 16385 11104
rect 16419 11101 16431 11135
rect 16373 11095 16431 11101
rect 19978 11092 19984 11144
rect 20036 11132 20042 11144
rect 20450 11135 20508 11141
rect 20450 11132 20462 11135
rect 20036 11104 20462 11132
rect 20036 11092 20042 11104
rect 20450 11101 20462 11104
rect 20496 11101 20508 11135
rect 20450 11095 20508 11101
rect 17865 11067 17923 11073
rect 17865 11033 17877 11067
rect 17911 11064 17923 11067
rect 17911 11036 18000 11064
rect 17911 11033 17923 11036
rect 17865 11027 17923 11033
rect 12345 10999 12403 11005
rect 12345 10996 12357 10999
rect 12308 10968 12357 10996
rect 12308 10956 12314 10968
rect 12345 10965 12357 10968
rect 12391 10965 12403 10999
rect 12345 10959 12403 10965
rect 14185 10999 14243 11005
rect 14185 10965 14197 10999
rect 14231 10996 14243 10999
rect 14458 10996 14464 11008
rect 14231 10968 14464 10996
rect 14231 10965 14243 10968
rect 14185 10959 14243 10965
rect 14458 10956 14464 10968
rect 14516 10956 14522 11008
rect 16298 10956 16304 11008
rect 16356 10956 16362 11008
rect 17972 10996 18000 11036
rect 18141 10999 18199 11005
rect 18141 10996 18153 10999
rect 17972 10968 18153 10996
rect 18141 10965 18153 10968
rect 18187 10996 18199 10999
rect 18322 10996 18328 11008
rect 18187 10968 18328 10996
rect 18187 10965 18199 10968
rect 18141 10959 18199 10965
rect 18322 10956 18328 10968
rect 18380 10996 18386 11008
rect 18509 10999 18567 11005
rect 18509 10996 18521 10999
rect 18380 10968 18521 10996
rect 18380 10956 18386 10968
rect 18509 10965 18521 10968
rect 18555 10996 18567 10999
rect 19794 10996 19800 11008
rect 18555 10968 19800 10996
rect 18555 10965 18567 10968
rect 18509 10959 18567 10965
rect 19794 10956 19800 10968
rect 19852 10956 19858 11008
rect 1104 10906 22056 10928
rect 1104 10854 6148 10906
rect 6200 10854 6212 10906
rect 6264 10854 6276 10906
rect 6328 10854 6340 10906
rect 6392 10854 6404 10906
rect 6456 10854 11346 10906
rect 11398 10854 11410 10906
rect 11462 10854 11474 10906
rect 11526 10854 11538 10906
rect 11590 10854 11602 10906
rect 11654 10854 16544 10906
rect 16596 10854 16608 10906
rect 16660 10854 16672 10906
rect 16724 10854 16736 10906
rect 16788 10854 16800 10906
rect 16852 10854 21742 10906
rect 21794 10854 21806 10906
rect 21858 10854 21870 10906
rect 21922 10854 21934 10906
rect 21986 10854 21998 10906
rect 22050 10854 22056 10906
rect 1104 10832 22056 10854
rect 1949 10795 2007 10801
rect 1949 10761 1961 10795
rect 1995 10792 2007 10795
rect 2130 10792 2136 10804
rect 1995 10764 2136 10792
rect 1995 10761 2007 10764
rect 1949 10755 2007 10761
rect 2130 10752 2136 10764
rect 2188 10752 2194 10804
rect 2317 10795 2375 10801
rect 2317 10761 2329 10795
rect 2363 10792 2375 10795
rect 2774 10792 2780 10804
rect 2363 10764 2780 10792
rect 2363 10761 2375 10764
rect 2317 10755 2375 10761
rect 2774 10752 2780 10764
rect 2832 10752 2838 10804
rect 3878 10792 3884 10804
rect 3839 10764 3884 10792
rect 3878 10752 3884 10764
rect 3936 10752 3942 10804
rect 4249 10795 4307 10801
rect 4249 10761 4261 10795
rect 4295 10792 4307 10795
rect 4890 10792 4896 10804
rect 4295 10764 4896 10792
rect 4295 10761 4307 10764
rect 4249 10755 4307 10761
rect 4890 10752 4896 10764
rect 4948 10752 4954 10804
rect 5445 10795 5503 10801
rect 5445 10761 5457 10795
rect 5491 10792 5503 10795
rect 7193 10795 7251 10801
rect 7193 10792 7205 10795
rect 5491 10764 7205 10792
rect 5491 10761 5503 10764
rect 5445 10755 5503 10761
rect 7193 10761 7205 10764
rect 7239 10761 7251 10795
rect 7193 10755 7251 10761
rect 7466 10752 7472 10804
rect 7524 10792 7530 10804
rect 8941 10795 8999 10801
rect 8941 10792 8953 10795
rect 7524 10764 8953 10792
rect 7524 10752 7530 10764
rect 8941 10761 8953 10764
rect 8987 10761 8999 10795
rect 10042 10792 10048 10804
rect 10003 10764 10048 10792
rect 8941 10755 8999 10761
rect 10042 10752 10048 10764
rect 10100 10792 10106 10804
rect 10778 10792 10784 10804
rect 10100 10764 10784 10792
rect 10100 10752 10106 10764
rect 10778 10752 10784 10764
rect 10836 10752 10842 10804
rect 16298 10792 16304 10804
rect 12406 10764 16304 10792
rect 2409 10727 2467 10733
rect 2409 10693 2421 10727
rect 2455 10724 2467 10727
rect 2498 10724 2504 10736
rect 2455 10696 2504 10724
rect 2455 10693 2467 10696
rect 2409 10687 2467 10693
rect 2498 10684 2504 10696
rect 2556 10684 2562 10736
rect 3142 10684 3148 10736
rect 3200 10724 3206 10736
rect 3789 10727 3847 10733
rect 3789 10724 3801 10727
rect 3200 10696 3801 10724
rect 3200 10684 3206 10696
rect 3789 10693 3801 10696
rect 3835 10693 3847 10727
rect 5718 10724 5724 10736
rect 3789 10687 3847 10693
rect 4724 10696 5724 10724
rect 2593 10591 2651 10597
rect 2593 10557 2605 10591
rect 2639 10588 2651 10591
rect 2682 10588 2688 10600
rect 2639 10560 2688 10588
rect 2639 10557 2651 10560
rect 2593 10551 2651 10557
rect 2682 10548 2688 10560
rect 2740 10548 2746 10600
rect 3697 10591 3755 10597
rect 3697 10557 3709 10591
rect 3743 10588 3755 10591
rect 4724 10588 4752 10696
rect 5718 10684 5724 10696
rect 5776 10684 5782 10736
rect 8202 10684 8208 10736
rect 8260 10724 8266 10736
rect 8570 10724 8576 10736
rect 8260 10696 8576 10724
rect 8260 10684 8266 10696
rect 8570 10684 8576 10696
rect 8628 10684 8634 10736
rect 12406 10724 12434 10764
rect 16298 10752 16304 10764
rect 16356 10792 16362 10804
rect 16669 10795 16727 10801
rect 16669 10792 16681 10795
rect 16356 10764 16681 10792
rect 16356 10752 16362 10764
rect 16669 10761 16681 10764
rect 16715 10761 16727 10795
rect 16669 10755 16727 10761
rect 18325 10795 18383 10801
rect 18325 10761 18337 10795
rect 18371 10792 18383 10795
rect 18598 10792 18604 10804
rect 18371 10764 18604 10792
rect 18371 10761 18383 10764
rect 18325 10755 18383 10761
rect 18598 10752 18604 10764
rect 18656 10752 18662 10804
rect 8680 10696 12434 10724
rect 14216 10727 14274 10733
rect 5077 10659 5135 10665
rect 5077 10625 5089 10659
rect 5123 10625 5135 10659
rect 5077 10619 5135 10625
rect 7285 10659 7343 10665
rect 7285 10625 7297 10659
rect 7331 10656 7343 10659
rect 7929 10659 7987 10665
rect 7929 10656 7941 10659
rect 7331 10628 7941 10656
rect 7331 10625 7343 10628
rect 7285 10619 7343 10625
rect 7929 10625 7941 10628
rect 7975 10625 7987 10659
rect 7929 10619 7987 10625
rect 4890 10588 4896 10600
rect 3743 10560 4752 10588
rect 4851 10560 4896 10588
rect 3743 10557 3755 10560
rect 3697 10551 3755 10557
rect 4890 10548 4896 10560
rect 4948 10548 4954 10600
rect 4985 10591 5043 10597
rect 4985 10557 4997 10591
rect 5031 10557 5043 10591
rect 4985 10551 5043 10557
rect 3237 10523 3295 10529
rect 3237 10489 3249 10523
rect 3283 10520 3295 10523
rect 4522 10520 4528 10532
rect 3283 10492 4528 10520
rect 3283 10489 3295 10492
rect 3237 10483 3295 10489
rect 4522 10480 4528 10492
rect 4580 10520 4586 10532
rect 5000 10520 5028 10551
rect 4580 10492 5028 10520
rect 4580 10480 4586 10492
rect 3418 10412 3424 10464
rect 3476 10452 3482 10464
rect 5092 10452 5120 10619
rect 7101 10591 7159 10597
rect 7101 10557 7113 10591
rect 7147 10588 7159 10591
rect 8680 10588 8708 10696
rect 14216 10693 14228 10727
rect 14262 10724 14274 10727
rect 15654 10724 15660 10736
rect 14262 10696 15660 10724
rect 14262 10693 14274 10696
rect 14216 10687 14274 10693
rect 15654 10684 15660 10696
rect 15712 10684 15718 10736
rect 19794 10724 19800 10736
rect 18064 10696 19800 10724
rect 8938 10656 8944 10668
rect 8851 10628 8944 10656
rect 8864 10597 8892 10628
rect 8938 10616 8944 10628
rect 8996 10656 9002 10668
rect 9585 10659 9643 10665
rect 9585 10656 9597 10659
rect 8996 10628 9597 10656
rect 8996 10616 9002 10628
rect 9585 10625 9597 10628
rect 9631 10625 9643 10659
rect 15470 10656 15476 10668
rect 9585 10619 9643 10625
rect 12406 10628 15476 10656
rect 7147 10560 8708 10588
rect 8757 10591 8815 10597
rect 7147 10557 7159 10560
rect 7101 10551 7159 10557
rect 8757 10557 8769 10591
rect 8803 10557 8815 10591
rect 8757 10551 8815 10557
rect 8849 10591 8907 10597
rect 8849 10557 8861 10591
rect 8895 10557 8907 10591
rect 12406 10588 12434 10628
rect 15470 10616 15476 10628
rect 15528 10616 15534 10668
rect 15562 10616 15568 10668
rect 15620 10656 15626 10668
rect 15850 10659 15908 10665
rect 15850 10656 15862 10659
rect 15620 10628 15862 10656
rect 15620 10616 15626 10628
rect 15850 10625 15862 10628
rect 15896 10625 15908 10659
rect 15850 10619 15908 10625
rect 16942 10616 16948 10668
rect 17000 10656 17006 10668
rect 18064 10665 18092 10696
rect 17782 10659 17840 10665
rect 17782 10656 17794 10659
rect 17000 10628 17794 10656
rect 17000 10616 17006 10628
rect 17782 10625 17794 10628
rect 17828 10625 17840 10659
rect 17782 10619 17840 10625
rect 18049 10659 18107 10665
rect 18049 10625 18061 10659
rect 18095 10625 18107 10659
rect 19426 10656 19432 10668
rect 19484 10665 19490 10668
rect 19720 10665 19748 10696
rect 19794 10684 19800 10696
rect 19852 10724 19858 10736
rect 19852 10696 21404 10724
rect 19852 10684 19858 10696
rect 21376 10668 21404 10696
rect 19396 10628 19432 10656
rect 18049 10619 18107 10625
rect 19426 10616 19432 10628
rect 19484 10619 19496 10665
rect 19705 10659 19763 10665
rect 19705 10625 19717 10659
rect 19751 10625 19763 10659
rect 19705 10619 19763 10625
rect 19484 10616 19490 10619
rect 20622 10616 20628 10668
rect 20680 10656 20686 10668
rect 21094 10659 21152 10665
rect 21094 10656 21106 10659
rect 20680 10628 21106 10656
rect 20680 10616 20686 10628
rect 21094 10625 21106 10628
rect 21140 10625 21152 10659
rect 21358 10656 21364 10668
rect 21319 10628 21364 10656
rect 21094 10619 21152 10625
rect 21358 10616 21364 10628
rect 21416 10616 21422 10668
rect 14458 10588 14464 10600
rect 8849 10551 8907 10557
rect 8956 10560 12434 10588
rect 14419 10560 14464 10588
rect 5534 10480 5540 10532
rect 5592 10520 5598 10532
rect 8386 10520 8392 10532
rect 5592 10492 8392 10520
rect 5592 10480 5598 10492
rect 8386 10480 8392 10492
rect 8444 10480 8450 10532
rect 8772 10520 8800 10551
rect 8956 10520 8984 10560
rect 14458 10548 14464 10560
rect 14516 10548 14522 10600
rect 16114 10588 16120 10600
rect 16075 10560 16120 10588
rect 16114 10548 16120 10560
rect 16172 10548 16178 10600
rect 8772 10492 8984 10520
rect 9309 10523 9367 10529
rect 9309 10489 9321 10523
rect 9355 10520 9367 10523
rect 9858 10520 9864 10532
rect 9355 10492 9864 10520
rect 9355 10489 9367 10492
rect 9309 10483 9367 10489
rect 9858 10480 9864 10492
rect 9916 10480 9922 10532
rect 9950 10480 9956 10532
rect 10008 10520 10014 10532
rect 12618 10520 12624 10532
rect 10008 10492 12624 10520
rect 10008 10480 10014 10492
rect 12618 10480 12624 10492
rect 12676 10520 12682 10532
rect 19978 10520 19984 10532
rect 12676 10492 13308 10520
rect 19939 10492 19984 10520
rect 12676 10480 12682 10492
rect 5718 10452 5724 10464
rect 3476 10424 5120 10452
rect 5679 10424 5724 10452
rect 3476 10412 3482 10424
rect 5718 10412 5724 10424
rect 5776 10412 5782 10464
rect 5810 10412 5816 10464
rect 5868 10452 5874 10464
rect 6549 10455 6607 10461
rect 6549 10452 6561 10455
rect 5868 10424 6561 10452
rect 5868 10412 5874 10424
rect 6549 10421 6561 10424
rect 6595 10452 6607 10455
rect 7374 10452 7380 10464
rect 6595 10424 7380 10452
rect 6595 10421 6607 10424
rect 6549 10415 6607 10421
rect 7374 10412 7380 10424
rect 7432 10412 7438 10464
rect 7653 10455 7711 10461
rect 7653 10421 7665 10455
rect 7699 10452 7711 10455
rect 7926 10452 7932 10464
rect 7699 10424 7932 10452
rect 7699 10421 7711 10424
rect 7653 10415 7711 10421
rect 7926 10412 7932 10424
rect 7984 10412 7990 10464
rect 12253 10455 12311 10461
rect 12253 10421 12265 10455
rect 12299 10452 12311 10455
rect 12434 10452 12440 10464
rect 12299 10424 12440 10452
rect 12299 10421 12311 10424
rect 12253 10415 12311 10421
rect 12434 10412 12440 10424
rect 12492 10412 12498 10464
rect 13078 10452 13084 10464
rect 13039 10424 13084 10452
rect 13078 10412 13084 10424
rect 13136 10412 13142 10464
rect 13280 10452 13308 10492
rect 19978 10480 19984 10492
rect 20036 10480 20042 10532
rect 14737 10455 14795 10461
rect 14737 10452 14749 10455
rect 13280 10424 14749 10452
rect 14737 10421 14749 10424
rect 14783 10421 14795 10455
rect 14737 10415 14795 10421
rect 1104 10362 21896 10384
rect 1104 10310 3549 10362
rect 3601 10310 3613 10362
rect 3665 10310 3677 10362
rect 3729 10310 3741 10362
rect 3793 10310 3805 10362
rect 3857 10310 8747 10362
rect 8799 10310 8811 10362
rect 8863 10310 8875 10362
rect 8927 10310 8939 10362
rect 8991 10310 9003 10362
rect 9055 10310 13945 10362
rect 13997 10310 14009 10362
rect 14061 10310 14073 10362
rect 14125 10310 14137 10362
rect 14189 10310 14201 10362
rect 14253 10310 19143 10362
rect 19195 10310 19207 10362
rect 19259 10310 19271 10362
rect 19323 10310 19335 10362
rect 19387 10310 19399 10362
rect 19451 10310 21896 10362
rect 1104 10288 21896 10310
rect 2685 10251 2743 10257
rect 2685 10217 2697 10251
rect 2731 10248 2743 10251
rect 2866 10248 2872 10260
rect 2731 10220 2872 10248
rect 2731 10217 2743 10220
rect 2685 10211 2743 10217
rect 2866 10208 2872 10220
rect 2924 10208 2930 10260
rect 3418 10248 3424 10260
rect 3379 10220 3424 10248
rect 3418 10208 3424 10220
rect 3476 10208 3482 10260
rect 5810 10248 5816 10260
rect 4816 10220 5816 10248
rect 3694 10072 3700 10124
rect 3752 10112 3758 10124
rect 4816 10112 4844 10220
rect 5810 10208 5816 10220
rect 5868 10208 5874 10260
rect 5994 10208 6000 10260
rect 6052 10248 6058 10260
rect 6181 10251 6239 10257
rect 6181 10248 6193 10251
rect 6052 10220 6193 10248
rect 6052 10208 6058 10220
rect 6181 10217 6193 10220
rect 6227 10217 6239 10251
rect 7466 10248 7472 10260
rect 7427 10220 7472 10248
rect 6181 10211 6239 10217
rect 7466 10208 7472 10220
rect 7524 10208 7530 10260
rect 8294 10208 8300 10260
rect 8352 10248 8358 10260
rect 8941 10251 8999 10257
rect 8941 10248 8953 10251
rect 8352 10220 8953 10248
rect 8352 10208 8358 10220
rect 8941 10217 8953 10220
rect 8987 10217 8999 10251
rect 12434 10248 12440 10260
rect 8941 10211 8999 10217
rect 10796 10220 12440 10248
rect 7742 10180 7748 10192
rect 5552 10152 7748 10180
rect 3752 10084 4844 10112
rect 3752 10072 3758 10084
rect 2866 10004 2872 10056
rect 2924 10044 2930 10056
rect 4816 10053 4844 10084
rect 5077 10115 5135 10121
rect 5077 10081 5089 10115
rect 5123 10112 5135 10115
rect 5258 10112 5264 10124
rect 5123 10084 5264 10112
rect 5123 10081 5135 10084
rect 5077 10075 5135 10081
rect 5258 10072 5264 10084
rect 5316 10072 5322 10124
rect 5552 10121 5580 10152
rect 7742 10140 7748 10152
rect 7800 10140 7806 10192
rect 8018 10140 8024 10192
rect 8076 10180 8082 10192
rect 8076 10152 8432 10180
rect 8076 10140 8082 10152
rect 5537 10115 5595 10121
rect 5537 10081 5549 10115
rect 5583 10081 5595 10115
rect 5537 10075 5595 10081
rect 5626 10072 5632 10124
rect 5684 10112 5690 10124
rect 8404 10121 8432 10152
rect 8389 10115 8447 10121
rect 5684 10084 8340 10112
rect 5684 10072 5690 10084
rect 3789 10047 3847 10053
rect 3789 10044 3801 10047
rect 2924 10016 3801 10044
rect 2924 10004 2930 10016
rect 3789 10013 3801 10016
rect 3835 10013 3847 10047
rect 3789 10007 3847 10013
rect 4801 10047 4859 10053
rect 4801 10013 4813 10047
rect 4847 10013 4859 10047
rect 4801 10007 4859 10013
rect 5721 10047 5779 10053
rect 5721 10013 5733 10047
rect 5767 10044 5779 10047
rect 5810 10044 5816 10056
rect 5767 10016 5816 10044
rect 5767 10013 5779 10016
rect 5721 10007 5779 10013
rect 5810 10004 5816 10016
rect 5868 10004 5874 10056
rect 7834 10044 7840 10056
rect 6748 10016 7840 10044
rect 3050 9936 3056 9988
rect 3108 9976 3114 9988
rect 6748 9985 6776 10016
rect 7834 10004 7840 10016
rect 7892 10044 7898 10056
rect 8205 10047 8263 10053
rect 8205 10044 8217 10047
rect 7892 10016 8217 10044
rect 7892 10004 7898 10016
rect 8205 10013 8217 10016
rect 8251 10013 8263 10047
rect 8312 10044 8340 10084
rect 8389 10081 8401 10115
rect 8435 10081 8447 10115
rect 9490 10112 9496 10124
rect 9451 10084 9496 10112
rect 8389 10075 8447 10081
rect 9490 10072 9496 10084
rect 9548 10072 9554 10124
rect 9674 10072 9680 10124
rect 9732 10112 9738 10124
rect 10796 10121 10824 10220
rect 12434 10208 12440 10220
rect 12492 10248 12498 10260
rect 13262 10248 13268 10260
rect 12492 10220 13268 10248
rect 12492 10208 12498 10220
rect 13262 10208 13268 10220
rect 13320 10208 13326 10260
rect 14458 10208 14464 10260
rect 14516 10248 14522 10260
rect 14645 10251 14703 10257
rect 14645 10248 14657 10251
rect 14516 10220 14657 10248
rect 14516 10208 14522 10220
rect 14645 10217 14657 10220
rect 14691 10248 14703 10251
rect 16114 10248 16120 10260
rect 14691 10220 16120 10248
rect 14691 10217 14703 10220
rect 14645 10211 14703 10217
rect 16114 10208 16120 10220
rect 16172 10248 16178 10260
rect 16209 10251 16267 10257
rect 16209 10248 16221 10251
rect 16172 10220 16221 10248
rect 16172 10208 16178 10220
rect 16209 10217 16221 10220
rect 16255 10217 16267 10251
rect 16209 10211 16267 10217
rect 17126 10208 17132 10260
rect 17184 10248 17190 10260
rect 17313 10251 17371 10257
rect 17313 10248 17325 10251
rect 17184 10220 17325 10248
rect 17184 10208 17190 10220
rect 17313 10217 17325 10220
rect 17359 10217 17371 10251
rect 17313 10211 17371 10217
rect 20993 10251 21051 10257
rect 20993 10217 21005 10251
rect 21039 10248 21051 10251
rect 21358 10248 21364 10260
rect 21039 10220 21364 10248
rect 21039 10217 21051 10220
rect 20993 10211 21051 10217
rect 21358 10208 21364 10220
rect 21416 10208 21422 10260
rect 10321 10115 10379 10121
rect 10321 10112 10333 10115
rect 9732 10084 10333 10112
rect 9732 10072 9738 10084
rect 10321 10081 10333 10084
rect 10367 10081 10379 10115
rect 10321 10075 10379 10081
rect 10781 10115 10839 10121
rect 10781 10081 10793 10115
rect 10827 10081 10839 10115
rect 10781 10075 10839 10081
rect 8312 10016 9904 10044
rect 8205 10007 8263 10013
rect 6733 9979 6791 9985
rect 6733 9976 6745 9979
rect 3108 9948 6745 9976
rect 3108 9936 3114 9948
rect 6733 9945 6745 9948
rect 6779 9945 6791 9979
rect 8297 9979 8355 9985
rect 8297 9976 8309 9979
rect 6733 9939 6791 9945
rect 7116 9948 8309 9976
rect 2961 9911 3019 9917
rect 2961 9877 2973 9911
rect 3007 9908 3019 9911
rect 3602 9908 3608 9920
rect 3007 9880 3608 9908
rect 3007 9877 3019 9880
rect 2961 9871 3019 9877
rect 3602 9868 3608 9880
rect 3660 9868 3666 9920
rect 3973 9911 4031 9917
rect 3973 9877 3985 9911
rect 4019 9908 4031 9911
rect 4062 9908 4068 9920
rect 4019 9880 4068 9908
rect 4019 9877 4031 9880
rect 3973 9871 4031 9877
rect 4062 9868 4068 9880
rect 4120 9868 4126 9920
rect 4430 9908 4436 9920
rect 4391 9880 4436 9908
rect 4430 9868 4436 9880
rect 4488 9868 4494 9920
rect 4614 9868 4620 9920
rect 4672 9908 4678 9920
rect 4893 9911 4951 9917
rect 4893 9908 4905 9911
rect 4672 9880 4905 9908
rect 4672 9868 4678 9880
rect 4893 9877 4905 9880
rect 4939 9908 4951 9911
rect 5534 9908 5540 9920
rect 4939 9880 5540 9908
rect 4939 9877 4951 9880
rect 4893 9871 4951 9877
rect 5534 9868 5540 9880
rect 5592 9868 5598 9920
rect 5718 9868 5724 9920
rect 5776 9908 5782 9920
rect 5813 9911 5871 9917
rect 5813 9908 5825 9911
rect 5776 9880 5825 9908
rect 5776 9868 5782 9880
rect 5813 9877 5825 9880
rect 5859 9877 5871 9911
rect 5813 9871 5871 9877
rect 6822 9868 6828 9920
rect 6880 9908 6886 9920
rect 7116 9917 7144 9948
rect 8297 9945 8309 9948
rect 8343 9945 8355 9979
rect 9876 9976 9904 10016
rect 10870 10004 10876 10056
rect 10928 10044 10934 10056
rect 18693 10047 18751 10053
rect 10928 10016 18552 10044
rect 10928 10004 10934 10016
rect 11054 9985 11060 9988
rect 11048 9976 11060 9985
rect 9876 9948 10456 9976
rect 10967 9948 11060 9976
rect 8297 9939 8355 9945
rect 7101 9911 7159 9917
rect 7101 9908 7113 9911
rect 6880 9880 7113 9908
rect 6880 9868 6886 9880
rect 7101 9877 7113 9880
rect 7147 9877 7159 9911
rect 7834 9908 7840 9920
rect 7795 9880 7840 9908
rect 7101 9871 7159 9877
rect 7834 9868 7840 9880
rect 7892 9868 7898 9920
rect 9122 9868 9128 9920
rect 9180 9908 9186 9920
rect 9309 9911 9367 9917
rect 9309 9908 9321 9911
rect 9180 9880 9321 9908
rect 9180 9868 9186 9880
rect 9309 9877 9321 9880
rect 9355 9877 9367 9911
rect 9309 9871 9367 9877
rect 9398 9868 9404 9920
rect 9456 9908 9462 9920
rect 9953 9911 10011 9917
rect 9953 9908 9965 9911
rect 9456 9880 9965 9908
rect 9456 9868 9462 9880
rect 9953 9877 9965 9880
rect 9999 9877 10011 9911
rect 10428 9908 10456 9948
rect 11048 9939 11060 9948
rect 11112 9976 11118 9988
rect 11882 9976 11888 9988
rect 11112 9948 11888 9976
rect 11054 9936 11060 9939
rect 11112 9936 11118 9948
rect 11882 9936 11888 9948
rect 11940 9936 11946 9988
rect 12710 9936 12716 9988
rect 12768 9976 12774 9988
rect 18414 9976 18420 9988
rect 18472 9985 18478 9988
rect 12768 9948 18420 9976
rect 12768 9936 12774 9948
rect 18414 9936 18420 9948
rect 18472 9939 18484 9985
rect 18524 9976 18552 10016
rect 18693 10013 18705 10047
rect 18739 10044 18751 10047
rect 19245 10047 19303 10053
rect 19245 10044 19257 10047
rect 18739 10016 19257 10044
rect 18739 10013 18751 10016
rect 18693 10007 18751 10013
rect 19245 10013 19257 10016
rect 19291 10044 19303 10047
rect 19334 10044 19340 10056
rect 19291 10016 19340 10044
rect 19291 10013 19303 10016
rect 19245 10007 19303 10013
rect 19334 10004 19340 10016
rect 19392 10044 19398 10056
rect 19794 10044 19800 10056
rect 19392 10016 19800 10044
rect 19392 10004 19398 10016
rect 19794 10004 19800 10016
rect 19852 10004 19858 10056
rect 19426 9976 19432 9988
rect 18524 9948 19432 9976
rect 18472 9936 18478 9939
rect 19426 9936 19432 9948
rect 19484 9985 19490 9988
rect 19484 9979 19548 9985
rect 19484 9945 19502 9979
rect 19536 9945 19548 9979
rect 19484 9939 19548 9945
rect 19484 9936 19490 9939
rect 12161 9911 12219 9917
rect 12161 9908 12173 9911
rect 10428 9880 12173 9908
rect 9953 9871 10011 9877
rect 12161 9877 12173 9880
rect 12207 9908 12219 9911
rect 12250 9908 12256 9920
rect 12207 9880 12256 9908
rect 12207 9877 12219 9880
rect 12161 9871 12219 9877
rect 12250 9868 12256 9880
rect 12308 9868 12314 9920
rect 20622 9908 20628 9920
rect 20583 9880 20628 9908
rect 20622 9868 20628 9880
rect 20680 9908 20686 9920
rect 21082 9908 21088 9920
rect 20680 9880 21088 9908
rect 20680 9868 20686 9880
rect 21082 9868 21088 9880
rect 21140 9868 21146 9920
rect 1104 9818 22056 9840
rect 1104 9766 6148 9818
rect 6200 9766 6212 9818
rect 6264 9766 6276 9818
rect 6328 9766 6340 9818
rect 6392 9766 6404 9818
rect 6456 9766 11346 9818
rect 11398 9766 11410 9818
rect 11462 9766 11474 9818
rect 11526 9766 11538 9818
rect 11590 9766 11602 9818
rect 11654 9766 16544 9818
rect 16596 9766 16608 9818
rect 16660 9766 16672 9818
rect 16724 9766 16736 9818
rect 16788 9766 16800 9818
rect 16852 9766 21742 9818
rect 21794 9766 21806 9818
rect 21858 9766 21870 9818
rect 21922 9766 21934 9818
rect 21986 9766 21998 9818
rect 22050 9766 22056 9818
rect 1104 9744 22056 9766
rect 3234 9664 3240 9716
rect 3292 9704 3298 9716
rect 3418 9704 3424 9716
rect 3292 9676 3424 9704
rect 3292 9664 3298 9676
rect 3418 9664 3424 9676
rect 3476 9664 3482 9716
rect 3602 9664 3608 9716
rect 3660 9704 3666 9716
rect 4614 9704 4620 9716
rect 3660 9676 4620 9704
rect 3660 9664 3666 9676
rect 4614 9664 4620 9676
rect 4672 9664 4678 9716
rect 6365 9707 6423 9713
rect 6365 9673 6377 9707
rect 6411 9673 6423 9707
rect 6365 9667 6423 9673
rect 3970 9596 3976 9648
rect 4028 9636 4034 9648
rect 6380 9636 6408 9667
rect 9674 9664 9680 9716
rect 9732 9704 9738 9716
rect 10873 9707 10931 9713
rect 10873 9704 10885 9707
rect 9732 9676 10885 9704
rect 9732 9664 9738 9676
rect 10873 9673 10885 9676
rect 10919 9673 10931 9707
rect 10873 9667 10931 9673
rect 11517 9707 11575 9713
rect 11517 9673 11529 9707
rect 11563 9704 11575 9707
rect 11698 9704 11704 9716
rect 11563 9676 11704 9704
rect 11563 9673 11575 9676
rect 11517 9667 11575 9673
rect 11698 9664 11704 9676
rect 11756 9664 11762 9716
rect 19337 9707 19395 9713
rect 19337 9673 19349 9707
rect 19383 9704 19395 9707
rect 19426 9704 19432 9716
rect 19383 9676 19432 9704
rect 19383 9673 19395 9676
rect 19337 9667 19395 9673
rect 19426 9664 19432 9676
rect 19484 9664 19490 9716
rect 21358 9704 21364 9716
rect 21319 9676 21364 9704
rect 21358 9664 21364 9676
rect 21416 9664 21422 9716
rect 4028 9608 6408 9636
rect 6825 9639 6883 9645
rect 4028 9596 4034 9608
rect 6825 9605 6837 9639
rect 6871 9636 6883 9639
rect 7834 9636 7840 9648
rect 6871 9608 7840 9636
rect 6871 9605 6883 9608
rect 6825 9599 6883 9605
rect 7834 9596 7840 9608
rect 7892 9596 7898 9648
rect 9858 9636 9864 9648
rect 9819 9608 9864 9636
rect 9858 9596 9864 9608
rect 9916 9596 9922 9648
rect 12526 9636 12532 9648
rect 9968 9608 12532 9636
rect 3234 9528 3240 9580
rect 3292 9568 3298 9580
rect 3881 9571 3939 9577
rect 3881 9568 3893 9571
rect 3292 9540 3893 9568
rect 3292 9528 3298 9540
rect 3881 9537 3893 9540
rect 3927 9537 3939 9571
rect 3881 9531 3939 9537
rect 4246 9528 4252 9580
rect 4304 9568 4310 9580
rect 4985 9571 5043 9577
rect 4985 9568 4997 9571
rect 4304 9540 4997 9568
rect 4304 9528 4310 9540
rect 4985 9537 4997 9540
rect 5031 9568 5043 9571
rect 5718 9568 5724 9580
rect 5031 9540 5724 9568
rect 5031 9537 5043 9540
rect 4985 9531 5043 9537
rect 5718 9528 5724 9540
rect 5776 9528 5782 9580
rect 6730 9568 6736 9580
rect 6691 9540 6736 9568
rect 6730 9528 6736 9540
rect 6788 9528 6794 9580
rect 7745 9571 7803 9577
rect 7745 9537 7757 9571
rect 7791 9568 7803 9571
rect 8389 9571 8447 9577
rect 8389 9568 8401 9571
rect 7791 9540 8401 9568
rect 7791 9537 7803 9540
rect 7745 9531 7803 9537
rect 8389 9537 8401 9540
rect 8435 9537 8447 9571
rect 8389 9531 8447 9537
rect 9125 9571 9183 9577
rect 9125 9537 9137 9571
rect 9171 9568 9183 9571
rect 9769 9571 9827 9577
rect 9769 9568 9781 9571
rect 9171 9540 9781 9568
rect 9171 9537 9183 9540
rect 9125 9531 9183 9537
rect 9769 9537 9781 9540
rect 9815 9537 9827 9571
rect 9769 9531 9827 9537
rect 2222 9460 2228 9512
rect 2280 9500 2286 9512
rect 3602 9500 3608 9512
rect 2280 9472 3608 9500
rect 2280 9460 2286 9472
rect 3602 9460 3608 9472
rect 3660 9460 3666 9512
rect 3970 9500 3976 9512
rect 3931 9472 3976 9500
rect 3970 9460 3976 9472
rect 4028 9460 4034 9512
rect 4062 9460 4068 9512
rect 4120 9500 4126 9512
rect 5074 9500 5080 9512
rect 4120 9472 4165 9500
rect 5035 9472 5080 9500
rect 4120 9460 4126 9472
rect 5074 9460 5080 9472
rect 5132 9460 5138 9512
rect 5258 9500 5264 9512
rect 5219 9472 5264 9500
rect 5258 9460 5264 9472
rect 5316 9460 5322 9512
rect 6546 9460 6552 9512
rect 6604 9500 6610 9512
rect 6917 9503 6975 9509
rect 6917 9500 6929 9503
rect 6604 9472 6929 9500
rect 6604 9460 6610 9472
rect 6917 9469 6929 9472
rect 6963 9469 6975 9503
rect 6917 9463 6975 9469
rect 7837 9503 7895 9509
rect 7837 9469 7849 9503
rect 7883 9469 7895 9503
rect 7837 9463 7895 9469
rect 8021 9503 8079 9509
rect 8021 9469 8033 9503
rect 8067 9500 8079 9503
rect 9968 9500 9996 9608
rect 12526 9596 12532 9608
rect 12584 9596 12590 9648
rect 12618 9596 12624 9648
rect 12676 9645 12682 9648
rect 12676 9636 12688 9645
rect 13262 9636 13268 9648
rect 12676 9608 12721 9636
rect 13004 9608 13268 9636
rect 12676 9599 12688 9608
rect 12676 9596 12682 9599
rect 10778 9568 10784 9580
rect 10739 9540 10784 9568
rect 10778 9528 10784 9540
rect 10836 9528 10842 9580
rect 10962 9528 10968 9580
rect 11020 9568 11026 9580
rect 11698 9568 11704 9580
rect 11020 9540 11704 9568
rect 11020 9528 11026 9540
rect 11698 9528 11704 9540
rect 11756 9528 11762 9580
rect 8067 9472 9996 9500
rect 10045 9503 10103 9509
rect 8067 9469 8079 9472
rect 8021 9463 8079 9469
rect 10045 9469 10057 9503
rect 10091 9469 10103 9503
rect 11054 9500 11060 9512
rect 11015 9472 11060 9500
rect 10045 9463 10103 9469
rect 1854 9392 1860 9444
rect 1912 9432 1918 9444
rect 3513 9435 3571 9441
rect 3513 9432 3525 9435
rect 1912 9404 3525 9432
rect 1912 9392 1918 9404
rect 3513 9401 3525 9404
rect 3559 9401 3571 9435
rect 3513 9395 3571 9401
rect 3786 9392 3792 9444
rect 3844 9432 3850 9444
rect 3844 9404 7052 9432
rect 3844 9392 3850 9404
rect 2866 9324 2872 9376
rect 2924 9364 2930 9376
rect 3145 9367 3203 9373
rect 3145 9364 3157 9367
rect 2924 9336 3157 9364
rect 2924 9324 2930 9336
rect 3145 9333 3157 9336
rect 3191 9364 3203 9367
rect 3694 9364 3700 9376
rect 3191 9336 3700 9364
rect 3191 9333 3203 9336
rect 3145 9327 3203 9333
rect 3694 9324 3700 9336
rect 3752 9324 3758 9376
rect 4617 9367 4675 9373
rect 4617 9333 4629 9367
rect 4663 9364 4675 9367
rect 4706 9364 4712 9376
rect 4663 9336 4712 9364
rect 4663 9333 4675 9336
rect 4617 9327 4675 9333
rect 4706 9324 4712 9336
rect 4764 9324 4770 9376
rect 5810 9324 5816 9376
rect 5868 9364 5874 9376
rect 5905 9367 5963 9373
rect 5905 9364 5917 9367
rect 5868 9336 5917 9364
rect 5868 9324 5874 9336
rect 5905 9333 5917 9336
rect 5951 9333 5963 9367
rect 7024 9364 7052 9404
rect 7190 9392 7196 9444
rect 7248 9432 7254 9444
rect 7377 9435 7435 9441
rect 7377 9432 7389 9435
rect 7248 9404 7389 9432
rect 7248 9392 7254 9404
rect 7377 9401 7389 9404
rect 7423 9401 7435 9435
rect 7852 9432 7880 9463
rect 10060 9432 10088 9463
rect 11054 9460 11060 9472
rect 11112 9460 11118 9512
rect 12897 9503 12955 9509
rect 12897 9469 12909 9503
rect 12943 9500 12955 9503
rect 13004 9500 13032 9608
rect 13262 9596 13268 9608
rect 13320 9596 13326 9648
rect 18046 9596 18052 9648
rect 18104 9596 18110 9648
rect 19978 9596 19984 9648
rect 20036 9636 20042 9648
rect 20450 9639 20508 9645
rect 20450 9636 20462 9639
rect 20036 9608 20462 9636
rect 20036 9596 20042 9608
rect 20450 9605 20462 9608
rect 20496 9605 20508 9639
rect 20450 9599 20508 9605
rect 18064 9568 18092 9596
rect 18150 9571 18208 9577
rect 18150 9568 18162 9571
rect 12943 9472 13032 9500
rect 13096 9540 18162 9568
rect 12943 9469 12955 9472
rect 12897 9463 12955 9469
rect 7852 9404 9904 9432
rect 10060 9404 11652 9432
rect 7377 9395 7435 9401
rect 8386 9364 8392 9376
rect 7024 9336 8392 9364
rect 5905 9327 5963 9333
rect 8386 9324 8392 9336
rect 8444 9324 8450 9376
rect 9214 9324 9220 9376
rect 9272 9364 9278 9376
rect 9401 9367 9459 9373
rect 9401 9364 9413 9367
rect 9272 9336 9413 9364
rect 9272 9324 9278 9336
rect 9401 9333 9413 9336
rect 9447 9333 9459 9367
rect 9876 9364 9904 9404
rect 10413 9367 10471 9373
rect 10413 9364 10425 9367
rect 9876 9336 10425 9364
rect 9401 9327 9459 9333
rect 10413 9333 10425 9336
rect 10459 9333 10471 9367
rect 11624 9364 11652 9404
rect 13096 9364 13124 9540
rect 18150 9537 18162 9540
rect 18196 9537 18208 9571
rect 18150 9531 18208 9537
rect 18417 9571 18475 9577
rect 18417 9537 18429 9571
rect 18463 9568 18475 9571
rect 18785 9571 18843 9577
rect 18785 9568 18797 9571
rect 18463 9540 18797 9568
rect 18463 9537 18475 9540
rect 18417 9531 18475 9537
rect 18785 9537 18797 9540
rect 18831 9568 18843 9571
rect 19334 9568 19340 9580
rect 18831 9540 19340 9568
rect 18831 9537 18843 9540
rect 18785 9531 18843 9537
rect 19334 9528 19340 9540
rect 19392 9528 19398 9580
rect 20717 9571 20775 9577
rect 20717 9537 20729 9571
rect 20763 9568 20775 9571
rect 21376 9568 21404 9664
rect 20763 9540 21404 9568
rect 20763 9537 20775 9540
rect 20717 9531 20775 9537
rect 17034 9432 17040 9444
rect 16995 9404 17040 9432
rect 17034 9392 17040 9404
rect 17092 9392 17098 9444
rect 13262 9364 13268 9376
rect 11624 9336 13124 9364
rect 13223 9336 13268 9364
rect 10413 9327 10471 9333
rect 13262 9324 13268 9336
rect 13320 9324 13326 9376
rect 1104 9274 21896 9296
rect 1104 9222 3549 9274
rect 3601 9222 3613 9274
rect 3665 9222 3677 9274
rect 3729 9222 3741 9274
rect 3793 9222 3805 9274
rect 3857 9222 8747 9274
rect 8799 9222 8811 9274
rect 8863 9222 8875 9274
rect 8927 9222 8939 9274
rect 8991 9222 9003 9274
rect 9055 9222 13945 9274
rect 13997 9222 14009 9274
rect 14061 9222 14073 9274
rect 14125 9222 14137 9274
rect 14189 9222 14201 9274
rect 14253 9222 19143 9274
rect 19195 9222 19207 9274
rect 19259 9222 19271 9274
rect 19323 9222 19335 9274
rect 19387 9222 19399 9274
rect 19451 9222 21896 9274
rect 1104 9200 21896 9222
rect 3234 9160 3240 9172
rect 3195 9132 3240 9160
rect 3234 9120 3240 9132
rect 3292 9120 3298 9172
rect 3970 9120 3976 9172
rect 4028 9160 4034 9172
rect 4249 9163 4307 9169
rect 4249 9160 4261 9163
rect 4028 9132 4261 9160
rect 4028 9120 4034 9132
rect 4249 9129 4261 9132
rect 4295 9129 4307 9163
rect 4249 9123 4307 9129
rect 4890 9120 4896 9172
rect 4948 9160 4954 9172
rect 15933 9163 15991 9169
rect 15933 9160 15945 9163
rect 4948 9132 15945 9160
rect 4948 9120 4954 9132
rect 15933 9129 15945 9132
rect 15979 9160 15991 9163
rect 16942 9160 16948 9172
rect 15979 9132 16948 9160
rect 15979 9129 15991 9132
rect 15933 9123 15991 9129
rect 16942 9120 16948 9132
rect 17000 9120 17006 9172
rect 18414 9120 18420 9172
rect 18472 9160 18478 9172
rect 19705 9163 19763 9169
rect 19705 9160 19717 9163
rect 18472 9132 19717 9160
rect 18472 9120 18478 9132
rect 19705 9129 19717 9132
rect 19751 9129 19763 9163
rect 19705 9123 19763 9129
rect 2225 9095 2283 9101
rect 2225 9061 2237 9095
rect 2271 9092 2283 9095
rect 2774 9092 2780 9104
rect 2271 9064 2780 9092
rect 2271 9061 2283 9064
rect 2225 9055 2283 9061
rect 2608 8956 2636 9064
rect 2774 9052 2780 9064
rect 2832 9092 2838 9104
rect 3142 9092 3148 9104
rect 2832 9064 3148 9092
rect 2832 9052 2838 9064
rect 3142 9052 3148 9064
rect 3200 9052 3206 9104
rect 4540 9064 4936 9092
rect 2685 9027 2743 9033
rect 2685 8993 2697 9027
rect 2731 9024 2743 9027
rect 4540 9024 4568 9064
rect 4706 9024 4712 9036
rect 2731 8996 4568 9024
rect 4667 8996 4712 9024
rect 2731 8993 2743 8996
rect 2685 8987 2743 8993
rect 4706 8984 4712 8996
rect 4764 8984 4770 9036
rect 4908 9033 4936 9064
rect 5718 9052 5724 9104
rect 5776 9092 5782 9104
rect 6089 9095 6147 9101
rect 6089 9092 6101 9095
rect 5776 9064 6101 9092
rect 5776 9052 5782 9064
rect 6089 9061 6101 9064
rect 6135 9092 6147 9095
rect 6135 9064 7696 9092
rect 6135 9061 6147 9064
rect 6089 9055 6147 9061
rect 4893 9027 4951 9033
rect 4893 8993 4905 9027
rect 4939 9024 4951 9027
rect 4982 9024 4988 9036
rect 4939 8996 4988 9024
rect 4939 8993 4951 8996
rect 4893 8987 4951 8993
rect 4982 8984 4988 8996
rect 5040 8984 5046 9036
rect 6730 8984 6736 9036
rect 6788 9024 6794 9036
rect 6917 9027 6975 9033
rect 6917 9024 6929 9027
rect 6788 8996 6929 9024
rect 6788 8984 6794 8996
rect 6917 8993 6929 8996
rect 6963 8993 6975 9027
rect 6917 8987 6975 8993
rect 2777 8959 2835 8965
rect 2777 8956 2789 8959
rect 2608 8928 2789 8956
rect 2777 8925 2789 8928
rect 2823 8925 2835 8959
rect 4246 8956 4252 8968
rect 2777 8919 2835 8925
rect 3896 8928 4252 8956
rect 1210 8848 1216 8900
rect 1268 8888 1274 8900
rect 3896 8897 3924 8928
rect 4246 8916 4252 8928
rect 4304 8916 4310 8968
rect 4430 8916 4436 8968
rect 4488 8956 4494 8968
rect 4617 8959 4675 8965
rect 4617 8956 4629 8959
rect 4488 8928 4629 8956
rect 4488 8916 4494 8928
rect 4617 8925 4629 8928
rect 4663 8925 4675 8959
rect 7466 8956 7472 8968
rect 4617 8919 4675 8925
rect 5644 8928 7472 8956
rect 3881 8891 3939 8897
rect 3881 8888 3893 8891
rect 1268 8860 3893 8888
rect 1268 8848 1274 8860
rect 3881 8857 3893 8860
rect 3927 8857 3939 8891
rect 3881 8851 3939 8857
rect 4062 8848 4068 8900
rect 4120 8888 4126 8900
rect 5644 8888 5672 8928
rect 7466 8916 7472 8928
rect 7524 8916 7530 8968
rect 7668 8956 7696 9064
rect 12986 9052 12992 9104
rect 13044 9092 13050 9104
rect 14550 9092 14556 9104
rect 13044 9064 14556 9092
rect 13044 9052 13050 9064
rect 14550 9052 14556 9064
rect 14608 9052 14614 9104
rect 8021 9027 8079 9033
rect 8021 8993 8033 9027
rect 8067 9024 8079 9027
rect 9766 9024 9772 9036
rect 8067 8996 9772 9024
rect 8067 8993 8079 8996
rect 8021 8987 8079 8993
rect 9766 8984 9772 8996
rect 9824 8984 9830 9036
rect 12894 8984 12900 9036
rect 12952 9024 12958 9036
rect 21085 9027 21143 9033
rect 12952 8996 13400 9024
rect 12952 8984 12958 8996
rect 7745 8959 7803 8965
rect 7745 8956 7757 8959
rect 7668 8928 7757 8956
rect 7745 8925 7757 8928
rect 7791 8956 7803 8959
rect 8941 8959 8999 8965
rect 8941 8956 8953 8959
rect 7791 8928 8953 8956
rect 7791 8925 7803 8928
rect 7745 8919 7803 8925
rect 8941 8925 8953 8928
rect 8987 8956 8999 8959
rect 9122 8956 9128 8968
rect 8987 8928 9128 8956
rect 8987 8925 8999 8928
rect 8941 8919 8999 8925
rect 9122 8916 9128 8928
rect 9180 8916 9186 8968
rect 10318 8916 10324 8968
rect 10376 8956 10382 8968
rect 10870 8956 10876 8968
rect 10928 8965 10934 8968
rect 10376 8928 10876 8956
rect 10376 8916 10382 8928
rect 10870 8916 10876 8928
rect 10928 8919 10940 8965
rect 11146 8956 11152 8968
rect 11059 8928 11152 8956
rect 10928 8916 10934 8919
rect 11146 8916 11152 8928
rect 11204 8956 11210 8968
rect 12805 8959 12863 8965
rect 12805 8956 12817 8959
rect 11204 8928 12817 8956
rect 11204 8916 11210 8928
rect 12805 8925 12817 8928
rect 12851 8956 12863 8959
rect 12851 8928 13216 8956
rect 12851 8925 12863 8928
rect 12805 8919 12863 8925
rect 4120 8860 5672 8888
rect 4120 8848 4126 8860
rect 7006 8848 7012 8900
rect 7064 8888 7070 8900
rect 7837 8891 7895 8897
rect 7837 8888 7849 8891
rect 7064 8860 7849 8888
rect 7064 8848 7070 8860
rect 7837 8857 7849 8860
rect 7883 8857 7895 8891
rect 7837 8851 7895 8857
rect 2774 8780 2780 8832
rect 2832 8820 2838 8832
rect 2869 8823 2927 8829
rect 2869 8820 2881 8823
rect 2832 8792 2881 8820
rect 2832 8780 2838 8792
rect 2869 8789 2881 8792
rect 2915 8789 2927 8823
rect 2869 8783 2927 8789
rect 5258 8780 5264 8832
rect 5316 8820 5322 8832
rect 5353 8823 5411 8829
rect 5353 8820 5365 8823
rect 5316 8792 5365 8820
rect 5316 8780 5322 8792
rect 5353 8789 5365 8792
rect 5399 8789 5411 8823
rect 6638 8820 6644 8832
rect 6599 8792 6644 8820
rect 5353 8783 5411 8789
rect 6638 8780 6644 8792
rect 6696 8780 6702 8832
rect 7374 8820 7380 8832
rect 7335 8792 7380 8820
rect 7374 8780 7380 8792
rect 7432 8780 7438 8832
rect 7852 8820 7880 8851
rect 8294 8848 8300 8900
rect 8352 8888 8358 8900
rect 8352 8860 11560 8888
rect 8352 8848 8358 8860
rect 8389 8823 8447 8829
rect 8389 8820 8401 8823
rect 7852 8792 8401 8820
rect 8389 8789 8401 8792
rect 8435 8789 8447 8823
rect 9490 8820 9496 8832
rect 9451 8792 9496 8820
rect 8389 8783 8447 8789
rect 9490 8780 9496 8792
rect 9548 8780 9554 8832
rect 9766 8820 9772 8832
rect 9727 8792 9772 8820
rect 9766 8780 9772 8792
rect 9824 8780 9830 8832
rect 10870 8780 10876 8832
rect 10928 8820 10934 8832
rect 11425 8823 11483 8829
rect 11425 8820 11437 8823
rect 10928 8792 11437 8820
rect 10928 8780 10934 8792
rect 11425 8789 11437 8792
rect 11471 8789 11483 8823
rect 11532 8820 11560 8860
rect 11974 8848 11980 8900
rect 12032 8888 12038 8900
rect 12538 8891 12596 8897
rect 12538 8888 12550 8891
rect 12032 8860 12550 8888
rect 12032 8848 12038 8860
rect 12538 8857 12550 8860
rect 12584 8857 12596 8891
rect 12538 8851 12596 8857
rect 12986 8820 12992 8832
rect 11532 8792 12992 8820
rect 11425 8783 11483 8789
rect 12986 8780 12992 8792
rect 13044 8780 13050 8832
rect 13188 8829 13216 8928
rect 13372 8888 13400 8996
rect 21085 8993 21097 9027
rect 21131 9024 21143 9027
rect 21358 9024 21364 9036
rect 21131 8996 21364 9024
rect 21131 8993 21143 8996
rect 21085 8987 21143 8993
rect 13446 8916 13452 8968
rect 13504 8956 13510 8968
rect 15298 8959 15356 8965
rect 15298 8956 15310 8959
rect 13504 8928 15310 8956
rect 13504 8916 13510 8928
rect 15298 8925 15310 8928
rect 15344 8925 15356 8959
rect 15298 8919 15356 8925
rect 15565 8959 15623 8965
rect 15565 8925 15577 8959
rect 15611 8956 15623 8959
rect 15746 8956 15752 8968
rect 15611 8928 15752 8956
rect 15611 8925 15623 8928
rect 15565 8919 15623 8925
rect 15746 8916 15752 8928
rect 15804 8956 15810 8968
rect 17313 8959 17371 8965
rect 17313 8956 17325 8959
rect 15804 8928 17325 8956
rect 15804 8916 15810 8928
rect 17313 8925 17325 8928
rect 17359 8956 17371 8959
rect 17681 8959 17739 8965
rect 17681 8956 17693 8959
rect 17359 8928 17693 8956
rect 17359 8925 17371 8928
rect 17313 8919 17371 8925
rect 17681 8925 17693 8928
rect 17727 8956 17739 8959
rect 18233 8959 18291 8965
rect 18233 8956 18245 8959
rect 17727 8928 18245 8956
rect 17727 8925 17739 8928
rect 17681 8919 17739 8925
rect 18233 8925 18245 8928
rect 18279 8956 18291 8959
rect 18322 8956 18328 8968
rect 18279 8928 18328 8956
rect 18279 8925 18291 8928
rect 18233 8919 18291 8925
rect 18322 8916 18328 8928
rect 18380 8956 18386 8968
rect 18601 8959 18659 8965
rect 18601 8956 18613 8959
rect 18380 8928 18613 8956
rect 18380 8916 18386 8928
rect 18601 8925 18613 8928
rect 18647 8956 18659 8959
rect 19429 8959 19487 8965
rect 19429 8956 19441 8959
rect 18647 8928 19441 8956
rect 18647 8925 18659 8928
rect 18601 8919 18659 8925
rect 19429 8925 19441 8928
rect 19475 8956 19487 8959
rect 19978 8956 19984 8968
rect 19475 8928 19984 8956
rect 19475 8925 19487 8928
rect 19429 8919 19487 8925
rect 19978 8916 19984 8928
rect 20036 8956 20042 8968
rect 21100 8956 21128 8987
rect 21358 8984 21364 8996
rect 21416 8984 21422 9036
rect 20036 8928 21128 8956
rect 20036 8916 20042 8928
rect 16942 8888 16948 8900
rect 13372 8860 16948 8888
rect 16942 8848 16948 8860
rect 17000 8848 17006 8900
rect 17068 8891 17126 8897
rect 17068 8857 17080 8891
rect 17114 8888 17126 8891
rect 18046 8888 18052 8900
rect 17114 8860 18052 8888
rect 17114 8857 17126 8860
rect 17068 8851 17126 8857
rect 18046 8848 18052 8860
rect 18104 8848 18110 8900
rect 20714 8848 20720 8900
rect 20772 8888 20778 8900
rect 20818 8891 20876 8897
rect 20818 8888 20830 8891
rect 20772 8860 20830 8888
rect 20772 8848 20778 8860
rect 20818 8857 20830 8860
rect 20864 8857 20876 8891
rect 20818 8851 20876 8857
rect 13173 8823 13231 8829
rect 13173 8789 13185 8823
rect 13219 8820 13231 8823
rect 13262 8820 13268 8832
rect 13219 8792 13268 8820
rect 13219 8789 13231 8792
rect 13173 8783 13231 8789
rect 13262 8780 13268 8792
rect 13320 8780 13326 8832
rect 14185 8823 14243 8829
rect 14185 8789 14197 8823
rect 14231 8820 14243 8823
rect 14366 8820 14372 8832
rect 14231 8792 14372 8820
rect 14231 8789 14243 8792
rect 14185 8783 14243 8789
rect 14366 8780 14372 8792
rect 14424 8780 14430 8832
rect 14550 8780 14556 8832
rect 14608 8820 14614 8832
rect 18966 8820 18972 8832
rect 14608 8792 18972 8820
rect 14608 8780 14614 8792
rect 18966 8780 18972 8792
rect 19024 8780 19030 8832
rect 1104 8730 22056 8752
rect 1104 8678 6148 8730
rect 6200 8678 6212 8730
rect 6264 8678 6276 8730
rect 6328 8678 6340 8730
rect 6392 8678 6404 8730
rect 6456 8678 11346 8730
rect 11398 8678 11410 8730
rect 11462 8678 11474 8730
rect 11526 8678 11538 8730
rect 11590 8678 11602 8730
rect 11654 8678 16544 8730
rect 16596 8678 16608 8730
rect 16660 8678 16672 8730
rect 16724 8678 16736 8730
rect 16788 8678 16800 8730
rect 16852 8678 21742 8730
rect 21794 8678 21806 8730
rect 21858 8678 21870 8730
rect 21922 8678 21934 8730
rect 21986 8678 21998 8730
rect 22050 8678 22056 8730
rect 1104 8656 22056 8678
rect 2774 8576 2780 8628
rect 2832 8616 2838 8628
rect 2832 8588 2877 8616
rect 2832 8576 2838 8588
rect 3326 8576 3332 8628
rect 3384 8616 3390 8628
rect 3513 8619 3571 8625
rect 3513 8616 3525 8619
rect 3384 8588 3525 8616
rect 3384 8576 3390 8588
rect 3513 8585 3525 8588
rect 3559 8616 3571 8619
rect 5258 8616 5264 8628
rect 3559 8588 4568 8616
rect 5219 8588 5264 8616
rect 3559 8585 3571 8588
rect 3513 8579 3571 8585
rect 2314 8508 2320 8560
rect 2372 8548 2378 8560
rect 4540 8548 4568 8588
rect 5258 8576 5264 8588
rect 5316 8576 5322 8628
rect 6638 8576 6644 8628
rect 6696 8616 6702 8628
rect 7469 8619 7527 8625
rect 7469 8616 7481 8619
rect 6696 8588 7481 8616
rect 6696 8576 6702 8588
rect 7469 8585 7481 8588
rect 7515 8585 7527 8619
rect 7469 8579 7527 8585
rect 9490 8576 9496 8628
rect 9548 8616 9554 8628
rect 9769 8619 9827 8625
rect 9769 8616 9781 8619
rect 9548 8588 9781 8616
rect 9548 8576 9554 8588
rect 9769 8585 9781 8588
rect 9815 8585 9827 8619
rect 11146 8616 11152 8628
rect 11107 8588 11152 8616
rect 9769 8579 9827 8585
rect 11146 8576 11152 8588
rect 11204 8576 11210 8628
rect 13354 8616 13360 8628
rect 11256 8588 13032 8616
rect 13315 8588 13360 8616
rect 5353 8551 5411 8557
rect 5353 8548 5365 8551
rect 2372 8520 4476 8548
rect 4540 8520 5365 8548
rect 2372 8508 2378 8520
rect 3418 8440 3424 8492
rect 3476 8480 3482 8492
rect 3970 8480 3976 8492
rect 3476 8452 3976 8480
rect 3476 8440 3482 8452
rect 3970 8440 3976 8452
rect 4028 8440 4034 8492
rect 4246 8480 4252 8492
rect 4207 8452 4252 8480
rect 4246 8440 4252 8452
rect 4304 8440 4310 8492
rect 4338 8412 4344 8424
rect 4299 8384 4344 8412
rect 4338 8372 4344 8384
rect 4396 8372 4402 8424
rect 4448 8421 4476 8520
rect 5353 8517 5365 8520
rect 5399 8517 5411 8551
rect 5353 8511 5411 8517
rect 6825 8483 6883 8489
rect 6825 8449 6837 8483
rect 6871 8480 6883 8483
rect 8481 8483 8539 8489
rect 8481 8480 8493 8483
rect 6871 8452 8493 8480
rect 6871 8449 6883 8452
rect 6825 8443 6883 8449
rect 8481 8449 8493 8452
rect 8527 8449 8539 8483
rect 11256 8480 11284 8588
rect 12894 8548 12900 8560
rect 8481 8443 8539 8449
rect 8772 8452 11284 8480
rect 11440 8520 12900 8548
rect 4433 8415 4491 8421
rect 4433 8381 4445 8415
rect 4479 8381 4491 8415
rect 4433 8375 4491 8381
rect 5445 8415 5503 8421
rect 5445 8381 5457 8415
rect 5491 8412 5503 8415
rect 5626 8412 5632 8424
rect 5491 8384 5632 8412
rect 5491 8381 5503 8384
rect 5445 8375 5503 8381
rect 5626 8372 5632 8384
rect 5684 8372 5690 8424
rect 7558 8412 7564 8424
rect 7519 8384 7564 8412
rect 7558 8372 7564 8384
rect 7616 8372 7622 8424
rect 7650 8372 7656 8424
rect 7708 8412 7714 8424
rect 8570 8412 8576 8424
rect 7708 8384 7753 8412
rect 8531 8384 8576 8412
rect 7708 8372 7714 8384
rect 8570 8372 8576 8384
rect 8628 8372 8634 8424
rect 8772 8421 8800 8452
rect 8757 8415 8815 8421
rect 8757 8381 8769 8415
rect 8803 8381 8815 8415
rect 9858 8412 9864 8424
rect 9819 8384 9864 8412
rect 8757 8375 8815 8381
rect 9858 8372 9864 8384
rect 9916 8372 9922 8424
rect 10045 8415 10103 8421
rect 10045 8381 10057 8415
rect 10091 8412 10103 8415
rect 11440 8412 11468 8520
rect 12894 8508 12900 8520
rect 12952 8508 12958 8560
rect 12250 8440 12256 8492
rect 12308 8480 12314 8492
rect 12814 8483 12872 8489
rect 12814 8480 12826 8483
rect 12308 8452 12826 8480
rect 12308 8440 12314 8452
rect 12814 8449 12826 8452
rect 12860 8449 12872 8483
rect 13004 8480 13032 8588
rect 13354 8576 13360 8588
rect 13412 8576 13418 8628
rect 15746 8616 15752 8628
rect 15707 8588 15752 8616
rect 15746 8576 15752 8588
rect 15804 8576 15810 8628
rect 17954 8576 17960 8628
rect 18012 8616 18018 8628
rect 18049 8619 18107 8625
rect 18049 8616 18061 8619
rect 18012 8588 18061 8616
rect 18012 8576 18018 8588
rect 18049 8585 18061 8588
rect 18095 8585 18107 8619
rect 18049 8579 18107 8585
rect 21361 8619 21419 8625
rect 21361 8585 21373 8619
rect 21407 8616 21419 8619
rect 21450 8616 21456 8628
rect 21407 8588 21456 8616
rect 21407 8585 21419 8588
rect 21361 8579 21419 8585
rect 13078 8508 13084 8560
rect 13136 8548 13142 8560
rect 13136 8520 14688 8548
rect 13136 8508 13142 8520
rect 14182 8480 14188 8492
rect 13004 8452 14188 8480
rect 12814 8443 12872 8449
rect 14182 8440 14188 8452
rect 14240 8440 14246 8492
rect 14458 8440 14464 8492
rect 14516 8489 14522 8492
rect 14516 8480 14528 8489
rect 14516 8452 14561 8480
rect 14516 8443 14528 8452
rect 14516 8440 14522 8443
rect 10091 8384 11468 8412
rect 13081 8415 13139 8421
rect 10091 8381 10103 8384
rect 10045 8375 10103 8381
rect 13081 8381 13093 8415
rect 13127 8412 13139 8415
rect 13262 8412 13268 8424
rect 13127 8384 13268 8412
rect 13127 8381 13139 8384
rect 13081 8375 13139 8381
rect 13262 8372 13268 8384
rect 13320 8372 13326 8424
rect 14660 8412 14688 8520
rect 14737 8483 14795 8489
rect 14737 8449 14749 8483
rect 14783 8480 14795 8483
rect 15105 8483 15163 8489
rect 15105 8480 15117 8483
rect 14783 8452 15117 8480
rect 14783 8449 14795 8452
rect 14737 8443 14795 8449
rect 15105 8449 15117 8452
rect 15151 8480 15163 8483
rect 15764 8480 15792 8576
rect 18064 8548 18092 8579
rect 21450 8576 21456 8588
rect 21508 8576 21514 8628
rect 20226 8551 20284 8557
rect 20226 8548 20238 8551
rect 18064 8520 20238 8548
rect 20226 8517 20238 8520
rect 20272 8517 20284 8551
rect 20226 8511 20284 8517
rect 16669 8483 16727 8489
rect 16669 8480 16681 8483
rect 15151 8452 16681 8480
rect 15151 8449 15163 8452
rect 15105 8443 15163 8449
rect 16669 8449 16681 8452
rect 16715 8449 16727 8483
rect 16925 8483 16983 8489
rect 16925 8480 16937 8483
rect 16669 8443 16727 8449
rect 16776 8452 16937 8480
rect 16776 8412 16804 8452
rect 16925 8449 16937 8452
rect 16971 8449 16983 8483
rect 18322 8480 18328 8492
rect 18283 8452 18328 8480
rect 16925 8443 16983 8449
rect 18322 8440 18328 8452
rect 18380 8440 18386 8492
rect 18414 8440 18420 8492
rect 18472 8480 18478 8492
rect 18581 8483 18639 8489
rect 18581 8480 18593 8483
rect 18472 8452 18593 8480
rect 18472 8440 18478 8452
rect 18581 8449 18593 8452
rect 18627 8449 18639 8483
rect 19978 8480 19984 8492
rect 19939 8452 19984 8480
rect 18581 8443 18639 8449
rect 19978 8440 19984 8452
rect 20036 8440 20042 8492
rect 14660 8384 16804 8412
rect 3881 8347 3939 8353
rect 3881 8313 3893 8347
rect 3927 8344 3939 8347
rect 4154 8344 4160 8356
rect 3927 8316 4160 8344
rect 3927 8313 3939 8316
rect 3881 8307 3939 8313
rect 4154 8304 4160 8316
rect 4212 8304 4218 8356
rect 5074 8304 5080 8356
rect 5132 8344 5138 8356
rect 5905 8347 5963 8353
rect 5905 8344 5917 8347
rect 5132 8316 5917 8344
rect 5132 8304 5138 8316
rect 5905 8313 5917 8316
rect 5951 8313 5963 8347
rect 5905 8307 5963 8313
rect 7101 8347 7159 8353
rect 7101 8313 7113 8347
rect 7147 8344 7159 8347
rect 7190 8344 7196 8356
rect 7147 8316 7196 8344
rect 7147 8313 7159 8316
rect 7101 8307 7159 8313
rect 7190 8304 7196 8316
rect 7248 8304 7254 8356
rect 7742 8304 7748 8356
rect 7800 8344 7806 8356
rect 8113 8347 8171 8353
rect 8113 8344 8125 8347
rect 7800 8316 8125 8344
rect 7800 8304 7806 8316
rect 8113 8313 8125 8316
rect 8159 8313 8171 8347
rect 8113 8307 8171 8313
rect 11701 8347 11759 8353
rect 11701 8313 11713 8347
rect 11747 8344 11759 8347
rect 11974 8344 11980 8356
rect 11747 8316 11980 8344
rect 11747 8313 11759 8316
rect 11701 8307 11759 8313
rect 11974 8304 11980 8316
rect 12032 8304 12038 8356
rect 19705 8347 19763 8353
rect 19705 8313 19717 8347
rect 19751 8313 19763 8347
rect 19705 8307 19763 8313
rect 4890 8276 4896 8288
rect 4851 8248 4896 8276
rect 4890 8236 4896 8248
rect 4948 8236 4954 8288
rect 9398 8276 9404 8288
rect 9359 8248 9404 8276
rect 9398 8236 9404 8248
rect 9456 8236 9462 8288
rect 18506 8236 18512 8288
rect 18564 8276 18570 8288
rect 19720 8276 19748 8307
rect 20714 8276 20720 8288
rect 18564 8248 20720 8276
rect 18564 8236 18570 8248
rect 20714 8236 20720 8248
rect 20772 8236 20778 8288
rect 1104 8186 21896 8208
rect 1104 8134 3549 8186
rect 3601 8134 3613 8186
rect 3665 8134 3677 8186
rect 3729 8134 3741 8186
rect 3793 8134 3805 8186
rect 3857 8134 8747 8186
rect 8799 8134 8811 8186
rect 8863 8134 8875 8186
rect 8927 8134 8939 8186
rect 8991 8134 9003 8186
rect 9055 8134 13945 8186
rect 13997 8134 14009 8186
rect 14061 8134 14073 8186
rect 14125 8134 14137 8186
rect 14189 8134 14201 8186
rect 14253 8134 19143 8186
rect 19195 8134 19207 8186
rect 19259 8134 19271 8186
rect 19323 8134 19335 8186
rect 19387 8134 19399 8186
rect 19451 8134 21896 8186
rect 1104 8112 21896 8134
rect 4157 8075 4215 8081
rect 4157 8041 4169 8075
rect 4203 8072 4215 8075
rect 4246 8072 4252 8084
rect 4203 8044 4252 8072
rect 4203 8041 4215 8044
rect 4157 8035 4215 8041
rect 4246 8032 4252 8044
rect 4304 8032 4310 8084
rect 5258 8032 5264 8084
rect 5316 8072 5322 8084
rect 6825 8075 6883 8081
rect 6825 8072 6837 8075
rect 5316 8044 6837 8072
rect 5316 8032 5322 8044
rect 6825 8041 6837 8044
rect 6871 8041 6883 8075
rect 6825 8035 6883 8041
rect 7193 8075 7251 8081
rect 7193 8041 7205 8075
rect 7239 8072 7251 8075
rect 7558 8072 7564 8084
rect 7239 8044 7564 8072
rect 7239 8041 7251 8044
rect 7193 8035 7251 8041
rect 6546 8004 6552 8016
rect 4816 7976 6552 8004
rect 3234 7896 3240 7948
rect 3292 7936 3298 7948
rect 4614 7936 4620 7948
rect 3292 7908 4620 7936
rect 3292 7896 3298 7908
rect 4614 7896 4620 7908
rect 4672 7896 4678 7948
rect 4816 7945 4844 7976
rect 6546 7964 6552 7976
rect 6604 7964 6610 8016
rect 4801 7939 4859 7945
rect 4801 7905 4813 7939
rect 4847 7905 4859 7939
rect 4801 7899 4859 7905
rect 5353 7939 5411 7945
rect 5353 7905 5365 7939
rect 5399 7936 5411 7939
rect 5534 7936 5540 7948
rect 5399 7908 5540 7936
rect 5399 7905 5411 7908
rect 5353 7899 5411 7905
rect 5534 7896 5540 7908
rect 5592 7896 5598 7948
rect 6840 7936 6868 8035
rect 7558 8032 7564 8044
rect 7616 8032 7622 8084
rect 8386 8032 8392 8084
rect 8444 8072 8450 8084
rect 8481 8075 8539 8081
rect 8481 8072 8493 8075
rect 8444 8044 8493 8072
rect 8444 8032 8450 8044
rect 8481 8041 8493 8044
rect 8527 8072 8539 8075
rect 8527 8044 8708 8072
rect 8527 8041 8539 8044
rect 8481 8035 8539 8041
rect 7653 7939 7711 7945
rect 7653 7936 7665 7939
rect 6840 7908 7665 7936
rect 7653 7905 7665 7908
rect 7699 7905 7711 7939
rect 7834 7936 7840 7948
rect 7795 7908 7840 7936
rect 7653 7899 7711 7905
rect 7834 7896 7840 7908
rect 7892 7896 7898 7948
rect 3878 7828 3884 7880
rect 3936 7868 3942 7880
rect 6457 7871 6515 7877
rect 6457 7868 6469 7871
rect 3936 7840 6469 7868
rect 3936 7828 3942 7840
rect 6457 7837 6469 7840
rect 6503 7868 6515 7871
rect 7561 7871 7619 7877
rect 7561 7868 7573 7871
rect 6503 7840 7573 7868
rect 6503 7837 6515 7840
rect 6457 7831 6515 7837
rect 7561 7837 7573 7840
rect 7607 7837 7619 7871
rect 8570 7868 8576 7880
rect 7561 7831 7619 7837
rect 7668 7840 8576 7868
rect 3418 7800 3424 7812
rect 3331 7772 3424 7800
rect 3418 7760 3424 7772
rect 3476 7800 3482 7812
rect 5537 7803 5595 7809
rect 5537 7800 5549 7803
rect 3476 7772 5549 7800
rect 3476 7760 3482 7772
rect 5537 7769 5549 7772
rect 5583 7769 5595 7803
rect 5537 7763 5595 7769
rect 3053 7735 3111 7741
rect 3053 7701 3065 7735
rect 3099 7732 3111 7735
rect 3234 7732 3240 7744
rect 3099 7704 3240 7732
rect 3099 7701 3111 7704
rect 3053 7695 3111 7701
rect 3234 7692 3240 7704
rect 3292 7692 3298 7744
rect 3878 7732 3884 7744
rect 3839 7704 3884 7732
rect 3878 7692 3884 7704
rect 3936 7732 3942 7744
rect 4525 7735 4583 7741
rect 4525 7732 4537 7735
rect 3936 7704 4537 7732
rect 3936 7692 3942 7704
rect 4525 7701 4537 7704
rect 4571 7732 4583 7735
rect 5258 7732 5264 7744
rect 4571 7704 5264 7732
rect 4571 7701 4583 7704
rect 4525 7695 4583 7701
rect 5258 7692 5264 7704
rect 5316 7692 5322 7744
rect 5442 7732 5448 7744
rect 5403 7704 5448 7732
rect 5442 7692 5448 7704
rect 5500 7692 5506 7744
rect 5905 7735 5963 7741
rect 5905 7701 5917 7735
rect 5951 7732 5963 7735
rect 7668 7732 7696 7840
rect 8570 7828 8576 7840
rect 8628 7828 8634 7880
rect 8680 7868 8708 8044
rect 9858 8032 9864 8084
rect 9916 8072 9922 8084
rect 10045 8075 10103 8081
rect 10045 8072 10057 8075
rect 9916 8044 10057 8072
rect 9916 8032 9922 8044
rect 10045 8041 10057 8044
rect 10091 8041 10103 8075
rect 11330 8072 11336 8084
rect 11243 8044 11336 8072
rect 10045 8035 10103 8041
rect 11330 8032 11336 8044
rect 11388 8072 11394 8084
rect 15470 8072 15476 8084
rect 11388 8044 15476 8072
rect 11388 8032 11394 8044
rect 15470 8032 15476 8044
rect 15528 8032 15534 8084
rect 15654 8072 15660 8084
rect 15615 8044 15660 8072
rect 15654 8032 15660 8044
rect 15712 8072 15718 8084
rect 15712 8044 16896 8072
rect 15712 8032 15718 8044
rect 16868 8004 16896 8044
rect 16942 8032 16948 8084
rect 17000 8072 17006 8084
rect 17313 8075 17371 8081
rect 17313 8072 17325 8075
rect 17000 8044 17325 8072
rect 17000 8032 17006 8044
rect 17313 8041 17325 8044
rect 17359 8041 17371 8075
rect 17313 8035 17371 8041
rect 17681 8075 17739 8081
rect 17681 8041 17693 8075
rect 17727 8072 17739 8075
rect 18322 8072 18328 8084
rect 17727 8044 18328 8072
rect 17727 8041 17739 8044
rect 17681 8035 17739 8041
rect 18322 8032 18328 8044
rect 18380 8032 18386 8084
rect 19978 8072 19984 8084
rect 19260 8044 19984 8072
rect 18141 8007 18199 8013
rect 18141 8004 18153 8007
rect 16868 7976 18153 8004
rect 18141 7973 18153 7976
rect 18187 8004 18199 8007
rect 18414 8004 18420 8016
rect 18187 7976 18420 8004
rect 18187 7973 18199 7976
rect 18141 7967 18199 7973
rect 18414 7964 18420 7976
rect 18472 7964 18478 8016
rect 9493 7939 9551 7945
rect 9493 7905 9505 7939
rect 9539 7936 9551 7939
rect 9539 7908 11008 7936
rect 9539 7905 9551 7908
rect 9493 7899 9551 7905
rect 9677 7871 9735 7877
rect 9677 7868 9689 7871
rect 8680 7840 9689 7868
rect 9677 7837 9689 7840
rect 9723 7837 9735 7871
rect 10980 7868 11008 7908
rect 15746 7896 15752 7948
rect 15804 7936 15810 7948
rect 19260 7945 19288 8044
rect 19978 8032 19984 8044
rect 20036 8072 20042 8084
rect 20901 8075 20959 8081
rect 20901 8072 20913 8075
rect 20036 8044 20913 8072
rect 20036 8032 20042 8044
rect 20901 8041 20913 8044
rect 20947 8072 20959 8075
rect 21082 8072 21088 8084
rect 20947 8044 21088 8072
rect 20947 8041 20959 8044
rect 20901 8035 20959 8041
rect 21082 8032 21088 8044
rect 21140 8072 21146 8084
rect 21269 8075 21327 8081
rect 21269 8072 21281 8075
rect 21140 8044 21281 8072
rect 21140 8032 21146 8044
rect 21269 8041 21281 8044
rect 21315 8041 21327 8075
rect 21269 8035 21327 8041
rect 15933 7939 15991 7945
rect 15933 7936 15945 7939
rect 15804 7908 15945 7936
rect 15804 7896 15810 7908
rect 15933 7905 15945 7908
rect 15979 7905 15991 7939
rect 15933 7899 15991 7905
rect 19245 7939 19303 7945
rect 19245 7905 19257 7939
rect 19291 7905 19303 7939
rect 19245 7899 19303 7905
rect 12713 7871 12771 7877
rect 10980 7840 12434 7868
rect 9677 7831 9735 7837
rect 8202 7760 8208 7812
rect 8260 7800 8266 7812
rect 11330 7800 11336 7812
rect 8260 7772 11336 7800
rect 8260 7760 8266 7772
rect 11330 7760 11336 7772
rect 11388 7760 11394 7812
rect 5951 7704 7696 7732
rect 5951 7701 5963 7704
rect 5905 7695 5963 7701
rect 8018 7692 8024 7744
rect 8076 7732 8082 7744
rect 9033 7735 9091 7741
rect 9033 7732 9045 7735
rect 8076 7704 9045 7732
rect 8076 7692 8082 7704
rect 9033 7701 9045 7704
rect 9079 7732 9091 7735
rect 9585 7735 9643 7741
rect 9585 7732 9597 7735
rect 9079 7704 9597 7732
rect 9079 7701 9091 7704
rect 9033 7695 9091 7701
rect 9585 7701 9597 7704
rect 9631 7701 9643 7735
rect 12406 7732 12434 7840
rect 12713 7837 12725 7871
rect 12759 7868 12771 7871
rect 13262 7868 13268 7880
rect 12759 7840 13268 7868
rect 12759 7837 12771 7840
rect 12713 7831 12771 7837
rect 13262 7828 13268 7840
rect 13320 7868 13326 7880
rect 13633 7871 13691 7877
rect 13633 7868 13645 7871
rect 13320 7840 13645 7868
rect 13320 7828 13326 7840
rect 13633 7837 13645 7840
rect 13679 7868 13691 7871
rect 13722 7868 13728 7880
rect 13679 7840 13728 7868
rect 13679 7837 13691 7840
rect 13633 7831 13691 7837
rect 13722 7828 13728 7840
rect 13780 7868 13786 7880
rect 14277 7871 14335 7877
rect 14277 7868 14289 7871
rect 13780 7840 14289 7868
rect 13780 7828 13786 7840
rect 14277 7837 14289 7840
rect 14323 7868 14335 7871
rect 15764 7868 15792 7896
rect 14323 7840 15792 7868
rect 14323 7837 14335 7840
rect 14277 7831 14335 7837
rect 12526 7809 12532 7812
rect 12468 7803 12532 7809
rect 12468 7769 12480 7803
rect 12514 7769 12532 7803
rect 12468 7763 12532 7769
rect 12526 7760 12532 7763
rect 12584 7760 12590 7812
rect 13814 7760 13820 7812
rect 13872 7800 13878 7812
rect 16206 7809 16212 7812
rect 14522 7803 14580 7809
rect 14522 7800 14534 7803
rect 13872 7772 14534 7800
rect 13872 7760 13878 7772
rect 14522 7769 14534 7772
rect 14568 7769 14580 7803
rect 16200 7800 16212 7809
rect 14522 7763 14580 7769
rect 14752 7772 16212 7800
rect 14752 7732 14780 7772
rect 16200 7763 16212 7772
rect 16206 7760 16212 7763
rect 16264 7760 16270 7812
rect 19512 7803 19570 7809
rect 19512 7769 19524 7803
rect 19558 7800 19570 7803
rect 19610 7800 19616 7812
rect 19558 7772 19616 7800
rect 19558 7769 19570 7772
rect 19512 7763 19570 7769
rect 19610 7760 19616 7772
rect 19668 7760 19674 7812
rect 12406 7704 14780 7732
rect 9585 7695 9643 7701
rect 17402 7692 17408 7744
rect 17460 7732 17466 7744
rect 19426 7732 19432 7744
rect 17460 7704 19432 7732
rect 17460 7692 17466 7704
rect 19426 7692 19432 7704
rect 19484 7692 19490 7744
rect 20622 7732 20628 7744
rect 20583 7704 20628 7732
rect 20622 7692 20628 7704
rect 20680 7692 20686 7744
rect 1104 7642 22056 7664
rect 1104 7590 6148 7642
rect 6200 7590 6212 7642
rect 6264 7590 6276 7642
rect 6328 7590 6340 7642
rect 6392 7590 6404 7642
rect 6456 7590 11346 7642
rect 11398 7590 11410 7642
rect 11462 7590 11474 7642
rect 11526 7590 11538 7642
rect 11590 7590 11602 7642
rect 11654 7590 16544 7642
rect 16596 7590 16608 7642
rect 16660 7590 16672 7642
rect 16724 7590 16736 7642
rect 16788 7590 16800 7642
rect 16852 7590 21742 7642
rect 21794 7590 21806 7642
rect 21858 7590 21870 7642
rect 21922 7590 21934 7642
rect 21986 7590 21998 7642
rect 22050 7590 22056 7642
rect 1104 7568 22056 7590
rect 2409 7531 2467 7537
rect 2409 7497 2421 7531
rect 2455 7528 2467 7531
rect 2958 7528 2964 7540
rect 2455 7500 2964 7528
rect 2455 7497 2467 7500
rect 2409 7491 2467 7497
rect 1857 7395 1915 7401
rect 1857 7361 1869 7395
rect 1903 7392 1915 7395
rect 2424 7392 2452 7491
rect 2958 7488 2964 7500
rect 3016 7488 3022 7540
rect 4338 7488 4344 7540
rect 4396 7528 4402 7540
rect 4433 7531 4491 7537
rect 4433 7528 4445 7531
rect 4396 7500 4445 7528
rect 4396 7488 4402 7500
rect 4433 7497 4445 7500
rect 4479 7497 4491 7531
rect 4433 7491 4491 7497
rect 4890 7488 4896 7540
rect 4948 7528 4954 7540
rect 5077 7531 5135 7537
rect 5077 7528 5089 7531
rect 4948 7500 5089 7528
rect 4948 7488 4954 7500
rect 5077 7497 5089 7500
rect 5123 7497 5135 7531
rect 7098 7528 7104 7540
rect 7059 7500 7104 7528
rect 5077 7491 5135 7497
rect 7098 7488 7104 7500
rect 7156 7488 7162 7540
rect 7374 7488 7380 7540
rect 7432 7528 7438 7540
rect 7561 7531 7619 7537
rect 7561 7528 7573 7531
rect 7432 7500 7573 7528
rect 7432 7488 7438 7500
rect 7561 7497 7573 7500
rect 7607 7497 7619 7531
rect 7561 7491 7619 7497
rect 11146 7488 11152 7540
rect 11204 7528 11210 7540
rect 11517 7531 11575 7537
rect 11517 7528 11529 7531
rect 11204 7500 11529 7528
rect 11204 7488 11210 7500
rect 11517 7497 11529 7500
rect 11563 7528 11575 7531
rect 12618 7528 12624 7540
rect 11563 7500 12624 7528
rect 11563 7497 11575 7500
rect 11517 7491 11575 7497
rect 12618 7488 12624 7500
rect 12676 7488 12682 7540
rect 14458 7488 14464 7540
rect 14516 7528 14522 7540
rect 15289 7531 15347 7537
rect 15289 7528 15301 7531
rect 14516 7500 15301 7528
rect 14516 7488 14522 7500
rect 15289 7497 15301 7500
rect 15335 7497 15347 7531
rect 15746 7528 15752 7540
rect 15707 7500 15752 7528
rect 15289 7491 15347 7497
rect 15746 7488 15752 7500
rect 15804 7528 15810 7540
rect 16117 7531 16175 7537
rect 16117 7528 16129 7531
rect 15804 7500 16129 7528
rect 15804 7488 15810 7500
rect 16117 7497 16129 7500
rect 16163 7497 16175 7531
rect 17402 7528 17408 7540
rect 17363 7500 17408 7528
rect 16117 7491 16175 7497
rect 17402 7488 17408 7500
rect 17460 7488 17466 7540
rect 18046 7488 18052 7540
rect 18104 7528 18110 7540
rect 19061 7531 19119 7537
rect 19061 7528 19073 7531
rect 18104 7500 19073 7528
rect 18104 7488 18110 7500
rect 19061 7497 19073 7500
rect 19107 7497 19119 7531
rect 20714 7528 20720 7540
rect 20675 7500 20720 7528
rect 19061 7491 19119 7497
rect 20714 7488 20720 7500
rect 20772 7488 20778 7540
rect 21082 7528 21088 7540
rect 21043 7500 21088 7528
rect 21082 7488 21088 7500
rect 21140 7488 21146 7540
rect 2682 7420 2688 7472
rect 2740 7460 2746 7472
rect 3421 7463 3479 7469
rect 3421 7460 3433 7463
rect 2740 7432 3433 7460
rect 2740 7420 2746 7432
rect 3421 7429 3433 7432
rect 3467 7460 3479 7463
rect 3973 7463 4031 7469
rect 3973 7460 3985 7463
rect 3467 7432 3985 7460
rect 3467 7429 3479 7432
rect 3421 7423 3479 7429
rect 3973 7429 3985 7432
rect 4019 7460 4031 7463
rect 4522 7460 4528 7472
rect 4019 7432 4528 7460
rect 4019 7429 4031 7432
rect 3973 7423 4031 7429
rect 4522 7420 4528 7432
rect 4580 7460 4586 7472
rect 5442 7460 5448 7472
rect 4580 7432 5448 7460
rect 4580 7420 4586 7432
rect 5442 7420 5448 7432
rect 5500 7460 5506 7472
rect 5721 7463 5779 7469
rect 5721 7460 5733 7463
rect 5500 7432 5733 7460
rect 5500 7420 5506 7432
rect 5721 7429 5733 7432
rect 5767 7429 5779 7463
rect 5721 7423 5779 7429
rect 10962 7420 10968 7472
rect 11020 7460 11026 7472
rect 13354 7460 13360 7472
rect 11020 7432 13360 7460
rect 11020 7420 11026 7432
rect 13354 7420 13360 7432
rect 13412 7460 13418 7472
rect 14154 7463 14212 7469
rect 14154 7460 14166 7463
rect 13412 7432 14166 7460
rect 13412 7420 13418 7432
rect 14154 7429 14166 7432
rect 14200 7429 14212 7463
rect 14154 7423 14212 7429
rect 1903 7364 2452 7392
rect 1903 7361 1915 7364
rect 1857 7355 1915 7361
rect 2958 7352 2964 7404
rect 3016 7392 3022 7404
rect 4065 7395 4123 7401
rect 4065 7392 4077 7395
rect 3016 7364 4077 7392
rect 3016 7352 3022 7364
rect 4065 7361 4077 7364
rect 4111 7361 4123 7395
rect 4065 7355 4123 7361
rect 4614 7352 4620 7404
rect 4672 7392 4678 7404
rect 6825 7395 6883 7401
rect 4672 7364 6776 7392
rect 4672 7352 4678 7364
rect 3881 7327 3939 7333
rect 3881 7293 3893 7327
rect 3927 7293 3939 7327
rect 4798 7324 4804 7336
rect 4759 7296 4804 7324
rect 3881 7287 3939 7293
rect 2038 7256 2044 7268
rect 1999 7228 2044 7256
rect 2038 7216 2044 7228
rect 2096 7216 2102 7268
rect 3896 7256 3924 7287
rect 4798 7284 4804 7296
rect 4856 7284 4862 7336
rect 4982 7324 4988 7336
rect 4943 7296 4988 7324
rect 4982 7284 4988 7296
rect 5040 7284 5046 7336
rect 6748 7324 6776 7364
rect 6825 7361 6837 7395
rect 6871 7392 6883 7395
rect 7469 7395 7527 7401
rect 7469 7392 7481 7395
rect 6871 7364 7481 7392
rect 6871 7361 6883 7364
rect 6825 7355 6883 7361
rect 7469 7361 7481 7364
rect 7515 7361 7527 7395
rect 8570 7392 8576 7404
rect 8531 7364 8576 7392
rect 7469 7355 7527 7361
rect 8570 7352 8576 7364
rect 8628 7352 8634 7404
rect 12342 7352 12348 7404
rect 12400 7392 12406 7404
rect 12630 7395 12688 7401
rect 12630 7392 12642 7395
rect 12400 7364 12642 7392
rect 12400 7352 12406 7364
rect 12630 7361 12642 7364
rect 12676 7361 12688 7395
rect 12630 7355 12688 7361
rect 12897 7395 12955 7401
rect 12897 7361 12909 7395
rect 12943 7392 12955 7395
rect 13265 7395 13323 7401
rect 13265 7392 13277 7395
rect 12943 7364 13277 7392
rect 12943 7361 12955 7364
rect 12897 7355 12955 7361
rect 13265 7361 13277 7364
rect 13311 7392 13323 7395
rect 13722 7392 13728 7404
rect 13311 7364 13728 7392
rect 13311 7361 13323 7364
rect 13265 7355 13323 7361
rect 13722 7352 13728 7364
rect 13780 7392 13786 7404
rect 13909 7395 13967 7401
rect 13909 7392 13921 7395
rect 13780 7364 13921 7392
rect 13780 7352 13786 7364
rect 13909 7361 13921 7364
rect 13955 7361 13967 7395
rect 17420 7392 17448 7488
rect 18322 7420 18328 7472
rect 18380 7460 18386 7472
rect 18380 7432 18828 7460
rect 18380 7420 18386 7432
rect 13909 7355 13967 7361
rect 14016 7364 17448 7392
rect 6914 7324 6920 7336
rect 6748 7296 6920 7324
rect 6914 7284 6920 7296
rect 6972 7284 6978 7336
rect 7745 7327 7803 7333
rect 7745 7293 7757 7327
rect 7791 7293 7803 7327
rect 7745 7287 7803 7293
rect 6546 7256 6552 7268
rect 3896 7228 6552 7256
rect 6546 7216 6552 7228
rect 6604 7216 6610 7268
rect 2958 7188 2964 7200
rect 2919 7160 2964 7188
rect 2958 7148 2964 7160
rect 3016 7148 3022 7200
rect 5442 7188 5448 7200
rect 5403 7160 5448 7188
rect 5442 7148 5448 7160
rect 5500 7148 5506 7200
rect 7760 7188 7788 7287
rect 8202 7284 8208 7336
rect 8260 7324 8266 7336
rect 8297 7327 8355 7333
rect 8297 7324 8309 7327
rect 8260 7296 8309 7324
rect 8260 7284 8266 7296
rect 8297 7293 8309 7296
rect 8343 7293 8355 7327
rect 14016 7324 14044 7364
rect 18506 7352 18512 7404
rect 18564 7401 18570 7404
rect 18800 7401 18828 7432
rect 18564 7392 18576 7401
rect 18785 7395 18843 7401
rect 18564 7364 18609 7392
rect 18564 7355 18576 7364
rect 18785 7361 18797 7395
rect 18831 7361 18843 7395
rect 20174 7395 20232 7401
rect 20174 7392 20186 7395
rect 18785 7355 18843 7361
rect 19444 7364 20186 7392
rect 18564 7352 18570 7355
rect 8297 7287 8355 7293
rect 13096 7296 14044 7324
rect 9582 7216 9588 7268
rect 9640 7256 9646 7268
rect 9640 7228 11652 7256
rect 9640 7216 9646 7228
rect 9858 7188 9864 7200
rect 7760 7160 9864 7188
rect 9858 7148 9864 7160
rect 9916 7148 9922 7200
rect 11624 7188 11652 7228
rect 13096 7188 13124 7296
rect 19444 7256 19472 7364
rect 20174 7361 20186 7364
rect 20220 7361 20232 7395
rect 20174 7355 20232 7361
rect 20441 7395 20499 7401
rect 20441 7361 20453 7395
rect 20487 7392 20499 7395
rect 21100 7392 21128 7488
rect 20487 7364 21128 7392
rect 20487 7361 20499 7364
rect 20441 7355 20499 7361
rect 15212 7228 17908 7256
rect 11624 7160 13124 7188
rect 13170 7148 13176 7200
rect 13228 7188 13234 7200
rect 15212 7188 15240 7228
rect 13228 7160 15240 7188
rect 17880 7188 17908 7228
rect 18984 7228 19564 7256
rect 18984 7188 19012 7228
rect 19536 7200 19564 7228
rect 17880 7160 19012 7188
rect 13228 7148 13234 7160
rect 19518 7148 19524 7200
rect 19576 7148 19582 7200
rect 1104 7098 21896 7120
rect 1104 7046 3549 7098
rect 3601 7046 3613 7098
rect 3665 7046 3677 7098
rect 3729 7046 3741 7098
rect 3793 7046 3805 7098
rect 3857 7046 8747 7098
rect 8799 7046 8811 7098
rect 8863 7046 8875 7098
rect 8927 7046 8939 7098
rect 8991 7046 9003 7098
rect 9055 7046 13945 7098
rect 13997 7046 14009 7098
rect 14061 7046 14073 7098
rect 14125 7046 14137 7098
rect 14189 7046 14201 7098
rect 14253 7046 19143 7098
rect 19195 7046 19207 7098
rect 19259 7046 19271 7098
rect 19323 7046 19335 7098
rect 19387 7046 19399 7098
rect 19451 7046 21896 7098
rect 1104 7024 21896 7046
rect 4246 6984 4252 6996
rect 3896 6956 4252 6984
rect 2225 6851 2283 6857
rect 2225 6817 2237 6851
rect 2271 6848 2283 6851
rect 2314 6848 2320 6860
rect 2271 6820 2320 6848
rect 2271 6817 2283 6820
rect 2225 6811 2283 6817
rect 2314 6808 2320 6820
rect 2372 6808 2378 6860
rect 3896 6857 3924 6956
rect 4246 6944 4252 6956
rect 4304 6944 4310 6996
rect 4982 6944 4988 6996
rect 5040 6984 5046 6996
rect 5169 6987 5227 6993
rect 5169 6984 5181 6987
rect 5040 6956 5181 6984
rect 5040 6944 5046 6956
rect 5169 6953 5181 6956
rect 5215 6953 5227 6987
rect 8386 6984 8392 6996
rect 5169 6947 5227 6953
rect 5552 6956 8392 6984
rect 3970 6876 3976 6928
rect 4028 6916 4034 6928
rect 5552 6916 5580 6956
rect 8386 6944 8392 6956
rect 8444 6984 8450 6996
rect 8481 6987 8539 6993
rect 8481 6984 8493 6987
rect 8444 6956 8493 6984
rect 8444 6944 8450 6956
rect 8481 6953 8493 6956
rect 8527 6953 8539 6987
rect 8481 6947 8539 6953
rect 8570 6944 8576 6996
rect 8628 6984 8634 6996
rect 8941 6987 8999 6993
rect 8941 6984 8953 6987
rect 8628 6956 8953 6984
rect 8628 6944 8634 6956
rect 8941 6953 8953 6956
rect 8987 6953 8999 6987
rect 13170 6984 13176 6996
rect 8941 6947 8999 6953
rect 9048 6956 13176 6984
rect 4028 6888 5580 6916
rect 4028 6876 4034 6888
rect 5626 6876 5632 6928
rect 5684 6916 5690 6928
rect 9048 6916 9076 6956
rect 13170 6944 13176 6956
rect 13228 6944 13234 6996
rect 13354 6984 13360 6996
rect 13315 6956 13360 6984
rect 13354 6944 13360 6956
rect 13412 6944 13418 6996
rect 13722 6984 13728 6996
rect 13683 6956 13728 6984
rect 13722 6944 13728 6956
rect 13780 6944 13786 6996
rect 15746 6944 15752 6996
rect 15804 6984 15810 6996
rect 16301 6987 16359 6993
rect 16301 6984 16313 6987
rect 15804 6956 16313 6984
rect 15804 6944 15810 6956
rect 5684 6888 9076 6916
rect 5684 6876 5690 6888
rect 3881 6851 3939 6857
rect 3881 6817 3893 6851
rect 3927 6817 3939 6851
rect 3881 6811 3939 6817
rect 4065 6851 4123 6857
rect 4065 6817 4077 6851
rect 4111 6848 4123 6851
rect 4154 6848 4160 6860
rect 4111 6820 4160 6848
rect 4111 6817 4123 6820
rect 4065 6811 4123 6817
rect 4154 6808 4160 6820
rect 4212 6808 4218 6860
rect 5166 6808 5172 6860
rect 5224 6848 5230 6860
rect 5828 6857 5856 6888
rect 5813 6851 5871 6857
rect 5224 6820 5764 6848
rect 5224 6808 5230 6820
rect 3421 6783 3479 6789
rect 3421 6749 3433 6783
rect 3467 6780 3479 6783
rect 4338 6780 4344 6792
rect 3467 6752 4344 6780
rect 3467 6749 3479 6752
rect 3421 6743 3479 6749
rect 4338 6740 4344 6752
rect 4396 6780 4402 6792
rect 5258 6780 5264 6792
rect 4396 6752 5264 6780
rect 4396 6740 4402 6752
rect 5258 6740 5264 6752
rect 5316 6780 5322 6792
rect 5537 6783 5595 6789
rect 5537 6780 5549 6783
rect 5316 6752 5549 6780
rect 5316 6740 5322 6752
rect 5537 6749 5549 6752
rect 5583 6749 5595 6783
rect 5736 6780 5764 6820
rect 5813 6817 5825 6851
rect 5859 6817 5871 6851
rect 5813 6811 5871 6817
rect 5994 6808 6000 6860
rect 6052 6848 6058 6860
rect 6825 6851 6883 6857
rect 6825 6848 6837 6851
rect 6052 6820 6837 6848
rect 6052 6808 6058 6820
rect 6825 6817 6837 6820
rect 6871 6848 6883 6851
rect 9122 6848 9128 6860
rect 6871 6820 9128 6848
rect 6871 6817 6883 6820
rect 6825 6811 6883 6817
rect 9122 6808 9128 6820
rect 9180 6808 9186 6860
rect 9582 6848 9588 6860
rect 9543 6820 9588 6848
rect 9582 6808 9588 6820
rect 9640 6808 9646 6860
rect 16040 6857 16068 6956
rect 16301 6953 16313 6956
rect 16347 6953 16359 6987
rect 16301 6947 16359 6953
rect 18322 6944 18328 6996
rect 18380 6984 18386 6996
rect 18417 6987 18475 6993
rect 18417 6984 18429 6987
rect 18380 6956 18429 6984
rect 18380 6944 18386 6956
rect 18417 6953 18429 6956
rect 18463 6984 18475 6987
rect 19245 6987 19303 6993
rect 19245 6984 19257 6987
rect 18463 6956 19257 6984
rect 18463 6953 18475 6956
rect 18417 6947 18475 6953
rect 19245 6953 19257 6956
rect 19291 6953 19303 6987
rect 19245 6947 19303 6953
rect 19518 6944 19524 6996
rect 19576 6984 19582 6996
rect 19613 6987 19671 6993
rect 19613 6984 19625 6987
rect 19576 6956 19625 6984
rect 19576 6944 19582 6956
rect 19613 6953 19625 6956
rect 19659 6953 19671 6987
rect 19613 6947 19671 6953
rect 21082 6944 21088 6996
rect 21140 6984 21146 6996
rect 21269 6987 21327 6993
rect 21269 6984 21281 6987
rect 21140 6956 21281 6984
rect 21140 6944 21146 6956
rect 21269 6953 21281 6956
rect 21315 6953 21327 6987
rect 21269 6947 21327 6953
rect 16025 6851 16083 6857
rect 16025 6817 16037 6851
rect 16071 6817 16083 6851
rect 16025 6811 16083 6817
rect 18141 6851 18199 6857
rect 18141 6817 18153 6851
rect 18187 6848 18199 6851
rect 18340 6848 18368 6944
rect 18187 6820 18368 6848
rect 20993 6851 21051 6857
rect 18187 6817 18199 6820
rect 18141 6811 18199 6817
rect 20993 6817 21005 6851
rect 21039 6848 21051 6851
rect 21100 6848 21128 6944
rect 21039 6820 21128 6848
rect 21039 6817 21051 6820
rect 20993 6811 21051 6817
rect 7742 6780 7748 6792
rect 5736 6752 7604 6780
rect 7703 6752 7748 6780
rect 5537 6743 5595 6749
rect 4157 6715 4215 6721
rect 4157 6712 4169 6715
rect 2792 6684 4169 6712
rect 1670 6644 1676 6656
rect 1631 6616 1676 6644
rect 1670 6604 1676 6616
rect 1728 6644 1734 6656
rect 2317 6647 2375 6653
rect 2317 6644 2329 6647
rect 1728 6616 2329 6644
rect 1728 6604 1734 6616
rect 2317 6613 2329 6616
rect 2363 6613 2375 6647
rect 2317 6607 2375 6613
rect 2409 6647 2467 6653
rect 2409 6613 2421 6647
rect 2455 6644 2467 6647
rect 2498 6644 2504 6656
rect 2455 6616 2504 6644
rect 2455 6613 2467 6616
rect 2409 6607 2467 6613
rect 2498 6604 2504 6616
rect 2556 6604 2562 6656
rect 2792 6653 2820 6684
rect 4157 6681 4169 6684
rect 4203 6681 4215 6715
rect 4157 6675 4215 6681
rect 6641 6715 6699 6721
rect 6641 6681 6653 6715
rect 6687 6712 6699 6715
rect 7466 6712 7472 6724
rect 6687 6684 7052 6712
rect 7427 6684 7472 6712
rect 6687 6681 6699 6684
rect 6641 6675 6699 6681
rect 2777 6647 2835 6653
rect 2777 6613 2789 6647
rect 2823 6613 2835 6647
rect 4522 6644 4528 6656
rect 4483 6616 4528 6644
rect 2777 6607 2835 6613
rect 4522 6604 4528 6616
rect 4580 6604 4586 6656
rect 4893 6647 4951 6653
rect 4893 6613 4905 6647
rect 4939 6644 4951 6647
rect 5166 6644 5172 6656
rect 4939 6616 5172 6644
rect 4939 6613 4951 6616
rect 4893 6607 4951 6613
rect 5166 6604 5172 6616
rect 5224 6644 5230 6656
rect 5629 6647 5687 6653
rect 5629 6644 5641 6647
rect 5224 6616 5641 6644
rect 5224 6604 5230 6616
rect 5629 6613 5641 6616
rect 5675 6613 5687 6647
rect 5629 6607 5687 6613
rect 5718 6604 5724 6656
rect 5776 6644 5782 6656
rect 6273 6647 6331 6653
rect 6273 6644 6285 6647
rect 5776 6616 6285 6644
rect 5776 6604 5782 6616
rect 6273 6613 6285 6616
rect 6319 6613 6331 6647
rect 6273 6607 6331 6613
rect 6730 6604 6736 6656
rect 6788 6644 6794 6656
rect 7024 6644 7052 6684
rect 7466 6672 7472 6684
rect 7524 6672 7530 6724
rect 7576 6712 7604 6752
rect 7742 6740 7748 6752
rect 7800 6740 7806 6792
rect 11977 6783 12035 6789
rect 8496 6752 10088 6780
rect 8496 6712 8524 6752
rect 7576 6684 8524 6712
rect 9309 6715 9367 6721
rect 9309 6681 9321 6715
rect 9355 6712 9367 6715
rect 9953 6715 10011 6721
rect 9953 6712 9965 6715
rect 9355 6684 9965 6712
rect 9355 6681 9367 6684
rect 9309 6675 9367 6681
rect 9953 6681 9965 6684
rect 9999 6681 10011 6715
rect 10060 6712 10088 6752
rect 11977 6749 11989 6783
rect 12023 6780 12035 6783
rect 13722 6780 13728 6792
rect 12023 6752 13728 6780
rect 12023 6749 12035 6752
rect 11977 6743 12035 6749
rect 13722 6740 13728 6752
rect 13780 6740 13786 6792
rect 15470 6740 15476 6792
rect 15528 6780 15534 6792
rect 15769 6783 15827 6789
rect 15769 6780 15781 6783
rect 15528 6752 15781 6780
rect 15528 6740 15534 6752
rect 15769 6749 15781 6752
rect 15815 6780 15827 6783
rect 18230 6780 18236 6792
rect 15815 6752 18236 6780
rect 15815 6749 15827 6752
rect 15769 6743 15827 6749
rect 18230 6740 18236 6752
rect 18288 6740 18294 6792
rect 19794 6740 19800 6792
rect 19852 6780 19858 6792
rect 20726 6783 20784 6789
rect 20726 6780 20738 6783
rect 19852 6752 20738 6780
rect 19852 6740 19858 6752
rect 20726 6749 20738 6752
rect 20772 6749 20784 6783
rect 20726 6743 20784 6749
rect 11146 6712 11152 6724
rect 10060 6684 11152 6712
rect 9953 6675 10011 6681
rect 11146 6672 11152 6684
rect 11204 6712 11210 6724
rect 12222 6715 12280 6721
rect 12222 6712 12234 6715
rect 11204 6684 12234 6712
rect 11204 6672 11210 6684
rect 12222 6681 12234 6684
rect 12268 6681 12280 6715
rect 12222 6675 12280 6681
rect 12434 6672 12440 6724
rect 12492 6712 12498 6724
rect 12492 6684 14872 6712
rect 12492 6672 12498 6684
rect 8021 6647 8079 6653
rect 8021 6644 8033 6647
rect 6788 6616 6833 6644
rect 7024 6616 8033 6644
rect 6788 6604 6794 6616
rect 8021 6613 8033 6616
rect 8067 6613 8079 6647
rect 8021 6607 8079 6613
rect 9030 6604 9036 6656
rect 9088 6644 9094 6656
rect 9401 6647 9459 6653
rect 9401 6644 9413 6647
rect 9088 6616 9413 6644
rect 9088 6604 9094 6616
rect 9401 6613 9413 6616
rect 9447 6613 9459 6647
rect 9401 6607 9459 6613
rect 10318 6604 10324 6656
rect 10376 6644 10382 6656
rect 12342 6644 12348 6656
rect 10376 6616 12348 6644
rect 10376 6604 10382 6616
rect 12342 6604 12348 6616
rect 12400 6604 12406 6656
rect 14274 6604 14280 6656
rect 14332 6644 14338 6656
rect 14645 6647 14703 6653
rect 14645 6644 14657 6647
rect 14332 6616 14657 6644
rect 14332 6604 14338 6616
rect 14645 6613 14657 6616
rect 14691 6613 14703 6647
rect 14844 6644 14872 6684
rect 17770 6672 17776 6724
rect 17828 6712 17834 6724
rect 17874 6715 17932 6721
rect 17874 6712 17886 6715
rect 17828 6684 17886 6712
rect 17828 6672 17834 6684
rect 17874 6681 17886 6684
rect 17920 6681 17932 6715
rect 17874 6675 17932 6681
rect 15378 6644 15384 6656
rect 14844 6616 15384 6644
rect 14645 6607 14703 6613
rect 15378 6604 15384 6616
rect 15436 6644 15442 6656
rect 16761 6647 16819 6653
rect 16761 6644 16773 6647
rect 15436 6616 16773 6644
rect 15436 6604 15442 6616
rect 16761 6613 16773 6616
rect 16807 6613 16819 6647
rect 16761 6607 16819 6613
rect 16942 6604 16948 6656
rect 17000 6644 17006 6656
rect 19702 6644 19708 6656
rect 17000 6616 19708 6644
rect 17000 6604 17006 6616
rect 19702 6604 19708 6616
rect 19760 6604 19766 6656
rect 1104 6554 22056 6576
rect 1104 6502 6148 6554
rect 6200 6502 6212 6554
rect 6264 6502 6276 6554
rect 6328 6502 6340 6554
rect 6392 6502 6404 6554
rect 6456 6502 11346 6554
rect 11398 6502 11410 6554
rect 11462 6502 11474 6554
rect 11526 6502 11538 6554
rect 11590 6502 11602 6554
rect 11654 6502 16544 6554
rect 16596 6502 16608 6554
rect 16660 6502 16672 6554
rect 16724 6502 16736 6554
rect 16788 6502 16800 6554
rect 16852 6502 21742 6554
rect 21794 6502 21806 6554
rect 21858 6502 21870 6554
rect 21922 6502 21934 6554
rect 21986 6502 21998 6554
rect 22050 6502 22056 6554
rect 1104 6480 22056 6502
rect 2498 6440 2504 6452
rect 2459 6412 2504 6440
rect 2498 6400 2504 6412
rect 2556 6400 2562 6452
rect 5629 6443 5687 6449
rect 5629 6409 5641 6443
rect 5675 6440 5687 6443
rect 5718 6440 5724 6452
rect 5675 6412 5724 6440
rect 5675 6409 5687 6412
rect 5629 6403 5687 6409
rect 5718 6400 5724 6412
rect 5776 6400 5782 6452
rect 6730 6440 6736 6452
rect 6691 6412 6736 6440
rect 6730 6400 6736 6412
rect 6788 6400 6794 6452
rect 8386 6400 8392 6452
rect 8444 6440 8450 6452
rect 8665 6443 8723 6449
rect 8665 6440 8677 6443
rect 8444 6412 8677 6440
rect 8444 6400 8450 6412
rect 8665 6409 8677 6412
rect 8711 6409 8723 6443
rect 9030 6440 9036 6452
rect 8991 6412 9036 6440
rect 8665 6403 8723 6409
rect 9030 6400 9036 6412
rect 9088 6400 9094 6452
rect 9122 6400 9128 6452
rect 9180 6440 9186 6452
rect 15473 6443 15531 6449
rect 9180 6412 15424 6440
rect 9180 6400 9186 6412
rect 5258 6332 5264 6384
rect 5316 6372 5322 6384
rect 6365 6375 6423 6381
rect 6365 6372 6377 6375
rect 5316 6344 6377 6372
rect 5316 6332 5322 6344
rect 6365 6341 6377 6344
rect 6411 6341 6423 6375
rect 6365 6335 6423 6341
rect 4522 6304 4528 6316
rect 4483 6276 4528 6304
rect 4522 6264 4528 6276
rect 4580 6264 4586 6316
rect 5534 6264 5540 6316
rect 5592 6304 5598 6316
rect 6270 6304 6276 6316
rect 5592 6276 6276 6304
rect 5592 6264 5598 6276
rect 6270 6264 6276 6276
rect 6328 6264 6334 6316
rect 1762 6196 1768 6248
rect 1820 6236 1826 6248
rect 2961 6239 3019 6245
rect 2961 6236 2973 6239
rect 1820 6208 2973 6236
rect 1820 6196 1826 6208
rect 2961 6205 2973 6208
rect 3007 6205 3019 6239
rect 2961 6199 3019 6205
rect 4614 6196 4620 6248
rect 4672 6236 4678 6248
rect 4709 6239 4767 6245
rect 4709 6236 4721 6239
rect 4672 6208 4721 6236
rect 4672 6196 4678 6208
rect 4709 6205 4721 6208
rect 4755 6205 4767 6239
rect 4709 6199 4767 6205
rect 5258 6196 5264 6248
rect 5316 6236 5322 6248
rect 5721 6239 5779 6245
rect 5721 6236 5733 6239
rect 5316 6208 5733 6236
rect 5316 6196 5322 6208
rect 5721 6205 5733 6208
rect 5767 6205 5779 6239
rect 5902 6236 5908 6248
rect 5863 6208 5908 6236
rect 5721 6199 5779 6205
rect 5902 6196 5908 6208
rect 5960 6196 5966 6248
rect 6380 6236 6408 6335
rect 6546 6332 6552 6384
rect 6604 6372 6610 6384
rect 10318 6372 10324 6384
rect 6604 6344 10324 6372
rect 6604 6332 6610 6344
rect 10318 6332 10324 6344
rect 10376 6332 10382 6384
rect 15396 6372 15424 6412
rect 15473 6409 15485 6443
rect 15519 6440 15531 6443
rect 15746 6440 15752 6452
rect 15519 6412 15752 6440
rect 15519 6409 15531 6412
rect 15473 6403 15531 6409
rect 15746 6400 15752 6412
rect 15804 6400 15810 6452
rect 18049 6443 18107 6449
rect 18049 6409 18061 6443
rect 18095 6409 18107 6443
rect 18322 6440 18328 6452
rect 18283 6412 18328 6440
rect 18049 6403 18107 6409
rect 18064 6372 18092 6403
rect 18322 6400 18328 6412
rect 18380 6440 18386 6452
rect 19061 6443 19119 6449
rect 19061 6440 19073 6443
rect 18380 6412 19073 6440
rect 18380 6400 18386 6412
rect 19061 6409 19073 6412
rect 19107 6409 19119 6443
rect 19061 6403 19119 6409
rect 12176 6344 15056 6372
rect 15396 6344 18092 6372
rect 6454 6264 6460 6316
rect 6512 6304 6518 6316
rect 7101 6307 7159 6313
rect 7101 6304 7113 6307
rect 6512 6276 7113 6304
rect 6512 6264 6518 6276
rect 7101 6273 7113 6276
rect 7147 6273 7159 6307
rect 10042 6304 10048 6316
rect 7101 6267 7159 6273
rect 7392 6276 10048 6304
rect 7193 6239 7251 6245
rect 7193 6236 7205 6239
rect 6380 6208 7205 6236
rect 7193 6205 7205 6208
rect 7239 6236 7251 6239
rect 7282 6236 7288 6248
rect 7239 6208 7288 6236
rect 7239 6205 7251 6208
rect 7193 6199 7251 6205
rect 7282 6196 7288 6208
rect 7340 6196 7346 6248
rect 7392 6245 7420 6276
rect 10042 6264 10048 6276
rect 10100 6304 10106 6316
rect 12176 6304 12204 6344
rect 12998 6307 13056 6313
rect 12998 6304 13010 6307
rect 10100 6276 12204 6304
rect 12268 6276 13010 6304
rect 10100 6264 10106 6276
rect 7377 6239 7435 6245
rect 7377 6205 7389 6239
rect 7423 6205 7435 6239
rect 7377 6199 7435 6205
rect 8481 6239 8539 6245
rect 8481 6205 8493 6239
rect 8527 6205 8539 6239
rect 8481 6199 8539 6205
rect 8573 6239 8631 6245
rect 8573 6205 8585 6239
rect 8619 6236 8631 6239
rect 8662 6236 8668 6248
rect 8619 6208 8668 6236
rect 8619 6205 8631 6208
rect 8573 6199 8631 6205
rect 4249 6171 4307 6177
rect 4249 6137 4261 6171
rect 4295 6168 4307 6171
rect 5920 6168 5948 6196
rect 7392 6168 7420 6199
rect 4295 6140 5948 6168
rect 6012 6140 7420 6168
rect 8496 6168 8524 6199
rect 8662 6196 8668 6208
rect 8720 6196 8726 6248
rect 9306 6236 9312 6248
rect 9267 6208 9312 6236
rect 9306 6196 9312 6208
rect 9364 6196 9370 6248
rect 11790 6196 11796 6248
rect 11848 6236 11854 6248
rect 12268 6236 12296 6276
rect 12998 6273 13010 6276
rect 13044 6273 13056 6307
rect 12998 6267 13056 6273
rect 13265 6307 13323 6313
rect 13265 6273 13277 6307
rect 13311 6304 13323 6307
rect 13722 6304 13728 6316
rect 13311 6276 13728 6304
rect 13311 6273 13323 6276
rect 13265 6267 13323 6273
rect 13722 6264 13728 6276
rect 13780 6264 13786 6316
rect 14274 6264 14280 6316
rect 14332 6304 14338 6316
rect 14838 6307 14896 6313
rect 14838 6304 14850 6307
rect 14332 6276 14850 6304
rect 14332 6264 14338 6276
rect 14838 6273 14850 6276
rect 14884 6273 14896 6307
rect 14838 6267 14896 6273
rect 11848 6208 12296 6236
rect 15028 6236 15056 6344
rect 15105 6307 15163 6313
rect 15105 6273 15117 6307
rect 15151 6304 15163 6307
rect 15746 6304 15752 6316
rect 15151 6276 15752 6304
rect 15151 6273 15163 6276
rect 15105 6267 15163 6273
rect 15746 6264 15752 6276
rect 15804 6304 15810 6316
rect 16669 6307 16727 6313
rect 16669 6304 16681 6307
rect 15804 6276 16681 6304
rect 15804 6264 15810 6276
rect 16669 6273 16681 6276
rect 16715 6273 16727 6307
rect 16925 6307 16983 6313
rect 16925 6304 16937 6307
rect 16669 6267 16727 6273
rect 16776 6276 16937 6304
rect 16776 6236 16804 6276
rect 16925 6273 16937 6276
rect 16971 6273 16983 6307
rect 16925 6267 16983 6273
rect 15028 6208 16804 6236
rect 18064 6236 18092 6344
rect 19076 6304 19104 6403
rect 19150 6400 19156 6452
rect 19208 6440 19214 6452
rect 20809 6443 20867 6449
rect 20809 6440 20821 6443
rect 19208 6412 20821 6440
rect 19208 6400 19214 6412
rect 20809 6409 20821 6412
rect 20855 6409 20867 6443
rect 21082 6440 21088 6452
rect 21043 6412 21088 6440
rect 20809 6403 20867 6409
rect 21082 6400 21088 6412
rect 21140 6400 21146 6452
rect 19429 6307 19487 6313
rect 19429 6304 19441 6307
rect 19076 6276 19441 6304
rect 19429 6273 19441 6276
rect 19475 6273 19487 6307
rect 19429 6267 19487 6273
rect 19518 6264 19524 6316
rect 19576 6264 19582 6316
rect 19702 6313 19708 6316
rect 19696 6304 19708 6313
rect 19663 6276 19708 6304
rect 19696 6267 19708 6276
rect 19702 6264 19708 6267
rect 19760 6264 19766 6316
rect 19536 6236 19564 6264
rect 18064 6208 19564 6236
rect 11848 6196 11854 6208
rect 8496 6140 12020 6168
rect 4295 6137 4307 6140
rect 4249 6131 4307 6137
rect 5074 6060 5080 6112
rect 5132 6100 5138 6112
rect 5261 6103 5319 6109
rect 5261 6100 5273 6103
rect 5132 6072 5273 6100
rect 5132 6060 5138 6072
rect 5261 6069 5273 6072
rect 5307 6069 5319 6103
rect 5261 6063 5319 6069
rect 5626 6060 5632 6112
rect 5684 6100 5690 6112
rect 6012 6100 6040 6140
rect 5684 6072 6040 6100
rect 5684 6060 5690 6072
rect 7006 6060 7012 6112
rect 7064 6100 7070 6112
rect 8021 6103 8079 6109
rect 8021 6100 8033 6103
rect 7064 6072 8033 6100
rect 7064 6060 7070 6072
rect 8021 6069 8033 6072
rect 8067 6100 8079 6103
rect 8662 6100 8668 6112
rect 8067 6072 8668 6100
rect 8067 6069 8079 6072
rect 8021 6063 8079 6069
rect 8662 6060 8668 6072
rect 8720 6060 8726 6112
rect 11882 6100 11888 6112
rect 11843 6072 11888 6100
rect 11882 6060 11888 6072
rect 11940 6060 11946 6112
rect 11992 6100 12020 6140
rect 13725 6103 13783 6109
rect 13725 6100 13737 6103
rect 11992 6072 13737 6100
rect 13725 6069 13737 6072
rect 13771 6100 13783 6103
rect 14734 6100 14740 6112
rect 13771 6072 14740 6100
rect 13771 6069 13783 6072
rect 13725 6063 13783 6069
rect 14734 6060 14740 6072
rect 14792 6060 14798 6112
rect 1104 6010 21896 6032
rect 1104 5958 3549 6010
rect 3601 5958 3613 6010
rect 3665 5958 3677 6010
rect 3729 5958 3741 6010
rect 3793 5958 3805 6010
rect 3857 5958 8747 6010
rect 8799 5958 8811 6010
rect 8863 5958 8875 6010
rect 8927 5958 8939 6010
rect 8991 5958 9003 6010
rect 9055 5958 13945 6010
rect 13997 5958 14009 6010
rect 14061 5958 14073 6010
rect 14125 5958 14137 6010
rect 14189 5958 14201 6010
rect 14253 5958 19143 6010
rect 19195 5958 19207 6010
rect 19259 5958 19271 6010
rect 19323 5958 19335 6010
rect 19387 5958 19399 6010
rect 19451 5958 21896 6010
rect 1104 5936 21896 5958
rect 3326 5856 3332 5908
rect 3384 5896 3390 5908
rect 3789 5899 3847 5905
rect 3789 5896 3801 5899
rect 3384 5868 3801 5896
rect 3384 5856 3390 5868
rect 3789 5865 3801 5868
rect 3835 5865 3847 5899
rect 5258 5896 5264 5908
rect 5219 5868 5264 5896
rect 3789 5859 3847 5865
rect 2498 5788 2504 5840
rect 2556 5828 2562 5840
rect 2958 5828 2964 5840
rect 2556 5800 2964 5828
rect 2556 5788 2562 5800
rect 2958 5788 2964 5800
rect 3016 5828 3022 5840
rect 3804 5828 3832 5859
rect 5258 5856 5264 5868
rect 5316 5856 5322 5908
rect 5902 5856 5908 5908
rect 5960 5896 5966 5908
rect 5960 5868 9536 5896
rect 5960 5856 5966 5868
rect 6914 5828 6920 5840
rect 3016 5800 3740 5828
rect 3804 5800 6316 5828
rect 6875 5800 6920 5828
rect 3016 5788 3022 5800
rect 1581 5763 1639 5769
rect 1581 5729 1593 5763
rect 1627 5760 1639 5763
rect 3053 5763 3111 5769
rect 3053 5760 3065 5763
rect 1627 5732 3065 5760
rect 1627 5729 1639 5732
rect 1581 5723 1639 5729
rect 3053 5729 3065 5732
rect 3099 5729 3111 5763
rect 3712 5760 3740 5800
rect 4157 5763 4215 5769
rect 4157 5760 4169 5763
rect 3712 5732 4169 5760
rect 3053 5723 3111 5729
rect 4157 5729 4169 5732
rect 4203 5760 4215 5763
rect 4522 5760 4528 5772
rect 4203 5732 4528 5760
rect 4203 5729 4215 5732
rect 4157 5723 4215 5729
rect 1670 5692 1676 5704
rect 1631 5664 1676 5692
rect 1670 5652 1676 5664
rect 1728 5652 1734 5704
rect 1762 5652 1768 5704
rect 1820 5692 1826 5704
rect 3068 5692 3096 5723
rect 4522 5720 4528 5732
rect 4580 5720 4586 5772
rect 4709 5763 4767 5769
rect 4709 5729 4721 5763
rect 4755 5760 4767 5763
rect 5994 5760 6000 5772
rect 4755 5732 6000 5760
rect 4755 5729 4767 5732
rect 4709 5723 4767 5729
rect 5994 5720 6000 5732
rect 6052 5720 6058 5772
rect 6089 5763 6147 5769
rect 6089 5729 6101 5763
rect 6135 5729 6147 5763
rect 6089 5723 6147 5729
rect 5902 5692 5908 5704
rect 1820 5664 1865 5692
rect 3068 5664 5908 5692
rect 1820 5652 1826 5664
rect 5902 5652 5908 5664
rect 5960 5652 5966 5704
rect 2777 5627 2835 5633
rect 2777 5593 2789 5627
rect 2823 5624 2835 5627
rect 3234 5624 3240 5636
rect 2823 5596 3240 5624
rect 2823 5593 2835 5596
rect 2777 5587 2835 5593
rect 3234 5584 3240 5596
rect 3292 5584 3298 5636
rect 4522 5584 4528 5636
rect 4580 5624 4586 5636
rect 6104 5624 6132 5723
rect 6288 5701 6316 5800
rect 6914 5788 6920 5800
rect 6972 5788 6978 5840
rect 8021 5831 8079 5837
rect 8021 5797 8033 5831
rect 8067 5828 8079 5831
rect 9508 5828 9536 5868
rect 9582 5856 9588 5908
rect 9640 5896 9646 5908
rect 9640 5868 13400 5896
rect 9640 5856 9646 5868
rect 8067 5800 9444 5828
rect 9508 5800 9720 5828
rect 8067 5797 8079 5800
rect 8021 5791 8079 5797
rect 7469 5763 7527 5769
rect 7469 5729 7481 5763
rect 7515 5760 7527 5763
rect 8294 5760 8300 5772
rect 7515 5732 8300 5760
rect 7515 5729 7527 5732
rect 7469 5723 7527 5729
rect 8294 5720 8300 5732
rect 8352 5720 8358 5772
rect 9416 5769 9444 5800
rect 9401 5763 9459 5769
rect 9401 5729 9413 5763
rect 9447 5729 9459 5763
rect 9582 5760 9588 5772
rect 9543 5732 9588 5760
rect 9401 5723 9459 5729
rect 9582 5720 9588 5732
rect 9640 5720 9646 5772
rect 6273 5695 6331 5701
rect 6273 5661 6285 5695
rect 6319 5661 6331 5695
rect 6273 5655 6331 5661
rect 7282 5652 7288 5704
rect 7340 5692 7346 5704
rect 7558 5692 7564 5704
rect 7340 5664 7564 5692
rect 7340 5652 7346 5664
rect 7558 5652 7564 5664
rect 7616 5652 7622 5704
rect 7650 5652 7656 5704
rect 7708 5692 7714 5704
rect 9306 5692 9312 5704
rect 7708 5664 7753 5692
rect 9267 5664 9312 5692
rect 7708 5652 7714 5664
rect 9306 5652 9312 5664
rect 9364 5652 9370 5704
rect 9692 5692 9720 5800
rect 11146 5788 11152 5840
rect 11204 5828 11210 5840
rect 11425 5831 11483 5837
rect 11425 5828 11437 5831
rect 11204 5800 11437 5828
rect 11204 5788 11210 5800
rect 11425 5797 11437 5800
rect 11471 5797 11483 5831
rect 13372 5828 13400 5868
rect 13446 5856 13452 5908
rect 13504 5896 13510 5908
rect 13722 5896 13728 5908
rect 13504 5868 13728 5896
rect 13504 5856 13510 5868
rect 13722 5856 13728 5868
rect 13780 5856 13786 5908
rect 15746 5896 15752 5908
rect 14568 5868 15608 5896
rect 15707 5868 15752 5896
rect 14568 5828 14596 5868
rect 13372 5800 14596 5828
rect 15580 5828 15608 5868
rect 15746 5856 15752 5868
rect 15804 5856 15810 5908
rect 17052 5868 18000 5896
rect 17052 5828 17080 5868
rect 15580 5800 17080 5828
rect 17972 5828 18000 5868
rect 18322 5856 18328 5908
rect 18380 5896 18386 5908
rect 18693 5899 18751 5905
rect 18693 5896 18705 5899
rect 18380 5868 18705 5896
rect 18380 5856 18386 5868
rect 18693 5865 18705 5868
rect 18739 5865 18751 5899
rect 18693 5859 18751 5865
rect 19337 5899 19395 5905
rect 19337 5865 19349 5899
rect 19383 5896 19395 5899
rect 19794 5896 19800 5908
rect 19383 5868 19800 5896
rect 19383 5865 19395 5868
rect 19337 5859 19395 5865
rect 19794 5856 19800 5868
rect 19852 5856 19858 5908
rect 21082 5896 21088 5908
rect 21043 5868 21088 5896
rect 21082 5856 21088 5868
rect 21140 5856 21146 5908
rect 18417 5831 18475 5837
rect 18417 5828 18429 5831
rect 17972 5800 18429 5828
rect 11425 5791 11483 5797
rect 18417 5797 18429 5800
rect 18463 5828 18475 5831
rect 19702 5828 19708 5840
rect 18463 5800 19708 5828
rect 18463 5797 18475 5800
rect 18417 5791 18475 5797
rect 19702 5788 19708 5800
rect 19760 5788 19766 5840
rect 12805 5763 12863 5769
rect 12805 5729 12817 5763
rect 12851 5760 12863 5763
rect 13446 5760 13452 5772
rect 12851 5732 13452 5760
rect 12851 5729 12863 5732
rect 12805 5723 12863 5729
rect 13446 5720 13452 5732
rect 13504 5720 13510 5772
rect 15473 5763 15531 5769
rect 13740 5732 14504 5760
rect 12250 5692 12256 5704
rect 9692 5664 12256 5692
rect 12250 5652 12256 5664
rect 12308 5652 12314 5704
rect 13740 5692 13768 5732
rect 12406 5664 13768 5692
rect 12406 5624 12434 5664
rect 4580 5596 5672 5624
rect 6104 5596 12434 5624
rect 12560 5627 12618 5633
rect 4580 5584 4586 5596
rect 2130 5556 2136 5568
rect 2091 5528 2136 5556
rect 2130 5516 2136 5528
rect 2188 5516 2194 5568
rect 2406 5556 2412 5568
rect 2367 5528 2412 5556
rect 2406 5516 2412 5528
rect 2464 5516 2470 5568
rect 2866 5516 2872 5568
rect 2924 5556 2930 5568
rect 4798 5556 4804 5568
rect 2924 5528 2969 5556
rect 4759 5528 4804 5556
rect 2924 5516 2930 5528
rect 4798 5516 4804 5528
rect 4856 5516 4862 5568
rect 4893 5559 4951 5565
rect 4893 5525 4905 5559
rect 4939 5556 4951 5559
rect 5166 5556 5172 5568
rect 4939 5528 5172 5556
rect 4939 5525 4951 5528
rect 4893 5519 4951 5525
rect 5166 5516 5172 5528
rect 5224 5516 5230 5568
rect 5534 5556 5540 5568
rect 5495 5528 5540 5556
rect 5534 5516 5540 5528
rect 5592 5516 5598 5568
rect 5644 5556 5672 5596
rect 12560 5593 12572 5627
rect 12606 5624 12618 5627
rect 14366 5624 14372 5636
rect 12606 5596 14372 5624
rect 12606 5593 12618 5596
rect 12560 5587 12618 5593
rect 14366 5584 14372 5596
rect 14424 5584 14430 5636
rect 14476 5624 14504 5732
rect 15473 5729 15485 5763
rect 15519 5760 15531 5763
rect 15746 5760 15752 5772
rect 15519 5732 15752 5760
rect 15519 5729 15531 5732
rect 15473 5723 15531 5729
rect 15746 5720 15752 5732
rect 15804 5760 15810 5772
rect 17037 5763 17095 5769
rect 17037 5760 17049 5763
rect 15804 5732 17049 5760
rect 15804 5720 15810 5732
rect 17037 5729 17049 5732
rect 17083 5729 17095 5763
rect 17037 5723 17095 5729
rect 20717 5763 20775 5769
rect 20717 5729 20729 5763
rect 20763 5760 20775 5763
rect 21100 5760 21128 5856
rect 20763 5732 21128 5760
rect 20763 5729 20775 5732
rect 20717 5723 20775 5729
rect 14734 5652 14740 5704
rect 14792 5692 14798 5704
rect 17293 5695 17351 5701
rect 17293 5692 17305 5695
rect 14792 5664 17305 5692
rect 14792 5652 14798 5664
rect 17293 5661 17305 5664
rect 17339 5661 17351 5695
rect 17293 5655 17351 5661
rect 19058 5652 19064 5704
rect 19116 5692 19122 5704
rect 20450 5695 20508 5701
rect 20450 5692 20462 5695
rect 19116 5664 20462 5692
rect 19116 5652 19122 5664
rect 20450 5661 20462 5664
rect 20496 5661 20508 5695
rect 20450 5655 20508 5661
rect 15228 5627 15286 5633
rect 15228 5624 15240 5627
rect 14476 5596 15240 5624
rect 15228 5593 15240 5596
rect 15274 5624 15286 5627
rect 16390 5624 16396 5636
rect 15274 5596 16396 5624
rect 15274 5593 15286 5596
rect 15228 5587 15286 5593
rect 16390 5584 16396 5596
rect 16448 5584 16454 5636
rect 17770 5584 17776 5636
rect 17828 5624 17834 5636
rect 19702 5624 19708 5636
rect 17828 5596 19708 5624
rect 17828 5584 17834 5596
rect 19702 5584 19708 5596
rect 19760 5584 19766 5636
rect 6181 5559 6239 5565
rect 6181 5556 6193 5559
rect 5644 5528 6193 5556
rect 6181 5525 6193 5528
rect 6227 5525 6239 5559
rect 6638 5556 6644 5568
rect 6599 5528 6644 5556
rect 6181 5519 6239 5525
rect 6638 5516 6644 5528
rect 6696 5516 6702 5568
rect 6914 5516 6920 5568
rect 6972 5556 6978 5568
rect 7561 5559 7619 5565
rect 7561 5556 7573 5559
rect 6972 5528 7573 5556
rect 6972 5516 6978 5528
rect 7561 5525 7573 5528
rect 7607 5525 7619 5559
rect 8570 5556 8576 5568
rect 8531 5528 8576 5556
rect 7561 5519 7619 5525
rect 8570 5516 8576 5528
rect 8628 5516 8634 5568
rect 8938 5556 8944 5568
rect 8899 5528 8944 5556
rect 8938 5516 8944 5528
rect 8996 5516 9002 5568
rect 9950 5556 9956 5568
rect 9911 5528 9956 5556
rect 9950 5516 9956 5528
rect 10008 5516 10014 5568
rect 11146 5556 11152 5568
rect 11107 5528 11152 5556
rect 11146 5516 11152 5528
rect 11204 5516 11210 5568
rect 14090 5556 14096 5568
rect 14051 5528 14096 5556
rect 14090 5516 14096 5528
rect 14148 5516 14154 5568
rect 1104 5466 22056 5488
rect 1104 5414 6148 5466
rect 6200 5414 6212 5466
rect 6264 5414 6276 5466
rect 6328 5414 6340 5466
rect 6392 5414 6404 5466
rect 6456 5414 11346 5466
rect 11398 5414 11410 5466
rect 11462 5414 11474 5466
rect 11526 5414 11538 5466
rect 11590 5414 11602 5466
rect 11654 5414 16544 5466
rect 16596 5414 16608 5466
rect 16660 5414 16672 5466
rect 16724 5414 16736 5466
rect 16788 5414 16800 5466
rect 16852 5414 21742 5466
rect 21794 5414 21806 5466
rect 21858 5414 21870 5466
rect 21922 5414 21934 5466
rect 21986 5414 21998 5466
rect 22050 5414 22056 5466
rect 1104 5392 22056 5414
rect 1489 5355 1547 5361
rect 1489 5321 1501 5355
rect 1535 5352 1547 5355
rect 1670 5352 1676 5364
rect 1535 5324 1676 5352
rect 1535 5321 1547 5324
rect 1489 5315 1547 5321
rect 1670 5312 1676 5324
rect 1728 5312 1734 5364
rect 2498 5312 2504 5364
rect 2556 5352 2562 5364
rect 2593 5355 2651 5361
rect 2593 5352 2605 5355
rect 2556 5324 2605 5352
rect 2556 5312 2562 5324
rect 2593 5321 2605 5324
rect 2639 5321 2651 5355
rect 2593 5315 2651 5321
rect 2866 5312 2872 5364
rect 2924 5352 2930 5364
rect 2961 5355 3019 5361
rect 2961 5352 2973 5355
rect 2924 5324 2973 5352
rect 2924 5312 2930 5324
rect 2961 5321 2973 5324
rect 3007 5321 3019 5355
rect 3234 5352 3240 5364
rect 3195 5324 3240 5352
rect 2961 5315 3019 5321
rect 3234 5312 3240 5324
rect 3292 5312 3298 5364
rect 3418 5312 3424 5364
rect 3476 5352 3482 5364
rect 3697 5355 3755 5361
rect 3697 5352 3709 5355
rect 3476 5324 3709 5352
rect 3476 5312 3482 5324
rect 3697 5321 3709 5324
rect 3743 5321 3755 5355
rect 3697 5315 3755 5321
rect 4709 5355 4767 5361
rect 4709 5321 4721 5355
rect 4755 5352 4767 5355
rect 4798 5352 4804 5364
rect 4755 5324 4804 5352
rect 4755 5321 4767 5324
rect 4709 5315 4767 5321
rect 4798 5312 4804 5324
rect 4856 5312 4862 5364
rect 4890 5312 4896 5364
rect 4948 5352 4954 5364
rect 5077 5355 5135 5361
rect 5077 5352 5089 5355
rect 4948 5324 5089 5352
rect 4948 5312 4954 5324
rect 5077 5321 5089 5324
rect 5123 5352 5135 5355
rect 6733 5355 6791 5361
rect 6733 5352 6745 5355
rect 5123 5324 6745 5352
rect 5123 5321 5135 5324
rect 5077 5315 5135 5321
rect 6733 5321 6745 5324
rect 6779 5352 6791 5355
rect 7006 5352 7012 5364
rect 6779 5324 7012 5352
rect 6779 5321 6791 5324
rect 6733 5315 6791 5321
rect 7006 5312 7012 5324
rect 7064 5312 7070 5364
rect 7469 5355 7527 5361
rect 7469 5321 7481 5355
rect 7515 5352 7527 5355
rect 7650 5352 7656 5364
rect 7515 5324 7656 5352
rect 7515 5321 7527 5324
rect 7469 5315 7527 5321
rect 7650 5312 7656 5324
rect 7708 5312 7714 5364
rect 8570 5312 8576 5364
rect 8628 5352 8634 5364
rect 9125 5355 9183 5361
rect 9125 5352 9137 5355
rect 8628 5324 9137 5352
rect 8628 5312 8634 5324
rect 9125 5321 9137 5324
rect 9171 5321 9183 5355
rect 13265 5355 13323 5361
rect 9125 5315 9183 5321
rect 9416 5324 12848 5352
rect 2516 5256 3924 5284
rect 2516 5216 2544 5256
rect 2424 5188 2544 5216
rect 3605 5219 3663 5225
rect 2424 5157 2452 5188
rect 3605 5185 3617 5219
rect 3651 5216 3663 5219
rect 3786 5216 3792 5228
rect 3651 5188 3792 5216
rect 3651 5185 3663 5188
rect 3605 5179 3663 5185
rect 2409 5151 2467 5157
rect 2409 5117 2421 5151
rect 2455 5117 2467 5151
rect 2409 5111 2467 5117
rect 2501 5151 2559 5157
rect 2501 5117 2513 5151
rect 2547 5148 2559 5151
rect 2682 5148 2688 5160
rect 2547 5120 2688 5148
rect 2547 5117 2559 5120
rect 2501 5111 2559 5117
rect 1762 4972 1768 5024
rect 1820 5012 1826 5024
rect 1857 5015 1915 5021
rect 1857 5012 1869 5015
rect 1820 4984 1869 5012
rect 1820 4972 1826 4984
rect 1857 4981 1869 4984
rect 1903 5012 1915 5015
rect 2516 5012 2544 5111
rect 2682 5108 2688 5120
rect 2740 5108 2746 5160
rect 3712 5080 3740 5188
rect 3786 5176 3792 5188
rect 3844 5176 3850 5228
rect 3896 5160 3924 5256
rect 4062 5244 4068 5296
rect 4120 5284 4126 5296
rect 5534 5284 5540 5296
rect 4120 5256 5540 5284
rect 4120 5244 4126 5256
rect 5534 5244 5540 5256
rect 5592 5244 5598 5296
rect 6638 5244 6644 5296
rect 6696 5284 6702 5296
rect 9217 5287 9275 5293
rect 9217 5284 9229 5287
rect 6696 5256 9229 5284
rect 6696 5244 6702 5256
rect 9217 5253 9229 5256
rect 9263 5253 9275 5287
rect 9217 5247 9275 5253
rect 4433 5219 4491 5225
rect 4433 5185 4445 5219
rect 4479 5216 4491 5219
rect 4890 5216 4896 5228
rect 4479 5188 4896 5216
rect 4479 5185 4491 5188
rect 4433 5179 4491 5185
rect 4890 5176 4896 5188
rect 4948 5176 4954 5228
rect 5169 5219 5227 5225
rect 5169 5185 5181 5219
rect 5215 5216 5227 5219
rect 5258 5216 5264 5228
rect 5215 5188 5264 5216
rect 5215 5185 5227 5188
rect 5169 5179 5227 5185
rect 5258 5176 5264 5188
rect 5316 5216 5322 5228
rect 5997 5219 6055 5225
rect 5997 5216 6009 5219
rect 5316 5188 6009 5216
rect 5316 5176 5322 5188
rect 5997 5185 6009 5188
rect 6043 5216 6055 5219
rect 6825 5219 6883 5225
rect 6825 5216 6837 5219
rect 6043 5188 6837 5216
rect 6043 5185 6055 5188
rect 5997 5179 6055 5185
rect 6825 5185 6837 5188
rect 6871 5216 6883 5219
rect 7006 5216 7012 5228
rect 6871 5188 7012 5216
rect 6871 5185 6883 5188
rect 6825 5179 6883 5185
rect 7006 5176 7012 5188
rect 7064 5176 7070 5228
rect 8205 5219 8263 5225
rect 8205 5185 8217 5219
rect 8251 5216 8263 5219
rect 8938 5216 8944 5228
rect 8251 5188 8944 5216
rect 8251 5185 8263 5188
rect 8205 5179 8263 5185
rect 8938 5176 8944 5188
rect 8996 5176 9002 5228
rect 3878 5148 3884 5160
rect 3839 5120 3884 5148
rect 3878 5108 3884 5120
rect 3936 5108 3942 5160
rect 5353 5151 5411 5157
rect 5353 5117 5365 5151
rect 5399 5148 5411 5151
rect 5626 5148 5632 5160
rect 5399 5120 5632 5148
rect 5399 5117 5411 5120
rect 5353 5111 5411 5117
rect 5626 5108 5632 5120
rect 5684 5148 5690 5160
rect 5902 5148 5908 5160
rect 5684 5120 5908 5148
rect 5684 5108 5690 5120
rect 5902 5108 5908 5120
rect 5960 5108 5966 5160
rect 6917 5151 6975 5157
rect 6917 5117 6929 5151
rect 6963 5117 6975 5151
rect 6917 5111 6975 5117
rect 4246 5080 4252 5092
rect 3712 5052 4252 5080
rect 4246 5040 4252 5052
rect 4304 5040 4310 5092
rect 6730 5040 6736 5092
rect 6788 5080 6794 5092
rect 6932 5080 6960 5111
rect 7374 5108 7380 5160
rect 7432 5148 7438 5160
rect 9416 5157 9444 5324
rect 9582 5244 9588 5296
rect 9640 5284 9646 5296
rect 12434 5284 12440 5296
rect 9640 5256 12440 5284
rect 9640 5244 9646 5256
rect 12434 5244 12440 5256
rect 12492 5244 12498 5296
rect 12618 5244 12624 5296
rect 12676 5293 12682 5296
rect 12676 5284 12688 5293
rect 12676 5256 12721 5284
rect 12676 5247 12688 5256
rect 12676 5244 12682 5247
rect 10870 5176 10876 5228
rect 10928 5225 10934 5228
rect 10928 5216 10940 5225
rect 11146 5216 11152 5228
rect 10928 5188 10973 5216
rect 11107 5188 11152 5216
rect 10928 5179 10940 5188
rect 10928 5176 10934 5179
rect 11146 5176 11152 5188
rect 11204 5176 11210 5228
rect 7929 5151 7987 5157
rect 7929 5148 7941 5151
rect 7432 5120 7941 5148
rect 7432 5108 7438 5120
rect 7929 5117 7941 5120
rect 7975 5117 7987 5151
rect 7929 5111 7987 5117
rect 9401 5151 9459 5157
rect 9401 5117 9413 5151
rect 9447 5117 9459 5151
rect 12820 5148 12848 5324
rect 13265 5321 13277 5355
rect 13311 5352 13323 5355
rect 13446 5352 13452 5364
rect 13311 5324 13452 5352
rect 13311 5321 13323 5324
rect 13265 5315 13323 5321
rect 12897 5219 12955 5225
rect 12897 5185 12909 5219
rect 12943 5216 12955 5219
rect 12986 5216 12992 5228
rect 12943 5188 12992 5216
rect 12943 5185 12955 5188
rect 12897 5179 12955 5185
rect 12986 5176 12992 5188
rect 13044 5216 13050 5228
rect 13280 5216 13308 5315
rect 13446 5312 13452 5324
rect 13504 5352 13510 5364
rect 13541 5355 13599 5361
rect 13541 5352 13553 5355
rect 13504 5324 13553 5352
rect 13504 5312 13510 5324
rect 13541 5321 13553 5324
rect 13587 5321 13599 5355
rect 13541 5315 13599 5321
rect 15746 5312 15752 5364
rect 15804 5352 15810 5364
rect 16209 5355 16267 5361
rect 16209 5352 16221 5355
rect 15804 5324 16221 5352
rect 15804 5312 15810 5324
rect 14090 5244 14096 5296
rect 14148 5284 14154 5296
rect 15666 5287 15724 5293
rect 15666 5284 15678 5287
rect 14148 5256 15678 5284
rect 14148 5244 14154 5256
rect 15666 5253 15678 5256
rect 15712 5253 15724 5287
rect 15666 5247 15724 5253
rect 13044 5188 13308 5216
rect 13044 5176 13050 5188
rect 14108 5148 14136 5244
rect 15948 5225 15976 5324
rect 16209 5321 16221 5324
rect 16255 5321 16267 5355
rect 18322 5352 18328 5364
rect 18283 5324 18328 5352
rect 16209 5315 16267 5321
rect 18322 5312 18328 5324
rect 18380 5352 18386 5364
rect 18969 5355 19027 5361
rect 18969 5352 18981 5355
rect 18380 5324 18981 5352
rect 18380 5312 18386 5324
rect 18969 5321 18981 5324
rect 19015 5352 19027 5355
rect 19337 5355 19395 5361
rect 19337 5352 19349 5355
rect 19015 5324 19349 5352
rect 19015 5321 19027 5324
rect 18969 5315 19027 5321
rect 19337 5321 19349 5324
rect 19383 5321 19395 5355
rect 19702 5352 19708 5364
rect 19663 5324 19708 5352
rect 19337 5315 19395 5321
rect 19702 5312 19708 5324
rect 19760 5312 19766 5364
rect 17034 5244 17040 5296
rect 17092 5284 17098 5296
rect 18598 5284 18604 5296
rect 17092 5256 18604 5284
rect 17092 5244 17098 5256
rect 18598 5244 18604 5256
rect 18656 5244 18662 5296
rect 20714 5244 20720 5296
rect 20772 5284 20778 5296
rect 20818 5287 20876 5293
rect 20818 5284 20830 5287
rect 20772 5256 20830 5284
rect 20772 5244 20778 5256
rect 20818 5253 20830 5256
rect 20864 5253 20876 5287
rect 20818 5247 20876 5253
rect 15933 5219 15991 5225
rect 15933 5185 15945 5219
rect 15979 5216 15991 5219
rect 16482 5216 16488 5228
rect 15979 5188 16488 5216
rect 15979 5185 15991 5188
rect 15933 5179 15991 5185
rect 16482 5176 16488 5188
rect 16540 5216 16546 5228
rect 16942 5225 16948 5228
rect 16669 5219 16727 5225
rect 16669 5216 16681 5219
rect 16540 5188 16681 5216
rect 16540 5176 16546 5188
rect 16669 5185 16681 5188
rect 16715 5185 16727 5219
rect 16669 5179 16727 5185
rect 16936 5179 16948 5225
rect 17000 5216 17006 5228
rect 21082 5216 21088 5228
rect 17000 5188 17036 5216
rect 21043 5188 21088 5216
rect 16942 5176 16948 5179
rect 17000 5176 17006 5188
rect 21082 5176 21088 5188
rect 21140 5176 21146 5228
rect 12820 5120 14136 5148
rect 9401 5111 9459 5117
rect 6788 5052 6960 5080
rect 9769 5083 9827 5089
rect 6788 5040 6794 5052
rect 9769 5049 9781 5083
rect 9815 5080 9827 5083
rect 10042 5080 10048 5092
rect 9815 5052 10048 5080
rect 9815 5049 9827 5052
rect 9769 5043 9827 5049
rect 10042 5040 10048 5052
rect 10100 5040 10106 5092
rect 11517 5083 11575 5089
rect 11517 5049 11529 5083
rect 11563 5080 11575 5083
rect 11790 5080 11796 5092
rect 11563 5052 11796 5080
rect 11563 5049 11575 5052
rect 11517 5043 11575 5049
rect 11790 5040 11796 5052
rect 11848 5040 11854 5092
rect 1903 4984 2544 5012
rect 1903 4981 1915 4984
rect 1857 4975 1915 4981
rect 3142 4972 3148 5024
rect 3200 5012 3206 5024
rect 3970 5012 3976 5024
rect 3200 4984 3976 5012
rect 3200 4972 3206 4984
rect 3970 4972 3976 4984
rect 4028 4972 4034 5024
rect 6362 5012 6368 5024
rect 6323 4984 6368 5012
rect 6362 4972 6368 4984
rect 6420 4972 6426 5024
rect 8570 4972 8576 5024
rect 8628 5012 8634 5024
rect 8757 5015 8815 5021
rect 8757 5012 8769 5015
rect 8628 4984 8769 5012
rect 8628 4972 8634 4984
rect 8757 4981 8769 4984
rect 8803 4981 8815 5015
rect 8757 4975 8815 4981
rect 9122 4972 9128 5024
rect 9180 5012 9186 5024
rect 9398 5012 9404 5024
rect 9180 4984 9404 5012
rect 9180 4972 9186 4984
rect 9398 4972 9404 4984
rect 9456 4972 9462 5024
rect 11606 4972 11612 5024
rect 11664 5012 11670 5024
rect 14553 5015 14611 5021
rect 14553 5012 14565 5015
rect 11664 4984 14565 5012
rect 11664 4972 11670 4984
rect 14553 4981 14565 4984
rect 14599 5012 14611 5015
rect 15194 5012 15200 5024
rect 14599 4984 15200 5012
rect 14599 4981 14611 4984
rect 14553 4975 14611 4981
rect 15194 4972 15200 4984
rect 15252 4972 15258 5024
rect 18049 5015 18107 5021
rect 18049 4981 18061 5015
rect 18095 5012 18107 5015
rect 18138 5012 18144 5024
rect 18095 4984 18144 5012
rect 18095 4981 18107 4984
rect 18049 4975 18107 4981
rect 18138 4972 18144 4984
rect 18196 4972 18202 5024
rect 1104 4922 21896 4944
rect 1104 4870 3549 4922
rect 3601 4870 3613 4922
rect 3665 4870 3677 4922
rect 3729 4870 3741 4922
rect 3793 4870 3805 4922
rect 3857 4870 8747 4922
rect 8799 4870 8811 4922
rect 8863 4870 8875 4922
rect 8927 4870 8939 4922
rect 8991 4870 9003 4922
rect 9055 4870 13945 4922
rect 13997 4870 14009 4922
rect 14061 4870 14073 4922
rect 14125 4870 14137 4922
rect 14189 4870 14201 4922
rect 14253 4870 19143 4922
rect 19195 4870 19207 4922
rect 19259 4870 19271 4922
rect 19323 4870 19335 4922
rect 19387 4870 19399 4922
rect 19451 4870 21896 4922
rect 1104 4848 21896 4870
rect 4522 4768 4528 4820
rect 4580 4808 4586 4820
rect 4617 4811 4675 4817
rect 4617 4808 4629 4811
rect 4580 4780 4629 4808
rect 4580 4768 4586 4780
rect 4617 4777 4629 4780
rect 4663 4808 4675 4811
rect 4890 4808 4896 4820
rect 4663 4780 4896 4808
rect 4663 4777 4675 4780
rect 4617 4771 4675 4777
rect 4890 4768 4896 4780
rect 4948 4768 4954 4820
rect 5169 4811 5227 4817
rect 5169 4777 5181 4811
rect 5215 4808 5227 4811
rect 5258 4808 5264 4820
rect 5215 4780 5264 4808
rect 5215 4777 5227 4780
rect 5169 4771 5227 4777
rect 5258 4768 5264 4780
rect 5316 4768 5322 4820
rect 5626 4768 5632 4820
rect 5684 4808 5690 4820
rect 8573 4811 8631 4817
rect 8573 4808 8585 4811
rect 5684 4780 8585 4808
rect 5684 4768 5690 4780
rect 8573 4777 8585 4780
rect 8619 4808 8631 4811
rect 10870 4808 10876 4820
rect 8619 4780 9628 4808
rect 10831 4780 10876 4808
rect 8619 4777 8631 4780
rect 8573 4771 8631 4777
rect 3329 4743 3387 4749
rect 3329 4709 3341 4743
rect 3375 4740 3387 4743
rect 3878 4740 3884 4752
rect 3375 4712 3884 4740
rect 3375 4709 3387 4712
rect 3329 4703 3387 4709
rect 3878 4700 3884 4712
rect 3936 4740 3942 4752
rect 4249 4743 4307 4749
rect 4249 4740 4261 4743
rect 3936 4712 4261 4740
rect 3936 4700 3942 4712
rect 4249 4709 4261 4712
rect 4295 4740 4307 4743
rect 4295 4712 9536 4740
rect 4295 4709 4307 4712
rect 4249 4703 4307 4709
rect 1854 4672 1860 4684
rect 1815 4644 1860 4672
rect 1854 4632 1860 4644
rect 1912 4632 1918 4684
rect 1949 4675 2007 4681
rect 1949 4641 1961 4675
rect 1995 4672 2007 4675
rect 2406 4672 2412 4684
rect 1995 4644 2412 4672
rect 1995 4641 2007 4644
rect 1949 4635 2007 4641
rect 2406 4632 2412 4644
rect 2464 4632 2470 4684
rect 5629 4675 5687 4681
rect 5629 4641 5641 4675
rect 5675 4641 5687 4675
rect 5629 4635 5687 4641
rect 5721 4675 5779 4681
rect 5721 4641 5733 4675
rect 5767 4672 5779 4675
rect 6362 4672 6368 4684
rect 5767 4644 6368 4672
rect 5767 4641 5779 4644
rect 5721 4635 5779 4641
rect 2041 4607 2099 4613
rect 2041 4573 2053 4607
rect 2087 4604 2099 4607
rect 2130 4604 2136 4616
rect 2087 4576 2136 4604
rect 2087 4573 2099 4576
rect 2041 4567 2099 4573
rect 2130 4564 2136 4576
rect 2188 4564 2194 4616
rect 5644 4604 5672 4635
rect 6362 4632 6368 4644
rect 6420 4632 6426 4684
rect 7098 4632 7104 4684
rect 7156 4632 7162 4684
rect 7282 4672 7288 4684
rect 7243 4644 7288 4672
rect 7282 4632 7288 4644
rect 7340 4632 7346 4684
rect 8386 4632 8392 4684
rect 8444 4672 8450 4684
rect 8444 4644 9444 4672
rect 8444 4632 8450 4644
rect 7006 4604 7012 4616
rect 5644 4576 7012 4604
rect 7006 4564 7012 4576
rect 7064 4564 7070 4616
rect 7116 4604 7144 4632
rect 8113 4607 8171 4613
rect 7116 4576 7328 4604
rect 7300 4548 7328 4576
rect 8113 4573 8125 4607
rect 8159 4604 8171 4607
rect 9122 4604 9128 4616
rect 8159 4576 9128 4604
rect 8159 4573 8171 4576
rect 8113 4567 8171 4573
rect 9122 4564 9128 4576
rect 9180 4564 9186 4616
rect 2498 4496 2504 4548
rect 2556 4536 2562 4548
rect 2869 4539 2927 4545
rect 2869 4536 2881 4539
rect 2556 4508 2881 4536
rect 2556 4496 2562 4508
rect 2869 4505 2881 4508
rect 2915 4505 2927 4539
rect 7101 4539 7159 4545
rect 7101 4536 7113 4539
rect 2869 4499 2927 4505
rect 6196 4508 7113 4536
rect 2409 4471 2467 4477
rect 2409 4437 2421 4471
rect 2455 4468 2467 4471
rect 2682 4468 2688 4480
rect 2455 4440 2688 4468
rect 2455 4437 2467 4440
rect 2409 4431 2467 4437
rect 2682 4428 2688 4440
rect 2740 4428 2746 4480
rect 3881 4471 3939 4477
rect 3881 4437 3893 4471
rect 3927 4468 3939 4471
rect 4246 4468 4252 4480
rect 3927 4440 4252 4468
rect 3927 4437 3939 4440
rect 3881 4431 3939 4437
rect 4246 4428 4252 4440
rect 4304 4428 4310 4480
rect 5810 4428 5816 4480
rect 5868 4468 5874 4480
rect 6196 4477 6224 4508
rect 7101 4505 7113 4508
rect 7147 4505 7159 4539
rect 7101 4499 7159 4505
rect 7282 4496 7288 4548
rect 7340 4496 7346 4548
rect 7837 4539 7895 4545
rect 7837 4505 7849 4539
rect 7883 4536 7895 4539
rect 9306 4536 9312 4548
rect 7883 4508 9312 4536
rect 7883 4505 7895 4508
rect 7837 4499 7895 4505
rect 9306 4496 9312 4508
rect 9364 4496 9370 4548
rect 6181 4471 6239 4477
rect 5868 4440 5913 4468
rect 5868 4428 5874 4440
rect 6181 4437 6193 4471
rect 6227 4437 6239 4471
rect 6181 4431 6239 4437
rect 6641 4471 6699 4477
rect 6641 4437 6653 4471
rect 6687 4468 6699 4471
rect 6822 4468 6828 4480
rect 6687 4440 6828 4468
rect 6687 4437 6699 4440
rect 6641 4431 6699 4437
rect 6822 4428 6828 4440
rect 6880 4428 6886 4480
rect 7006 4468 7012 4480
rect 6967 4440 7012 4468
rect 7006 4428 7012 4440
rect 7064 4428 7070 4480
rect 9122 4468 9128 4480
rect 9083 4440 9128 4468
rect 9122 4428 9128 4440
rect 9180 4428 9186 4480
rect 9416 4468 9444 4644
rect 9508 4536 9536 4712
rect 9600 4681 9628 4780
rect 10870 4768 10876 4780
rect 10928 4768 10934 4820
rect 11606 4808 11612 4820
rect 11072 4780 11612 4808
rect 9585 4675 9643 4681
rect 9585 4641 9597 4675
rect 9631 4641 9643 4675
rect 9585 4635 9643 4641
rect 9769 4675 9827 4681
rect 9769 4641 9781 4675
rect 9815 4672 9827 4675
rect 11072 4672 11100 4780
rect 11606 4768 11612 4780
rect 11664 4768 11670 4820
rect 12526 4768 12532 4820
rect 12584 4808 12590 4820
rect 12621 4811 12679 4817
rect 12621 4808 12633 4811
rect 12584 4780 12633 4808
rect 12584 4768 12590 4780
rect 12621 4777 12633 4780
rect 12667 4777 12679 4811
rect 12986 4808 12992 4820
rect 12947 4780 12992 4808
rect 12621 4771 12679 4777
rect 12986 4768 12992 4780
rect 13044 4808 13050 4820
rect 13630 4808 13636 4820
rect 13044 4780 13636 4808
rect 13044 4768 13050 4780
rect 13630 4768 13636 4780
rect 13688 4808 13694 4820
rect 14093 4811 14151 4817
rect 14093 4808 14105 4811
rect 13688 4780 14105 4808
rect 13688 4768 13694 4780
rect 14093 4777 14105 4780
rect 14139 4777 14151 4811
rect 16482 4808 16488 4820
rect 14093 4771 14151 4777
rect 16132 4780 16488 4808
rect 12434 4700 12440 4752
rect 12492 4740 12498 4752
rect 15102 4740 15108 4752
rect 12492 4712 15108 4740
rect 12492 4700 12498 4712
rect 15102 4700 15108 4712
rect 15160 4700 15166 4752
rect 16132 4684 16160 4780
rect 16482 4768 16488 4780
rect 16540 4808 16546 4820
rect 17129 4811 17187 4817
rect 17129 4808 17141 4811
rect 16540 4780 17141 4808
rect 16540 4768 16546 4780
rect 17129 4777 17141 4780
rect 17175 4808 17187 4811
rect 20993 4811 21051 4817
rect 17175 4780 18920 4808
rect 17175 4777 17187 4780
rect 17129 4771 17187 4777
rect 16206 4700 16212 4752
rect 16264 4740 16270 4752
rect 17497 4743 17555 4749
rect 17497 4740 17509 4743
rect 16264 4712 17509 4740
rect 16264 4700 16270 4712
rect 17497 4709 17509 4712
rect 17543 4709 17555 4743
rect 17497 4703 17555 4709
rect 9815 4644 11100 4672
rect 9815 4641 9827 4644
rect 9769 4635 9827 4641
rect 11146 4632 11152 4684
rect 11204 4672 11210 4684
rect 11241 4675 11299 4681
rect 11241 4672 11253 4675
rect 11204 4644 11253 4672
rect 11204 4632 11210 4644
rect 11241 4641 11253 4644
rect 11287 4641 11299 4675
rect 11241 4635 11299 4641
rect 16114 4632 16120 4684
rect 16172 4672 16178 4684
rect 18892 4681 18920 4780
rect 20993 4777 21005 4811
rect 21039 4808 21051 4811
rect 21082 4808 21088 4820
rect 21039 4780 21088 4808
rect 21039 4777 21051 4780
rect 20993 4771 21051 4777
rect 18877 4675 18935 4681
rect 16172 4644 16265 4672
rect 16172 4632 16178 4644
rect 18877 4641 18889 4675
rect 18923 4672 18935 4675
rect 19610 4672 19616 4684
rect 18923 4644 19616 4672
rect 18923 4641 18935 4644
rect 18877 4635 18935 4641
rect 19610 4632 19616 4644
rect 19668 4632 19674 4684
rect 20625 4675 20683 4681
rect 20625 4641 20637 4675
rect 20671 4672 20683 4675
rect 21008 4672 21036 4771
rect 21082 4768 21088 4780
rect 21140 4808 21146 4820
rect 21269 4811 21327 4817
rect 21269 4808 21281 4811
rect 21140 4780 21281 4808
rect 21140 4768 21146 4780
rect 21269 4777 21281 4780
rect 21315 4777 21327 4811
rect 21269 4771 21327 4777
rect 20671 4644 21036 4672
rect 20671 4641 20683 4644
rect 20625 4635 20683 4641
rect 15850 4607 15908 4613
rect 15850 4604 15862 4607
rect 9646 4576 15862 4604
rect 9646 4536 9674 4576
rect 15850 4573 15862 4576
rect 15896 4604 15908 4607
rect 16761 4607 16819 4613
rect 16761 4604 16773 4607
rect 15896 4576 16773 4604
rect 15896 4573 15908 4576
rect 15850 4567 15908 4573
rect 16761 4573 16773 4576
rect 16807 4604 16819 4607
rect 19978 4604 19984 4616
rect 16807 4576 19984 4604
rect 16807 4573 16819 4576
rect 16761 4567 16819 4573
rect 19978 4564 19984 4576
rect 20036 4564 20042 4616
rect 9508 4508 9674 4536
rect 11054 4496 11060 4548
rect 11112 4536 11118 4548
rect 11486 4539 11544 4545
rect 11486 4536 11498 4539
rect 11112 4508 11498 4536
rect 11112 4496 11118 4508
rect 11486 4505 11498 4508
rect 11532 4505 11544 4539
rect 18610 4539 18668 4545
rect 18610 4536 18622 4539
rect 11486 4499 11544 4505
rect 17972 4508 18622 4536
rect 9493 4471 9551 4477
rect 9493 4468 9505 4471
rect 9416 4440 9505 4468
rect 9493 4437 9505 4440
rect 9539 4468 9551 4471
rect 10137 4471 10195 4477
rect 10137 4468 10149 4471
rect 9539 4440 10149 4468
rect 9539 4437 9551 4440
rect 9493 4431 9551 4437
rect 10137 4437 10149 4440
rect 10183 4437 10195 4471
rect 10137 4431 10195 4437
rect 10226 4428 10232 4480
rect 10284 4468 10290 4480
rect 10870 4468 10876 4480
rect 10284 4440 10876 4468
rect 10284 4428 10290 4440
rect 10870 4428 10876 4440
rect 10928 4428 10934 4480
rect 12434 4428 12440 4480
rect 12492 4468 12498 4480
rect 14737 4471 14795 4477
rect 14737 4468 14749 4471
rect 12492 4440 14749 4468
rect 12492 4428 12498 4440
rect 14737 4437 14749 4440
rect 14783 4437 14795 4471
rect 14737 4431 14795 4437
rect 15102 4428 15108 4480
rect 15160 4468 15166 4480
rect 17034 4468 17040 4480
rect 15160 4440 17040 4468
rect 15160 4428 15166 4440
rect 17034 4428 17040 4440
rect 17092 4468 17098 4480
rect 17972 4468 18000 4508
rect 18610 4505 18622 4508
rect 18656 4505 18668 4539
rect 18610 4499 18668 4505
rect 19518 4496 19524 4548
rect 19576 4536 19582 4548
rect 20358 4539 20416 4545
rect 20358 4536 20370 4539
rect 19576 4508 20370 4536
rect 19576 4496 19582 4508
rect 20358 4505 20370 4508
rect 20404 4505 20416 4539
rect 20358 4499 20416 4505
rect 17092 4440 18000 4468
rect 17092 4428 17098 4440
rect 18046 4428 18052 4480
rect 18104 4468 18110 4480
rect 19245 4471 19303 4477
rect 19245 4468 19257 4471
rect 18104 4440 19257 4468
rect 18104 4428 18110 4440
rect 19245 4437 19257 4440
rect 19291 4437 19303 4471
rect 19245 4431 19303 4437
rect 1104 4378 22056 4400
rect 1104 4326 6148 4378
rect 6200 4326 6212 4378
rect 6264 4326 6276 4378
rect 6328 4326 6340 4378
rect 6392 4326 6404 4378
rect 6456 4326 11346 4378
rect 11398 4326 11410 4378
rect 11462 4326 11474 4378
rect 11526 4326 11538 4378
rect 11590 4326 11602 4378
rect 11654 4326 16544 4378
rect 16596 4326 16608 4378
rect 16660 4326 16672 4378
rect 16724 4326 16736 4378
rect 16788 4326 16800 4378
rect 16852 4326 21742 4378
rect 21794 4326 21806 4378
rect 21858 4326 21870 4378
rect 21922 4326 21934 4378
rect 21986 4326 21998 4378
rect 22050 4326 22056 4378
rect 1104 4304 22056 4326
rect 5537 4267 5595 4273
rect 5537 4233 5549 4267
rect 5583 4264 5595 4267
rect 6178 4264 6184 4276
rect 5583 4236 6184 4264
rect 5583 4233 5595 4236
rect 5537 4227 5595 4233
rect 2682 4128 2688 4140
rect 2643 4100 2688 4128
rect 2682 4088 2688 4100
rect 2740 4088 2746 4140
rect 4154 4088 4160 4140
rect 4212 4128 4218 4140
rect 4798 4128 4804 4140
rect 4212 4100 4804 4128
rect 4212 4088 4218 4100
rect 4798 4088 4804 4100
rect 4856 4088 4862 4140
rect 2961 4063 3019 4069
rect 2961 4029 2973 4063
rect 3007 4060 3019 4063
rect 4890 4060 4896 4072
rect 3007 4032 4896 4060
rect 3007 4029 3019 4032
rect 2961 4023 3019 4029
rect 4890 4020 4896 4032
rect 4948 4020 4954 4072
rect 5552 4060 5580 4227
rect 6178 4224 6184 4236
rect 6236 4264 6242 4276
rect 8018 4264 8024 4276
rect 6236 4236 8024 4264
rect 6236 4224 6242 4236
rect 8018 4224 8024 4236
rect 8076 4224 8082 4276
rect 9122 4224 9128 4276
rect 9180 4264 9186 4276
rect 9401 4267 9459 4273
rect 9401 4264 9413 4267
rect 9180 4236 9413 4264
rect 9180 4224 9186 4236
rect 9401 4233 9413 4236
rect 9447 4233 9459 4267
rect 11146 4264 11152 4276
rect 11107 4236 11152 4264
rect 9401 4227 9459 4233
rect 11146 4224 11152 4236
rect 11204 4224 11210 4276
rect 16025 4267 16083 4273
rect 13096 4236 14136 4264
rect 6914 4156 6920 4208
rect 6972 4196 6978 4208
rect 9309 4199 9367 4205
rect 6972 4168 7512 4196
rect 6972 4156 6978 4168
rect 5626 4088 5632 4140
rect 5684 4128 5690 4140
rect 6822 4128 6828 4140
rect 5684 4100 5729 4128
rect 6783 4100 6828 4128
rect 5684 4088 5690 4100
rect 6822 4088 6828 4100
rect 6880 4088 6886 4140
rect 7377 4131 7435 4137
rect 7377 4097 7389 4131
rect 7423 4097 7435 4131
rect 7484 4128 7512 4168
rect 8588 4168 9076 4196
rect 8588 4128 8616 4168
rect 7484 4100 8616 4128
rect 8665 4131 8723 4137
rect 7377 4091 7435 4097
rect 8665 4097 8677 4131
rect 8711 4128 8723 4131
rect 9048 4128 9076 4168
rect 9309 4165 9321 4199
rect 9355 4196 9367 4199
rect 9950 4196 9956 4208
rect 9355 4168 9956 4196
rect 9355 4165 9367 4168
rect 9309 4159 9367 4165
rect 9950 4156 9956 4168
rect 10008 4156 10014 4208
rect 10042 4128 10048 4140
rect 8711 4100 8984 4128
rect 9048 4100 10048 4128
rect 8711 4097 8723 4100
rect 8665 4091 8723 4097
rect 5000 4032 5580 4060
rect 5813 4063 5871 4069
rect 3418 3952 3424 4004
rect 3476 3992 3482 4004
rect 4157 3995 4215 4001
rect 4157 3992 4169 3995
rect 3476 3964 4169 3992
rect 3476 3952 3482 3964
rect 4157 3961 4169 3964
rect 4203 3961 4215 3995
rect 5000 3992 5028 4032
rect 5813 4029 5825 4063
rect 5859 4060 5871 4063
rect 5902 4060 5908 4072
rect 5859 4032 5908 4060
rect 5859 4029 5871 4032
rect 5813 4023 5871 4029
rect 5902 4020 5908 4032
rect 5960 4020 5966 4072
rect 6638 4060 6644 4072
rect 6599 4032 6644 4060
rect 6638 4020 6644 4032
rect 6696 4020 6702 4072
rect 5166 3992 5172 4004
rect 4157 3955 4215 3961
rect 4448 3964 5028 3992
rect 5127 3964 5172 3992
rect 3789 3927 3847 3933
rect 3789 3893 3801 3927
rect 3835 3924 3847 3927
rect 3878 3924 3884 3936
rect 3835 3896 3884 3924
rect 3835 3893 3847 3896
rect 3789 3887 3847 3893
rect 3878 3884 3884 3896
rect 3936 3924 3942 3936
rect 4448 3924 4476 3964
rect 5166 3952 5172 3964
rect 5224 3952 5230 4004
rect 5442 3952 5448 4004
rect 5500 3992 5506 4004
rect 7392 3992 7420 4091
rect 7653 4063 7711 4069
rect 7653 4029 7665 4063
rect 7699 4029 7711 4063
rect 7653 4023 7711 4029
rect 5500 3964 7420 3992
rect 5500 3952 5506 3964
rect 3936 3896 4476 3924
rect 4525 3927 4583 3933
rect 3936 3884 3942 3896
rect 4525 3893 4537 3927
rect 4571 3924 4583 3927
rect 5626 3924 5632 3936
rect 4571 3896 5632 3924
rect 4571 3893 4583 3896
rect 4525 3887 4583 3893
rect 5626 3884 5632 3896
rect 5684 3884 5690 3936
rect 7668 3924 7696 4023
rect 8018 4020 8024 4072
rect 8076 4060 8082 4072
rect 8389 4063 8447 4069
rect 8389 4060 8401 4063
rect 8076 4032 8401 4060
rect 8076 4020 8082 4032
rect 8389 4029 8401 4032
rect 8435 4029 8447 4063
rect 8389 4023 8447 4029
rect 8956 4001 8984 4100
rect 10042 4088 10048 4100
rect 10100 4088 10106 4140
rect 11698 4088 11704 4140
rect 11756 4128 11762 4140
rect 13096 4128 13124 4236
rect 13630 4156 13636 4208
rect 13688 4196 13694 4208
rect 13688 4168 14044 4196
rect 13688 4156 13694 4168
rect 11756 4100 13124 4128
rect 11756 4088 11762 4100
rect 13170 4088 13176 4140
rect 13228 4128 13234 4140
rect 14016 4137 14044 4168
rect 13734 4131 13792 4137
rect 13734 4128 13746 4131
rect 13228 4100 13746 4128
rect 13228 4088 13234 4100
rect 13734 4097 13746 4100
rect 13780 4097 13792 4131
rect 13734 4091 13792 4097
rect 14001 4131 14059 4137
rect 14001 4097 14013 4131
rect 14047 4097 14059 4131
rect 14001 4091 14059 4097
rect 9582 4060 9588 4072
rect 9543 4032 9588 4060
rect 9582 4020 9588 4032
rect 9640 4020 9646 4072
rect 12802 4060 12808 4072
rect 9692 4032 12808 4060
rect 8941 3995 8999 4001
rect 8941 3961 8953 3995
rect 8987 3961 8999 3995
rect 8941 3955 8999 3961
rect 9122 3952 9128 4004
rect 9180 3992 9186 4004
rect 9692 3992 9720 4032
rect 12802 4020 12808 4032
rect 12860 4020 12866 4072
rect 9180 3964 9720 3992
rect 9968 3964 13124 3992
rect 9180 3952 9186 3964
rect 9968 3924 9996 3964
rect 7668 3896 9996 3924
rect 10042 3884 10048 3936
rect 10100 3924 10106 3936
rect 12618 3924 12624 3936
rect 10100 3896 12624 3924
rect 10100 3884 10106 3896
rect 12618 3884 12624 3896
rect 12676 3884 12682 3936
rect 13096 3924 13124 3964
rect 13722 3924 13728 3936
rect 13096 3896 13728 3924
rect 13722 3884 13728 3896
rect 13780 3884 13786 3936
rect 14108 3924 14136 4236
rect 16025 4233 16037 4267
rect 16071 4264 16083 4267
rect 16114 4264 16120 4276
rect 16071 4236 16120 4264
rect 16071 4233 16083 4236
rect 16025 4227 16083 4233
rect 15378 4088 15384 4140
rect 15436 4137 15442 4140
rect 15436 4128 15448 4137
rect 15657 4131 15715 4137
rect 15436 4100 15481 4128
rect 15436 4091 15448 4100
rect 15657 4097 15669 4131
rect 15703 4128 15715 4131
rect 16040 4128 16068 4227
rect 16114 4224 16120 4236
rect 16172 4224 16178 4276
rect 18049 4267 18107 4273
rect 18049 4233 18061 4267
rect 18095 4264 18107 4267
rect 18782 4264 18788 4276
rect 18095 4236 18788 4264
rect 18095 4233 18107 4236
rect 18049 4227 18107 4233
rect 18782 4224 18788 4236
rect 18840 4224 18846 4276
rect 19978 4264 19984 4276
rect 19939 4236 19984 4264
rect 19978 4224 19984 4236
rect 20036 4224 20042 4276
rect 19720 4168 21404 4196
rect 16669 4131 16727 4137
rect 16669 4128 16681 4131
rect 15703 4100 16681 4128
rect 15703 4097 15715 4100
rect 15657 4091 15715 4097
rect 16669 4097 16681 4100
rect 16715 4097 16727 4131
rect 16669 4091 16727 4097
rect 15436 4088 15442 4091
rect 16758 4088 16764 4140
rect 16816 4128 16822 4140
rect 16925 4131 16983 4137
rect 16925 4128 16937 4131
rect 16816 4100 16937 4128
rect 16816 4088 16822 4100
rect 16925 4097 16937 4100
rect 16971 4097 16983 4131
rect 16925 4091 16983 4097
rect 19058 4088 19064 4140
rect 19116 4128 19122 4140
rect 19438 4131 19496 4137
rect 19438 4128 19450 4131
rect 19116 4100 19450 4128
rect 19116 4088 19122 4100
rect 19438 4097 19450 4100
rect 19484 4097 19496 4131
rect 19438 4091 19496 4097
rect 19610 4088 19616 4140
rect 19668 4128 19674 4140
rect 19720 4137 19748 4168
rect 19705 4131 19763 4137
rect 19705 4128 19717 4131
rect 19668 4100 19717 4128
rect 19668 4088 19674 4100
rect 19705 4097 19717 4100
rect 19751 4097 19763 4131
rect 20806 4128 20812 4140
rect 19705 4091 19763 4097
rect 19812 4100 20812 4128
rect 14274 3992 14280 4004
rect 14235 3964 14280 3992
rect 14274 3952 14280 3964
rect 14332 3952 14338 4004
rect 17954 3952 17960 4004
rect 18012 3992 18018 4004
rect 18012 3964 18184 3992
rect 18012 3952 18018 3964
rect 16942 3924 16948 3936
rect 14108 3896 16948 3924
rect 16942 3884 16948 3896
rect 17000 3884 17006 3936
rect 18156 3924 18184 3964
rect 18230 3952 18236 4004
rect 18288 3992 18294 4004
rect 18325 3995 18383 4001
rect 18325 3992 18337 3995
rect 18288 3964 18337 3992
rect 18288 3952 18294 3964
rect 18325 3961 18337 3964
rect 18371 3961 18383 3995
rect 18325 3955 18383 3961
rect 19812 3924 19840 4100
rect 20806 4088 20812 4100
rect 20864 4128 20870 4140
rect 21376 4137 21404 4168
rect 21094 4131 21152 4137
rect 21094 4128 21106 4131
rect 20864 4100 21106 4128
rect 20864 4088 20870 4100
rect 21094 4097 21106 4100
rect 21140 4097 21152 4131
rect 21094 4091 21152 4097
rect 21361 4131 21419 4137
rect 21361 4097 21373 4131
rect 21407 4097 21419 4131
rect 21361 4091 21419 4097
rect 18156 3896 19840 3924
rect 1104 3834 21896 3856
rect 1104 3782 3549 3834
rect 3601 3782 3613 3834
rect 3665 3782 3677 3834
rect 3729 3782 3741 3834
rect 3793 3782 3805 3834
rect 3857 3782 8747 3834
rect 8799 3782 8811 3834
rect 8863 3782 8875 3834
rect 8927 3782 8939 3834
rect 8991 3782 9003 3834
rect 9055 3782 13945 3834
rect 13997 3782 14009 3834
rect 14061 3782 14073 3834
rect 14125 3782 14137 3834
rect 14189 3782 14201 3834
rect 14253 3782 19143 3834
rect 19195 3782 19207 3834
rect 19259 3782 19271 3834
rect 19323 3782 19335 3834
rect 19387 3782 19399 3834
rect 19451 3782 21896 3834
rect 1104 3760 21896 3782
rect 2406 3680 2412 3732
rect 2464 3720 2470 3732
rect 4338 3720 4344 3732
rect 2464 3692 2774 3720
rect 4299 3692 4344 3720
rect 2464 3680 2470 3692
rect 2746 3652 2774 3692
rect 4338 3680 4344 3692
rect 4396 3680 4402 3732
rect 5810 3720 5816 3732
rect 5771 3692 5816 3720
rect 5810 3680 5816 3692
rect 5868 3680 5874 3732
rect 5902 3680 5908 3732
rect 5960 3720 5966 3732
rect 9122 3720 9128 3732
rect 5960 3692 9128 3720
rect 5960 3680 5966 3692
rect 9122 3680 9128 3692
rect 9180 3680 9186 3732
rect 9582 3680 9588 3732
rect 9640 3720 9646 3732
rect 12710 3720 12716 3732
rect 9640 3692 12716 3720
rect 9640 3680 9646 3692
rect 12710 3680 12716 3692
rect 12768 3680 12774 3732
rect 12986 3720 12992 3732
rect 12947 3692 12992 3720
rect 12986 3680 12992 3692
rect 13044 3680 13050 3732
rect 15841 3723 15899 3729
rect 15841 3689 15853 3723
rect 15887 3720 15899 3723
rect 16114 3720 16120 3732
rect 15887 3692 16120 3720
rect 15887 3689 15899 3692
rect 15841 3683 15899 3689
rect 4522 3652 4528 3664
rect 2746 3624 4528 3652
rect 4522 3612 4528 3624
rect 4580 3612 4586 3664
rect 5442 3612 5448 3664
rect 5500 3652 5506 3664
rect 7466 3652 7472 3664
rect 5500 3624 7472 3652
rect 5500 3612 5506 3624
rect 7466 3612 7472 3624
rect 7524 3612 7530 3664
rect 7650 3612 7656 3664
rect 7708 3652 7714 3664
rect 9217 3655 9275 3661
rect 7708 3624 9168 3652
rect 7708 3612 7714 3624
rect 3142 3544 3148 3596
rect 3200 3584 3206 3596
rect 3973 3587 4031 3593
rect 3973 3584 3985 3587
rect 3200 3556 3985 3584
rect 3200 3544 3206 3556
rect 3973 3553 3985 3556
rect 4019 3584 4031 3587
rect 5626 3584 5632 3596
rect 4019 3556 5632 3584
rect 4019 3553 4031 3556
rect 3973 3547 4031 3553
rect 5626 3544 5632 3556
rect 5684 3584 5690 3596
rect 6273 3587 6331 3593
rect 6273 3584 6285 3587
rect 5684 3556 6285 3584
rect 5684 3544 5690 3556
rect 6273 3553 6285 3556
rect 6319 3553 6331 3587
rect 6273 3547 6331 3553
rect 6457 3587 6515 3593
rect 6457 3553 6469 3587
rect 6503 3584 6515 3587
rect 6730 3584 6736 3596
rect 6503 3556 6736 3584
rect 6503 3553 6515 3556
rect 6457 3547 6515 3553
rect 6730 3544 6736 3556
rect 6788 3584 6794 3596
rect 7742 3584 7748 3596
rect 6788 3556 7748 3584
rect 6788 3544 6794 3556
rect 7742 3544 7748 3556
rect 7800 3544 7806 3596
rect 9140 3584 9168 3624
rect 9217 3621 9229 3655
rect 9263 3652 9275 3655
rect 9950 3652 9956 3664
rect 9263 3624 9956 3652
rect 9263 3621 9275 3624
rect 9217 3615 9275 3621
rect 9950 3612 9956 3624
rect 10008 3612 10014 3664
rect 11241 3655 11299 3661
rect 11241 3621 11253 3655
rect 11287 3621 11299 3655
rect 13004 3652 13032 3680
rect 11241 3615 11299 3621
rect 12636 3624 13032 3652
rect 9674 3584 9680 3596
rect 9140 3556 9680 3584
rect 9674 3544 9680 3556
rect 9732 3544 9738 3596
rect 10965 3587 11023 3593
rect 10965 3553 10977 3587
rect 11011 3584 11023 3587
rect 11146 3584 11152 3596
rect 11011 3556 11152 3584
rect 11011 3553 11023 3556
rect 10965 3547 11023 3553
rect 11146 3544 11152 3556
rect 11204 3544 11210 3596
rect 11256 3584 11284 3615
rect 11606 3584 11612 3596
rect 11256 3556 11612 3584
rect 11606 3544 11612 3556
rect 11664 3544 11670 3596
rect 12636 3593 12664 3624
rect 12621 3587 12679 3593
rect 12621 3553 12633 3587
rect 12667 3553 12679 3587
rect 12621 3547 12679 3553
rect 15473 3587 15531 3593
rect 15473 3553 15485 3587
rect 15519 3584 15531 3587
rect 15856 3584 15884 3683
rect 16114 3680 16120 3692
rect 16172 3680 16178 3732
rect 16945 3723 17003 3729
rect 16945 3689 16957 3723
rect 16991 3720 17003 3723
rect 17034 3720 17040 3732
rect 16991 3692 17040 3720
rect 16991 3689 17003 3692
rect 16945 3683 17003 3689
rect 17034 3680 17040 3692
rect 17092 3680 17098 3732
rect 18693 3723 18751 3729
rect 18693 3689 18705 3723
rect 18739 3720 18751 3723
rect 19610 3720 19616 3732
rect 18739 3692 19616 3720
rect 18739 3689 18751 3692
rect 18693 3683 18751 3689
rect 15519 3556 15884 3584
rect 15519 3553 15531 3556
rect 15473 3547 15531 3553
rect 5074 3516 5080 3528
rect 5035 3488 5080 3516
rect 5074 3476 5080 3488
rect 5132 3476 5138 3528
rect 5353 3519 5411 3525
rect 5353 3485 5365 3519
rect 5399 3516 5411 3519
rect 8570 3516 8576 3528
rect 5399 3488 8432 3516
rect 8531 3488 8576 3516
rect 5399 3485 5411 3488
rect 5353 3479 5411 3485
rect 6178 3448 6184 3460
rect 6139 3420 6184 3448
rect 6178 3408 6184 3420
rect 6236 3408 6242 3460
rect 7466 3448 7472 3460
rect 7427 3420 7472 3448
rect 7466 3408 7472 3420
rect 7524 3408 7530 3460
rect 7558 3408 7564 3460
rect 7616 3448 7622 3460
rect 8294 3448 8300 3460
rect 7616 3420 7661 3448
rect 8255 3420 8300 3448
rect 7616 3408 7622 3420
rect 8294 3408 8300 3420
rect 8352 3408 8358 3460
rect 8404 3448 8432 3488
rect 8570 3476 8576 3488
rect 8628 3476 8634 3528
rect 9033 3519 9091 3525
rect 9033 3485 9045 3519
rect 9079 3485 9091 3519
rect 9033 3479 9091 3485
rect 9048 3448 9076 3479
rect 10410 3476 10416 3528
rect 10468 3516 10474 3528
rect 10698 3519 10756 3525
rect 10698 3516 10710 3519
rect 10468 3488 10710 3516
rect 10468 3476 10474 3488
rect 10698 3485 10710 3488
rect 10744 3485 10756 3519
rect 11164 3516 11192 3544
rect 12636 3516 12664 3547
rect 18322 3544 18328 3596
rect 18380 3584 18386 3596
rect 18708 3584 18736 3683
rect 19610 3680 19616 3692
rect 19668 3720 19674 3732
rect 20901 3723 20959 3729
rect 20901 3720 20913 3723
rect 19668 3692 20913 3720
rect 19668 3680 19674 3692
rect 20640 3596 20668 3692
rect 20901 3689 20913 3692
rect 20947 3720 20959 3723
rect 21269 3723 21327 3729
rect 21269 3720 21281 3723
rect 20947 3692 21281 3720
rect 20947 3689 20959 3692
rect 20901 3683 20959 3689
rect 21269 3689 21281 3692
rect 21315 3689 21327 3723
rect 21269 3683 21327 3689
rect 18380 3556 18736 3584
rect 18380 3544 18386 3556
rect 20622 3544 20628 3596
rect 20680 3584 20686 3596
rect 20680 3556 20773 3584
rect 20680 3544 20686 3556
rect 11164 3488 12664 3516
rect 10698 3479 10756 3485
rect 12802 3476 12808 3528
rect 12860 3516 12866 3528
rect 14274 3516 14280 3528
rect 12860 3488 14280 3516
rect 12860 3476 12866 3488
rect 14274 3476 14280 3488
rect 14332 3476 14338 3528
rect 15194 3476 15200 3528
rect 15252 3525 15258 3528
rect 15252 3516 15264 3525
rect 15252 3488 15297 3516
rect 15252 3479 15264 3488
rect 15252 3476 15258 3479
rect 18046 3476 18052 3528
rect 18104 3525 18110 3528
rect 18104 3516 18116 3525
rect 18104 3488 18149 3516
rect 18104 3479 18116 3488
rect 18104 3476 18110 3479
rect 19794 3476 19800 3528
rect 19852 3516 19858 3528
rect 20358 3519 20416 3525
rect 20358 3516 20370 3519
rect 19852 3488 20370 3516
rect 19852 3476 19858 3488
rect 20358 3485 20370 3488
rect 20404 3485 20416 3519
rect 20358 3479 20416 3485
rect 8404 3420 9076 3448
rect 9674 3408 9680 3460
rect 9732 3448 9738 3460
rect 12342 3448 12348 3460
rect 12400 3457 12406 3460
rect 9732 3420 11376 3448
rect 12312 3420 12348 3448
rect 9732 3408 9738 3420
rect 4798 3380 4804 3392
rect 4759 3352 4804 3380
rect 4798 3340 4804 3352
rect 4856 3340 4862 3392
rect 6914 3340 6920 3392
rect 6972 3380 6978 3392
rect 7101 3383 7159 3389
rect 7101 3380 7113 3383
rect 6972 3352 7113 3380
rect 6972 3340 6978 3352
rect 7101 3349 7113 3352
rect 7147 3349 7159 3383
rect 7101 3343 7159 3349
rect 8662 3340 8668 3392
rect 8720 3380 8726 3392
rect 9582 3380 9588 3392
rect 8720 3352 9588 3380
rect 8720 3340 8726 3352
rect 9582 3340 9588 3352
rect 9640 3340 9646 3392
rect 11348 3380 11376 3420
rect 12342 3408 12348 3420
rect 12400 3411 12412 3457
rect 12400 3408 12406 3411
rect 12710 3408 12716 3460
rect 12768 3448 12774 3460
rect 19518 3448 19524 3460
rect 12768 3420 19524 3448
rect 12768 3408 12774 3420
rect 13446 3380 13452 3392
rect 11348 3352 13452 3380
rect 13446 3340 13452 3352
rect 13504 3340 13510 3392
rect 14108 3389 14136 3420
rect 19518 3408 19524 3420
rect 19576 3408 19582 3460
rect 14093 3383 14151 3389
rect 14093 3349 14105 3383
rect 14139 3349 14151 3383
rect 14093 3343 14151 3349
rect 14642 3340 14648 3392
rect 14700 3380 14706 3392
rect 16390 3380 16396 3392
rect 14700 3352 16396 3380
rect 14700 3340 14706 3352
rect 16390 3340 16396 3352
rect 16448 3340 16454 3392
rect 16482 3340 16488 3392
rect 16540 3380 16546 3392
rect 19245 3383 19303 3389
rect 19245 3380 19257 3383
rect 16540 3352 19257 3380
rect 16540 3340 16546 3352
rect 19245 3349 19257 3352
rect 19291 3349 19303 3383
rect 19245 3343 19303 3349
rect 1104 3290 22056 3312
rect 1104 3238 6148 3290
rect 6200 3238 6212 3290
rect 6264 3238 6276 3290
rect 6328 3238 6340 3290
rect 6392 3238 6404 3290
rect 6456 3238 11346 3290
rect 11398 3238 11410 3290
rect 11462 3238 11474 3290
rect 11526 3238 11538 3290
rect 11590 3238 11602 3290
rect 11654 3238 16544 3290
rect 16596 3238 16608 3290
rect 16660 3238 16672 3290
rect 16724 3238 16736 3290
rect 16788 3238 16800 3290
rect 16852 3238 21742 3290
rect 21794 3238 21806 3290
rect 21858 3238 21870 3290
rect 21922 3238 21934 3290
rect 21986 3238 21998 3290
rect 22050 3238 22056 3290
rect 1104 3216 22056 3238
rect 1486 3176 1492 3188
rect 1447 3148 1492 3176
rect 1486 3136 1492 3148
rect 1544 3136 1550 3188
rect 5261 3179 5319 3185
rect 5261 3145 5273 3179
rect 5307 3176 5319 3179
rect 5902 3176 5908 3188
rect 5307 3148 5908 3176
rect 5307 3145 5319 3148
rect 5261 3139 5319 3145
rect 5902 3136 5908 3148
rect 5960 3136 5966 3188
rect 6914 3176 6920 3188
rect 6875 3148 6920 3176
rect 6914 3136 6920 3148
rect 6972 3136 6978 3188
rect 7006 3136 7012 3188
rect 7064 3176 7070 3188
rect 7377 3179 7435 3185
rect 7377 3176 7389 3179
rect 7064 3148 7389 3176
rect 7064 3136 7070 3148
rect 7377 3145 7389 3148
rect 7423 3145 7435 3179
rect 7377 3139 7435 3145
rect 7926 3136 7932 3188
rect 7984 3176 7990 3188
rect 9030 3176 9036 3188
rect 7984 3148 9036 3176
rect 7984 3136 7990 3148
rect 9030 3136 9036 3148
rect 9088 3136 9094 3188
rect 9769 3179 9827 3185
rect 9769 3145 9781 3179
rect 9815 3176 9827 3179
rect 9858 3176 9864 3188
rect 9815 3148 9864 3176
rect 9815 3145 9827 3148
rect 9769 3139 9827 3145
rect 9858 3136 9864 3148
rect 9916 3176 9922 3188
rect 11422 3176 11428 3188
rect 9916 3148 11428 3176
rect 9916 3136 9922 3148
rect 11422 3136 11428 3148
rect 11480 3136 11486 3188
rect 12802 3136 12808 3188
rect 12860 3176 12866 3188
rect 12897 3179 12955 3185
rect 12897 3176 12909 3179
rect 12860 3148 12909 3176
rect 12860 3136 12866 3148
rect 12897 3145 12909 3148
rect 12943 3176 12955 3179
rect 13170 3176 13176 3188
rect 12943 3148 13176 3176
rect 12943 3145 12955 3148
rect 12897 3139 12955 3145
rect 13170 3136 13176 3148
rect 13228 3136 13234 3188
rect 13357 3179 13415 3185
rect 13357 3145 13369 3179
rect 13403 3176 13415 3179
rect 14642 3176 14648 3188
rect 13403 3148 14648 3176
rect 13403 3145 13415 3148
rect 13357 3139 13415 3145
rect 14642 3136 14648 3148
rect 14700 3136 14706 3188
rect 16669 3179 16727 3185
rect 16669 3176 16681 3179
rect 14936 3148 16681 3176
rect 1504 3040 1532 3136
rect 4798 3068 4804 3120
rect 4856 3108 4862 3120
rect 9309 3111 9367 3117
rect 4856 3080 7052 3108
rect 4856 3068 4862 3080
rect 1857 3043 1915 3049
rect 1857 3040 1869 3043
rect 1504 3012 1869 3040
rect 1857 3009 1869 3012
rect 1903 3009 1915 3043
rect 1857 3003 1915 3009
rect 2409 3043 2467 3049
rect 2409 3009 2421 3043
rect 2455 3040 2467 3043
rect 2961 3043 3019 3049
rect 2961 3040 2973 3043
rect 2455 3012 2973 3040
rect 2455 3009 2467 3012
rect 2409 3003 2467 3009
rect 2961 3009 2973 3012
rect 3007 3040 3019 3043
rect 4430 3040 4436 3052
rect 3007 3012 4436 3040
rect 3007 3009 3019 3012
rect 2961 3003 3019 3009
rect 4430 3000 4436 3012
rect 4488 3000 4494 3052
rect 4614 3040 4620 3052
rect 4575 3012 4620 3040
rect 4614 3000 4620 3012
rect 4672 3000 4678 3052
rect 5442 3040 5448 3052
rect 5403 3012 5448 3040
rect 5442 3000 5448 3012
rect 5500 3000 5506 3052
rect 7024 3049 7052 3080
rect 9309 3077 9321 3111
rect 9355 3108 9367 3111
rect 13078 3108 13084 3120
rect 9355 3080 13084 3108
rect 9355 3077 9367 3080
rect 9309 3071 9367 3077
rect 13078 3068 13084 3080
rect 13136 3068 13142 3120
rect 5997 3043 6055 3049
rect 5997 3009 6009 3043
rect 6043 3009 6055 3043
rect 5997 3003 6055 3009
rect 7009 3043 7067 3049
rect 7009 3009 7021 3043
rect 7055 3009 7067 3043
rect 8018 3040 8024 3052
rect 7979 3012 8024 3040
rect 7009 3003 7067 3009
rect 4801 2907 4859 2913
rect 4801 2873 4813 2907
rect 4847 2904 4859 2907
rect 5810 2904 5816 2916
rect 4847 2876 5672 2904
rect 5771 2876 5816 2904
rect 4847 2873 4859 2876
rect 4801 2867 4859 2873
rect 2038 2836 2044 2848
rect 1999 2808 2044 2836
rect 2038 2796 2044 2808
rect 2096 2796 2102 2848
rect 2590 2836 2596 2848
rect 2551 2808 2596 2836
rect 2590 2796 2596 2808
rect 2648 2796 2654 2848
rect 5644 2836 5672 2876
rect 5810 2864 5816 2876
rect 5868 2864 5874 2916
rect 6012 2904 6040 3003
rect 8018 3000 8024 3012
rect 8076 3000 8082 3052
rect 8754 3040 8760 3052
rect 8715 3012 8760 3040
rect 8754 3000 8760 3012
rect 8812 3000 8818 3052
rect 9030 3040 9036 3052
rect 8991 3012 9036 3040
rect 9030 3000 9036 3012
rect 9088 3000 9094 3052
rect 9766 3000 9772 3052
rect 9824 3040 9830 3052
rect 10882 3043 10940 3049
rect 10882 3040 10894 3043
rect 9824 3012 10894 3040
rect 9824 3000 9830 3012
rect 10882 3009 10894 3012
rect 10928 3009 10940 3043
rect 11146 3040 11152 3052
rect 11107 3012 11152 3040
rect 10882 3003 10940 3009
rect 11146 3000 11152 3012
rect 11204 3040 11210 3052
rect 11517 3043 11575 3049
rect 11517 3040 11529 3043
rect 11204 3012 11529 3040
rect 11204 3000 11210 3012
rect 11517 3009 11529 3012
rect 11563 3009 11575 3043
rect 11773 3043 11831 3049
rect 11773 3040 11785 3043
rect 11517 3003 11575 3009
rect 11624 3012 11785 3040
rect 6825 2975 6883 2981
rect 6825 2941 6837 2975
rect 6871 2972 6883 2975
rect 6914 2972 6920 2984
rect 6871 2944 6920 2972
rect 6871 2941 6883 2944
rect 6825 2935 6883 2941
rect 6914 2932 6920 2944
rect 6972 2972 6978 2984
rect 7098 2972 7104 2984
rect 6972 2944 7104 2972
rect 6972 2932 6978 2944
rect 7098 2932 7104 2944
rect 7156 2932 7162 2984
rect 8573 2975 8631 2981
rect 8573 2941 8585 2975
rect 8619 2972 8631 2975
rect 9582 2972 9588 2984
rect 8619 2944 9588 2972
rect 8619 2941 8631 2944
rect 8573 2935 8631 2941
rect 9582 2932 9588 2944
rect 9640 2932 9646 2984
rect 11422 2932 11428 2984
rect 11480 2972 11486 2984
rect 11624 2972 11652 3012
rect 11773 3009 11785 3012
rect 11819 3009 11831 3043
rect 13170 3040 13176 3052
rect 13131 3012 13176 3040
rect 11773 3003 11831 3009
rect 13170 3000 13176 3012
rect 13228 3000 13234 3052
rect 13722 3040 13728 3052
rect 13683 3012 13728 3040
rect 13722 3000 13728 3012
rect 13780 3000 13786 3052
rect 14642 3040 14648 3052
rect 13832 3012 14648 3040
rect 13832 2972 13860 3012
rect 14642 3000 14648 3012
rect 14700 3000 14706 3052
rect 14737 3043 14795 3049
rect 14737 3009 14749 3043
rect 14783 3040 14795 3043
rect 14936 3040 14964 3148
rect 16669 3145 16681 3148
rect 16715 3145 16727 3179
rect 17126 3176 17132 3188
rect 17087 3148 17132 3176
rect 16669 3139 16727 3145
rect 17126 3136 17132 3148
rect 17184 3136 17190 3188
rect 18233 3179 18291 3185
rect 17236 3148 18184 3176
rect 15746 3068 15752 3120
rect 15804 3108 15810 3120
rect 15804 3080 17172 3108
rect 15804 3068 15810 3080
rect 14783 3012 14964 3040
rect 15013 3043 15071 3049
rect 14783 3009 14795 3012
rect 14737 3003 14795 3009
rect 15013 3009 15025 3043
rect 15059 3009 15071 3043
rect 15562 3040 15568 3052
rect 15523 3012 15568 3040
rect 15013 3003 15071 3009
rect 11480 2944 11652 2972
rect 12820 2944 13860 2972
rect 14553 2975 14611 2981
rect 11480 2932 11486 2944
rect 7374 2904 7380 2916
rect 6012 2876 7380 2904
rect 7374 2864 7380 2876
rect 7432 2864 7438 2916
rect 7837 2907 7895 2913
rect 7837 2873 7849 2907
rect 7883 2904 7895 2907
rect 7883 2876 10180 2904
rect 7883 2873 7895 2876
rect 7837 2867 7895 2873
rect 9674 2836 9680 2848
rect 5644 2808 9680 2836
rect 9674 2796 9680 2808
rect 9732 2796 9738 2848
rect 10152 2836 10180 2876
rect 12820 2836 12848 2944
rect 14553 2941 14565 2975
rect 14599 2972 14611 2975
rect 15028 2972 15056 3003
rect 15562 3000 15568 3012
rect 15620 3000 15626 3052
rect 16301 3043 16359 3049
rect 16301 3009 16313 3043
rect 16347 3040 16359 3043
rect 17037 3043 17095 3049
rect 17037 3040 17049 3043
rect 16347 3012 17049 3040
rect 16347 3009 16359 3012
rect 16301 3003 16359 3009
rect 17037 3009 17049 3012
rect 17083 3009 17095 3043
rect 17037 3003 17095 3009
rect 14599 2944 15056 2972
rect 14599 2941 14611 2944
rect 14553 2935 14611 2941
rect 13814 2864 13820 2916
rect 13872 2904 13878 2916
rect 15197 2907 15255 2913
rect 15197 2904 15209 2907
rect 13872 2876 15209 2904
rect 13872 2864 13878 2876
rect 15197 2873 15209 2876
rect 15243 2873 15255 2907
rect 15197 2867 15255 2873
rect 15749 2907 15807 2913
rect 15749 2873 15761 2907
rect 15795 2904 15807 2907
rect 17034 2904 17040 2916
rect 15795 2876 17040 2904
rect 15795 2873 15807 2876
rect 15749 2867 15807 2873
rect 17034 2864 17040 2876
rect 17092 2864 17098 2916
rect 10152 2808 12848 2836
rect 13909 2839 13967 2845
rect 13909 2805 13921 2839
rect 13955 2836 13967 2839
rect 16942 2836 16948 2848
rect 13955 2808 16948 2836
rect 13955 2805 13967 2808
rect 13909 2799 13967 2805
rect 16942 2796 16948 2808
rect 17000 2796 17006 2848
rect 17144 2836 17172 3080
rect 17236 2981 17264 3148
rect 17865 3111 17923 3117
rect 17865 3077 17877 3111
rect 17911 3108 17923 3111
rect 17954 3108 17960 3120
rect 17911 3080 17960 3108
rect 17911 3077 17923 3080
rect 17865 3071 17923 3077
rect 17954 3068 17960 3080
rect 18012 3068 18018 3120
rect 18156 3108 18184 3148
rect 18233 3145 18245 3179
rect 18279 3176 18291 3179
rect 18322 3176 18328 3188
rect 18279 3148 18328 3176
rect 18279 3145 18291 3148
rect 18233 3139 18291 3145
rect 18322 3136 18328 3148
rect 18380 3136 18386 3188
rect 19889 3179 19947 3185
rect 19889 3145 19901 3179
rect 19935 3145 19947 3179
rect 19889 3139 19947 3145
rect 19058 3108 19064 3120
rect 18156 3080 19064 3108
rect 19058 3068 19064 3080
rect 19116 3108 19122 3120
rect 19904 3108 19932 3139
rect 19116 3080 19932 3108
rect 19116 3068 19122 3080
rect 17770 3000 17776 3052
rect 17828 3040 17834 3052
rect 18322 3040 18328 3052
rect 17828 3012 18328 3040
rect 17828 3000 17834 3012
rect 18322 3000 18328 3012
rect 18380 3040 18386 3052
rect 18782 3049 18788 3052
rect 18509 3043 18567 3049
rect 18509 3040 18521 3043
rect 18380 3012 18521 3040
rect 18380 3000 18386 3012
rect 18509 3009 18521 3012
rect 18555 3009 18567 3043
rect 18776 3040 18788 3049
rect 18743 3012 18788 3040
rect 18509 3003 18567 3009
rect 18776 3003 18788 3012
rect 18782 3000 18788 3003
rect 18840 3000 18846 3052
rect 20346 3040 20352 3052
rect 20307 3012 20352 3040
rect 20346 3000 20352 3012
rect 20404 3040 20410 3052
rect 20806 3040 20812 3052
rect 20404 3012 20812 3040
rect 20404 3000 20410 3012
rect 20806 3000 20812 3012
rect 20864 3000 20870 3052
rect 17221 2975 17279 2981
rect 17221 2941 17233 2975
rect 17267 2941 17279 2975
rect 20622 2972 20628 2984
rect 20583 2944 20628 2972
rect 17221 2935 17279 2941
rect 20622 2932 20628 2944
rect 20680 2932 20686 2984
rect 19794 2836 19800 2848
rect 17144 2808 19800 2836
rect 19794 2796 19800 2808
rect 19852 2796 19858 2848
rect 1104 2746 21896 2768
rect 1104 2694 3549 2746
rect 3601 2694 3613 2746
rect 3665 2694 3677 2746
rect 3729 2694 3741 2746
rect 3793 2694 3805 2746
rect 3857 2694 8747 2746
rect 8799 2694 8811 2746
rect 8863 2694 8875 2746
rect 8927 2694 8939 2746
rect 8991 2694 9003 2746
rect 9055 2694 13945 2746
rect 13997 2694 14009 2746
rect 14061 2694 14073 2746
rect 14125 2694 14137 2746
rect 14189 2694 14201 2746
rect 14253 2694 19143 2746
rect 19195 2694 19207 2746
rect 19259 2694 19271 2746
rect 19323 2694 19335 2746
rect 19387 2694 19399 2746
rect 19451 2694 21896 2746
rect 1104 2672 21896 2694
rect 6638 2592 6644 2644
rect 6696 2632 6702 2644
rect 10318 2632 10324 2644
rect 6696 2604 8432 2632
rect 6696 2592 6702 2604
rect 6730 2564 6736 2576
rect 6691 2536 6736 2564
rect 6730 2524 6736 2536
rect 6788 2524 6794 2576
rect 8294 2564 8300 2576
rect 7024 2536 8300 2564
rect 1946 2428 1952 2440
rect 1907 2400 1952 2428
rect 1946 2388 1952 2400
rect 2004 2428 2010 2440
rect 2501 2431 2559 2437
rect 2501 2428 2513 2431
rect 2004 2400 2513 2428
rect 2004 2388 2010 2400
rect 2501 2397 2513 2400
rect 2547 2397 2559 2431
rect 2501 2391 2559 2397
rect 4890 2388 4896 2440
rect 4948 2428 4954 2440
rect 5169 2431 5227 2437
rect 5169 2428 5181 2431
rect 4948 2400 5181 2428
rect 4948 2388 4954 2400
rect 5169 2397 5181 2400
rect 5215 2397 5227 2431
rect 5169 2391 5227 2397
rect 5997 2431 6055 2437
rect 5997 2397 6009 2431
rect 6043 2428 6055 2431
rect 6917 2431 6975 2437
rect 6043 2400 6868 2428
rect 6043 2397 6055 2400
rect 5997 2391 6055 2397
rect 3050 2320 3056 2372
rect 3108 2360 3114 2372
rect 6840 2360 6868 2400
rect 6917 2397 6929 2431
rect 6963 2428 6975 2431
rect 7024 2428 7052 2536
rect 8294 2524 8300 2536
rect 8352 2524 8358 2576
rect 8202 2496 8208 2508
rect 7392 2468 8208 2496
rect 7190 2428 7196 2440
rect 6963 2400 7052 2428
rect 7151 2400 7196 2428
rect 6963 2397 6975 2400
rect 6917 2391 6975 2397
rect 7190 2388 7196 2400
rect 7248 2388 7254 2440
rect 7392 2360 7420 2468
rect 8202 2456 8208 2468
rect 8260 2456 8266 2508
rect 8404 2496 8432 2604
rect 9646 2604 10324 2632
rect 8481 2567 8539 2573
rect 8481 2533 8493 2567
rect 8527 2533 8539 2567
rect 8481 2527 8539 2533
rect 8312 2468 8432 2496
rect 8312 2437 8340 2468
rect 8297 2431 8355 2437
rect 8297 2397 8309 2431
rect 8343 2397 8355 2431
rect 8496 2428 8524 2527
rect 9490 2524 9496 2576
rect 9548 2564 9554 2576
rect 9646 2564 9674 2604
rect 10318 2592 10324 2604
rect 10376 2592 10382 2644
rect 11146 2632 11152 2644
rect 11107 2604 11152 2632
rect 11146 2592 11152 2604
rect 11204 2592 11210 2644
rect 17126 2632 17132 2644
rect 11624 2604 17132 2632
rect 9950 2564 9956 2576
rect 9548 2536 9674 2564
rect 9876 2536 9956 2564
rect 9548 2524 9554 2536
rect 9030 2456 9036 2508
rect 9088 2496 9094 2508
rect 9401 2499 9459 2505
rect 9088 2468 9352 2496
rect 9088 2456 9094 2468
rect 9324 2428 9352 2468
rect 9401 2465 9413 2499
rect 9447 2496 9459 2499
rect 9876 2496 9904 2536
rect 9950 2524 9956 2536
rect 10008 2524 10014 2576
rect 10045 2567 10103 2573
rect 10045 2533 10057 2567
rect 10091 2564 10103 2567
rect 10091 2536 10640 2564
rect 10091 2533 10103 2536
rect 10045 2527 10103 2533
rect 9447 2468 9904 2496
rect 10612 2496 10640 2536
rect 11054 2524 11060 2576
rect 11112 2564 11118 2576
rect 11517 2567 11575 2573
rect 11517 2564 11529 2567
rect 11112 2536 11529 2564
rect 11112 2524 11118 2536
rect 11517 2533 11529 2536
rect 11563 2533 11575 2567
rect 11517 2527 11575 2533
rect 11624 2496 11652 2604
rect 17126 2592 17132 2604
rect 17184 2592 17190 2644
rect 17589 2635 17647 2641
rect 17589 2601 17601 2635
rect 17635 2632 17647 2635
rect 17770 2632 17776 2644
rect 17635 2604 17776 2632
rect 17635 2601 17647 2604
rect 17589 2595 17647 2601
rect 17770 2592 17776 2604
rect 17828 2592 17834 2644
rect 17957 2635 18015 2641
rect 17957 2601 17969 2635
rect 18003 2632 18015 2635
rect 20346 2632 20352 2644
rect 18003 2604 20352 2632
rect 18003 2601 18015 2604
rect 17957 2595 18015 2601
rect 20346 2592 20352 2604
rect 20404 2592 20410 2644
rect 20622 2592 20628 2644
rect 20680 2632 20686 2644
rect 21085 2635 21143 2641
rect 21085 2632 21097 2635
rect 20680 2604 21097 2632
rect 20680 2592 20686 2604
rect 21085 2601 21097 2604
rect 21131 2601 21143 2635
rect 21085 2595 21143 2601
rect 20714 2524 20720 2576
rect 20772 2564 20778 2576
rect 20809 2567 20867 2573
rect 20809 2564 20821 2567
rect 20772 2536 20821 2564
rect 20772 2524 20778 2536
rect 20809 2533 20821 2536
rect 20855 2533 20867 2567
rect 20809 2527 20867 2533
rect 12894 2496 12900 2508
rect 10612 2468 11652 2496
rect 12855 2468 12900 2496
rect 9447 2465 9459 2468
rect 9401 2459 9459 2465
rect 12894 2456 12900 2468
rect 12952 2496 12958 2508
rect 13173 2499 13231 2505
rect 13173 2496 13185 2499
rect 12952 2468 13185 2496
rect 12952 2456 12958 2468
rect 13173 2465 13185 2468
rect 13219 2496 13231 2499
rect 13541 2499 13599 2505
rect 13541 2496 13553 2499
rect 13219 2468 13553 2496
rect 13219 2465 13231 2468
rect 13173 2459 13231 2465
rect 13541 2465 13553 2468
rect 13587 2465 13599 2499
rect 13541 2459 13599 2465
rect 9585 2431 9643 2437
rect 9585 2428 9597 2431
rect 8496 2400 9168 2428
rect 9324 2400 9597 2428
rect 8297 2391 8355 2397
rect 3108 2332 5948 2360
rect 6840 2332 7420 2360
rect 7469 2363 7527 2369
rect 3108 2320 3114 2332
rect 2130 2292 2136 2304
rect 2091 2264 2136 2292
rect 2130 2252 2136 2264
rect 2188 2252 2194 2304
rect 3878 2252 3884 2304
rect 3936 2292 3942 2304
rect 4801 2295 4859 2301
rect 4801 2292 4813 2295
rect 3936 2264 4813 2292
rect 3936 2252 3942 2264
rect 4801 2261 4813 2264
rect 4847 2261 4859 2295
rect 4801 2255 4859 2261
rect 5353 2295 5411 2301
rect 5353 2261 5365 2295
rect 5399 2292 5411 2295
rect 5534 2292 5540 2304
rect 5399 2264 5540 2292
rect 5399 2261 5411 2264
rect 5353 2255 5411 2261
rect 5534 2252 5540 2264
rect 5592 2252 5598 2304
rect 5810 2292 5816 2304
rect 5771 2264 5816 2292
rect 5810 2252 5816 2264
rect 5868 2252 5874 2304
rect 5920 2292 5948 2332
rect 7469 2329 7481 2363
rect 7515 2360 7527 2363
rect 8202 2360 8208 2372
rect 7515 2332 8208 2360
rect 7515 2329 7527 2332
rect 7469 2323 7527 2329
rect 8202 2320 8208 2332
rect 8260 2320 8266 2372
rect 9030 2360 9036 2372
rect 8991 2332 9036 2360
rect 9030 2320 9036 2332
rect 9088 2320 9094 2372
rect 9140 2360 9168 2400
rect 9585 2397 9597 2400
rect 9631 2397 9643 2431
rect 9585 2391 9643 2397
rect 10318 2388 10324 2440
rect 10376 2437 10382 2440
rect 10376 2428 10385 2437
rect 10376 2400 10421 2428
rect 10376 2391 10385 2400
rect 10376 2388 10382 2391
rect 10594 2388 10600 2440
rect 10652 2428 10658 2440
rect 15105 2431 15163 2437
rect 15105 2428 15117 2431
rect 10652 2400 15117 2428
rect 10652 2388 10658 2400
rect 15105 2397 15117 2400
rect 15151 2397 15163 2431
rect 15105 2391 15163 2397
rect 18325 2431 18383 2437
rect 18325 2397 18337 2431
rect 18371 2428 18383 2431
rect 18601 2431 18659 2437
rect 18601 2428 18613 2431
rect 18371 2400 18613 2428
rect 18371 2397 18383 2400
rect 18325 2391 18383 2397
rect 18601 2397 18613 2400
rect 18647 2428 18659 2431
rect 19334 2428 19340 2440
rect 18647 2400 19340 2428
rect 18647 2397 18659 2400
rect 18601 2391 18659 2397
rect 19334 2388 19340 2400
rect 19392 2388 19398 2440
rect 19429 2431 19487 2437
rect 19429 2397 19441 2431
rect 19475 2428 19487 2431
rect 20622 2428 20628 2440
rect 19475 2400 20628 2428
rect 19475 2397 19487 2400
rect 19429 2391 19487 2397
rect 20622 2388 20628 2400
rect 20680 2388 20686 2440
rect 9140 2332 12434 2360
rect 7929 2295 7987 2301
rect 7929 2292 7941 2295
rect 5920 2264 7941 2292
rect 7929 2261 7941 2264
rect 7975 2292 7987 2295
rect 9214 2292 9220 2304
rect 7975 2264 9220 2292
rect 7975 2261 7987 2264
rect 7929 2255 7987 2261
rect 9214 2252 9220 2264
rect 9272 2252 9278 2304
rect 9490 2252 9496 2304
rect 9548 2292 9554 2304
rect 9677 2295 9735 2301
rect 9677 2292 9689 2295
rect 9548 2264 9689 2292
rect 9548 2252 9554 2264
rect 9677 2261 9689 2264
rect 9723 2261 9735 2295
rect 9677 2255 9735 2261
rect 10505 2295 10563 2301
rect 10505 2261 10517 2295
rect 10551 2292 10563 2295
rect 11698 2292 11704 2304
rect 10551 2264 11704 2292
rect 10551 2261 10563 2264
rect 10505 2255 10563 2261
rect 11698 2252 11704 2264
rect 11756 2252 11762 2304
rect 12406 2292 12434 2332
rect 12618 2320 12624 2372
rect 12676 2369 12682 2372
rect 12676 2360 12688 2369
rect 12676 2332 12721 2360
rect 12676 2323 12688 2332
rect 12676 2320 12682 2323
rect 18138 2320 18144 2372
rect 18196 2360 18202 2372
rect 19674 2363 19732 2369
rect 19674 2360 19686 2363
rect 18196 2332 19686 2360
rect 18196 2320 18202 2332
rect 19674 2329 19686 2332
rect 19720 2329 19732 2363
rect 19674 2323 19732 2329
rect 13078 2292 13084 2304
rect 12406 2264 13084 2292
rect 13078 2252 13084 2264
rect 13136 2252 13142 2304
rect 15289 2295 15347 2301
rect 15289 2261 15301 2295
rect 15335 2292 15347 2295
rect 17494 2292 17500 2304
rect 15335 2264 17500 2292
rect 15335 2261 15347 2264
rect 15289 2255 15347 2261
rect 17494 2252 17500 2264
rect 17552 2252 17558 2304
rect 18785 2295 18843 2301
rect 18785 2261 18797 2295
rect 18831 2292 18843 2295
rect 20438 2292 20444 2304
rect 18831 2264 20444 2292
rect 18831 2261 18843 2264
rect 18785 2255 18843 2261
rect 20438 2252 20444 2264
rect 20496 2252 20502 2304
rect 1104 2202 22056 2224
rect 1104 2150 6148 2202
rect 6200 2150 6212 2202
rect 6264 2150 6276 2202
rect 6328 2150 6340 2202
rect 6392 2150 6404 2202
rect 6456 2150 11346 2202
rect 11398 2150 11410 2202
rect 11462 2150 11474 2202
rect 11526 2150 11538 2202
rect 11590 2150 11602 2202
rect 11654 2150 16544 2202
rect 16596 2150 16608 2202
rect 16660 2150 16672 2202
rect 16724 2150 16736 2202
rect 16788 2150 16800 2202
rect 16852 2150 21742 2202
rect 21794 2150 21806 2202
rect 21858 2150 21870 2202
rect 21922 2150 21934 2202
rect 21986 2150 21998 2202
rect 22050 2150 22056 2202
rect 1104 2128 22056 2150
rect 6454 2048 6460 2100
rect 6512 2088 6518 2100
rect 7282 2088 7288 2100
rect 6512 2060 7288 2088
rect 6512 2048 6518 2060
rect 7282 2048 7288 2060
rect 7340 2048 7346 2100
rect 9950 2048 9956 2100
rect 10008 2088 10014 2100
rect 18782 2088 18788 2100
rect 10008 2060 18788 2088
rect 10008 2048 10014 2060
rect 18782 2048 18788 2060
rect 18840 2048 18846 2100
rect 19334 1980 19340 2032
rect 19392 2020 19398 2032
rect 20070 2020 20076 2032
rect 19392 1992 20076 2020
rect 19392 1980 19398 1992
rect 20070 1980 20076 1992
rect 20128 1980 20134 2032
rect 8202 1912 8208 1964
rect 8260 1952 8266 1964
rect 13170 1952 13176 1964
rect 8260 1924 13176 1952
rect 8260 1912 8266 1924
rect 13170 1912 13176 1924
rect 13228 1912 13234 1964
rect 11698 1844 11704 1896
rect 11756 1884 11762 1896
rect 16022 1884 16028 1896
rect 11756 1856 16028 1884
rect 11756 1844 11762 1856
rect 16022 1844 16028 1856
rect 16080 1844 16086 1896
rect 6730 1708 6736 1760
rect 6788 1748 6794 1760
rect 14918 1748 14924 1760
rect 6788 1720 14924 1748
rect 6788 1708 6794 1720
rect 14918 1708 14924 1720
rect 14976 1708 14982 1760
rect 5534 1640 5540 1692
rect 5592 1680 5598 1692
rect 12710 1680 12716 1692
rect 5592 1652 12716 1680
rect 5592 1640 5598 1652
rect 12710 1640 12716 1652
rect 12768 1640 12774 1692
rect 9030 1572 9036 1624
rect 9088 1612 9094 1624
rect 15746 1612 15752 1624
rect 9088 1584 15752 1612
rect 9088 1572 9094 1584
rect 15746 1572 15752 1584
rect 15804 1572 15810 1624
rect 5810 1504 5816 1556
rect 5868 1544 5874 1556
rect 14550 1544 14556 1556
rect 5868 1516 14556 1544
rect 5868 1504 5874 1516
rect 14550 1504 14556 1516
rect 14608 1504 14614 1556
rect 7558 1368 7564 1420
rect 7616 1408 7622 1420
rect 8110 1408 8116 1420
rect 7616 1380 8116 1408
rect 7616 1368 7622 1380
rect 8110 1368 8116 1380
rect 8168 1368 8174 1420
rect 11974 1232 11980 1284
rect 12032 1232 12038 1284
rect 11992 1080 12020 1232
rect 11974 1028 11980 1080
rect 12032 1028 12038 1080
rect 9766 892 9772 944
rect 9824 932 9830 944
rect 10686 932 10692 944
rect 9824 904 10692 932
rect 9824 892 9830 904
rect 10686 892 10692 904
rect 10744 892 10750 944
<< via1 >>
rect 2964 20952 3016 21004
rect 5908 20952 5960 21004
rect 3884 20748 3936 20800
rect 5632 20748 5684 20800
rect 6148 20646 6200 20698
rect 6212 20646 6264 20698
rect 6276 20646 6328 20698
rect 6340 20646 6392 20698
rect 6404 20646 6456 20698
rect 11346 20646 11398 20698
rect 11410 20646 11462 20698
rect 11474 20646 11526 20698
rect 11538 20646 11590 20698
rect 11602 20646 11654 20698
rect 16544 20646 16596 20698
rect 16608 20646 16660 20698
rect 16672 20646 16724 20698
rect 16736 20646 16788 20698
rect 16800 20646 16852 20698
rect 21742 20646 21794 20698
rect 21806 20646 21858 20698
rect 21870 20646 21922 20698
rect 21934 20646 21986 20698
rect 21998 20646 22050 20698
rect 3549 20102 3601 20154
rect 3613 20102 3665 20154
rect 3677 20102 3729 20154
rect 3741 20102 3793 20154
rect 3805 20102 3857 20154
rect 8747 20102 8799 20154
rect 8811 20102 8863 20154
rect 8875 20102 8927 20154
rect 8939 20102 8991 20154
rect 9003 20102 9055 20154
rect 13945 20102 13997 20154
rect 14009 20102 14061 20154
rect 14073 20102 14125 20154
rect 14137 20102 14189 20154
rect 14201 20102 14253 20154
rect 19143 20102 19195 20154
rect 19207 20102 19259 20154
rect 19271 20102 19323 20154
rect 19335 20102 19387 20154
rect 19399 20102 19451 20154
rect 4068 20000 4120 20052
rect 5632 20043 5684 20052
rect 5632 20009 5641 20043
rect 5641 20009 5675 20043
rect 5675 20009 5684 20043
rect 5632 20000 5684 20009
rect 5816 19839 5868 19848
rect 5816 19805 5825 19839
rect 5825 19805 5859 19839
rect 5859 19805 5868 19839
rect 5816 19796 5868 19805
rect 10416 19796 10468 19848
rect 6148 19558 6200 19610
rect 6212 19558 6264 19610
rect 6276 19558 6328 19610
rect 6340 19558 6392 19610
rect 6404 19558 6456 19610
rect 11346 19558 11398 19610
rect 11410 19558 11462 19610
rect 11474 19558 11526 19610
rect 11538 19558 11590 19610
rect 11602 19558 11654 19610
rect 16544 19558 16596 19610
rect 16608 19558 16660 19610
rect 16672 19558 16724 19610
rect 16736 19558 16788 19610
rect 16800 19558 16852 19610
rect 21742 19558 21794 19610
rect 21806 19558 21858 19610
rect 21870 19558 21922 19610
rect 21934 19558 21986 19610
rect 21998 19558 22050 19610
rect 3240 19456 3292 19508
rect 5816 19388 5868 19440
rect 4712 19363 4764 19372
rect 4712 19329 4721 19363
rect 4721 19329 4755 19363
rect 4755 19329 4764 19363
rect 4712 19320 4764 19329
rect 9128 19320 9180 19372
rect 3549 19014 3601 19066
rect 3613 19014 3665 19066
rect 3677 19014 3729 19066
rect 3741 19014 3793 19066
rect 3805 19014 3857 19066
rect 8747 19014 8799 19066
rect 8811 19014 8863 19066
rect 8875 19014 8927 19066
rect 8939 19014 8991 19066
rect 9003 19014 9055 19066
rect 13945 19014 13997 19066
rect 14009 19014 14061 19066
rect 14073 19014 14125 19066
rect 14137 19014 14189 19066
rect 14201 19014 14253 19066
rect 19143 19014 19195 19066
rect 19207 19014 19259 19066
rect 19271 19014 19323 19066
rect 19335 19014 19387 19066
rect 19399 19014 19451 19066
rect 4160 18912 4212 18964
rect 5816 18708 5868 18760
rect 6148 18470 6200 18522
rect 6212 18470 6264 18522
rect 6276 18470 6328 18522
rect 6340 18470 6392 18522
rect 6404 18470 6456 18522
rect 11346 18470 11398 18522
rect 11410 18470 11462 18522
rect 11474 18470 11526 18522
rect 11538 18470 11590 18522
rect 11602 18470 11654 18522
rect 16544 18470 16596 18522
rect 16608 18470 16660 18522
rect 16672 18470 16724 18522
rect 16736 18470 16788 18522
rect 16800 18470 16852 18522
rect 21742 18470 21794 18522
rect 21806 18470 21858 18522
rect 21870 18470 21922 18522
rect 21934 18470 21986 18522
rect 21998 18470 22050 18522
rect 4068 18368 4120 18420
rect 7656 18232 7708 18284
rect 3549 17926 3601 17978
rect 3613 17926 3665 17978
rect 3677 17926 3729 17978
rect 3741 17926 3793 17978
rect 3805 17926 3857 17978
rect 8747 17926 8799 17978
rect 8811 17926 8863 17978
rect 8875 17926 8927 17978
rect 8939 17926 8991 17978
rect 9003 17926 9055 17978
rect 13945 17926 13997 17978
rect 14009 17926 14061 17978
rect 14073 17926 14125 17978
rect 14137 17926 14189 17978
rect 14201 17926 14253 17978
rect 19143 17926 19195 17978
rect 19207 17926 19259 17978
rect 19271 17926 19323 17978
rect 19335 17926 19387 17978
rect 19399 17926 19451 17978
rect 1952 17867 2004 17876
rect 1952 17833 1961 17867
rect 1961 17833 1995 17867
rect 1995 17833 2004 17867
rect 1952 17824 2004 17833
rect 3976 17867 4028 17876
rect 3976 17833 3985 17867
rect 3985 17833 4019 17867
rect 4019 17833 4028 17867
rect 3976 17824 4028 17833
rect 4160 17824 4212 17876
rect 5816 17688 5868 17740
rect 2228 17620 2280 17672
rect 6736 17620 6788 17672
rect 9404 17620 9456 17672
rect 6000 17552 6052 17604
rect 6148 17382 6200 17434
rect 6212 17382 6264 17434
rect 6276 17382 6328 17434
rect 6340 17382 6392 17434
rect 6404 17382 6456 17434
rect 11346 17382 11398 17434
rect 11410 17382 11462 17434
rect 11474 17382 11526 17434
rect 11538 17382 11590 17434
rect 11602 17382 11654 17434
rect 16544 17382 16596 17434
rect 16608 17382 16660 17434
rect 16672 17382 16724 17434
rect 16736 17382 16788 17434
rect 16800 17382 16852 17434
rect 21742 17382 21794 17434
rect 21806 17382 21858 17434
rect 21870 17382 21922 17434
rect 21934 17382 21986 17434
rect 21998 17382 22050 17434
rect 1584 17323 1636 17332
rect 1584 17289 1593 17323
rect 1593 17289 1627 17323
rect 1627 17289 1636 17323
rect 1584 17280 1636 17289
rect 3700 17323 3752 17332
rect 3700 17289 3709 17323
rect 3709 17289 3743 17323
rect 3743 17289 3752 17323
rect 3700 17280 3752 17289
rect 2228 17255 2280 17264
rect 2228 17221 2237 17255
rect 2237 17221 2271 17255
rect 2271 17221 2280 17255
rect 2228 17212 2280 17221
rect 4712 17212 4764 17264
rect 6644 17144 6696 17196
rect 12164 17144 12216 17196
rect 4252 17076 4304 17128
rect 4436 17008 4488 17060
rect 3549 16838 3601 16890
rect 3613 16838 3665 16890
rect 3677 16838 3729 16890
rect 3741 16838 3793 16890
rect 3805 16838 3857 16890
rect 8747 16838 8799 16890
rect 8811 16838 8863 16890
rect 8875 16838 8927 16890
rect 8939 16838 8991 16890
rect 9003 16838 9055 16890
rect 13945 16838 13997 16890
rect 14009 16838 14061 16890
rect 14073 16838 14125 16890
rect 14137 16838 14189 16890
rect 14201 16838 14253 16890
rect 19143 16838 19195 16890
rect 19207 16838 19259 16890
rect 19271 16838 19323 16890
rect 19335 16838 19387 16890
rect 19399 16838 19451 16890
rect 10876 16668 10928 16720
rect 21456 16600 21508 16652
rect 4436 16575 4488 16584
rect 4436 16541 4445 16575
rect 4445 16541 4479 16575
rect 4479 16541 4488 16575
rect 4436 16532 4488 16541
rect 5816 16532 5868 16584
rect 6000 16532 6052 16584
rect 6828 16532 6880 16584
rect 7196 16575 7248 16584
rect 7196 16541 7205 16575
rect 7205 16541 7239 16575
rect 7239 16541 7248 16575
rect 7196 16532 7248 16541
rect 7656 16575 7708 16584
rect 7656 16541 7665 16575
rect 7665 16541 7699 16575
rect 7699 16541 7708 16575
rect 7656 16532 7708 16541
rect 8576 16532 8628 16584
rect 6736 16464 6788 16516
rect 9128 16396 9180 16448
rect 6148 16294 6200 16346
rect 6212 16294 6264 16346
rect 6276 16294 6328 16346
rect 6340 16294 6392 16346
rect 6404 16294 6456 16346
rect 11346 16294 11398 16346
rect 11410 16294 11462 16346
rect 11474 16294 11526 16346
rect 11538 16294 11590 16346
rect 11602 16294 11654 16346
rect 16544 16294 16596 16346
rect 16608 16294 16660 16346
rect 16672 16294 16724 16346
rect 16736 16294 16788 16346
rect 16800 16294 16852 16346
rect 21742 16294 21794 16346
rect 21806 16294 21858 16346
rect 21870 16294 21922 16346
rect 21934 16294 21986 16346
rect 21998 16294 22050 16346
rect 1952 16235 2004 16244
rect 1952 16201 1961 16235
rect 1961 16201 1995 16235
rect 1995 16201 2004 16235
rect 1952 16192 2004 16201
rect 5356 16056 5408 16108
rect 5172 15895 5224 15904
rect 5172 15861 5181 15895
rect 5181 15861 5215 15895
rect 5215 15861 5224 15895
rect 5172 15852 5224 15861
rect 3549 15750 3601 15802
rect 3613 15750 3665 15802
rect 3677 15750 3729 15802
rect 3741 15750 3793 15802
rect 3805 15750 3857 15802
rect 8747 15750 8799 15802
rect 8811 15750 8863 15802
rect 8875 15750 8927 15802
rect 8939 15750 8991 15802
rect 9003 15750 9055 15802
rect 13945 15750 13997 15802
rect 14009 15750 14061 15802
rect 14073 15750 14125 15802
rect 14137 15750 14189 15802
rect 14201 15750 14253 15802
rect 19143 15750 19195 15802
rect 19207 15750 19259 15802
rect 19271 15750 19323 15802
rect 19335 15750 19387 15802
rect 19399 15750 19451 15802
rect 1676 15691 1728 15700
rect 1676 15657 1685 15691
rect 1685 15657 1719 15691
rect 1719 15657 1728 15691
rect 1676 15648 1728 15657
rect 2780 15691 2832 15700
rect 2780 15657 2789 15691
rect 2789 15657 2823 15691
rect 2823 15657 2832 15691
rect 2780 15648 2832 15657
rect 5908 15691 5960 15700
rect 5908 15657 5917 15691
rect 5917 15657 5951 15691
rect 5951 15657 5960 15691
rect 5908 15648 5960 15657
rect 6644 15648 6696 15700
rect 2228 15623 2280 15632
rect 2228 15589 2237 15623
rect 2237 15589 2271 15623
rect 2271 15589 2280 15623
rect 2228 15580 2280 15589
rect 5356 15555 5408 15564
rect 5356 15521 5365 15555
rect 5365 15521 5399 15555
rect 5399 15521 5408 15555
rect 5356 15512 5408 15521
rect 11796 15512 11848 15564
rect 2872 15444 2924 15496
rect 3700 15444 3752 15496
rect 7748 15444 7800 15496
rect 6000 15376 6052 15428
rect 9312 15308 9364 15360
rect 6148 15206 6200 15258
rect 6212 15206 6264 15258
rect 6276 15206 6328 15258
rect 6340 15206 6392 15258
rect 6404 15206 6456 15258
rect 11346 15206 11398 15258
rect 11410 15206 11462 15258
rect 11474 15206 11526 15258
rect 11538 15206 11590 15258
rect 11602 15206 11654 15258
rect 16544 15206 16596 15258
rect 16608 15206 16660 15258
rect 16672 15206 16724 15258
rect 16736 15206 16788 15258
rect 16800 15206 16852 15258
rect 21742 15206 21794 15258
rect 21806 15206 21858 15258
rect 21870 15206 21922 15258
rect 21934 15206 21986 15258
rect 21998 15206 22050 15258
rect 4252 15147 4304 15156
rect 4252 15113 4261 15147
rect 4261 15113 4295 15147
rect 4295 15113 4304 15147
rect 4252 15104 4304 15113
rect 5816 15104 5868 15156
rect 2872 15036 2924 15088
rect 3700 15079 3752 15088
rect 3700 15045 3709 15079
rect 3709 15045 3743 15079
rect 3743 15045 3752 15079
rect 3700 15036 3752 15045
rect 2136 15011 2188 15020
rect 2136 14977 2145 15011
rect 2145 14977 2179 15011
rect 2179 14977 2188 15011
rect 2136 14968 2188 14977
rect 3884 14968 3936 15020
rect 7104 15036 7156 15088
rect 4896 14968 4948 15020
rect 5908 14968 5960 15020
rect 5172 14900 5224 14952
rect 5724 14943 5776 14952
rect 5724 14909 5733 14943
rect 5733 14909 5767 14943
rect 5767 14909 5776 14943
rect 5724 14900 5776 14909
rect 7380 14943 7432 14952
rect 1952 14807 2004 14816
rect 1952 14773 1961 14807
rect 1961 14773 1995 14807
rect 1995 14773 2004 14807
rect 1952 14764 2004 14773
rect 5540 14764 5592 14816
rect 7380 14909 7389 14943
rect 7389 14909 7423 14943
rect 7423 14909 7432 14943
rect 7380 14900 7432 14909
rect 15568 14900 15620 14952
rect 3549 14662 3601 14714
rect 3613 14662 3665 14714
rect 3677 14662 3729 14714
rect 3741 14662 3793 14714
rect 3805 14662 3857 14714
rect 8747 14662 8799 14714
rect 8811 14662 8863 14714
rect 8875 14662 8927 14714
rect 8939 14662 8991 14714
rect 9003 14662 9055 14714
rect 13945 14662 13997 14714
rect 14009 14662 14061 14714
rect 14073 14662 14125 14714
rect 14137 14662 14189 14714
rect 14201 14662 14253 14714
rect 19143 14662 19195 14714
rect 19207 14662 19259 14714
rect 19271 14662 19323 14714
rect 19335 14662 19387 14714
rect 19399 14662 19451 14714
rect 1492 14603 1544 14612
rect 1492 14569 1501 14603
rect 1501 14569 1535 14603
rect 1535 14569 1544 14603
rect 1492 14560 1544 14569
rect 9312 14603 9364 14612
rect 9312 14569 9321 14603
rect 9321 14569 9355 14603
rect 9355 14569 9364 14603
rect 9312 14560 9364 14569
rect 2136 14467 2188 14476
rect 2136 14433 2145 14467
rect 2145 14433 2179 14467
rect 2179 14433 2188 14467
rect 2136 14424 2188 14433
rect 7840 14492 7892 14544
rect 11888 14492 11940 14544
rect 3332 14356 3384 14408
rect 8392 14356 8444 14408
rect 10600 14424 10652 14476
rect 10324 14356 10376 14408
rect 11152 14356 11204 14408
rect 12348 14356 12400 14408
rect 8208 14288 8260 14340
rect 4068 14220 4120 14272
rect 4252 14263 4304 14272
rect 4252 14229 4261 14263
rect 4261 14229 4295 14263
rect 4295 14229 4304 14263
rect 4804 14263 4856 14272
rect 4252 14220 4304 14229
rect 4804 14229 4813 14263
rect 4813 14229 4847 14263
rect 4847 14229 4856 14263
rect 4804 14220 4856 14229
rect 5724 14220 5776 14272
rect 6552 14220 6604 14272
rect 8484 14263 8536 14272
rect 8484 14229 8493 14263
rect 8493 14229 8527 14263
rect 8527 14229 8536 14263
rect 9680 14263 9732 14272
rect 8484 14220 8536 14229
rect 9680 14229 9689 14263
rect 9689 14229 9723 14263
rect 9723 14229 9732 14263
rect 9680 14220 9732 14229
rect 10784 14220 10836 14272
rect 11888 14220 11940 14272
rect 12900 14220 12952 14272
rect 6148 14118 6200 14170
rect 6212 14118 6264 14170
rect 6276 14118 6328 14170
rect 6340 14118 6392 14170
rect 6404 14118 6456 14170
rect 11346 14118 11398 14170
rect 11410 14118 11462 14170
rect 11474 14118 11526 14170
rect 11538 14118 11590 14170
rect 11602 14118 11654 14170
rect 16544 14118 16596 14170
rect 16608 14118 16660 14170
rect 16672 14118 16724 14170
rect 16736 14118 16788 14170
rect 16800 14118 16852 14170
rect 21742 14118 21794 14170
rect 21806 14118 21858 14170
rect 21870 14118 21922 14170
rect 21934 14118 21986 14170
rect 21998 14118 22050 14170
rect 1952 14059 2004 14068
rect 1952 14025 1961 14059
rect 1961 14025 1995 14059
rect 1995 14025 2004 14059
rect 1952 14016 2004 14025
rect 2780 14016 2832 14068
rect 4068 14059 4120 14068
rect 4068 14025 4077 14059
rect 4077 14025 4111 14059
rect 4111 14025 4120 14059
rect 4068 14016 4120 14025
rect 4896 14059 4948 14068
rect 4896 14025 4905 14059
rect 4905 14025 4939 14059
rect 4939 14025 4948 14059
rect 4896 14016 4948 14025
rect 7380 14016 7432 14068
rect 8208 14016 8260 14068
rect 9404 14059 9456 14068
rect 9404 14025 9413 14059
rect 9413 14025 9447 14059
rect 9447 14025 9456 14059
rect 9404 14016 9456 14025
rect 10416 14059 10468 14068
rect 10416 14025 10425 14059
rect 10425 14025 10459 14059
rect 10459 14025 10468 14059
rect 10416 14016 10468 14025
rect 10784 14059 10836 14068
rect 10784 14025 10793 14059
rect 10793 14025 10827 14059
rect 10827 14025 10836 14059
rect 10784 14016 10836 14025
rect 2412 13923 2464 13932
rect 2412 13889 2421 13923
rect 2421 13889 2455 13923
rect 2455 13889 2464 13923
rect 2412 13880 2464 13889
rect 4804 13948 4856 14000
rect 6184 13948 6236 14000
rect 7656 13991 7708 14000
rect 7656 13957 7665 13991
rect 7665 13957 7699 13991
rect 7699 13957 7708 13991
rect 7656 13948 7708 13957
rect 3148 13812 3200 13864
rect 5264 13923 5316 13932
rect 5264 13889 5273 13923
rect 5273 13889 5307 13923
rect 5307 13889 5316 13923
rect 5264 13880 5316 13889
rect 9772 13923 9824 13932
rect 9772 13889 9781 13923
rect 9781 13889 9815 13923
rect 9815 13889 9824 13923
rect 9772 13880 9824 13889
rect 12900 14059 12952 14068
rect 12900 14025 12909 14059
rect 12909 14025 12943 14059
rect 12943 14025 12952 14059
rect 12900 14016 12952 14025
rect 11888 13991 11940 14000
rect 11888 13957 11897 13991
rect 11897 13957 11931 13991
rect 11931 13957 11940 13991
rect 11888 13948 11940 13957
rect 12348 13948 12400 14000
rect 5540 13855 5592 13864
rect 5540 13821 5549 13855
rect 5549 13821 5583 13855
rect 5583 13821 5592 13855
rect 5540 13812 5592 13821
rect 6644 13855 6696 13864
rect 6644 13821 6653 13855
rect 6653 13821 6687 13855
rect 6687 13821 6696 13855
rect 6644 13812 6696 13821
rect 9036 13855 9088 13864
rect 2136 13676 2188 13728
rect 4804 13744 4856 13796
rect 9036 13821 9045 13855
rect 9045 13821 9079 13855
rect 9079 13821 9088 13855
rect 9036 13812 9088 13821
rect 11980 13855 12032 13864
rect 9956 13744 10008 13796
rect 10140 13744 10192 13796
rect 11980 13821 11989 13855
rect 11989 13821 12023 13855
rect 12023 13821 12032 13855
rect 11980 13812 12032 13821
rect 3240 13676 3292 13728
rect 8484 13676 8536 13728
rect 13084 13676 13136 13728
rect 19984 13744 20036 13796
rect 15660 13676 15712 13728
rect 3549 13574 3601 13626
rect 3613 13574 3665 13626
rect 3677 13574 3729 13626
rect 3741 13574 3793 13626
rect 3805 13574 3857 13626
rect 8747 13574 8799 13626
rect 8811 13574 8863 13626
rect 8875 13574 8927 13626
rect 8939 13574 8991 13626
rect 9003 13574 9055 13626
rect 13945 13574 13997 13626
rect 14009 13574 14061 13626
rect 14073 13574 14125 13626
rect 14137 13574 14189 13626
rect 14201 13574 14253 13626
rect 19143 13574 19195 13626
rect 19207 13574 19259 13626
rect 19271 13574 19323 13626
rect 19335 13574 19387 13626
rect 19399 13574 19451 13626
rect 4252 13472 4304 13524
rect 7196 13472 7248 13524
rect 10876 13472 10928 13524
rect 1952 13379 2004 13388
rect 1952 13345 1961 13379
rect 1961 13345 1995 13379
rect 1995 13345 2004 13379
rect 1952 13336 2004 13345
rect 1492 13200 1544 13252
rect 2136 13243 2188 13252
rect 2136 13209 2145 13243
rect 2145 13209 2179 13243
rect 2179 13209 2188 13243
rect 2136 13200 2188 13209
rect 1584 13132 1636 13184
rect 3148 13379 3200 13388
rect 3148 13345 3157 13379
rect 3157 13345 3191 13379
rect 3191 13345 3200 13379
rect 3148 13336 3200 13345
rect 4804 13379 4856 13388
rect 4804 13345 4813 13379
rect 4813 13345 4847 13379
rect 4847 13345 4856 13379
rect 4804 13336 4856 13345
rect 5264 13336 5316 13388
rect 7656 13404 7708 13456
rect 6552 13336 6604 13388
rect 8300 13379 8352 13388
rect 8300 13345 8309 13379
rect 8309 13345 8343 13379
rect 8343 13345 8352 13379
rect 9772 13379 9824 13388
rect 8300 13336 8352 13345
rect 9772 13345 9781 13379
rect 9781 13345 9815 13379
rect 9815 13345 9824 13379
rect 9772 13336 9824 13345
rect 10876 13379 10928 13388
rect 10876 13345 10885 13379
rect 10885 13345 10919 13379
rect 10919 13345 10928 13379
rect 10876 13336 10928 13345
rect 17960 13336 18012 13388
rect 4528 13268 4580 13320
rect 6184 13311 6236 13320
rect 6184 13277 6193 13311
rect 6193 13277 6227 13311
rect 6227 13277 6236 13311
rect 6184 13268 6236 13277
rect 10692 13268 10744 13320
rect 11704 13268 11756 13320
rect 4068 13200 4120 13252
rect 2504 13175 2556 13184
rect 2504 13141 2513 13175
rect 2513 13141 2547 13175
rect 2547 13141 2556 13175
rect 2504 13132 2556 13141
rect 5908 13200 5960 13252
rect 10508 13200 10560 13252
rect 11980 13200 12032 13252
rect 4988 13132 5040 13184
rect 5816 13175 5868 13184
rect 5816 13141 5825 13175
rect 5825 13141 5859 13175
rect 5859 13141 5868 13175
rect 5816 13132 5868 13141
rect 7932 13132 7984 13184
rect 10692 13175 10744 13184
rect 10692 13141 10701 13175
rect 10701 13141 10735 13175
rect 10735 13141 10744 13175
rect 10692 13132 10744 13141
rect 12072 13132 12124 13184
rect 6148 13030 6200 13082
rect 6212 13030 6264 13082
rect 6276 13030 6328 13082
rect 6340 13030 6392 13082
rect 6404 13030 6456 13082
rect 11346 13030 11398 13082
rect 11410 13030 11462 13082
rect 11474 13030 11526 13082
rect 11538 13030 11590 13082
rect 11602 13030 11654 13082
rect 16544 13030 16596 13082
rect 16608 13030 16660 13082
rect 16672 13030 16724 13082
rect 16736 13030 16788 13082
rect 16800 13030 16852 13082
rect 21742 13030 21794 13082
rect 21806 13030 21858 13082
rect 21870 13030 21922 13082
rect 21934 13030 21986 13082
rect 21998 13030 22050 13082
rect 2780 12928 2832 12980
rect 7656 12928 7708 12980
rect 7840 12928 7892 12980
rect 2412 12860 2464 12912
rect 4804 12860 4856 12912
rect 9680 12928 9732 12980
rect 11704 12971 11756 12980
rect 11704 12937 11713 12971
rect 11713 12937 11747 12971
rect 11747 12937 11756 12971
rect 11704 12928 11756 12937
rect 12164 12971 12216 12980
rect 12164 12937 12173 12971
rect 12173 12937 12207 12971
rect 12207 12937 12216 12971
rect 12164 12928 12216 12937
rect 11980 12860 12032 12912
rect 1768 12835 1820 12844
rect 1768 12801 1777 12835
rect 1777 12801 1811 12835
rect 1811 12801 1820 12835
rect 1768 12792 1820 12801
rect 2320 12792 2372 12844
rect 4344 12792 4396 12844
rect 7932 12792 7984 12844
rect 3240 12767 3292 12776
rect 3240 12733 3249 12767
rect 3249 12733 3283 12767
rect 3283 12733 3292 12767
rect 3240 12724 3292 12733
rect 5724 12767 5776 12776
rect 5724 12733 5733 12767
rect 5733 12733 5767 12767
rect 5767 12733 5776 12767
rect 5724 12724 5776 12733
rect 7104 12767 7156 12776
rect 5632 12656 5684 12708
rect 7104 12733 7113 12767
rect 7113 12733 7147 12767
rect 7147 12733 7156 12767
rect 7104 12724 7156 12733
rect 8024 12767 8076 12776
rect 8024 12733 8033 12767
rect 8033 12733 8067 12767
rect 8067 12733 8076 12767
rect 8024 12724 8076 12733
rect 9128 12792 9180 12844
rect 10232 12724 10284 12776
rect 1492 12631 1544 12640
rect 1492 12597 1501 12631
rect 1501 12597 1535 12631
rect 1535 12597 1544 12631
rect 1492 12588 1544 12597
rect 4988 12631 5040 12640
rect 4988 12597 4997 12631
rect 4997 12597 5031 12631
rect 5031 12597 5040 12631
rect 4988 12588 5040 12597
rect 5264 12631 5316 12640
rect 5264 12597 5273 12631
rect 5273 12597 5307 12631
rect 5307 12597 5316 12631
rect 5264 12588 5316 12597
rect 6368 12588 6420 12640
rect 7656 12588 7708 12640
rect 8116 12588 8168 12640
rect 9128 12631 9180 12640
rect 9128 12597 9137 12631
rect 9137 12597 9171 12631
rect 9171 12597 9180 12631
rect 9128 12588 9180 12597
rect 17132 12724 17184 12776
rect 12716 12588 12768 12640
rect 3549 12486 3601 12538
rect 3613 12486 3665 12538
rect 3677 12486 3729 12538
rect 3741 12486 3793 12538
rect 3805 12486 3857 12538
rect 8747 12486 8799 12538
rect 8811 12486 8863 12538
rect 8875 12486 8927 12538
rect 8939 12486 8991 12538
rect 9003 12486 9055 12538
rect 13945 12486 13997 12538
rect 14009 12486 14061 12538
rect 14073 12486 14125 12538
rect 14137 12486 14189 12538
rect 14201 12486 14253 12538
rect 19143 12486 19195 12538
rect 19207 12486 19259 12538
rect 19271 12486 19323 12538
rect 19335 12486 19387 12538
rect 19399 12486 19451 12538
rect 1676 12427 1728 12436
rect 1676 12393 1685 12427
rect 1685 12393 1719 12427
rect 1719 12393 1728 12427
rect 1676 12384 1728 12393
rect 4344 12427 4396 12436
rect 4344 12393 4353 12427
rect 4353 12393 4387 12427
rect 4387 12393 4396 12427
rect 4344 12384 4396 12393
rect 5172 12384 5224 12436
rect 5448 12384 5500 12436
rect 5724 12384 5776 12436
rect 6368 12384 6420 12436
rect 6828 12427 6880 12436
rect 6828 12393 6837 12427
rect 6837 12393 6871 12427
rect 6871 12393 6880 12427
rect 6828 12384 6880 12393
rect 2688 12316 2740 12368
rect 1952 12248 2004 12300
rect 2412 12248 2464 12300
rect 5172 12248 5224 12300
rect 6552 12316 6604 12368
rect 8024 12384 8076 12436
rect 8300 12316 8352 12368
rect 8576 12384 8628 12436
rect 9956 12384 10008 12436
rect 13176 12384 13228 12436
rect 7472 12291 7524 12300
rect 7472 12257 7481 12291
rect 7481 12257 7515 12291
rect 7515 12257 7524 12291
rect 7472 12248 7524 12257
rect 8024 12248 8076 12300
rect 8208 12248 8260 12300
rect 8576 12248 8628 12300
rect 9588 12248 9640 12300
rect 10416 12248 10468 12300
rect 10876 12291 10928 12300
rect 10876 12257 10885 12291
rect 10885 12257 10919 12291
rect 10919 12257 10928 12291
rect 10876 12248 10928 12257
rect 3240 12180 3292 12232
rect 5264 12180 5316 12232
rect 5908 12180 5960 12232
rect 7104 12180 7156 12232
rect 8116 12180 8168 12232
rect 10048 12180 10100 12232
rect 10140 12180 10192 12232
rect 11796 12223 11848 12232
rect 11796 12189 11805 12223
rect 11805 12189 11839 12223
rect 11839 12189 11848 12223
rect 11796 12180 11848 12189
rect 7656 12112 7708 12164
rect 11704 12112 11756 12164
rect 12348 12112 12400 12164
rect 1400 12044 1452 12096
rect 2688 12044 2740 12096
rect 2872 12087 2924 12096
rect 2872 12053 2881 12087
rect 2881 12053 2915 12087
rect 2915 12053 2924 12087
rect 2872 12044 2924 12053
rect 3056 12044 3108 12096
rect 3976 12087 4028 12096
rect 3976 12053 3985 12087
rect 3985 12053 4019 12087
rect 4019 12053 4028 12087
rect 3976 12044 4028 12053
rect 4712 12087 4764 12096
rect 4712 12053 4721 12087
rect 4721 12053 4755 12087
rect 4755 12053 4764 12087
rect 4712 12044 4764 12053
rect 5356 12087 5408 12096
rect 5356 12053 5365 12087
rect 5365 12053 5399 12087
rect 5399 12053 5408 12087
rect 5356 12044 5408 12053
rect 6644 12044 6696 12096
rect 7380 12044 7432 12096
rect 8208 12087 8260 12096
rect 8208 12053 8217 12087
rect 8217 12053 8251 12087
rect 8251 12053 8260 12087
rect 8208 12044 8260 12053
rect 10416 12044 10468 12096
rect 13176 12087 13228 12096
rect 13176 12053 13185 12087
rect 13185 12053 13219 12087
rect 13219 12053 13228 12087
rect 13176 12044 13228 12053
rect 13728 12044 13780 12096
rect 15660 12087 15712 12096
rect 15660 12053 15669 12087
rect 15669 12053 15703 12087
rect 15703 12053 15712 12087
rect 15660 12044 15712 12053
rect 17132 12112 17184 12164
rect 17040 12044 17092 12096
rect 18328 12044 18380 12096
rect 21364 12087 21416 12096
rect 21364 12053 21373 12087
rect 21373 12053 21407 12087
rect 21407 12053 21416 12087
rect 21364 12044 21416 12053
rect 6148 11942 6200 11994
rect 6212 11942 6264 11994
rect 6276 11942 6328 11994
rect 6340 11942 6392 11994
rect 6404 11942 6456 11994
rect 11346 11942 11398 11994
rect 11410 11942 11462 11994
rect 11474 11942 11526 11994
rect 11538 11942 11590 11994
rect 11602 11942 11654 11994
rect 16544 11942 16596 11994
rect 16608 11942 16660 11994
rect 16672 11942 16724 11994
rect 16736 11942 16788 11994
rect 16800 11942 16852 11994
rect 21742 11942 21794 11994
rect 21806 11942 21858 11994
rect 21870 11942 21922 11994
rect 21934 11942 21986 11994
rect 21998 11942 22050 11994
rect 2872 11840 2924 11892
rect 3976 11840 4028 11892
rect 4712 11840 4764 11892
rect 5356 11883 5408 11892
rect 5356 11849 5365 11883
rect 5365 11849 5399 11883
rect 5399 11849 5408 11883
rect 5356 11840 5408 11849
rect 5816 11840 5868 11892
rect 6000 11840 6052 11892
rect 7380 11840 7432 11892
rect 7748 11883 7800 11892
rect 7748 11849 7757 11883
rect 7757 11849 7791 11883
rect 7791 11849 7800 11883
rect 7748 11840 7800 11849
rect 2320 11772 2372 11824
rect 2412 11772 2464 11824
rect 1860 11747 1912 11756
rect 1860 11713 1869 11747
rect 1869 11713 1903 11747
rect 1903 11713 1912 11747
rect 1860 11704 1912 11713
rect 2688 11679 2740 11688
rect 2688 11645 2697 11679
rect 2697 11645 2731 11679
rect 2731 11645 2740 11679
rect 2688 11636 2740 11645
rect 8392 11772 8444 11824
rect 11704 11840 11756 11892
rect 13176 11840 13228 11892
rect 15568 11883 15620 11892
rect 6736 11747 6788 11756
rect 6736 11713 6745 11747
rect 6745 11713 6779 11747
rect 6779 11713 6788 11747
rect 6736 11704 6788 11713
rect 8668 11704 8720 11756
rect 5632 11679 5684 11688
rect 5632 11645 5641 11679
rect 5641 11645 5675 11679
rect 5675 11645 5684 11679
rect 5632 11636 5684 11645
rect 10784 11772 10836 11824
rect 11336 11772 11388 11824
rect 9128 11747 9180 11756
rect 9128 11713 9137 11747
rect 9137 11713 9171 11747
rect 9171 11713 9180 11747
rect 9128 11704 9180 11713
rect 5356 11568 5408 11620
rect 9312 11636 9364 11688
rect 11704 11704 11756 11756
rect 9956 11568 10008 11620
rect 2228 11500 2280 11552
rect 7380 11543 7432 11552
rect 7380 11509 7389 11543
rect 7389 11509 7423 11543
rect 7423 11509 7432 11543
rect 7380 11500 7432 11509
rect 7932 11500 7984 11552
rect 9128 11500 9180 11552
rect 10784 11500 10836 11552
rect 11796 11636 11848 11688
rect 12348 11747 12400 11756
rect 12348 11713 12382 11747
rect 12382 11713 12400 11747
rect 12348 11704 12400 11713
rect 13728 11704 13780 11756
rect 15568 11849 15577 11883
rect 15577 11849 15611 11883
rect 15611 11849 15620 11883
rect 15568 11840 15620 11849
rect 19984 11883 20036 11892
rect 19984 11849 19993 11883
rect 19993 11849 20027 11883
rect 20027 11849 20036 11883
rect 19984 11840 20036 11849
rect 16488 11772 16540 11824
rect 18604 11815 18656 11824
rect 18604 11781 18638 11815
rect 18638 11781 18656 11815
rect 18604 11772 18656 11781
rect 16120 11704 16172 11756
rect 21088 11747 21140 11756
rect 21088 11713 21106 11747
rect 21106 11713 21140 11747
rect 21364 11747 21416 11756
rect 21088 11704 21140 11713
rect 21364 11713 21373 11747
rect 21373 11713 21407 11747
rect 21407 11713 21416 11747
rect 21364 11704 21416 11713
rect 18328 11679 18380 11688
rect 18328 11645 18337 11679
rect 18337 11645 18371 11679
rect 18371 11645 18380 11679
rect 18328 11636 18380 11645
rect 11336 11500 11388 11552
rect 13452 11543 13504 11552
rect 13452 11509 13461 11543
rect 13461 11509 13495 11543
rect 13495 11509 13504 11543
rect 13728 11543 13780 11552
rect 13452 11500 13504 11509
rect 13728 11509 13737 11543
rect 13737 11509 13771 11543
rect 13771 11509 13780 11543
rect 13728 11500 13780 11509
rect 18052 11543 18104 11552
rect 18052 11509 18061 11543
rect 18061 11509 18095 11543
rect 18095 11509 18104 11543
rect 18052 11500 18104 11509
rect 20628 11500 20680 11552
rect 3549 11398 3601 11450
rect 3613 11398 3665 11450
rect 3677 11398 3729 11450
rect 3741 11398 3793 11450
rect 3805 11398 3857 11450
rect 8747 11398 8799 11450
rect 8811 11398 8863 11450
rect 8875 11398 8927 11450
rect 8939 11398 8991 11450
rect 9003 11398 9055 11450
rect 13945 11398 13997 11450
rect 14009 11398 14061 11450
rect 14073 11398 14125 11450
rect 14137 11398 14189 11450
rect 14201 11398 14253 11450
rect 19143 11398 19195 11450
rect 19207 11398 19259 11450
rect 19271 11398 19323 11450
rect 19335 11398 19387 11450
rect 19399 11398 19451 11450
rect 1768 11339 1820 11348
rect 1768 11305 1777 11339
rect 1777 11305 1811 11339
rect 1811 11305 1820 11339
rect 1768 11296 1820 11305
rect 3148 11296 3200 11348
rect 4528 11339 4580 11348
rect 4528 11305 4537 11339
rect 4537 11305 4571 11339
rect 4571 11305 4580 11339
rect 4528 11296 4580 11305
rect 8208 11296 8260 11348
rect 8392 11296 8444 11348
rect 2228 11203 2280 11212
rect 2228 11169 2237 11203
rect 2237 11169 2271 11203
rect 2271 11169 2280 11203
rect 2228 11160 2280 11169
rect 2412 11203 2464 11212
rect 2412 11169 2421 11203
rect 2421 11169 2455 11203
rect 2455 11169 2464 11203
rect 2412 11160 2464 11169
rect 5632 11160 5684 11212
rect 5724 11160 5776 11212
rect 6184 11203 6236 11212
rect 6184 11169 6193 11203
rect 6193 11169 6227 11203
rect 6227 11169 6236 11203
rect 6184 11160 6236 11169
rect 6736 11203 6788 11212
rect 6736 11169 6745 11203
rect 6745 11169 6779 11203
rect 6779 11169 6788 11203
rect 6736 11160 6788 11169
rect 4068 11092 4120 11144
rect 1400 11067 1452 11076
rect 1400 11033 1409 11067
rect 1409 11033 1443 11067
rect 1443 11033 1452 11067
rect 1400 11024 1452 11033
rect 3424 11024 3476 11076
rect 4344 11024 4396 11076
rect 7932 11228 7984 11280
rect 8392 11203 8444 11212
rect 8392 11169 8401 11203
rect 8401 11169 8435 11203
rect 8435 11169 8444 11203
rect 8392 11160 8444 11169
rect 8668 11160 8720 11212
rect 11888 11296 11940 11348
rect 13820 11296 13872 11348
rect 15476 11296 15528 11348
rect 16488 11296 16540 11348
rect 19524 11296 19576 11348
rect 20720 11296 20772 11348
rect 14464 11271 14516 11280
rect 14464 11237 14473 11271
rect 14473 11237 14507 11271
rect 14507 11237 14516 11271
rect 14464 11228 14516 11237
rect 10048 11092 10100 11144
rect 10784 11092 10836 11144
rect 21364 11296 21416 11348
rect 13728 11135 13780 11144
rect 13728 11101 13737 11135
rect 13737 11101 13771 11135
rect 13771 11101 13780 11135
rect 13728 11092 13780 11101
rect 7472 11024 7524 11076
rect 8392 11024 8444 11076
rect 9312 11024 9364 11076
rect 10140 11067 10192 11076
rect 10140 11033 10149 11067
rect 10149 11033 10183 11067
rect 10183 11033 10192 11067
rect 10140 11024 10192 11033
rect 10600 11024 10652 11076
rect 13360 11024 13412 11076
rect 2136 10999 2188 11008
rect 2136 10965 2145 10999
rect 2145 10965 2179 10999
rect 2179 10965 2188 10999
rect 2136 10956 2188 10965
rect 2780 10999 2832 11008
rect 2780 10965 2789 10999
rect 2789 10965 2823 10999
rect 2823 10965 2832 10999
rect 3884 10999 3936 11008
rect 2780 10956 2832 10965
rect 3884 10965 3893 10999
rect 3893 10965 3927 10999
rect 3927 10965 3936 10999
rect 3884 10956 3936 10965
rect 4896 10999 4948 11008
rect 4896 10965 4905 10999
rect 4905 10965 4939 10999
rect 4939 10965 4948 10999
rect 4896 10956 4948 10965
rect 6000 10999 6052 11008
rect 6000 10965 6009 10999
rect 6009 10965 6043 10999
rect 6043 10965 6052 10999
rect 6000 10956 6052 10965
rect 6184 10956 6236 11008
rect 11060 10956 11112 11008
rect 12256 10956 12308 11008
rect 16120 11135 16172 11144
rect 16120 11101 16129 11135
rect 16129 11101 16163 11135
rect 16163 11101 16172 11135
rect 16120 11092 16172 11101
rect 15568 11067 15620 11076
rect 15568 11033 15586 11067
rect 15586 11033 15620 11067
rect 15568 11024 15620 11033
rect 19984 11092 20036 11144
rect 14464 10956 14516 11008
rect 16304 10956 16356 11008
rect 18328 10956 18380 11008
rect 19800 10956 19852 11008
rect 6148 10854 6200 10906
rect 6212 10854 6264 10906
rect 6276 10854 6328 10906
rect 6340 10854 6392 10906
rect 6404 10854 6456 10906
rect 11346 10854 11398 10906
rect 11410 10854 11462 10906
rect 11474 10854 11526 10906
rect 11538 10854 11590 10906
rect 11602 10854 11654 10906
rect 16544 10854 16596 10906
rect 16608 10854 16660 10906
rect 16672 10854 16724 10906
rect 16736 10854 16788 10906
rect 16800 10854 16852 10906
rect 21742 10854 21794 10906
rect 21806 10854 21858 10906
rect 21870 10854 21922 10906
rect 21934 10854 21986 10906
rect 21998 10854 22050 10906
rect 2136 10752 2188 10804
rect 2780 10752 2832 10804
rect 3884 10795 3936 10804
rect 3884 10761 3893 10795
rect 3893 10761 3927 10795
rect 3927 10761 3936 10795
rect 3884 10752 3936 10761
rect 4896 10752 4948 10804
rect 7472 10752 7524 10804
rect 10048 10795 10100 10804
rect 10048 10761 10057 10795
rect 10057 10761 10091 10795
rect 10091 10761 10100 10795
rect 10048 10752 10100 10761
rect 10784 10752 10836 10804
rect 2504 10684 2556 10736
rect 3148 10684 3200 10736
rect 2688 10548 2740 10600
rect 5724 10684 5776 10736
rect 8208 10684 8260 10736
rect 8576 10684 8628 10736
rect 16304 10752 16356 10804
rect 18604 10752 18656 10804
rect 4896 10591 4948 10600
rect 4896 10557 4905 10591
rect 4905 10557 4939 10591
rect 4939 10557 4948 10591
rect 4896 10548 4948 10557
rect 4528 10480 4580 10532
rect 3424 10412 3476 10464
rect 15660 10684 15712 10736
rect 8944 10616 8996 10668
rect 15476 10616 15528 10668
rect 15568 10616 15620 10668
rect 16948 10616 17000 10668
rect 19432 10659 19484 10668
rect 19800 10684 19852 10736
rect 19432 10625 19450 10659
rect 19450 10625 19484 10659
rect 19432 10616 19484 10625
rect 20628 10616 20680 10668
rect 21364 10659 21416 10668
rect 21364 10625 21373 10659
rect 21373 10625 21407 10659
rect 21407 10625 21416 10659
rect 21364 10616 21416 10625
rect 14464 10591 14516 10600
rect 5540 10480 5592 10532
rect 8392 10480 8444 10532
rect 14464 10557 14473 10591
rect 14473 10557 14507 10591
rect 14507 10557 14516 10591
rect 14464 10548 14516 10557
rect 16120 10591 16172 10600
rect 16120 10557 16129 10591
rect 16129 10557 16163 10591
rect 16163 10557 16172 10591
rect 16120 10548 16172 10557
rect 9864 10480 9916 10532
rect 9956 10480 10008 10532
rect 12624 10480 12676 10532
rect 19984 10523 20036 10532
rect 5724 10455 5776 10464
rect 5724 10421 5733 10455
rect 5733 10421 5767 10455
rect 5767 10421 5776 10455
rect 5724 10412 5776 10421
rect 5816 10412 5868 10464
rect 7380 10412 7432 10464
rect 7932 10412 7984 10464
rect 12440 10412 12492 10464
rect 13084 10455 13136 10464
rect 13084 10421 13093 10455
rect 13093 10421 13127 10455
rect 13127 10421 13136 10455
rect 13084 10412 13136 10421
rect 19984 10489 19993 10523
rect 19993 10489 20027 10523
rect 20027 10489 20036 10523
rect 19984 10480 20036 10489
rect 3549 10310 3601 10362
rect 3613 10310 3665 10362
rect 3677 10310 3729 10362
rect 3741 10310 3793 10362
rect 3805 10310 3857 10362
rect 8747 10310 8799 10362
rect 8811 10310 8863 10362
rect 8875 10310 8927 10362
rect 8939 10310 8991 10362
rect 9003 10310 9055 10362
rect 13945 10310 13997 10362
rect 14009 10310 14061 10362
rect 14073 10310 14125 10362
rect 14137 10310 14189 10362
rect 14201 10310 14253 10362
rect 19143 10310 19195 10362
rect 19207 10310 19259 10362
rect 19271 10310 19323 10362
rect 19335 10310 19387 10362
rect 19399 10310 19451 10362
rect 2872 10208 2924 10260
rect 3424 10251 3476 10260
rect 3424 10217 3433 10251
rect 3433 10217 3467 10251
rect 3467 10217 3476 10251
rect 3424 10208 3476 10217
rect 3700 10072 3752 10124
rect 5816 10208 5868 10260
rect 6000 10208 6052 10260
rect 7472 10251 7524 10260
rect 7472 10217 7481 10251
rect 7481 10217 7515 10251
rect 7515 10217 7524 10251
rect 7472 10208 7524 10217
rect 8300 10208 8352 10260
rect 12440 10251 12492 10260
rect 2872 10004 2924 10056
rect 5264 10072 5316 10124
rect 7748 10140 7800 10192
rect 8024 10140 8076 10192
rect 5632 10072 5684 10124
rect 5816 10004 5868 10056
rect 3056 9936 3108 9988
rect 7840 10004 7892 10056
rect 9496 10115 9548 10124
rect 9496 10081 9505 10115
rect 9505 10081 9539 10115
rect 9539 10081 9548 10115
rect 9496 10072 9548 10081
rect 9680 10072 9732 10124
rect 12440 10217 12449 10251
rect 12449 10217 12483 10251
rect 12483 10217 12492 10251
rect 12440 10208 12492 10217
rect 13268 10208 13320 10260
rect 14464 10208 14516 10260
rect 16120 10208 16172 10260
rect 17132 10208 17184 10260
rect 21364 10251 21416 10260
rect 21364 10217 21373 10251
rect 21373 10217 21407 10251
rect 21407 10217 21416 10251
rect 21364 10208 21416 10217
rect 3608 9868 3660 9920
rect 4068 9868 4120 9920
rect 4436 9911 4488 9920
rect 4436 9877 4445 9911
rect 4445 9877 4479 9911
rect 4479 9877 4488 9911
rect 4436 9868 4488 9877
rect 4620 9868 4672 9920
rect 5540 9868 5592 9920
rect 5724 9868 5776 9920
rect 6828 9868 6880 9920
rect 10876 10004 10928 10056
rect 11060 9979 11112 9988
rect 7840 9911 7892 9920
rect 7840 9877 7849 9911
rect 7849 9877 7883 9911
rect 7883 9877 7892 9911
rect 7840 9868 7892 9877
rect 9128 9868 9180 9920
rect 9404 9911 9456 9920
rect 9404 9877 9413 9911
rect 9413 9877 9447 9911
rect 9447 9877 9456 9911
rect 9404 9868 9456 9877
rect 11060 9945 11094 9979
rect 11094 9945 11112 9979
rect 11060 9936 11112 9945
rect 11888 9936 11940 9988
rect 12716 9936 12768 9988
rect 18420 9979 18472 9988
rect 18420 9945 18438 9979
rect 18438 9945 18472 9979
rect 18420 9936 18472 9945
rect 19340 10004 19392 10056
rect 19800 10004 19852 10056
rect 19432 9936 19484 9988
rect 12256 9868 12308 9920
rect 20628 9911 20680 9920
rect 20628 9877 20637 9911
rect 20637 9877 20671 9911
rect 20671 9877 20680 9911
rect 20628 9868 20680 9877
rect 21088 9868 21140 9920
rect 6148 9766 6200 9818
rect 6212 9766 6264 9818
rect 6276 9766 6328 9818
rect 6340 9766 6392 9818
rect 6404 9766 6456 9818
rect 11346 9766 11398 9818
rect 11410 9766 11462 9818
rect 11474 9766 11526 9818
rect 11538 9766 11590 9818
rect 11602 9766 11654 9818
rect 16544 9766 16596 9818
rect 16608 9766 16660 9818
rect 16672 9766 16724 9818
rect 16736 9766 16788 9818
rect 16800 9766 16852 9818
rect 21742 9766 21794 9818
rect 21806 9766 21858 9818
rect 21870 9766 21922 9818
rect 21934 9766 21986 9818
rect 21998 9766 22050 9818
rect 3240 9664 3292 9716
rect 3424 9664 3476 9716
rect 3608 9664 3660 9716
rect 4620 9664 4672 9716
rect 3976 9596 4028 9648
rect 9680 9664 9732 9716
rect 11704 9664 11756 9716
rect 19432 9664 19484 9716
rect 21364 9707 21416 9716
rect 21364 9673 21373 9707
rect 21373 9673 21407 9707
rect 21407 9673 21416 9707
rect 21364 9664 21416 9673
rect 7840 9596 7892 9648
rect 9864 9639 9916 9648
rect 9864 9605 9873 9639
rect 9873 9605 9907 9639
rect 9907 9605 9916 9639
rect 9864 9596 9916 9605
rect 3240 9528 3292 9580
rect 4252 9528 4304 9580
rect 5724 9528 5776 9580
rect 6736 9571 6788 9580
rect 6736 9537 6745 9571
rect 6745 9537 6779 9571
rect 6779 9537 6788 9571
rect 6736 9528 6788 9537
rect 2228 9460 2280 9512
rect 3608 9460 3660 9512
rect 3976 9503 4028 9512
rect 3976 9469 3985 9503
rect 3985 9469 4019 9503
rect 4019 9469 4028 9503
rect 3976 9460 4028 9469
rect 4068 9503 4120 9512
rect 4068 9469 4077 9503
rect 4077 9469 4111 9503
rect 4111 9469 4120 9503
rect 5080 9503 5132 9512
rect 4068 9460 4120 9469
rect 5080 9469 5089 9503
rect 5089 9469 5123 9503
rect 5123 9469 5132 9503
rect 5080 9460 5132 9469
rect 5264 9503 5316 9512
rect 5264 9469 5273 9503
rect 5273 9469 5307 9503
rect 5307 9469 5316 9503
rect 5264 9460 5316 9469
rect 6552 9460 6604 9512
rect 12532 9596 12584 9648
rect 12624 9639 12676 9648
rect 12624 9605 12642 9639
rect 12642 9605 12676 9639
rect 12624 9596 12676 9605
rect 10784 9571 10836 9580
rect 10784 9537 10793 9571
rect 10793 9537 10827 9571
rect 10827 9537 10836 9571
rect 10784 9528 10836 9537
rect 10968 9528 11020 9580
rect 11704 9528 11756 9580
rect 11060 9503 11112 9512
rect 1860 9392 1912 9444
rect 3792 9392 3844 9444
rect 2872 9324 2924 9376
rect 3700 9324 3752 9376
rect 4712 9324 4764 9376
rect 5816 9324 5868 9376
rect 7196 9392 7248 9444
rect 11060 9469 11069 9503
rect 11069 9469 11103 9503
rect 11103 9469 11112 9503
rect 11060 9460 11112 9469
rect 13268 9596 13320 9648
rect 18052 9596 18104 9648
rect 19984 9596 20036 9648
rect 8392 9324 8444 9376
rect 9220 9324 9272 9376
rect 19340 9528 19392 9580
rect 17040 9435 17092 9444
rect 17040 9401 17049 9435
rect 17049 9401 17083 9435
rect 17083 9401 17092 9435
rect 17040 9392 17092 9401
rect 13268 9367 13320 9376
rect 13268 9333 13277 9367
rect 13277 9333 13311 9367
rect 13311 9333 13320 9367
rect 13268 9324 13320 9333
rect 3549 9222 3601 9274
rect 3613 9222 3665 9274
rect 3677 9222 3729 9274
rect 3741 9222 3793 9274
rect 3805 9222 3857 9274
rect 8747 9222 8799 9274
rect 8811 9222 8863 9274
rect 8875 9222 8927 9274
rect 8939 9222 8991 9274
rect 9003 9222 9055 9274
rect 13945 9222 13997 9274
rect 14009 9222 14061 9274
rect 14073 9222 14125 9274
rect 14137 9222 14189 9274
rect 14201 9222 14253 9274
rect 19143 9222 19195 9274
rect 19207 9222 19259 9274
rect 19271 9222 19323 9274
rect 19335 9222 19387 9274
rect 19399 9222 19451 9274
rect 3240 9163 3292 9172
rect 3240 9129 3249 9163
rect 3249 9129 3283 9163
rect 3283 9129 3292 9163
rect 3240 9120 3292 9129
rect 3976 9120 4028 9172
rect 4896 9120 4948 9172
rect 16948 9120 17000 9172
rect 18420 9120 18472 9172
rect 2780 9052 2832 9104
rect 3148 9052 3200 9104
rect 4712 9027 4764 9036
rect 4712 8993 4721 9027
rect 4721 8993 4755 9027
rect 4755 8993 4764 9027
rect 4712 8984 4764 8993
rect 5724 9052 5776 9104
rect 4988 8984 5040 9036
rect 6736 8984 6788 9036
rect 1216 8848 1268 8900
rect 4252 8916 4304 8968
rect 4436 8916 4488 8968
rect 4068 8848 4120 8900
rect 7472 8916 7524 8968
rect 12992 9052 13044 9104
rect 14556 9052 14608 9104
rect 9772 8984 9824 9036
rect 12900 8984 12952 9036
rect 9128 8916 9180 8968
rect 10324 8916 10376 8968
rect 10876 8959 10928 8968
rect 10876 8925 10894 8959
rect 10894 8925 10928 8959
rect 10876 8916 10928 8925
rect 11152 8959 11204 8968
rect 11152 8925 11161 8959
rect 11161 8925 11195 8959
rect 11195 8925 11204 8959
rect 11152 8916 11204 8925
rect 7012 8848 7064 8900
rect 2780 8780 2832 8832
rect 5264 8780 5316 8832
rect 6644 8823 6696 8832
rect 6644 8789 6653 8823
rect 6653 8789 6687 8823
rect 6687 8789 6696 8823
rect 6644 8780 6696 8789
rect 7380 8823 7432 8832
rect 7380 8789 7389 8823
rect 7389 8789 7423 8823
rect 7423 8789 7432 8823
rect 7380 8780 7432 8789
rect 8300 8848 8352 8900
rect 9496 8823 9548 8832
rect 9496 8789 9505 8823
rect 9505 8789 9539 8823
rect 9539 8789 9548 8823
rect 9496 8780 9548 8789
rect 9772 8823 9824 8832
rect 9772 8789 9781 8823
rect 9781 8789 9815 8823
rect 9815 8789 9824 8823
rect 9772 8780 9824 8789
rect 10876 8780 10928 8832
rect 11980 8848 12032 8900
rect 12992 8780 13044 8832
rect 13452 8916 13504 8968
rect 15752 8916 15804 8968
rect 18328 8916 18380 8968
rect 19984 8916 20036 8968
rect 21364 8984 21416 9036
rect 16948 8848 17000 8900
rect 18052 8848 18104 8900
rect 20720 8848 20772 8900
rect 13268 8780 13320 8832
rect 14372 8780 14424 8832
rect 14556 8780 14608 8832
rect 18972 8780 19024 8832
rect 6148 8678 6200 8730
rect 6212 8678 6264 8730
rect 6276 8678 6328 8730
rect 6340 8678 6392 8730
rect 6404 8678 6456 8730
rect 11346 8678 11398 8730
rect 11410 8678 11462 8730
rect 11474 8678 11526 8730
rect 11538 8678 11590 8730
rect 11602 8678 11654 8730
rect 16544 8678 16596 8730
rect 16608 8678 16660 8730
rect 16672 8678 16724 8730
rect 16736 8678 16788 8730
rect 16800 8678 16852 8730
rect 21742 8678 21794 8730
rect 21806 8678 21858 8730
rect 21870 8678 21922 8730
rect 21934 8678 21986 8730
rect 21998 8678 22050 8730
rect 2780 8619 2832 8628
rect 2780 8585 2789 8619
rect 2789 8585 2823 8619
rect 2823 8585 2832 8619
rect 2780 8576 2832 8585
rect 3332 8576 3384 8628
rect 5264 8619 5316 8628
rect 2320 8508 2372 8560
rect 5264 8585 5273 8619
rect 5273 8585 5307 8619
rect 5307 8585 5316 8619
rect 5264 8576 5316 8585
rect 6644 8576 6696 8628
rect 9496 8576 9548 8628
rect 11152 8619 11204 8628
rect 11152 8585 11161 8619
rect 11161 8585 11195 8619
rect 11195 8585 11204 8619
rect 11152 8576 11204 8585
rect 13360 8619 13412 8628
rect 3424 8440 3476 8492
rect 3976 8440 4028 8492
rect 4252 8483 4304 8492
rect 4252 8449 4261 8483
rect 4261 8449 4295 8483
rect 4295 8449 4304 8483
rect 4252 8440 4304 8449
rect 4344 8415 4396 8424
rect 4344 8381 4353 8415
rect 4353 8381 4387 8415
rect 4387 8381 4396 8415
rect 4344 8372 4396 8381
rect 5632 8372 5684 8424
rect 7564 8415 7616 8424
rect 7564 8381 7573 8415
rect 7573 8381 7607 8415
rect 7607 8381 7616 8415
rect 7564 8372 7616 8381
rect 7656 8415 7708 8424
rect 7656 8381 7665 8415
rect 7665 8381 7699 8415
rect 7699 8381 7708 8415
rect 8576 8415 8628 8424
rect 7656 8372 7708 8381
rect 8576 8381 8585 8415
rect 8585 8381 8619 8415
rect 8619 8381 8628 8415
rect 8576 8372 8628 8381
rect 9864 8415 9916 8424
rect 9864 8381 9873 8415
rect 9873 8381 9907 8415
rect 9907 8381 9916 8415
rect 9864 8372 9916 8381
rect 12900 8508 12952 8560
rect 12256 8440 12308 8492
rect 13360 8585 13369 8619
rect 13369 8585 13403 8619
rect 13403 8585 13412 8619
rect 13360 8576 13412 8585
rect 15752 8619 15804 8628
rect 15752 8585 15761 8619
rect 15761 8585 15795 8619
rect 15795 8585 15804 8619
rect 15752 8576 15804 8585
rect 17960 8576 18012 8628
rect 13084 8508 13136 8560
rect 14188 8440 14240 8492
rect 14464 8483 14516 8492
rect 14464 8449 14482 8483
rect 14482 8449 14516 8483
rect 14464 8440 14516 8449
rect 13268 8372 13320 8424
rect 21456 8576 21508 8628
rect 18328 8483 18380 8492
rect 18328 8449 18337 8483
rect 18337 8449 18371 8483
rect 18371 8449 18380 8483
rect 18328 8440 18380 8449
rect 18420 8440 18472 8492
rect 19984 8483 20036 8492
rect 19984 8449 19993 8483
rect 19993 8449 20027 8483
rect 20027 8449 20036 8483
rect 19984 8440 20036 8449
rect 4160 8304 4212 8356
rect 5080 8304 5132 8356
rect 7196 8304 7248 8356
rect 7748 8304 7800 8356
rect 11980 8304 12032 8356
rect 4896 8279 4948 8288
rect 4896 8245 4905 8279
rect 4905 8245 4939 8279
rect 4939 8245 4948 8279
rect 4896 8236 4948 8245
rect 9404 8279 9456 8288
rect 9404 8245 9413 8279
rect 9413 8245 9447 8279
rect 9447 8245 9456 8279
rect 9404 8236 9456 8245
rect 18512 8236 18564 8288
rect 20720 8236 20772 8288
rect 3549 8134 3601 8186
rect 3613 8134 3665 8186
rect 3677 8134 3729 8186
rect 3741 8134 3793 8186
rect 3805 8134 3857 8186
rect 8747 8134 8799 8186
rect 8811 8134 8863 8186
rect 8875 8134 8927 8186
rect 8939 8134 8991 8186
rect 9003 8134 9055 8186
rect 13945 8134 13997 8186
rect 14009 8134 14061 8186
rect 14073 8134 14125 8186
rect 14137 8134 14189 8186
rect 14201 8134 14253 8186
rect 19143 8134 19195 8186
rect 19207 8134 19259 8186
rect 19271 8134 19323 8186
rect 19335 8134 19387 8186
rect 19399 8134 19451 8186
rect 4252 8032 4304 8084
rect 5264 8032 5316 8084
rect 3240 7896 3292 7948
rect 4620 7939 4672 7948
rect 4620 7905 4629 7939
rect 4629 7905 4663 7939
rect 4663 7905 4672 7939
rect 4620 7896 4672 7905
rect 6552 7964 6604 8016
rect 5540 7896 5592 7948
rect 7564 8032 7616 8084
rect 8392 8032 8444 8084
rect 7840 7939 7892 7948
rect 7840 7905 7849 7939
rect 7849 7905 7883 7939
rect 7883 7905 7892 7939
rect 7840 7896 7892 7905
rect 3884 7828 3936 7880
rect 3424 7803 3476 7812
rect 3424 7769 3433 7803
rect 3433 7769 3467 7803
rect 3467 7769 3476 7803
rect 3424 7760 3476 7769
rect 3240 7692 3292 7744
rect 3884 7735 3936 7744
rect 3884 7701 3893 7735
rect 3893 7701 3927 7735
rect 3927 7701 3936 7735
rect 3884 7692 3936 7701
rect 5264 7692 5316 7744
rect 5448 7735 5500 7744
rect 5448 7701 5457 7735
rect 5457 7701 5491 7735
rect 5491 7701 5500 7735
rect 5448 7692 5500 7701
rect 8576 7828 8628 7880
rect 9864 8032 9916 8084
rect 11336 8075 11388 8084
rect 11336 8041 11345 8075
rect 11345 8041 11379 8075
rect 11379 8041 11388 8075
rect 11336 8032 11388 8041
rect 15476 8032 15528 8084
rect 15660 8075 15712 8084
rect 15660 8041 15669 8075
rect 15669 8041 15703 8075
rect 15703 8041 15712 8075
rect 15660 8032 15712 8041
rect 16948 8032 17000 8084
rect 18328 8032 18380 8084
rect 18420 7964 18472 8016
rect 15752 7896 15804 7948
rect 19984 8032 20036 8084
rect 21088 8032 21140 8084
rect 8208 7760 8260 7812
rect 11336 7760 11388 7812
rect 8024 7692 8076 7744
rect 13268 7871 13320 7880
rect 13268 7837 13277 7871
rect 13277 7837 13311 7871
rect 13311 7837 13320 7871
rect 13268 7828 13320 7837
rect 13728 7828 13780 7880
rect 12532 7760 12584 7812
rect 13820 7760 13872 7812
rect 16212 7803 16264 7812
rect 16212 7769 16246 7803
rect 16246 7769 16264 7803
rect 16212 7760 16264 7769
rect 19616 7760 19668 7812
rect 17408 7692 17460 7744
rect 19432 7692 19484 7744
rect 20628 7735 20680 7744
rect 20628 7701 20637 7735
rect 20637 7701 20671 7735
rect 20671 7701 20680 7735
rect 20628 7692 20680 7701
rect 6148 7590 6200 7642
rect 6212 7590 6264 7642
rect 6276 7590 6328 7642
rect 6340 7590 6392 7642
rect 6404 7590 6456 7642
rect 11346 7590 11398 7642
rect 11410 7590 11462 7642
rect 11474 7590 11526 7642
rect 11538 7590 11590 7642
rect 11602 7590 11654 7642
rect 16544 7590 16596 7642
rect 16608 7590 16660 7642
rect 16672 7590 16724 7642
rect 16736 7590 16788 7642
rect 16800 7590 16852 7642
rect 21742 7590 21794 7642
rect 21806 7590 21858 7642
rect 21870 7590 21922 7642
rect 21934 7590 21986 7642
rect 21998 7590 22050 7642
rect 2964 7488 3016 7540
rect 4344 7488 4396 7540
rect 4896 7488 4948 7540
rect 7104 7531 7156 7540
rect 7104 7497 7113 7531
rect 7113 7497 7147 7531
rect 7147 7497 7156 7531
rect 7104 7488 7156 7497
rect 7380 7488 7432 7540
rect 11152 7488 11204 7540
rect 12624 7488 12676 7540
rect 14464 7488 14516 7540
rect 15752 7531 15804 7540
rect 15752 7497 15761 7531
rect 15761 7497 15795 7531
rect 15795 7497 15804 7531
rect 15752 7488 15804 7497
rect 17408 7531 17460 7540
rect 17408 7497 17417 7531
rect 17417 7497 17451 7531
rect 17451 7497 17460 7531
rect 17408 7488 17460 7497
rect 18052 7488 18104 7540
rect 20720 7531 20772 7540
rect 20720 7497 20729 7531
rect 20729 7497 20763 7531
rect 20763 7497 20772 7531
rect 20720 7488 20772 7497
rect 21088 7531 21140 7540
rect 21088 7497 21097 7531
rect 21097 7497 21131 7531
rect 21131 7497 21140 7531
rect 21088 7488 21140 7497
rect 2688 7420 2740 7472
rect 4528 7420 4580 7472
rect 5448 7420 5500 7472
rect 10968 7420 11020 7472
rect 13360 7420 13412 7472
rect 2964 7352 3016 7404
rect 4620 7352 4672 7404
rect 4804 7327 4856 7336
rect 2044 7259 2096 7268
rect 2044 7225 2053 7259
rect 2053 7225 2087 7259
rect 2087 7225 2096 7259
rect 2044 7216 2096 7225
rect 4804 7293 4813 7327
rect 4813 7293 4847 7327
rect 4847 7293 4856 7327
rect 4804 7284 4856 7293
rect 4988 7327 5040 7336
rect 4988 7293 4997 7327
rect 4997 7293 5031 7327
rect 5031 7293 5040 7327
rect 4988 7284 5040 7293
rect 8576 7395 8628 7404
rect 8576 7361 8585 7395
rect 8585 7361 8619 7395
rect 8619 7361 8628 7395
rect 8576 7352 8628 7361
rect 12348 7352 12400 7404
rect 13728 7352 13780 7404
rect 18328 7420 18380 7472
rect 6920 7284 6972 7336
rect 6552 7216 6604 7268
rect 2964 7191 3016 7200
rect 2964 7157 2973 7191
rect 2973 7157 3007 7191
rect 3007 7157 3016 7191
rect 2964 7148 3016 7157
rect 5448 7191 5500 7200
rect 5448 7157 5457 7191
rect 5457 7157 5491 7191
rect 5491 7157 5500 7191
rect 5448 7148 5500 7157
rect 8208 7284 8260 7336
rect 18512 7395 18564 7404
rect 18512 7361 18530 7395
rect 18530 7361 18564 7395
rect 18512 7352 18564 7361
rect 9588 7216 9640 7268
rect 9864 7148 9916 7200
rect 13176 7148 13228 7200
rect 19524 7148 19576 7200
rect 3549 7046 3601 7098
rect 3613 7046 3665 7098
rect 3677 7046 3729 7098
rect 3741 7046 3793 7098
rect 3805 7046 3857 7098
rect 8747 7046 8799 7098
rect 8811 7046 8863 7098
rect 8875 7046 8927 7098
rect 8939 7046 8991 7098
rect 9003 7046 9055 7098
rect 13945 7046 13997 7098
rect 14009 7046 14061 7098
rect 14073 7046 14125 7098
rect 14137 7046 14189 7098
rect 14201 7046 14253 7098
rect 19143 7046 19195 7098
rect 19207 7046 19259 7098
rect 19271 7046 19323 7098
rect 19335 7046 19387 7098
rect 19399 7046 19451 7098
rect 2320 6808 2372 6860
rect 4252 6944 4304 6996
rect 4988 6944 5040 6996
rect 3976 6876 4028 6928
rect 8392 6944 8444 6996
rect 8576 6944 8628 6996
rect 5632 6876 5684 6928
rect 13176 6944 13228 6996
rect 13360 6987 13412 6996
rect 13360 6953 13369 6987
rect 13369 6953 13403 6987
rect 13403 6953 13412 6987
rect 13360 6944 13412 6953
rect 13728 6987 13780 6996
rect 13728 6953 13737 6987
rect 13737 6953 13771 6987
rect 13771 6953 13780 6987
rect 13728 6944 13780 6953
rect 15752 6944 15804 6996
rect 4160 6808 4212 6860
rect 5172 6808 5224 6860
rect 4344 6740 4396 6792
rect 5264 6740 5316 6792
rect 6000 6808 6052 6860
rect 9128 6808 9180 6860
rect 9588 6851 9640 6860
rect 9588 6817 9597 6851
rect 9597 6817 9631 6851
rect 9631 6817 9640 6851
rect 9588 6808 9640 6817
rect 18328 6944 18380 6996
rect 19524 6944 19576 6996
rect 21088 6944 21140 6996
rect 7748 6783 7800 6792
rect 1676 6647 1728 6656
rect 1676 6613 1685 6647
rect 1685 6613 1719 6647
rect 1719 6613 1728 6647
rect 1676 6604 1728 6613
rect 2504 6604 2556 6656
rect 7472 6715 7524 6724
rect 4528 6647 4580 6656
rect 4528 6613 4537 6647
rect 4537 6613 4571 6647
rect 4571 6613 4580 6647
rect 4528 6604 4580 6613
rect 5172 6604 5224 6656
rect 5724 6604 5776 6656
rect 6736 6647 6788 6656
rect 6736 6613 6745 6647
rect 6745 6613 6779 6647
rect 6779 6613 6788 6647
rect 7472 6681 7481 6715
rect 7481 6681 7515 6715
rect 7515 6681 7524 6715
rect 7472 6672 7524 6681
rect 7748 6749 7757 6783
rect 7757 6749 7791 6783
rect 7791 6749 7800 6783
rect 7748 6740 7800 6749
rect 13728 6740 13780 6792
rect 15476 6740 15528 6792
rect 18236 6740 18288 6792
rect 19800 6740 19852 6792
rect 11152 6672 11204 6724
rect 12440 6672 12492 6724
rect 6736 6604 6788 6613
rect 9036 6604 9088 6656
rect 10324 6604 10376 6656
rect 12348 6604 12400 6656
rect 14280 6604 14332 6656
rect 17776 6672 17828 6724
rect 15384 6604 15436 6656
rect 16948 6604 17000 6656
rect 19708 6604 19760 6656
rect 6148 6502 6200 6554
rect 6212 6502 6264 6554
rect 6276 6502 6328 6554
rect 6340 6502 6392 6554
rect 6404 6502 6456 6554
rect 11346 6502 11398 6554
rect 11410 6502 11462 6554
rect 11474 6502 11526 6554
rect 11538 6502 11590 6554
rect 11602 6502 11654 6554
rect 16544 6502 16596 6554
rect 16608 6502 16660 6554
rect 16672 6502 16724 6554
rect 16736 6502 16788 6554
rect 16800 6502 16852 6554
rect 21742 6502 21794 6554
rect 21806 6502 21858 6554
rect 21870 6502 21922 6554
rect 21934 6502 21986 6554
rect 21998 6502 22050 6554
rect 2504 6443 2556 6452
rect 2504 6409 2513 6443
rect 2513 6409 2547 6443
rect 2547 6409 2556 6443
rect 2504 6400 2556 6409
rect 5724 6400 5776 6452
rect 6736 6443 6788 6452
rect 6736 6409 6745 6443
rect 6745 6409 6779 6443
rect 6779 6409 6788 6443
rect 6736 6400 6788 6409
rect 8392 6400 8444 6452
rect 9036 6443 9088 6452
rect 9036 6409 9045 6443
rect 9045 6409 9079 6443
rect 9079 6409 9088 6443
rect 9036 6400 9088 6409
rect 9128 6400 9180 6452
rect 5264 6332 5316 6384
rect 4528 6307 4580 6316
rect 4528 6273 4537 6307
rect 4537 6273 4571 6307
rect 4571 6273 4580 6307
rect 4528 6264 4580 6273
rect 5540 6264 5592 6316
rect 6276 6264 6328 6316
rect 1768 6196 1820 6248
rect 4620 6196 4672 6248
rect 5264 6196 5316 6248
rect 5908 6239 5960 6248
rect 5908 6205 5917 6239
rect 5917 6205 5951 6239
rect 5951 6205 5960 6239
rect 5908 6196 5960 6205
rect 6552 6332 6604 6384
rect 10324 6332 10376 6384
rect 15752 6400 15804 6452
rect 18328 6443 18380 6452
rect 18328 6409 18337 6443
rect 18337 6409 18371 6443
rect 18371 6409 18380 6443
rect 18328 6400 18380 6409
rect 6460 6264 6512 6316
rect 7288 6196 7340 6248
rect 10048 6264 10100 6316
rect 8668 6196 8720 6248
rect 9312 6239 9364 6248
rect 9312 6205 9321 6239
rect 9321 6205 9355 6239
rect 9355 6205 9364 6239
rect 9312 6196 9364 6205
rect 11796 6196 11848 6248
rect 13728 6264 13780 6316
rect 14280 6264 14332 6316
rect 15752 6264 15804 6316
rect 19156 6400 19208 6452
rect 21088 6443 21140 6452
rect 21088 6409 21097 6443
rect 21097 6409 21131 6443
rect 21131 6409 21140 6443
rect 21088 6400 21140 6409
rect 19524 6264 19576 6316
rect 19708 6307 19760 6316
rect 19708 6273 19742 6307
rect 19742 6273 19760 6307
rect 19708 6264 19760 6273
rect 5080 6060 5132 6112
rect 5632 6060 5684 6112
rect 7012 6060 7064 6112
rect 8668 6060 8720 6112
rect 11888 6103 11940 6112
rect 11888 6069 11897 6103
rect 11897 6069 11931 6103
rect 11931 6069 11940 6103
rect 11888 6060 11940 6069
rect 14740 6060 14792 6112
rect 3549 5958 3601 6010
rect 3613 5958 3665 6010
rect 3677 5958 3729 6010
rect 3741 5958 3793 6010
rect 3805 5958 3857 6010
rect 8747 5958 8799 6010
rect 8811 5958 8863 6010
rect 8875 5958 8927 6010
rect 8939 5958 8991 6010
rect 9003 5958 9055 6010
rect 13945 5958 13997 6010
rect 14009 5958 14061 6010
rect 14073 5958 14125 6010
rect 14137 5958 14189 6010
rect 14201 5958 14253 6010
rect 19143 5958 19195 6010
rect 19207 5958 19259 6010
rect 19271 5958 19323 6010
rect 19335 5958 19387 6010
rect 19399 5958 19451 6010
rect 3332 5856 3384 5908
rect 5264 5899 5316 5908
rect 2504 5788 2556 5840
rect 2964 5788 3016 5840
rect 5264 5865 5273 5899
rect 5273 5865 5307 5899
rect 5307 5865 5316 5899
rect 5264 5856 5316 5865
rect 5908 5856 5960 5908
rect 6920 5831 6972 5840
rect 1676 5695 1728 5704
rect 1676 5661 1685 5695
rect 1685 5661 1719 5695
rect 1719 5661 1728 5695
rect 1676 5652 1728 5661
rect 1768 5695 1820 5704
rect 1768 5661 1777 5695
rect 1777 5661 1811 5695
rect 1811 5661 1820 5695
rect 4528 5720 4580 5772
rect 6000 5720 6052 5772
rect 1768 5652 1820 5661
rect 5908 5652 5960 5704
rect 3240 5584 3292 5636
rect 4528 5584 4580 5636
rect 6920 5797 6929 5831
rect 6929 5797 6963 5831
rect 6963 5797 6972 5831
rect 6920 5788 6972 5797
rect 9588 5856 9640 5908
rect 8300 5720 8352 5772
rect 9588 5763 9640 5772
rect 9588 5729 9597 5763
rect 9597 5729 9631 5763
rect 9631 5729 9640 5763
rect 9588 5720 9640 5729
rect 7288 5652 7340 5704
rect 7564 5652 7616 5704
rect 7656 5695 7708 5704
rect 7656 5661 7665 5695
rect 7665 5661 7699 5695
rect 7699 5661 7708 5695
rect 9312 5695 9364 5704
rect 7656 5652 7708 5661
rect 9312 5661 9321 5695
rect 9321 5661 9355 5695
rect 9355 5661 9364 5695
rect 9312 5652 9364 5661
rect 11152 5788 11204 5840
rect 13452 5899 13504 5908
rect 13452 5865 13461 5899
rect 13461 5865 13495 5899
rect 13495 5865 13504 5899
rect 13452 5856 13504 5865
rect 13728 5856 13780 5908
rect 15752 5899 15804 5908
rect 15752 5865 15761 5899
rect 15761 5865 15795 5899
rect 15795 5865 15804 5899
rect 15752 5856 15804 5865
rect 18328 5856 18380 5908
rect 19800 5856 19852 5908
rect 21088 5899 21140 5908
rect 21088 5865 21097 5899
rect 21097 5865 21131 5899
rect 21131 5865 21140 5899
rect 21088 5856 21140 5865
rect 19708 5788 19760 5840
rect 13452 5720 13504 5772
rect 12256 5652 12308 5704
rect 2136 5559 2188 5568
rect 2136 5525 2145 5559
rect 2145 5525 2179 5559
rect 2179 5525 2188 5559
rect 2136 5516 2188 5525
rect 2412 5559 2464 5568
rect 2412 5525 2421 5559
rect 2421 5525 2455 5559
rect 2455 5525 2464 5559
rect 2412 5516 2464 5525
rect 2872 5559 2924 5568
rect 2872 5525 2881 5559
rect 2881 5525 2915 5559
rect 2915 5525 2924 5559
rect 4804 5559 4856 5568
rect 2872 5516 2924 5525
rect 4804 5525 4813 5559
rect 4813 5525 4847 5559
rect 4847 5525 4856 5559
rect 4804 5516 4856 5525
rect 5172 5516 5224 5568
rect 5540 5559 5592 5568
rect 5540 5525 5549 5559
rect 5549 5525 5583 5559
rect 5583 5525 5592 5559
rect 5540 5516 5592 5525
rect 14372 5584 14424 5636
rect 15752 5720 15804 5772
rect 14740 5652 14792 5704
rect 19064 5652 19116 5704
rect 16396 5584 16448 5636
rect 17776 5584 17828 5636
rect 19708 5584 19760 5636
rect 6644 5559 6696 5568
rect 6644 5525 6653 5559
rect 6653 5525 6687 5559
rect 6687 5525 6696 5559
rect 6644 5516 6696 5525
rect 6920 5516 6972 5568
rect 8576 5559 8628 5568
rect 8576 5525 8585 5559
rect 8585 5525 8619 5559
rect 8619 5525 8628 5559
rect 8576 5516 8628 5525
rect 8944 5559 8996 5568
rect 8944 5525 8953 5559
rect 8953 5525 8987 5559
rect 8987 5525 8996 5559
rect 8944 5516 8996 5525
rect 9956 5559 10008 5568
rect 9956 5525 9965 5559
rect 9965 5525 9999 5559
rect 9999 5525 10008 5559
rect 9956 5516 10008 5525
rect 11152 5559 11204 5568
rect 11152 5525 11161 5559
rect 11161 5525 11195 5559
rect 11195 5525 11204 5559
rect 11152 5516 11204 5525
rect 14096 5559 14148 5568
rect 14096 5525 14105 5559
rect 14105 5525 14139 5559
rect 14139 5525 14148 5559
rect 14096 5516 14148 5525
rect 6148 5414 6200 5466
rect 6212 5414 6264 5466
rect 6276 5414 6328 5466
rect 6340 5414 6392 5466
rect 6404 5414 6456 5466
rect 11346 5414 11398 5466
rect 11410 5414 11462 5466
rect 11474 5414 11526 5466
rect 11538 5414 11590 5466
rect 11602 5414 11654 5466
rect 16544 5414 16596 5466
rect 16608 5414 16660 5466
rect 16672 5414 16724 5466
rect 16736 5414 16788 5466
rect 16800 5414 16852 5466
rect 21742 5414 21794 5466
rect 21806 5414 21858 5466
rect 21870 5414 21922 5466
rect 21934 5414 21986 5466
rect 21998 5414 22050 5466
rect 1676 5312 1728 5364
rect 2504 5312 2556 5364
rect 2872 5312 2924 5364
rect 3240 5355 3292 5364
rect 3240 5321 3249 5355
rect 3249 5321 3283 5355
rect 3283 5321 3292 5355
rect 3240 5312 3292 5321
rect 3424 5312 3476 5364
rect 4804 5312 4856 5364
rect 4896 5312 4948 5364
rect 7012 5312 7064 5364
rect 7656 5312 7708 5364
rect 8576 5312 8628 5364
rect 1768 4972 1820 5024
rect 2688 5108 2740 5160
rect 3792 5176 3844 5228
rect 4068 5244 4120 5296
rect 5540 5244 5592 5296
rect 6644 5244 6696 5296
rect 4896 5176 4948 5228
rect 5264 5176 5316 5228
rect 7012 5176 7064 5228
rect 8944 5176 8996 5228
rect 3884 5151 3936 5160
rect 3884 5117 3893 5151
rect 3893 5117 3927 5151
rect 3927 5117 3936 5151
rect 3884 5108 3936 5117
rect 5632 5108 5684 5160
rect 5908 5108 5960 5160
rect 4252 5040 4304 5092
rect 6736 5040 6788 5092
rect 7380 5108 7432 5160
rect 9588 5244 9640 5296
rect 12440 5244 12492 5296
rect 12624 5287 12676 5296
rect 12624 5253 12642 5287
rect 12642 5253 12676 5287
rect 12624 5244 12676 5253
rect 10876 5219 10928 5228
rect 10876 5185 10894 5219
rect 10894 5185 10928 5219
rect 11152 5219 11204 5228
rect 10876 5176 10928 5185
rect 11152 5185 11161 5219
rect 11161 5185 11195 5219
rect 11195 5185 11204 5219
rect 11152 5176 11204 5185
rect 12992 5176 13044 5228
rect 13452 5312 13504 5364
rect 15752 5312 15804 5364
rect 14096 5244 14148 5296
rect 18328 5355 18380 5364
rect 18328 5321 18337 5355
rect 18337 5321 18371 5355
rect 18371 5321 18380 5355
rect 18328 5312 18380 5321
rect 19708 5355 19760 5364
rect 19708 5321 19717 5355
rect 19717 5321 19751 5355
rect 19751 5321 19760 5355
rect 19708 5312 19760 5321
rect 17040 5244 17092 5296
rect 18604 5244 18656 5296
rect 20720 5244 20772 5296
rect 16488 5176 16540 5228
rect 16948 5219 17000 5228
rect 16948 5185 16982 5219
rect 16982 5185 17000 5219
rect 21088 5219 21140 5228
rect 16948 5176 17000 5185
rect 21088 5185 21097 5219
rect 21097 5185 21131 5219
rect 21131 5185 21140 5219
rect 21088 5176 21140 5185
rect 10048 5040 10100 5092
rect 11796 5040 11848 5092
rect 3148 4972 3200 5024
rect 3976 4972 4028 5024
rect 6368 5015 6420 5024
rect 6368 4981 6377 5015
rect 6377 4981 6411 5015
rect 6411 4981 6420 5015
rect 6368 4972 6420 4981
rect 8576 4972 8628 5024
rect 9128 4972 9180 5024
rect 9404 4972 9456 5024
rect 11612 4972 11664 5024
rect 15200 4972 15252 5024
rect 18144 4972 18196 5024
rect 3549 4870 3601 4922
rect 3613 4870 3665 4922
rect 3677 4870 3729 4922
rect 3741 4870 3793 4922
rect 3805 4870 3857 4922
rect 8747 4870 8799 4922
rect 8811 4870 8863 4922
rect 8875 4870 8927 4922
rect 8939 4870 8991 4922
rect 9003 4870 9055 4922
rect 13945 4870 13997 4922
rect 14009 4870 14061 4922
rect 14073 4870 14125 4922
rect 14137 4870 14189 4922
rect 14201 4870 14253 4922
rect 19143 4870 19195 4922
rect 19207 4870 19259 4922
rect 19271 4870 19323 4922
rect 19335 4870 19387 4922
rect 19399 4870 19451 4922
rect 4528 4768 4580 4820
rect 4896 4768 4948 4820
rect 5264 4768 5316 4820
rect 5632 4768 5684 4820
rect 10876 4811 10928 4820
rect 3884 4700 3936 4752
rect 1860 4675 1912 4684
rect 1860 4641 1869 4675
rect 1869 4641 1903 4675
rect 1903 4641 1912 4675
rect 1860 4632 1912 4641
rect 2412 4632 2464 4684
rect 2136 4564 2188 4616
rect 6368 4632 6420 4684
rect 7104 4632 7156 4684
rect 7288 4675 7340 4684
rect 7288 4641 7297 4675
rect 7297 4641 7331 4675
rect 7331 4641 7340 4675
rect 7288 4632 7340 4641
rect 8392 4632 8444 4684
rect 7012 4564 7064 4616
rect 9128 4564 9180 4616
rect 2504 4496 2556 4548
rect 2688 4428 2740 4480
rect 4252 4428 4304 4480
rect 5816 4471 5868 4480
rect 5816 4437 5825 4471
rect 5825 4437 5859 4471
rect 5859 4437 5868 4471
rect 7288 4496 7340 4548
rect 9312 4496 9364 4548
rect 5816 4428 5868 4437
rect 6828 4428 6880 4480
rect 7012 4471 7064 4480
rect 7012 4437 7021 4471
rect 7021 4437 7055 4471
rect 7055 4437 7064 4471
rect 7012 4428 7064 4437
rect 9128 4471 9180 4480
rect 9128 4437 9137 4471
rect 9137 4437 9171 4471
rect 9171 4437 9180 4471
rect 9128 4428 9180 4437
rect 10876 4777 10885 4811
rect 10885 4777 10919 4811
rect 10919 4777 10928 4811
rect 10876 4768 10928 4777
rect 11612 4768 11664 4820
rect 12532 4768 12584 4820
rect 12992 4811 13044 4820
rect 12992 4777 13001 4811
rect 13001 4777 13035 4811
rect 13035 4777 13044 4811
rect 12992 4768 13044 4777
rect 13636 4768 13688 4820
rect 16488 4811 16540 4820
rect 12440 4700 12492 4752
rect 15108 4700 15160 4752
rect 16488 4777 16497 4811
rect 16497 4777 16531 4811
rect 16531 4777 16540 4811
rect 16488 4768 16540 4777
rect 16212 4700 16264 4752
rect 11152 4632 11204 4684
rect 16120 4675 16172 4684
rect 16120 4641 16129 4675
rect 16129 4641 16163 4675
rect 16163 4641 16172 4675
rect 16120 4632 16172 4641
rect 19616 4632 19668 4684
rect 21088 4768 21140 4820
rect 19984 4564 20036 4616
rect 11060 4496 11112 4548
rect 10232 4428 10284 4480
rect 10876 4428 10928 4480
rect 12440 4428 12492 4480
rect 15108 4428 15160 4480
rect 17040 4428 17092 4480
rect 19524 4496 19576 4548
rect 18052 4428 18104 4480
rect 6148 4326 6200 4378
rect 6212 4326 6264 4378
rect 6276 4326 6328 4378
rect 6340 4326 6392 4378
rect 6404 4326 6456 4378
rect 11346 4326 11398 4378
rect 11410 4326 11462 4378
rect 11474 4326 11526 4378
rect 11538 4326 11590 4378
rect 11602 4326 11654 4378
rect 16544 4326 16596 4378
rect 16608 4326 16660 4378
rect 16672 4326 16724 4378
rect 16736 4326 16788 4378
rect 16800 4326 16852 4378
rect 21742 4326 21794 4378
rect 21806 4326 21858 4378
rect 21870 4326 21922 4378
rect 21934 4326 21986 4378
rect 21998 4326 22050 4378
rect 2688 4131 2740 4140
rect 2688 4097 2697 4131
rect 2697 4097 2731 4131
rect 2731 4097 2740 4131
rect 2688 4088 2740 4097
rect 4160 4088 4212 4140
rect 4804 4131 4856 4140
rect 4804 4097 4813 4131
rect 4813 4097 4847 4131
rect 4847 4097 4856 4131
rect 4804 4088 4856 4097
rect 4896 4020 4948 4072
rect 6184 4224 6236 4276
rect 8024 4224 8076 4276
rect 9128 4224 9180 4276
rect 11152 4267 11204 4276
rect 11152 4233 11161 4267
rect 11161 4233 11195 4267
rect 11195 4233 11204 4267
rect 11152 4224 11204 4233
rect 6920 4156 6972 4208
rect 5632 4131 5684 4140
rect 5632 4097 5641 4131
rect 5641 4097 5675 4131
rect 5675 4097 5684 4131
rect 6828 4131 6880 4140
rect 5632 4088 5684 4097
rect 6828 4097 6837 4131
rect 6837 4097 6871 4131
rect 6871 4097 6880 4131
rect 6828 4088 6880 4097
rect 9956 4156 10008 4208
rect 3424 3952 3476 4004
rect 5908 4020 5960 4072
rect 6644 4063 6696 4072
rect 6644 4029 6653 4063
rect 6653 4029 6687 4063
rect 6687 4029 6696 4063
rect 6644 4020 6696 4029
rect 5172 3995 5224 4004
rect 3884 3884 3936 3936
rect 5172 3961 5181 3995
rect 5181 3961 5215 3995
rect 5215 3961 5224 3995
rect 5172 3952 5224 3961
rect 5448 3952 5500 4004
rect 5632 3884 5684 3936
rect 8024 4020 8076 4072
rect 10048 4088 10100 4140
rect 11704 4088 11756 4140
rect 13636 4156 13688 4208
rect 13176 4088 13228 4140
rect 9588 4063 9640 4072
rect 9588 4029 9597 4063
rect 9597 4029 9631 4063
rect 9631 4029 9640 4063
rect 9588 4020 9640 4029
rect 9128 3952 9180 4004
rect 12808 4020 12860 4072
rect 10048 3884 10100 3936
rect 12624 3927 12676 3936
rect 12624 3893 12633 3927
rect 12633 3893 12667 3927
rect 12667 3893 12676 3927
rect 12624 3884 12676 3893
rect 13728 3884 13780 3936
rect 15384 4131 15436 4140
rect 15384 4097 15402 4131
rect 15402 4097 15436 4131
rect 15384 4088 15436 4097
rect 16120 4224 16172 4276
rect 18788 4224 18840 4276
rect 19984 4267 20036 4276
rect 19984 4233 19993 4267
rect 19993 4233 20027 4267
rect 20027 4233 20036 4267
rect 19984 4224 20036 4233
rect 16764 4088 16816 4140
rect 19064 4088 19116 4140
rect 19616 4088 19668 4140
rect 14280 3995 14332 4004
rect 14280 3961 14289 3995
rect 14289 3961 14323 3995
rect 14323 3961 14332 3995
rect 14280 3952 14332 3961
rect 17960 3952 18012 4004
rect 16948 3884 17000 3936
rect 18236 3952 18288 4004
rect 20812 4088 20864 4140
rect 3549 3782 3601 3834
rect 3613 3782 3665 3834
rect 3677 3782 3729 3834
rect 3741 3782 3793 3834
rect 3805 3782 3857 3834
rect 8747 3782 8799 3834
rect 8811 3782 8863 3834
rect 8875 3782 8927 3834
rect 8939 3782 8991 3834
rect 9003 3782 9055 3834
rect 13945 3782 13997 3834
rect 14009 3782 14061 3834
rect 14073 3782 14125 3834
rect 14137 3782 14189 3834
rect 14201 3782 14253 3834
rect 19143 3782 19195 3834
rect 19207 3782 19259 3834
rect 19271 3782 19323 3834
rect 19335 3782 19387 3834
rect 19399 3782 19451 3834
rect 2412 3680 2464 3732
rect 4344 3723 4396 3732
rect 4344 3689 4353 3723
rect 4353 3689 4387 3723
rect 4387 3689 4396 3723
rect 4344 3680 4396 3689
rect 5816 3723 5868 3732
rect 5816 3689 5825 3723
rect 5825 3689 5859 3723
rect 5859 3689 5868 3723
rect 5816 3680 5868 3689
rect 5908 3680 5960 3732
rect 9128 3680 9180 3732
rect 9588 3680 9640 3732
rect 12716 3680 12768 3732
rect 12992 3723 13044 3732
rect 12992 3689 13001 3723
rect 13001 3689 13035 3723
rect 13035 3689 13044 3723
rect 12992 3680 13044 3689
rect 4528 3612 4580 3664
rect 5448 3612 5500 3664
rect 7472 3612 7524 3664
rect 7656 3612 7708 3664
rect 3148 3544 3200 3596
rect 5632 3544 5684 3596
rect 6736 3544 6788 3596
rect 7748 3587 7800 3596
rect 7748 3553 7757 3587
rect 7757 3553 7791 3587
rect 7791 3553 7800 3587
rect 7748 3544 7800 3553
rect 9956 3612 10008 3664
rect 9680 3544 9732 3596
rect 11152 3544 11204 3596
rect 11612 3544 11664 3596
rect 16120 3680 16172 3732
rect 17040 3680 17092 3732
rect 5080 3519 5132 3528
rect 5080 3485 5089 3519
rect 5089 3485 5123 3519
rect 5123 3485 5132 3519
rect 5080 3476 5132 3485
rect 8576 3519 8628 3528
rect 6184 3451 6236 3460
rect 6184 3417 6193 3451
rect 6193 3417 6227 3451
rect 6227 3417 6236 3451
rect 6184 3408 6236 3417
rect 7472 3451 7524 3460
rect 7472 3417 7481 3451
rect 7481 3417 7515 3451
rect 7515 3417 7524 3451
rect 7472 3408 7524 3417
rect 7564 3451 7616 3460
rect 7564 3417 7573 3451
rect 7573 3417 7607 3451
rect 7607 3417 7616 3451
rect 8300 3451 8352 3460
rect 7564 3408 7616 3417
rect 8300 3417 8309 3451
rect 8309 3417 8343 3451
rect 8343 3417 8352 3451
rect 8300 3408 8352 3417
rect 8576 3485 8585 3519
rect 8585 3485 8619 3519
rect 8619 3485 8628 3519
rect 8576 3476 8628 3485
rect 10416 3476 10468 3528
rect 18328 3587 18380 3596
rect 18328 3553 18337 3587
rect 18337 3553 18371 3587
rect 18371 3553 18380 3587
rect 19616 3680 19668 3732
rect 18328 3544 18380 3553
rect 20628 3587 20680 3596
rect 20628 3553 20637 3587
rect 20637 3553 20671 3587
rect 20671 3553 20680 3587
rect 20628 3544 20680 3553
rect 12808 3476 12860 3528
rect 14280 3476 14332 3528
rect 15200 3519 15252 3528
rect 15200 3485 15218 3519
rect 15218 3485 15252 3519
rect 15200 3476 15252 3485
rect 18052 3519 18104 3528
rect 18052 3485 18070 3519
rect 18070 3485 18104 3519
rect 18052 3476 18104 3485
rect 19800 3476 19852 3528
rect 9680 3408 9732 3460
rect 12348 3451 12400 3460
rect 4804 3383 4856 3392
rect 4804 3349 4813 3383
rect 4813 3349 4847 3383
rect 4847 3349 4856 3383
rect 4804 3340 4856 3349
rect 6920 3340 6972 3392
rect 8668 3340 8720 3392
rect 9588 3383 9640 3392
rect 9588 3349 9597 3383
rect 9597 3349 9631 3383
rect 9631 3349 9640 3383
rect 9588 3340 9640 3349
rect 12348 3417 12366 3451
rect 12366 3417 12400 3451
rect 12348 3408 12400 3417
rect 12716 3408 12768 3460
rect 13452 3340 13504 3392
rect 19524 3408 19576 3460
rect 14648 3340 14700 3392
rect 16396 3340 16448 3392
rect 16488 3340 16540 3392
rect 6148 3238 6200 3290
rect 6212 3238 6264 3290
rect 6276 3238 6328 3290
rect 6340 3238 6392 3290
rect 6404 3238 6456 3290
rect 11346 3238 11398 3290
rect 11410 3238 11462 3290
rect 11474 3238 11526 3290
rect 11538 3238 11590 3290
rect 11602 3238 11654 3290
rect 16544 3238 16596 3290
rect 16608 3238 16660 3290
rect 16672 3238 16724 3290
rect 16736 3238 16788 3290
rect 16800 3238 16852 3290
rect 21742 3238 21794 3290
rect 21806 3238 21858 3290
rect 21870 3238 21922 3290
rect 21934 3238 21986 3290
rect 21998 3238 22050 3290
rect 1492 3179 1544 3188
rect 1492 3145 1501 3179
rect 1501 3145 1535 3179
rect 1535 3145 1544 3179
rect 1492 3136 1544 3145
rect 5908 3136 5960 3188
rect 6920 3179 6972 3188
rect 6920 3145 6929 3179
rect 6929 3145 6963 3179
rect 6963 3145 6972 3179
rect 6920 3136 6972 3145
rect 7012 3136 7064 3188
rect 7932 3136 7984 3188
rect 9036 3136 9088 3188
rect 9864 3136 9916 3188
rect 11428 3136 11480 3188
rect 12808 3136 12860 3188
rect 13176 3136 13228 3188
rect 14648 3136 14700 3188
rect 4804 3068 4856 3120
rect 4436 3000 4488 3052
rect 4620 3043 4672 3052
rect 4620 3009 4629 3043
rect 4629 3009 4663 3043
rect 4663 3009 4672 3043
rect 4620 3000 4672 3009
rect 5448 3043 5500 3052
rect 5448 3009 5457 3043
rect 5457 3009 5491 3043
rect 5491 3009 5500 3043
rect 5448 3000 5500 3009
rect 13084 3068 13136 3120
rect 8024 3043 8076 3052
rect 5816 2907 5868 2916
rect 2044 2839 2096 2848
rect 2044 2805 2053 2839
rect 2053 2805 2087 2839
rect 2087 2805 2096 2839
rect 2044 2796 2096 2805
rect 2596 2839 2648 2848
rect 2596 2805 2605 2839
rect 2605 2805 2639 2839
rect 2639 2805 2648 2839
rect 2596 2796 2648 2805
rect 5816 2873 5825 2907
rect 5825 2873 5859 2907
rect 5859 2873 5868 2907
rect 5816 2864 5868 2873
rect 8024 3009 8033 3043
rect 8033 3009 8067 3043
rect 8067 3009 8076 3043
rect 8024 3000 8076 3009
rect 8760 3043 8812 3052
rect 8760 3009 8769 3043
rect 8769 3009 8803 3043
rect 8803 3009 8812 3043
rect 8760 3000 8812 3009
rect 9036 3043 9088 3052
rect 9036 3009 9045 3043
rect 9045 3009 9079 3043
rect 9079 3009 9088 3043
rect 9036 3000 9088 3009
rect 9772 3000 9824 3052
rect 11152 3043 11204 3052
rect 11152 3009 11161 3043
rect 11161 3009 11195 3043
rect 11195 3009 11204 3043
rect 11152 3000 11204 3009
rect 6920 2932 6972 2984
rect 7104 2932 7156 2984
rect 9588 2932 9640 2984
rect 11428 2932 11480 2984
rect 13176 3043 13228 3052
rect 13176 3009 13185 3043
rect 13185 3009 13219 3043
rect 13219 3009 13228 3043
rect 13176 3000 13228 3009
rect 13728 3043 13780 3052
rect 13728 3009 13737 3043
rect 13737 3009 13771 3043
rect 13771 3009 13780 3043
rect 13728 3000 13780 3009
rect 14648 3000 14700 3052
rect 17132 3179 17184 3188
rect 17132 3145 17141 3179
rect 17141 3145 17175 3179
rect 17175 3145 17184 3179
rect 17132 3136 17184 3145
rect 15752 3068 15804 3120
rect 15568 3043 15620 3052
rect 7380 2864 7432 2916
rect 9680 2796 9732 2848
rect 15568 3009 15577 3043
rect 15577 3009 15611 3043
rect 15611 3009 15620 3043
rect 15568 3000 15620 3009
rect 13820 2864 13872 2916
rect 17040 2864 17092 2916
rect 16948 2796 17000 2848
rect 17960 3068 18012 3120
rect 18328 3136 18380 3188
rect 19064 3068 19116 3120
rect 17776 3000 17828 3052
rect 18328 3000 18380 3052
rect 18788 3043 18840 3052
rect 18788 3009 18822 3043
rect 18822 3009 18840 3043
rect 18788 3000 18840 3009
rect 20352 3043 20404 3052
rect 20352 3009 20361 3043
rect 20361 3009 20395 3043
rect 20395 3009 20404 3043
rect 20352 3000 20404 3009
rect 20812 3000 20864 3052
rect 20628 2975 20680 2984
rect 20628 2941 20637 2975
rect 20637 2941 20671 2975
rect 20671 2941 20680 2975
rect 20628 2932 20680 2941
rect 19800 2796 19852 2848
rect 3549 2694 3601 2746
rect 3613 2694 3665 2746
rect 3677 2694 3729 2746
rect 3741 2694 3793 2746
rect 3805 2694 3857 2746
rect 8747 2694 8799 2746
rect 8811 2694 8863 2746
rect 8875 2694 8927 2746
rect 8939 2694 8991 2746
rect 9003 2694 9055 2746
rect 13945 2694 13997 2746
rect 14009 2694 14061 2746
rect 14073 2694 14125 2746
rect 14137 2694 14189 2746
rect 14201 2694 14253 2746
rect 19143 2694 19195 2746
rect 19207 2694 19259 2746
rect 19271 2694 19323 2746
rect 19335 2694 19387 2746
rect 19399 2694 19451 2746
rect 6644 2592 6696 2644
rect 6736 2567 6788 2576
rect 6736 2533 6745 2567
rect 6745 2533 6779 2567
rect 6779 2533 6788 2567
rect 6736 2524 6788 2533
rect 1952 2431 2004 2440
rect 1952 2397 1961 2431
rect 1961 2397 1995 2431
rect 1995 2397 2004 2431
rect 1952 2388 2004 2397
rect 4896 2388 4948 2440
rect 3056 2320 3108 2372
rect 8300 2524 8352 2576
rect 7196 2431 7248 2440
rect 7196 2397 7205 2431
rect 7205 2397 7239 2431
rect 7239 2397 7248 2431
rect 7196 2388 7248 2397
rect 8208 2456 8260 2508
rect 9496 2524 9548 2576
rect 10324 2592 10376 2644
rect 11152 2635 11204 2644
rect 11152 2601 11161 2635
rect 11161 2601 11195 2635
rect 11195 2601 11204 2635
rect 11152 2592 11204 2601
rect 9036 2456 9088 2508
rect 9956 2524 10008 2576
rect 11060 2524 11112 2576
rect 17132 2592 17184 2644
rect 17776 2592 17828 2644
rect 20352 2592 20404 2644
rect 20628 2592 20680 2644
rect 20720 2524 20772 2576
rect 12900 2499 12952 2508
rect 12900 2465 12909 2499
rect 12909 2465 12943 2499
rect 12943 2465 12952 2499
rect 12900 2456 12952 2465
rect 2136 2295 2188 2304
rect 2136 2261 2145 2295
rect 2145 2261 2179 2295
rect 2179 2261 2188 2295
rect 2136 2252 2188 2261
rect 3884 2252 3936 2304
rect 5540 2252 5592 2304
rect 5816 2295 5868 2304
rect 5816 2261 5825 2295
rect 5825 2261 5859 2295
rect 5859 2261 5868 2295
rect 5816 2252 5868 2261
rect 8208 2320 8260 2372
rect 9036 2363 9088 2372
rect 9036 2329 9045 2363
rect 9045 2329 9079 2363
rect 9079 2329 9088 2363
rect 9036 2320 9088 2329
rect 10324 2431 10376 2440
rect 10324 2397 10339 2431
rect 10339 2397 10373 2431
rect 10373 2397 10376 2431
rect 10324 2388 10376 2397
rect 10600 2388 10652 2440
rect 19340 2388 19392 2440
rect 20628 2388 20680 2440
rect 9220 2252 9272 2304
rect 9496 2252 9548 2304
rect 11704 2252 11756 2304
rect 12624 2363 12676 2372
rect 12624 2329 12642 2363
rect 12642 2329 12676 2363
rect 12624 2320 12676 2329
rect 18144 2320 18196 2372
rect 13084 2252 13136 2304
rect 17500 2252 17552 2304
rect 20444 2252 20496 2304
rect 6148 2150 6200 2202
rect 6212 2150 6264 2202
rect 6276 2150 6328 2202
rect 6340 2150 6392 2202
rect 6404 2150 6456 2202
rect 11346 2150 11398 2202
rect 11410 2150 11462 2202
rect 11474 2150 11526 2202
rect 11538 2150 11590 2202
rect 11602 2150 11654 2202
rect 16544 2150 16596 2202
rect 16608 2150 16660 2202
rect 16672 2150 16724 2202
rect 16736 2150 16788 2202
rect 16800 2150 16852 2202
rect 21742 2150 21794 2202
rect 21806 2150 21858 2202
rect 21870 2150 21922 2202
rect 21934 2150 21986 2202
rect 21998 2150 22050 2202
rect 6460 2048 6512 2100
rect 7288 2048 7340 2100
rect 9956 2048 10008 2100
rect 18788 2048 18840 2100
rect 19340 1980 19392 2032
rect 20076 1980 20128 2032
rect 8208 1912 8260 1964
rect 13176 1912 13228 1964
rect 11704 1844 11756 1896
rect 16028 1844 16080 1896
rect 6736 1708 6788 1760
rect 14924 1708 14976 1760
rect 5540 1640 5592 1692
rect 12716 1640 12768 1692
rect 9036 1572 9088 1624
rect 15752 1572 15804 1624
rect 5816 1504 5868 1556
rect 14556 1504 14608 1556
rect 7564 1368 7616 1420
rect 8116 1368 8168 1420
rect 11980 1232 12032 1284
rect 11980 1028 12032 1080
rect 9772 892 9824 944
rect 10692 892 10744 944
<< metal2 >>
rect 2962 21312 3018 21321
rect 2962 21247 3018 21256
rect 2976 21010 3004 21247
rect 2964 21004 3016 21010
rect 2964 20946 3016 20952
rect 5908 21004 5960 21010
rect 5908 20946 5960 20952
rect 3882 20904 3938 20913
rect 3882 20839 3938 20848
rect 3896 20806 3924 20839
rect 3884 20800 3936 20806
rect 3884 20742 3936 20748
rect 5632 20800 5684 20806
rect 5632 20742 5684 20748
rect 4066 20496 4122 20505
rect 4066 20431 4122 20440
rect 3549 20156 3857 20165
rect 3549 20154 3555 20156
rect 3611 20154 3635 20156
rect 3691 20154 3715 20156
rect 3771 20154 3795 20156
rect 3851 20154 3857 20156
rect 3611 20102 3613 20154
rect 3793 20102 3795 20154
rect 3549 20100 3555 20102
rect 3611 20100 3635 20102
rect 3691 20100 3715 20102
rect 3771 20100 3795 20102
rect 3851 20100 3857 20102
rect 3238 20088 3294 20097
rect 3549 20091 3857 20100
rect 4080 20058 4108 20431
rect 5644 20058 5672 20742
rect 3238 20023 3294 20032
rect 4068 20052 4120 20058
rect 3252 19514 3280 20023
rect 4068 19994 4120 20000
rect 5632 20052 5684 20058
rect 5632 19994 5684 20000
rect 5816 19848 5868 19854
rect 5816 19790 5868 19796
rect 4158 19680 4214 19689
rect 4158 19615 4214 19624
rect 3240 19508 3292 19514
rect 3240 19450 3292 19456
rect 4066 19272 4122 19281
rect 4066 19207 4122 19216
rect 3549 19068 3857 19077
rect 3549 19066 3555 19068
rect 3611 19066 3635 19068
rect 3691 19066 3715 19068
rect 3771 19066 3795 19068
rect 3851 19066 3857 19068
rect 3611 19014 3613 19066
rect 3793 19014 3795 19066
rect 3549 19012 3555 19014
rect 3611 19012 3635 19014
rect 3691 19012 3715 19014
rect 3771 19012 3795 19014
rect 3851 19012 3857 19014
rect 3549 19003 3857 19012
rect 3974 18456 4030 18465
rect 4080 18426 4108 19207
rect 4172 18970 4200 19615
rect 5828 19446 5856 19790
rect 5816 19440 5868 19446
rect 5816 19382 5868 19388
rect 4712 19372 4764 19378
rect 4712 19314 4764 19320
rect 4160 18964 4212 18970
rect 4160 18906 4212 18912
rect 4158 18864 4214 18873
rect 4158 18799 4214 18808
rect 3974 18391 4030 18400
rect 4068 18420 4120 18426
rect 1950 18048 2006 18057
rect 1950 17983 2006 17992
rect 1964 17882 1992 17983
rect 3549 17980 3857 17989
rect 3549 17978 3555 17980
rect 3611 17978 3635 17980
rect 3691 17978 3715 17980
rect 3771 17978 3795 17980
rect 3851 17978 3857 17980
rect 3611 17926 3613 17978
rect 3793 17926 3795 17978
rect 3549 17924 3555 17926
rect 3611 17924 3635 17926
rect 3691 17924 3715 17926
rect 3771 17924 3795 17926
rect 3851 17924 3857 17926
rect 3549 17915 3857 17924
rect 3988 17882 4016 18391
rect 4068 18362 4120 18368
rect 4172 17882 4200 18799
rect 1952 17876 2004 17882
rect 1952 17818 2004 17824
rect 3976 17876 4028 17882
rect 3976 17818 4028 17824
rect 4160 17876 4212 17882
rect 4160 17818 4212 17824
rect 2228 17672 2280 17678
rect 2228 17614 2280 17620
rect 3698 17640 3754 17649
rect 1584 17332 1636 17338
rect 1584 17274 1636 17280
rect 1596 17241 1624 17274
rect 2240 17270 2268 17614
rect 3698 17575 3754 17584
rect 3712 17338 3740 17575
rect 3700 17332 3752 17338
rect 3700 17274 3752 17280
rect 4724 17270 4752 19314
rect 5816 18760 5868 18766
rect 5816 18702 5868 18708
rect 5828 17746 5856 18702
rect 5816 17740 5868 17746
rect 5816 17682 5868 17688
rect 2228 17264 2280 17270
rect 1582 17232 1638 17241
rect 2228 17206 2280 17212
rect 4712 17264 4764 17270
rect 4712 17206 4764 17212
rect 1582 17167 1638 17176
rect 4252 17128 4304 17134
rect 4252 17070 4304 17076
rect 3549 16892 3857 16901
rect 3549 16890 3555 16892
rect 3611 16890 3635 16892
rect 3691 16890 3715 16892
rect 3771 16890 3795 16892
rect 3851 16890 3857 16892
rect 3611 16838 3613 16890
rect 3793 16838 3795 16890
rect 3549 16836 3555 16838
rect 3611 16836 3635 16838
rect 3691 16836 3715 16838
rect 3771 16836 3795 16838
rect 3851 16836 3857 16838
rect 1950 16824 2006 16833
rect 3549 16827 3857 16836
rect 1950 16759 2006 16768
rect 1674 16416 1730 16425
rect 1674 16351 1730 16360
rect 1688 15706 1716 16351
rect 1964 16250 1992 16759
rect 1952 16244 2004 16250
rect 1952 16186 2004 16192
rect 2778 16008 2834 16017
rect 2778 15943 2834 15952
rect 2792 15706 2820 15943
rect 3549 15804 3857 15813
rect 3549 15802 3555 15804
rect 3611 15802 3635 15804
rect 3691 15802 3715 15804
rect 3771 15802 3795 15804
rect 3851 15802 3857 15804
rect 3611 15750 3613 15802
rect 3793 15750 3795 15802
rect 3549 15748 3555 15750
rect 3611 15748 3635 15750
rect 3691 15748 3715 15750
rect 3771 15748 3795 15750
rect 3851 15748 3857 15750
rect 3549 15739 3857 15748
rect 1676 15700 1728 15706
rect 1676 15642 1728 15648
rect 2780 15700 2832 15706
rect 2780 15642 2832 15648
rect 2228 15632 2280 15638
rect 2226 15600 2228 15609
rect 2280 15600 2282 15609
rect 2226 15535 2282 15544
rect 2872 15496 2924 15502
rect 2872 15438 2924 15444
rect 3700 15496 3752 15502
rect 3700 15438 3752 15444
rect 1490 15192 1546 15201
rect 1490 15127 1546 15136
rect 1504 14618 1532 15127
rect 2884 15094 2912 15438
rect 3712 15094 3740 15438
rect 4264 15162 4292 17070
rect 4436 17060 4488 17066
rect 4436 17002 4488 17008
rect 4448 16590 4476 17002
rect 4436 16584 4488 16590
rect 4436 16526 4488 16532
rect 5816 16584 5868 16590
rect 5816 16526 5868 16532
rect 5356 16108 5408 16114
rect 5356 16050 5408 16056
rect 5172 15904 5224 15910
rect 5172 15846 5224 15852
rect 4252 15156 4304 15162
rect 4252 15098 4304 15104
rect 2872 15088 2924 15094
rect 2872 15030 2924 15036
rect 3700 15088 3752 15094
rect 3700 15030 3752 15036
rect 2136 15020 2188 15026
rect 2136 14962 2188 14968
rect 3884 15020 3936 15026
rect 3884 14962 3936 14968
rect 4896 15020 4948 15026
rect 4896 14962 4948 14968
rect 1952 14816 2004 14822
rect 1950 14784 1952 14793
rect 2004 14784 2006 14793
rect 1950 14719 2006 14728
rect 1492 14612 1544 14618
rect 1492 14554 1544 14560
rect 2148 14482 2176 14962
rect 3549 14716 3857 14725
rect 3549 14714 3555 14716
rect 3611 14714 3635 14716
rect 3691 14714 3715 14716
rect 3771 14714 3795 14716
rect 3851 14714 3857 14716
rect 3611 14662 3613 14714
rect 3793 14662 3795 14714
rect 3549 14660 3555 14662
rect 3611 14660 3635 14662
rect 3691 14660 3715 14662
rect 3771 14660 3795 14662
rect 3851 14660 3857 14662
rect 3549 14651 3857 14660
rect 2136 14476 2188 14482
rect 2136 14418 2188 14424
rect 3332 14408 3384 14414
rect 1950 14376 2006 14385
rect 3332 14350 3384 14356
rect 1950 14311 2006 14320
rect 1964 14074 1992 14311
rect 1952 14068 2004 14074
rect 1952 14010 2004 14016
rect 2780 14068 2832 14074
rect 2780 14010 2832 14016
rect 2792 13977 2820 14010
rect 2778 13968 2834 13977
rect 2412 13932 2464 13938
rect 2778 13903 2834 13912
rect 2412 13874 2464 13880
rect 2136 13728 2188 13734
rect 2136 13670 2188 13676
rect 1952 13388 2004 13394
rect 1952 13330 2004 13336
rect 1492 13252 1544 13258
rect 1492 13194 1544 13200
rect 1504 12646 1532 13194
rect 1584 13184 1636 13190
rect 1584 13126 1636 13132
rect 1674 13152 1730 13161
rect 1492 12640 1544 12646
rect 1492 12582 1544 12588
rect 1400 12096 1452 12102
rect 1400 12038 1452 12044
rect 1412 11082 1440 12038
rect 1400 11076 1452 11082
rect 1400 11018 1452 11024
rect 1216 8900 1268 8906
rect 1216 8842 1268 8848
rect 1228 1737 1256 8842
rect 1412 5250 1440 11018
rect 1320 5222 1440 5250
rect 1320 4468 1348 5222
rect 1504 5114 1532 12582
rect 1412 5086 1532 5114
rect 1412 4593 1440 5086
rect 1490 4992 1546 5001
rect 1490 4927 1546 4936
rect 1398 4584 1454 4593
rect 1398 4519 1454 4528
rect 1320 4440 1440 4468
rect 1412 2961 1440 4440
rect 1504 3194 1532 4927
rect 1596 3777 1624 13126
rect 1674 13087 1730 13096
rect 1688 12442 1716 13087
rect 1768 12844 1820 12850
rect 1768 12786 1820 12792
rect 1676 12436 1728 12442
rect 1676 12378 1728 12384
rect 1780 11354 1808 12786
rect 1964 12306 1992 13330
rect 2148 13258 2176 13670
rect 2136 13252 2188 13258
rect 2136 13194 2188 13200
rect 2424 12918 2452 13874
rect 3148 13864 3200 13870
rect 3148 13806 3200 13812
rect 2778 13560 2834 13569
rect 2778 13495 2834 13504
rect 2504 13184 2556 13190
rect 2504 13126 2556 13132
rect 2412 12912 2464 12918
rect 2412 12854 2464 12860
rect 2320 12844 2372 12850
rect 2320 12786 2372 12792
rect 1952 12300 2004 12306
rect 1952 12242 2004 12248
rect 1950 11928 2006 11937
rect 1950 11863 2006 11872
rect 1860 11756 1912 11762
rect 1860 11698 1912 11704
rect 1768 11348 1820 11354
rect 1768 11290 1820 11296
rect 1872 9450 1900 11698
rect 1860 9444 1912 9450
rect 1860 9386 1912 9392
rect 1676 6656 1728 6662
rect 1674 6624 1676 6633
rect 1728 6624 1730 6633
rect 1674 6559 1730 6568
rect 1768 6248 1820 6254
rect 1768 6190 1820 6196
rect 1674 5808 1730 5817
rect 1674 5743 1730 5752
rect 1688 5710 1716 5743
rect 1780 5710 1808 6190
rect 1676 5704 1728 5710
rect 1676 5646 1728 5652
rect 1768 5704 1820 5710
rect 1768 5646 1820 5652
rect 1688 5370 1716 5646
rect 1676 5364 1728 5370
rect 1676 5306 1728 5312
rect 1768 5024 1820 5030
rect 1768 4966 1820 4972
rect 1582 3768 1638 3777
rect 1582 3703 1638 3712
rect 1492 3188 1544 3194
rect 1492 3130 1544 3136
rect 1398 2952 1454 2961
rect 1398 2887 1454 2896
rect 1214 1728 1270 1737
rect 1214 1663 1270 1672
rect 1780 762 1808 4966
rect 1860 4684 1912 4690
rect 1860 4626 1912 4632
rect 1872 4593 1900 4626
rect 1858 4584 1914 4593
rect 1858 4519 1914 4528
rect 1964 2446 1992 11863
rect 2332 11830 2360 12786
rect 2412 12300 2464 12306
rect 2412 12242 2464 12248
rect 2424 11830 2452 12242
rect 2320 11824 2372 11830
rect 2320 11766 2372 11772
rect 2412 11824 2464 11830
rect 2412 11766 2464 11772
rect 2228 11552 2280 11558
rect 2228 11494 2280 11500
rect 2240 11218 2268 11494
rect 2228 11212 2280 11218
rect 2228 11154 2280 11160
rect 2412 11212 2464 11218
rect 2412 11154 2464 11160
rect 2136 11008 2188 11014
rect 2136 10950 2188 10956
rect 2148 10810 2176 10950
rect 2136 10804 2188 10810
rect 2136 10746 2188 10752
rect 2228 9512 2280 9518
rect 2228 9454 2280 9460
rect 2042 7304 2098 7313
rect 2042 7239 2044 7248
rect 2096 7239 2098 7248
rect 2044 7210 2096 7216
rect 2136 5568 2188 5574
rect 2136 5510 2188 5516
rect 2148 4622 2176 5510
rect 2136 4616 2188 4622
rect 2136 4558 2188 4564
rect 2044 2848 2096 2854
rect 2044 2790 2096 2796
rect 1952 2440 2004 2446
rect 1952 2382 2004 2388
rect 2056 1737 2084 2790
rect 2240 2553 2268 9454
rect 2320 8560 2372 8566
rect 2320 8502 2372 8508
rect 2332 6866 2360 8502
rect 2424 7993 2452 11154
rect 2516 10742 2544 13126
rect 2792 12986 2820 13495
rect 3160 13394 3188 13806
rect 3240 13728 3292 13734
rect 3240 13670 3292 13676
rect 3148 13388 3200 13394
rect 3148 13330 3200 13336
rect 2780 12980 2832 12986
rect 2780 12922 2832 12928
rect 3252 12866 3280 13670
rect 3160 12838 3280 12866
rect 2778 12744 2834 12753
rect 2778 12679 2834 12688
rect 2688 12368 2740 12374
rect 2688 12310 2740 12316
rect 2700 12102 2728 12310
rect 2688 12096 2740 12102
rect 2688 12038 2740 12044
rect 2686 11792 2742 11801
rect 2686 11727 2742 11736
rect 2700 11694 2728 11727
rect 2688 11688 2740 11694
rect 2688 11630 2740 11636
rect 2504 10736 2556 10742
rect 2504 10678 2556 10684
rect 2700 10606 2728 11630
rect 2792 11098 2820 12679
rect 2962 12336 3018 12345
rect 2962 12271 3018 12280
rect 2872 12096 2924 12102
rect 2872 12038 2924 12044
rect 2884 11898 2912 12038
rect 2872 11892 2924 11898
rect 2872 11834 2924 11840
rect 2792 11070 2912 11098
rect 2780 11008 2832 11014
rect 2780 10950 2832 10956
rect 2792 10810 2820 10950
rect 2780 10804 2832 10810
rect 2780 10746 2832 10752
rect 2688 10600 2740 10606
rect 2688 10542 2740 10548
rect 2884 10266 2912 11070
rect 2872 10260 2924 10266
rect 2872 10202 2924 10208
rect 2884 10062 2912 10202
rect 2872 10056 2924 10062
rect 2872 9998 2924 10004
rect 2872 9376 2924 9382
rect 2872 9318 2924 9324
rect 2780 9104 2832 9110
rect 2700 9052 2780 9058
rect 2700 9046 2832 9052
rect 2700 9030 2820 9046
rect 2700 8378 2728 9030
rect 2780 8832 2832 8838
rect 2780 8774 2832 8780
rect 2792 8634 2820 8774
rect 2780 8628 2832 8634
rect 2780 8570 2832 8576
rect 2700 8350 2820 8378
rect 2410 7984 2466 7993
rect 2410 7919 2466 7928
rect 2688 7472 2740 7478
rect 2688 7414 2740 7420
rect 2320 6860 2372 6866
rect 2320 6802 2372 6808
rect 2332 4049 2360 6802
rect 2504 6656 2556 6662
rect 2504 6598 2556 6604
rect 2516 6458 2544 6598
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 2504 5840 2556 5846
rect 2504 5782 2556 5788
rect 2412 5568 2464 5574
rect 2412 5510 2464 5516
rect 2424 4690 2452 5510
rect 2516 5370 2544 5782
rect 2504 5364 2556 5370
rect 2504 5306 2556 5312
rect 2412 4684 2464 4690
rect 2412 4626 2464 4632
rect 2516 4554 2544 5306
rect 2700 5166 2728 7414
rect 2688 5160 2740 5166
rect 2688 5102 2740 5108
rect 2504 4548 2556 4554
rect 2504 4490 2556 4496
rect 2318 4040 2374 4049
rect 2318 3975 2374 3984
rect 2412 3732 2464 3738
rect 2412 3674 2464 3680
rect 2226 2544 2282 2553
rect 2226 2479 2282 2488
rect 2134 2408 2190 2417
rect 2134 2343 2190 2352
rect 2148 2310 2176 2343
rect 2136 2304 2188 2310
rect 2136 2246 2188 2252
rect 2042 1728 2098 1737
rect 2042 1663 2098 1672
rect 1964 870 2084 898
rect 1964 762 1992 870
rect 2056 800 2084 870
rect 2424 800 2452 3674
rect 1780 734 1992 762
rect 2042 0 2098 800
rect 2410 0 2466 800
rect 2516 762 2544 4490
rect 2688 4480 2740 4486
rect 2688 4422 2740 4428
rect 2700 4146 2728 4422
rect 2792 4185 2820 8350
rect 2884 5681 2912 9318
rect 2976 7546 3004 12271
rect 3056 12096 3108 12102
rect 3056 12038 3108 12044
rect 3068 9994 3096 12038
rect 3160 11354 3188 12838
rect 3240 12776 3292 12782
rect 3240 12718 3292 12724
rect 3252 12238 3280 12718
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 3148 11348 3200 11354
rect 3148 11290 3200 11296
rect 3160 10742 3188 11290
rect 3148 10736 3200 10742
rect 3148 10678 3200 10684
rect 3056 9988 3108 9994
rect 3056 9930 3108 9936
rect 3068 8922 3096 9930
rect 3160 9110 3188 10678
rect 3344 10418 3372 14350
rect 3549 13628 3857 13637
rect 3549 13626 3555 13628
rect 3611 13626 3635 13628
rect 3691 13626 3715 13628
rect 3771 13626 3795 13628
rect 3851 13626 3857 13628
rect 3611 13574 3613 13626
rect 3793 13574 3795 13626
rect 3549 13572 3555 13574
rect 3611 13572 3635 13574
rect 3691 13572 3715 13574
rect 3771 13572 3795 13574
rect 3851 13572 3857 13574
rect 3549 13563 3857 13572
rect 3549 12540 3857 12549
rect 3549 12538 3555 12540
rect 3611 12538 3635 12540
rect 3691 12538 3715 12540
rect 3771 12538 3795 12540
rect 3851 12538 3857 12540
rect 3611 12486 3613 12538
rect 3793 12486 3795 12538
rect 3549 12484 3555 12486
rect 3611 12484 3635 12486
rect 3691 12484 3715 12486
rect 3771 12484 3795 12486
rect 3851 12484 3857 12486
rect 3549 12475 3857 12484
rect 3422 11520 3478 11529
rect 3422 11455 3478 11464
rect 3436 11082 3464 11455
rect 3549 11452 3857 11461
rect 3549 11450 3555 11452
rect 3611 11450 3635 11452
rect 3691 11450 3715 11452
rect 3771 11450 3795 11452
rect 3851 11450 3857 11452
rect 3611 11398 3613 11450
rect 3793 11398 3795 11450
rect 3549 11396 3555 11398
rect 3611 11396 3635 11398
rect 3691 11396 3715 11398
rect 3771 11396 3795 11398
rect 3851 11396 3857 11398
rect 3549 11387 3857 11396
rect 3896 11098 3924 14962
rect 4068 14272 4120 14278
rect 4068 14214 4120 14220
rect 4252 14272 4304 14278
rect 4252 14214 4304 14220
rect 4804 14272 4856 14278
rect 4804 14214 4856 14220
rect 4080 14074 4108 14214
rect 4068 14068 4120 14074
rect 4068 14010 4120 14016
rect 4264 13530 4292 14214
rect 4816 14006 4844 14214
rect 4908 14074 4936 14962
rect 5184 14958 5212 15846
rect 5368 15570 5396 16050
rect 5356 15564 5408 15570
rect 5356 15506 5408 15512
rect 5828 15162 5856 16526
rect 5920 15706 5948 20946
rect 6148 20700 6456 20709
rect 6148 20698 6154 20700
rect 6210 20698 6234 20700
rect 6290 20698 6314 20700
rect 6370 20698 6394 20700
rect 6450 20698 6456 20700
rect 6210 20646 6212 20698
rect 6392 20646 6394 20698
rect 6148 20644 6154 20646
rect 6210 20644 6234 20646
rect 6290 20644 6314 20646
rect 6370 20644 6394 20646
rect 6450 20644 6456 20646
rect 6148 20635 6456 20644
rect 11346 20700 11654 20709
rect 11346 20698 11352 20700
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11648 20698 11654 20700
rect 11408 20646 11410 20698
rect 11590 20646 11592 20698
rect 11346 20644 11352 20646
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11648 20644 11654 20646
rect 11346 20635 11654 20644
rect 16544 20700 16852 20709
rect 16544 20698 16550 20700
rect 16606 20698 16630 20700
rect 16686 20698 16710 20700
rect 16766 20698 16790 20700
rect 16846 20698 16852 20700
rect 16606 20646 16608 20698
rect 16788 20646 16790 20698
rect 16544 20644 16550 20646
rect 16606 20644 16630 20646
rect 16686 20644 16710 20646
rect 16766 20644 16790 20646
rect 16846 20644 16852 20646
rect 16544 20635 16852 20644
rect 21742 20700 22050 20709
rect 21742 20698 21748 20700
rect 21804 20698 21828 20700
rect 21884 20698 21908 20700
rect 21964 20698 21988 20700
rect 22044 20698 22050 20700
rect 21804 20646 21806 20698
rect 21986 20646 21988 20698
rect 21742 20644 21748 20646
rect 21804 20644 21828 20646
rect 21884 20644 21908 20646
rect 21964 20644 21988 20646
rect 22044 20644 22050 20646
rect 21742 20635 22050 20644
rect 8747 20156 9055 20165
rect 8747 20154 8753 20156
rect 8809 20154 8833 20156
rect 8889 20154 8913 20156
rect 8969 20154 8993 20156
rect 9049 20154 9055 20156
rect 8809 20102 8811 20154
rect 8991 20102 8993 20154
rect 8747 20100 8753 20102
rect 8809 20100 8833 20102
rect 8889 20100 8913 20102
rect 8969 20100 8993 20102
rect 9049 20100 9055 20102
rect 8747 20091 9055 20100
rect 13945 20156 14253 20165
rect 13945 20154 13951 20156
rect 14007 20154 14031 20156
rect 14087 20154 14111 20156
rect 14167 20154 14191 20156
rect 14247 20154 14253 20156
rect 14007 20102 14009 20154
rect 14189 20102 14191 20154
rect 13945 20100 13951 20102
rect 14007 20100 14031 20102
rect 14087 20100 14111 20102
rect 14167 20100 14191 20102
rect 14247 20100 14253 20102
rect 13945 20091 14253 20100
rect 19143 20156 19451 20165
rect 19143 20154 19149 20156
rect 19205 20154 19229 20156
rect 19285 20154 19309 20156
rect 19365 20154 19389 20156
rect 19445 20154 19451 20156
rect 19205 20102 19207 20154
rect 19387 20102 19389 20154
rect 19143 20100 19149 20102
rect 19205 20100 19229 20102
rect 19285 20100 19309 20102
rect 19365 20100 19389 20102
rect 19445 20100 19451 20102
rect 19143 20091 19451 20100
rect 10416 19848 10468 19854
rect 10416 19790 10468 19796
rect 6148 19612 6456 19621
rect 6148 19610 6154 19612
rect 6210 19610 6234 19612
rect 6290 19610 6314 19612
rect 6370 19610 6394 19612
rect 6450 19610 6456 19612
rect 6210 19558 6212 19610
rect 6392 19558 6394 19610
rect 6148 19556 6154 19558
rect 6210 19556 6234 19558
rect 6290 19556 6314 19558
rect 6370 19556 6394 19558
rect 6450 19556 6456 19558
rect 6148 19547 6456 19556
rect 9128 19372 9180 19378
rect 9128 19314 9180 19320
rect 8747 19068 9055 19077
rect 8747 19066 8753 19068
rect 8809 19066 8833 19068
rect 8889 19066 8913 19068
rect 8969 19066 8993 19068
rect 9049 19066 9055 19068
rect 8809 19014 8811 19066
rect 8991 19014 8993 19066
rect 8747 19012 8753 19014
rect 8809 19012 8833 19014
rect 8889 19012 8913 19014
rect 8969 19012 8993 19014
rect 9049 19012 9055 19014
rect 8747 19003 9055 19012
rect 6148 18524 6456 18533
rect 6148 18522 6154 18524
rect 6210 18522 6234 18524
rect 6290 18522 6314 18524
rect 6370 18522 6394 18524
rect 6450 18522 6456 18524
rect 6210 18470 6212 18522
rect 6392 18470 6394 18522
rect 6148 18468 6154 18470
rect 6210 18468 6234 18470
rect 6290 18468 6314 18470
rect 6370 18468 6394 18470
rect 6450 18468 6456 18470
rect 6148 18459 6456 18468
rect 7656 18284 7708 18290
rect 7656 18226 7708 18232
rect 6736 17672 6788 17678
rect 6736 17614 6788 17620
rect 6000 17604 6052 17610
rect 6000 17546 6052 17552
rect 6012 16590 6040 17546
rect 6148 17436 6456 17445
rect 6148 17434 6154 17436
rect 6210 17434 6234 17436
rect 6290 17434 6314 17436
rect 6370 17434 6394 17436
rect 6450 17434 6456 17436
rect 6210 17382 6212 17434
rect 6392 17382 6394 17434
rect 6148 17380 6154 17382
rect 6210 17380 6234 17382
rect 6290 17380 6314 17382
rect 6370 17380 6394 17382
rect 6450 17380 6456 17382
rect 6148 17371 6456 17380
rect 6644 17196 6696 17202
rect 6644 17138 6696 17144
rect 6000 16584 6052 16590
rect 6000 16526 6052 16532
rect 6148 16348 6456 16357
rect 6148 16346 6154 16348
rect 6210 16346 6234 16348
rect 6290 16346 6314 16348
rect 6370 16346 6394 16348
rect 6450 16346 6456 16348
rect 6210 16294 6212 16346
rect 6392 16294 6394 16346
rect 6148 16292 6154 16294
rect 6210 16292 6234 16294
rect 6290 16292 6314 16294
rect 6370 16292 6394 16294
rect 6450 16292 6456 16294
rect 6148 16283 6456 16292
rect 6656 15706 6684 17138
rect 6748 16522 6776 17614
rect 7668 16590 7696 18226
rect 8747 17980 9055 17989
rect 8747 17978 8753 17980
rect 8809 17978 8833 17980
rect 8889 17978 8913 17980
rect 8969 17978 8993 17980
rect 9049 17978 9055 17980
rect 8809 17926 8811 17978
rect 8991 17926 8993 17978
rect 8747 17924 8753 17926
rect 8809 17924 8833 17926
rect 8889 17924 8913 17926
rect 8969 17924 8993 17926
rect 9049 17924 9055 17926
rect 8747 17915 9055 17924
rect 8747 16892 9055 16901
rect 8747 16890 8753 16892
rect 8809 16890 8833 16892
rect 8889 16890 8913 16892
rect 8969 16890 8993 16892
rect 9049 16890 9055 16892
rect 8809 16838 8811 16890
rect 8991 16838 8993 16890
rect 8747 16836 8753 16838
rect 8809 16836 8833 16838
rect 8889 16836 8913 16838
rect 8969 16836 8993 16838
rect 9049 16836 9055 16838
rect 8747 16827 9055 16836
rect 6828 16584 6880 16590
rect 6828 16526 6880 16532
rect 7196 16584 7248 16590
rect 7196 16526 7248 16532
rect 7656 16584 7708 16590
rect 7656 16526 7708 16532
rect 8576 16584 8628 16590
rect 8576 16526 8628 16532
rect 6736 16516 6788 16522
rect 6736 16458 6788 16464
rect 5908 15700 5960 15706
rect 5908 15642 5960 15648
rect 6644 15700 6696 15706
rect 6644 15642 6696 15648
rect 5816 15156 5868 15162
rect 5816 15098 5868 15104
rect 5920 15026 5948 15642
rect 6000 15428 6052 15434
rect 6000 15370 6052 15376
rect 5908 15020 5960 15026
rect 5908 14962 5960 14968
rect 5172 14952 5224 14958
rect 5172 14894 5224 14900
rect 5724 14952 5776 14958
rect 5724 14894 5776 14900
rect 4896 14068 4948 14074
rect 4896 14010 4948 14016
rect 4804 14000 4856 14006
rect 4804 13942 4856 13948
rect 4804 13796 4856 13802
rect 4804 13738 4856 13744
rect 4252 13524 4304 13530
rect 4252 13466 4304 13472
rect 4816 13394 4844 13738
rect 4804 13388 4856 13394
rect 4804 13330 4856 13336
rect 4528 13320 4580 13326
rect 4528 13262 4580 13268
rect 4068 13252 4120 13258
rect 4068 13194 4120 13200
rect 3976 12096 4028 12102
rect 4080 12084 4108 13194
rect 4344 12844 4396 12850
rect 4344 12786 4396 12792
rect 4356 12442 4384 12786
rect 4344 12436 4396 12442
rect 4344 12378 4396 12384
rect 4028 12056 4108 12084
rect 3976 12038 4028 12044
rect 3988 11898 4016 12038
rect 3976 11892 4028 11898
rect 3976 11834 4028 11840
rect 4540 11354 4568 13262
rect 4816 12918 4844 13330
rect 4988 13184 5040 13190
rect 4988 13126 5040 13132
rect 4804 12912 4856 12918
rect 4804 12854 4856 12860
rect 5000 12646 5028 13126
rect 4988 12640 5040 12646
rect 4986 12608 4988 12617
rect 5040 12608 5042 12617
rect 4986 12543 5042 12552
rect 5184 12442 5212 14894
rect 5540 14816 5592 14822
rect 5540 14758 5592 14764
rect 5264 13932 5316 13938
rect 5264 13874 5316 13880
rect 5276 13394 5304 13874
rect 5552 13870 5580 14758
rect 5736 14278 5764 14894
rect 5724 14272 5776 14278
rect 5724 14214 5776 14220
rect 5540 13864 5592 13870
rect 5540 13806 5592 13812
rect 5264 13388 5316 13394
rect 5264 13330 5316 13336
rect 5264 12640 5316 12646
rect 5264 12582 5316 12588
rect 5172 12436 5224 12442
rect 5172 12378 5224 12384
rect 5172 12300 5224 12306
rect 5172 12242 5224 12248
rect 4712 12096 4764 12102
rect 4712 12038 4764 12044
rect 4724 11898 4752 12038
rect 4712 11892 4764 11898
rect 4712 11834 4764 11840
rect 4528 11348 4580 11354
rect 4528 11290 4580 11296
rect 4068 11144 4120 11150
rect 4066 11112 4068 11121
rect 4120 11112 4122 11121
rect 3424 11076 3476 11082
rect 3896 11070 4016 11098
rect 3424 11018 3476 11024
rect 3884 11008 3936 11014
rect 3884 10950 3936 10956
rect 3896 10810 3924 10950
rect 3884 10804 3936 10810
rect 3884 10746 3936 10752
rect 3422 10704 3478 10713
rect 3422 10639 3478 10648
rect 3436 10470 3464 10639
rect 3252 10390 3372 10418
rect 3424 10464 3476 10470
rect 3424 10406 3476 10412
rect 3252 9722 3280 10390
rect 3330 10296 3386 10305
rect 3436 10266 3464 10406
rect 3549 10364 3857 10373
rect 3549 10362 3555 10364
rect 3611 10362 3635 10364
rect 3691 10362 3715 10364
rect 3771 10362 3795 10364
rect 3851 10362 3857 10364
rect 3611 10310 3613 10362
rect 3793 10310 3795 10362
rect 3549 10308 3555 10310
rect 3611 10308 3635 10310
rect 3691 10308 3715 10310
rect 3771 10308 3795 10310
rect 3851 10308 3857 10310
rect 3549 10299 3857 10308
rect 3330 10231 3386 10240
rect 3424 10260 3476 10266
rect 3240 9716 3292 9722
rect 3240 9658 3292 9664
rect 3240 9580 3292 9586
rect 3240 9522 3292 9528
rect 3252 9178 3280 9522
rect 3240 9172 3292 9178
rect 3240 9114 3292 9120
rect 3148 9104 3200 9110
rect 3148 9046 3200 9052
rect 3068 8894 3188 8922
rect 2964 7540 3016 7546
rect 2964 7482 3016 7488
rect 2964 7404 3016 7410
rect 2964 7346 3016 7352
rect 2976 7206 3004 7346
rect 2964 7200 3016 7206
rect 2964 7142 3016 7148
rect 2976 5846 3004 7142
rect 3054 7032 3110 7041
rect 3054 6967 3110 6976
rect 2964 5840 3016 5846
rect 2964 5782 3016 5788
rect 2870 5672 2926 5681
rect 2870 5607 2926 5616
rect 2872 5568 2924 5574
rect 2872 5510 2924 5516
rect 2884 5370 2912 5510
rect 2872 5364 2924 5370
rect 2872 5306 2924 5312
rect 2778 4176 2834 4185
rect 2688 4140 2740 4146
rect 2778 4111 2834 4120
rect 2688 4082 2740 4088
rect 2596 2848 2648 2854
rect 2596 2790 2648 2796
rect 2608 1873 2636 2790
rect 3068 2378 3096 6967
rect 3160 5030 3188 8894
rect 3344 8634 3372 10231
rect 3424 10202 3476 10208
rect 3700 10124 3752 10130
rect 3700 10066 3752 10072
rect 3608 9920 3660 9926
rect 3608 9862 3660 9868
rect 3620 9722 3648 9862
rect 3424 9716 3476 9722
rect 3424 9658 3476 9664
rect 3608 9716 3660 9722
rect 3608 9658 3660 9664
rect 3332 8628 3384 8634
rect 3332 8570 3384 8576
rect 3436 8498 3464 9658
rect 3620 9518 3648 9658
rect 3608 9512 3660 9518
rect 3608 9454 3660 9460
rect 3712 9382 3740 10066
rect 3882 9888 3938 9897
rect 3882 9823 3938 9832
rect 3790 9480 3846 9489
rect 3790 9415 3792 9424
rect 3844 9415 3846 9424
rect 3792 9386 3844 9392
rect 3700 9376 3752 9382
rect 3700 9318 3752 9324
rect 3549 9276 3857 9285
rect 3549 9274 3555 9276
rect 3611 9274 3635 9276
rect 3691 9274 3715 9276
rect 3771 9274 3795 9276
rect 3851 9274 3857 9276
rect 3611 9222 3613 9274
rect 3793 9222 3795 9274
rect 3549 9220 3555 9222
rect 3611 9220 3635 9222
rect 3691 9220 3715 9222
rect 3771 9220 3795 9222
rect 3851 9220 3857 9222
rect 3549 9211 3857 9220
rect 3424 8492 3476 8498
rect 3424 8434 3476 8440
rect 3330 8256 3386 8265
rect 3330 8191 3386 8200
rect 3240 7948 3292 7954
rect 3240 7890 3292 7896
rect 3252 7750 3280 7890
rect 3240 7744 3292 7750
rect 3240 7686 3292 7692
rect 3252 5794 3280 7686
rect 3344 5914 3372 8191
rect 3549 8188 3857 8197
rect 3549 8186 3555 8188
rect 3611 8186 3635 8188
rect 3691 8186 3715 8188
rect 3771 8186 3795 8188
rect 3851 8186 3857 8188
rect 3611 8134 3613 8186
rect 3793 8134 3795 8186
rect 3549 8132 3555 8134
rect 3611 8132 3635 8134
rect 3691 8132 3715 8134
rect 3771 8132 3795 8134
rect 3851 8132 3857 8134
rect 3549 8123 3857 8132
rect 3896 7886 3924 9823
rect 3988 9654 4016 11070
rect 4066 11047 4122 11056
rect 4344 11076 4396 11082
rect 4344 11018 4396 11024
rect 4066 10024 4122 10033
rect 4066 9959 4122 9968
rect 4080 9926 4108 9959
rect 4068 9920 4120 9926
rect 4068 9862 4120 9868
rect 3976 9648 4028 9654
rect 3976 9590 4028 9596
rect 4252 9580 4304 9586
rect 4252 9522 4304 9528
rect 3976 9512 4028 9518
rect 4068 9512 4120 9518
rect 3976 9454 4028 9460
rect 4066 9480 4068 9489
rect 4120 9480 4122 9489
rect 3988 9178 4016 9454
rect 4066 9415 4122 9424
rect 3976 9172 4028 9178
rect 3976 9114 4028 9120
rect 4066 9072 4122 9081
rect 4066 9007 4122 9016
rect 4080 8906 4108 9007
rect 4264 8974 4292 9522
rect 4252 8968 4304 8974
rect 4252 8910 4304 8916
rect 4068 8900 4120 8906
rect 4068 8842 4120 8848
rect 4356 8514 4384 11018
rect 4896 11008 4948 11014
rect 4896 10950 4948 10956
rect 4908 10810 4936 10950
rect 4896 10804 4948 10810
rect 4896 10746 4948 10752
rect 4896 10600 4948 10606
rect 4896 10542 4948 10548
rect 4528 10532 4580 10538
rect 4528 10474 4580 10480
rect 4436 9920 4488 9926
rect 4436 9862 4488 9868
rect 4448 8974 4476 9862
rect 4436 8968 4488 8974
rect 4436 8910 4488 8916
rect 3976 8492 4028 8498
rect 3976 8434 4028 8440
rect 4252 8492 4304 8498
rect 4356 8486 4476 8514
rect 4252 8434 4304 8440
rect 3988 8265 4016 8434
rect 4160 8356 4212 8362
rect 4160 8298 4212 8304
rect 3974 8256 4030 8265
rect 3974 8191 4030 8200
rect 3884 7880 3936 7886
rect 3884 7822 3936 7828
rect 3974 7848 4030 7857
rect 3424 7812 3476 7818
rect 3974 7783 4030 7792
rect 3424 7754 3476 7760
rect 3436 7449 3464 7754
rect 3884 7744 3936 7750
rect 3884 7686 3936 7692
rect 3422 7440 3478 7449
rect 3422 7375 3478 7384
rect 3549 7100 3857 7109
rect 3549 7098 3555 7100
rect 3611 7098 3635 7100
rect 3691 7098 3715 7100
rect 3771 7098 3795 7100
rect 3851 7098 3857 7100
rect 3611 7046 3613 7098
rect 3793 7046 3795 7098
rect 3549 7044 3555 7046
rect 3611 7044 3635 7046
rect 3691 7044 3715 7046
rect 3771 7044 3795 7046
rect 3851 7044 3857 7046
rect 3549 7035 3857 7044
rect 3549 6012 3857 6021
rect 3549 6010 3555 6012
rect 3611 6010 3635 6012
rect 3691 6010 3715 6012
rect 3771 6010 3795 6012
rect 3851 6010 3857 6012
rect 3611 5958 3613 6010
rect 3793 5958 3795 6010
rect 3549 5956 3555 5958
rect 3611 5956 3635 5958
rect 3691 5956 3715 5958
rect 3771 5956 3795 5958
rect 3851 5956 3857 5958
rect 3549 5947 3857 5956
rect 3332 5908 3384 5914
rect 3896 5896 3924 7686
rect 3988 6934 4016 7783
rect 3976 6928 4028 6934
rect 3976 6870 4028 6876
rect 4172 6866 4200 8298
rect 4264 8090 4292 8434
rect 4344 8424 4396 8430
rect 4344 8366 4396 8372
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4356 7546 4384 8366
rect 4344 7540 4396 7546
rect 4344 7482 4396 7488
rect 4252 6996 4304 7002
rect 4252 6938 4304 6944
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 4158 6216 4214 6225
rect 4158 6151 4214 6160
rect 3332 5850 3384 5856
rect 3804 5868 3924 5896
rect 3252 5766 3464 5794
rect 3330 5672 3386 5681
rect 3240 5636 3292 5642
rect 3330 5607 3386 5616
rect 3240 5578 3292 5584
rect 3252 5370 3280 5578
rect 3240 5364 3292 5370
rect 3240 5306 3292 5312
rect 3148 5024 3200 5030
rect 3148 4966 3200 4972
rect 3148 3596 3200 3602
rect 3148 3538 3200 3544
rect 3056 2372 3108 2378
rect 3056 2314 3108 2320
rect 2594 1864 2650 1873
rect 2594 1799 2650 1808
rect 2700 870 2820 898
rect 2700 762 2728 870
rect 2792 800 2820 870
rect 3160 800 3188 3538
rect 3344 3369 3372 5607
rect 3436 5370 3464 5766
rect 3424 5364 3476 5370
rect 3424 5306 3476 5312
rect 3436 4010 3464 5306
rect 3804 5234 3832 5868
rect 4066 5400 4122 5409
rect 4066 5335 4122 5344
rect 4080 5302 4108 5335
rect 4068 5296 4120 5302
rect 4068 5238 4120 5244
rect 3792 5228 3844 5234
rect 3792 5170 3844 5176
rect 3884 5160 3936 5166
rect 3884 5102 3936 5108
rect 3549 4924 3857 4933
rect 3549 4922 3555 4924
rect 3611 4922 3635 4924
rect 3691 4922 3715 4924
rect 3771 4922 3795 4924
rect 3851 4922 3857 4924
rect 3611 4870 3613 4922
rect 3793 4870 3795 4922
rect 3549 4868 3555 4870
rect 3611 4868 3635 4870
rect 3691 4868 3715 4870
rect 3771 4868 3795 4870
rect 3851 4868 3857 4870
rect 3549 4859 3857 4868
rect 3896 4758 3924 5102
rect 3976 5024 4028 5030
rect 3976 4966 4028 4972
rect 3884 4752 3936 4758
rect 3884 4694 3936 4700
rect 3424 4004 3476 4010
rect 3424 3946 3476 3952
rect 3330 3360 3386 3369
rect 3330 3295 3386 3304
rect 3436 1442 3464 3946
rect 3884 3936 3936 3942
rect 3884 3878 3936 3884
rect 3549 3836 3857 3845
rect 3549 3834 3555 3836
rect 3611 3834 3635 3836
rect 3691 3834 3715 3836
rect 3771 3834 3795 3836
rect 3851 3834 3857 3836
rect 3611 3782 3613 3834
rect 3793 3782 3795 3834
rect 3549 3780 3555 3782
rect 3611 3780 3635 3782
rect 3691 3780 3715 3782
rect 3771 3780 3795 3782
rect 3851 3780 3857 3782
rect 3549 3771 3857 3780
rect 3549 2748 3857 2757
rect 3549 2746 3555 2748
rect 3611 2746 3635 2748
rect 3691 2746 3715 2748
rect 3771 2746 3795 2748
rect 3851 2746 3857 2748
rect 3611 2694 3613 2746
rect 3793 2694 3795 2746
rect 3549 2692 3555 2694
rect 3611 2692 3635 2694
rect 3691 2692 3715 2694
rect 3771 2692 3795 2694
rect 3851 2692 3857 2694
rect 3549 2683 3857 2692
rect 3896 2310 3924 3878
rect 3884 2304 3936 2310
rect 3884 2246 3936 2252
rect 3436 1414 3556 1442
rect 3528 800 3556 1414
rect 3896 800 3924 2246
rect 3988 2145 4016 4966
rect 4172 4146 4200 6151
rect 4264 5681 4292 6938
rect 4344 6792 4396 6798
rect 4344 6734 4396 6740
rect 4250 5672 4306 5681
rect 4250 5607 4306 5616
rect 4252 5092 4304 5098
rect 4252 5034 4304 5040
rect 4264 4486 4292 5034
rect 4252 4480 4304 4486
rect 4252 4422 4304 4428
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 3974 2136 4030 2145
rect 3974 2071 4030 2080
rect 4264 800 4292 4422
rect 4356 3738 4384 6734
rect 4344 3732 4396 3738
rect 4344 3674 4396 3680
rect 4356 2774 4384 3674
rect 4448 3058 4476 8486
rect 4540 7478 4568 10474
rect 4620 9920 4672 9926
rect 4620 9862 4672 9868
rect 4632 9722 4660 9862
rect 4620 9716 4672 9722
rect 4620 9658 4672 9664
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4724 9042 4752 9318
rect 4908 9178 4936 10542
rect 5080 9512 5132 9518
rect 5080 9454 5132 9460
rect 4896 9172 4948 9178
rect 4896 9114 4948 9120
rect 4712 9036 4764 9042
rect 4712 8978 4764 8984
rect 4988 9036 5040 9042
rect 4988 8978 5040 8984
rect 4896 8288 4948 8294
rect 4896 8230 4948 8236
rect 4620 7948 4672 7954
rect 4620 7890 4672 7896
rect 4528 7472 4580 7478
rect 4528 7414 4580 7420
rect 4632 7410 4660 7890
rect 4908 7546 4936 8230
rect 5000 7857 5028 8978
rect 5092 8362 5120 9454
rect 5184 9081 5212 12242
rect 5276 12238 5304 12582
rect 5448 12436 5500 12442
rect 5448 12378 5500 12384
rect 5264 12232 5316 12238
rect 5264 12174 5316 12180
rect 5356 12096 5408 12102
rect 5356 12038 5408 12044
rect 5368 11898 5396 12038
rect 5356 11892 5408 11898
rect 5356 11834 5408 11840
rect 5356 11620 5408 11626
rect 5356 11562 5408 11568
rect 5264 10124 5316 10130
rect 5264 10066 5316 10072
rect 5276 9518 5304 10066
rect 5264 9512 5316 9518
rect 5264 9454 5316 9460
rect 5170 9072 5226 9081
rect 5170 9007 5226 9016
rect 5276 8922 5304 9454
rect 5184 8894 5304 8922
rect 5080 8356 5132 8362
rect 5080 8298 5132 8304
rect 4986 7848 5042 7857
rect 4986 7783 5042 7792
rect 4896 7540 4948 7546
rect 4896 7482 4948 7488
rect 4802 7440 4858 7449
rect 4620 7404 4672 7410
rect 4802 7375 4858 7384
rect 4620 7346 4672 7352
rect 4816 7342 4844 7375
rect 4804 7336 4856 7342
rect 4804 7278 4856 7284
rect 4988 7336 5040 7342
rect 4988 7278 5040 7284
rect 5000 7002 5028 7278
rect 4988 6996 5040 7002
rect 4988 6938 5040 6944
rect 5092 6882 5120 8298
rect 5000 6854 5120 6882
rect 5184 6866 5212 8894
rect 5264 8832 5316 8838
rect 5264 8774 5316 8780
rect 5276 8634 5304 8774
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5264 8084 5316 8090
rect 5264 8026 5316 8032
rect 5276 7750 5304 8026
rect 5264 7744 5316 7750
rect 5264 7686 5316 7692
rect 5172 6860 5224 6866
rect 4528 6656 4580 6662
rect 4528 6598 4580 6604
rect 4540 6322 4568 6598
rect 4528 6316 4580 6322
rect 4528 6258 4580 6264
rect 4620 6248 4672 6254
rect 4620 6190 4672 6196
rect 4528 5772 4580 5778
rect 4528 5714 4580 5720
rect 4540 5642 4568 5714
rect 4528 5636 4580 5642
rect 4528 5578 4580 5584
rect 4528 4820 4580 4826
rect 4528 4762 4580 4768
rect 4540 3670 4568 4762
rect 4528 3664 4580 3670
rect 4528 3606 4580 3612
rect 4632 3058 4660 6190
rect 4804 5568 4856 5574
rect 4804 5510 4856 5516
rect 4816 5370 4844 5510
rect 4804 5364 4856 5370
rect 4804 5306 4856 5312
rect 4896 5364 4948 5370
rect 4896 5306 4948 5312
rect 4908 5234 4936 5306
rect 4896 5228 4948 5234
rect 4896 5170 4948 5176
rect 4908 4826 4936 5170
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 4816 3505 4844 4082
rect 4896 4072 4948 4078
rect 4896 4014 4948 4020
rect 4802 3496 4858 3505
rect 4802 3431 4858 3440
rect 4804 3392 4856 3398
rect 4804 3334 4856 3340
rect 4816 3126 4844 3334
rect 4804 3120 4856 3126
rect 4804 3062 4856 3068
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 4356 2746 4660 2774
rect 4632 800 4660 2746
rect 4908 2446 4936 4014
rect 4896 2440 4948 2446
rect 4896 2382 4948 2388
rect 5000 800 5028 6854
rect 5172 6802 5224 6808
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 5172 6656 5224 6662
rect 5172 6598 5224 6604
rect 5080 6112 5132 6118
rect 5080 6054 5132 6060
rect 5092 3534 5120 6054
rect 5184 5794 5212 6598
rect 5276 6390 5304 6734
rect 5264 6384 5316 6390
rect 5264 6326 5316 6332
rect 5264 6248 5316 6254
rect 5264 6190 5316 6196
rect 5276 5914 5304 6190
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 5184 5766 5304 5794
rect 5172 5568 5224 5574
rect 5172 5510 5224 5516
rect 5184 4010 5212 5510
rect 5276 5234 5304 5766
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 5276 4826 5304 5170
rect 5264 4820 5316 4826
rect 5264 4762 5316 4768
rect 5172 4004 5224 4010
rect 5172 3946 5224 3952
rect 5080 3528 5132 3534
rect 5080 3470 5132 3476
rect 5368 800 5396 11562
rect 5460 8537 5488 12378
rect 5552 11506 5580 13806
rect 5920 13258 5948 14962
rect 5908 13252 5960 13258
rect 5908 13194 5960 13200
rect 5816 13184 5868 13190
rect 5816 13126 5868 13132
rect 5724 12776 5776 12782
rect 5724 12718 5776 12724
rect 5632 12708 5684 12714
rect 5632 12650 5684 12656
rect 5644 11694 5672 12650
rect 5736 12442 5764 12718
rect 5724 12436 5776 12442
rect 5724 12378 5776 12384
rect 5828 11898 5856 13126
rect 5920 12238 5948 13194
rect 5908 12232 5960 12238
rect 5908 12174 5960 12180
rect 6012 11898 6040 15370
rect 6148 15260 6456 15269
rect 6148 15258 6154 15260
rect 6210 15258 6234 15260
rect 6290 15258 6314 15260
rect 6370 15258 6394 15260
rect 6450 15258 6456 15260
rect 6210 15206 6212 15258
rect 6392 15206 6394 15258
rect 6148 15204 6154 15206
rect 6210 15204 6234 15206
rect 6290 15204 6314 15206
rect 6370 15204 6394 15206
rect 6450 15204 6456 15206
rect 6148 15195 6456 15204
rect 6552 14272 6604 14278
rect 6552 14214 6604 14220
rect 6148 14172 6456 14181
rect 6148 14170 6154 14172
rect 6210 14170 6234 14172
rect 6290 14170 6314 14172
rect 6370 14170 6394 14172
rect 6450 14170 6456 14172
rect 6210 14118 6212 14170
rect 6392 14118 6394 14170
rect 6148 14116 6154 14118
rect 6210 14116 6234 14118
rect 6290 14116 6314 14118
rect 6370 14116 6394 14118
rect 6450 14116 6456 14118
rect 6148 14107 6456 14116
rect 6184 14000 6236 14006
rect 6564 13977 6592 14214
rect 6184 13942 6236 13948
rect 6550 13968 6606 13977
rect 6196 13326 6224 13942
rect 6550 13903 6606 13912
rect 6644 13864 6696 13870
rect 6644 13806 6696 13812
rect 6552 13388 6604 13394
rect 6552 13330 6604 13336
rect 6184 13320 6236 13326
rect 6184 13262 6236 13268
rect 6148 13084 6456 13093
rect 6148 13082 6154 13084
rect 6210 13082 6234 13084
rect 6290 13082 6314 13084
rect 6370 13082 6394 13084
rect 6450 13082 6456 13084
rect 6210 13030 6212 13082
rect 6392 13030 6394 13082
rect 6148 13028 6154 13030
rect 6210 13028 6234 13030
rect 6290 13028 6314 13030
rect 6370 13028 6394 13030
rect 6450 13028 6456 13030
rect 6148 13019 6456 13028
rect 6368 12640 6420 12646
rect 6368 12582 6420 12588
rect 6380 12442 6408 12582
rect 6368 12436 6420 12442
rect 6368 12378 6420 12384
rect 6564 12374 6592 13330
rect 6552 12368 6604 12374
rect 6552 12310 6604 12316
rect 6656 12102 6684 13806
rect 6840 12442 6868 16526
rect 7104 15088 7156 15094
rect 7104 15030 7156 15036
rect 7116 12866 7144 15030
rect 7208 13530 7236 16526
rect 7748 15496 7800 15502
rect 7748 15438 7800 15444
rect 7380 14952 7432 14958
rect 7380 14894 7432 14900
rect 7392 14074 7420 14894
rect 7380 14068 7432 14074
rect 7380 14010 7432 14016
rect 7656 14000 7708 14006
rect 7656 13942 7708 13948
rect 7196 13524 7248 13530
rect 7196 13466 7248 13472
rect 7668 13462 7696 13942
rect 7656 13456 7708 13462
rect 7656 13398 7708 13404
rect 7656 12980 7708 12986
rect 7656 12922 7708 12928
rect 7116 12838 7236 12866
rect 7104 12776 7156 12782
rect 7104 12718 7156 12724
rect 6828 12436 6880 12442
rect 6828 12378 6880 12384
rect 7116 12238 7144 12718
rect 7104 12232 7156 12238
rect 7104 12174 7156 12180
rect 6644 12096 6696 12102
rect 6644 12038 6696 12044
rect 6148 11996 6456 12005
rect 6148 11994 6154 11996
rect 6210 11994 6234 11996
rect 6290 11994 6314 11996
rect 6370 11994 6394 11996
rect 6450 11994 6456 11996
rect 6210 11942 6212 11994
rect 6392 11942 6394 11994
rect 6148 11940 6154 11942
rect 6210 11940 6234 11942
rect 6290 11940 6314 11942
rect 6370 11940 6394 11942
rect 6450 11940 6456 11942
rect 6148 11931 6456 11940
rect 5816 11892 5868 11898
rect 5816 11834 5868 11840
rect 6000 11892 6052 11898
rect 6000 11834 6052 11840
rect 5632 11688 5684 11694
rect 5630 11656 5632 11665
rect 5684 11656 5686 11665
rect 5630 11591 5686 11600
rect 5552 11478 5948 11506
rect 5632 11212 5684 11218
rect 5632 11154 5684 11160
rect 5724 11212 5776 11218
rect 5724 11154 5776 11160
rect 5540 10532 5592 10538
rect 5540 10474 5592 10480
rect 5552 9926 5580 10474
rect 5644 10130 5672 11154
rect 5736 10742 5764 11154
rect 5724 10736 5776 10742
rect 5724 10678 5776 10684
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 5816 10464 5868 10470
rect 5816 10406 5868 10412
rect 5632 10124 5684 10130
rect 5632 10066 5684 10072
rect 5736 9926 5764 10406
rect 5828 10266 5856 10406
rect 5816 10260 5868 10266
rect 5816 10202 5868 10208
rect 5816 10056 5868 10062
rect 5816 9998 5868 10004
rect 5540 9920 5592 9926
rect 5540 9862 5592 9868
rect 5724 9920 5776 9926
rect 5724 9862 5776 9868
rect 5736 9586 5764 9862
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 5736 9110 5764 9522
rect 5828 9382 5856 9998
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5724 9104 5776 9110
rect 5724 9046 5776 9052
rect 5538 8664 5594 8673
rect 5538 8599 5594 8608
rect 5446 8528 5502 8537
rect 5446 8463 5502 8472
rect 5552 8129 5580 8599
rect 5632 8424 5684 8430
rect 5632 8366 5684 8372
rect 5538 8120 5594 8129
rect 5538 8055 5594 8064
rect 5540 7948 5592 7954
rect 5540 7890 5592 7896
rect 5448 7744 5500 7750
rect 5448 7686 5500 7692
rect 5460 7478 5488 7686
rect 5448 7472 5500 7478
rect 5448 7414 5500 7420
rect 5448 7200 5500 7206
rect 5448 7142 5500 7148
rect 5460 4010 5488 7142
rect 5552 6769 5580 7890
rect 5644 6934 5672 8366
rect 5632 6928 5684 6934
rect 5632 6870 5684 6876
rect 5538 6760 5594 6769
rect 5538 6695 5594 6704
rect 5724 6656 5776 6662
rect 5724 6598 5776 6604
rect 5736 6458 5764 6598
rect 5724 6452 5776 6458
rect 5724 6394 5776 6400
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5552 5574 5580 6258
rect 5632 6112 5684 6118
rect 5828 6066 5856 9318
rect 5920 8401 5948 11478
rect 6184 11212 6236 11218
rect 6184 11154 6236 11160
rect 6196 11014 6224 11154
rect 6656 11121 6684 12038
rect 6736 11756 6788 11762
rect 6736 11698 6788 11704
rect 6748 11218 6776 11698
rect 6736 11212 6788 11218
rect 6736 11154 6788 11160
rect 6642 11112 6698 11121
rect 6642 11047 6698 11056
rect 6000 11008 6052 11014
rect 6000 10950 6052 10956
rect 6184 11008 6236 11014
rect 6184 10950 6236 10956
rect 6012 10266 6040 10950
rect 6148 10908 6456 10917
rect 6148 10906 6154 10908
rect 6210 10906 6234 10908
rect 6290 10906 6314 10908
rect 6370 10906 6394 10908
rect 6450 10906 6456 10908
rect 6210 10854 6212 10906
rect 6392 10854 6394 10906
rect 6148 10852 6154 10854
rect 6210 10852 6234 10854
rect 6290 10852 6314 10854
rect 6370 10852 6394 10854
rect 6450 10852 6456 10854
rect 6148 10843 6456 10852
rect 6000 10260 6052 10266
rect 6000 10202 6052 10208
rect 6828 9920 6880 9926
rect 6828 9862 6880 9868
rect 6148 9820 6456 9829
rect 6148 9818 6154 9820
rect 6210 9818 6234 9820
rect 6290 9818 6314 9820
rect 6370 9818 6394 9820
rect 6450 9818 6456 9820
rect 6210 9766 6212 9818
rect 6392 9766 6394 9818
rect 6148 9764 6154 9766
rect 6210 9764 6234 9766
rect 6290 9764 6314 9766
rect 6370 9764 6394 9766
rect 6450 9764 6456 9766
rect 6148 9755 6456 9764
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 6552 9512 6604 9518
rect 6552 9454 6604 9460
rect 6148 8732 6456 8741
rect 6148 8730 6154 8732
rect 6210 8730 6234 8732
rect 6290 8730 6314 8732
rect 6370 8730 6394 8732
rect 6450 8730 6456 8732
rect 6210 8678 6212 8730
rect 6392 8678 6394 8730
rect 6148 8676 6154 8678
rect 6210 8676 6234 8678
rect 6290 8676 6314 8678
rect 6370 8676 6394 8678
rect 6450 8676 6456 8678
rect 6148 8667 6456 8676
rect 6564 8514 6592 9454
rect 6748 9042 6776 9522
rect 6736 9036 6788 9042
rect 6736 8978 6788 8984
rect 6644 8832 6696 8838
rect 6644 8774 6696 8780
rect 6656 8634 6684 8774
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 6564 8486 6684 8514
rect 5906 8392 5962 8401
rect 5906 8327 5962 8336
rect 6552 8016 6604 8022
rect 6552 7958 6604 7964
rect 6148 7644 6456 7653
rect 6148 7642 6154 7644
rect 6210 7642 6234 7644
rect 6290 7642 6314 7644
rect 6370 7642 6394 7644
rect 6450 7642 6456 7644
rect 6210 7590 6212 7642
rect 6392 7590 6394 7642
rect 6148 7588 6154 7590
rect 6210 7588 6234 7590
rect 6290 7588 6314 7590
rect 6370 7588 6394 7590
rect 6450 7588 6456 7590
rect 6148 7579 6456 7588
rect 6564 7274 6592 7958
rect 6552 7268 6604 7274
rect 6552 7210 6604 7216
rect 5906 6896 5962 6905
rect 5906 6831 5962 6840
rect 6000 6860 6052 6866
rect 5920 6254 5948 6831
rect 6000 6802 6052 6808
rect 5908 6248 5960 6254
rect 5908 6190 5960 6196
rect 5632 6054 5684 6060
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 5552 5302 5580 5510
rect 5540 5296 5592 5302
rect 5540 5238 5592 5244
rect 5644 5166 5672 6054
rect 5736 6038 5856 6066
rect 5632 5160 5684 5166
rect 5632 5102 5684 5108
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 5644 4146 5672 4762
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 5448 4004 5500 4010
rect 5448 3946 5500 3952
rect 5644 3942 5672 4082
rect 5632 3936 5684 3942
rect 5632 3878 5684 3884
rect 5448 3664 5500 3670
rect 5448 3606 5500 3612
rect 5460 3058 5488 3606
rect 5644 3602 5672 3878
rect 5632 3596 5684 3602
rect 5632 3538 5684 3544
rect 5448 3052 5500 3058
rect 5448 2994 5500 3000
rect 5540 2304 5592 2310
rect 5540 2246 5592 2252
rect 5552 1698 5580 2246
rect 5540 1692 5592 1698
rect 5540 1634 5592 1640
rect 5736 800 5764 6038
rect 5908 5908 5960 5914
rect 5908 5850 5960 5856
rect 5920 5710 5948 5850
rect 6012 5778 6040 6802
rect 6148 6556 6456 6565
rect 6148 6554 6154 6556
rect 6210 6554 6234 6556
rect 6290 6554 6314 6556
rect 6370 6554 6394 6556
rect 6450 6554 6456 6556
rect 6210 6502 6212 6554
rect 6392 6502 6394 6554
rect 6148 6500 6154 6502
rect 6210 6500 6234 6502
rect 6290 6500 6314 6502
rect 6370 6500 6394 6502
rect 6450 6500 6456 6502
rect 6148 6491 6456 6500
rect 6564 6390 6592 7210
rect 6552 6384 6604 6390
rect 6288 6322 6500 6338
rect 6552 6326 6604 6332
rect 6276 6316 6512 6322
rect 6328 6310 6460 6316
rect 6276 6258 6328 6264
rect 6460 6258 6512 6264
rect 6550 6216 6606 6225
rect 6550 6151 6606 6160
rect 6000 5772 6052 5778
rect 6000 5714 6052 5720
rect 5908 5704 5960 5710
rect 5908 5646 5960 5652
rect 6148 5468 6456 5477
rect 6148 5466 6154 5468
rect 6210 5466 6234 5468
rect 6290 5466 6314 5468
rect 6370 5466 6394 5468
rect 6450 5466 6456 5468
rect 6210 5414 6212 5466
rect 6392 5414 6394 5466
rect 6148 5412 6154 5414
rect 6210 5412 6234 5414
rect 6290 5412 6314 5414
rect 6370 5412 6394 5414
rect 6450 5412 6456 5414
rect 6148 5403 6456 5412
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 5816 4480 5868 4486
rect 5816 4422 5868 4428
rect 5828 3738 5856 4422
rect 5920 4078 5948 5102
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 6380 4690 6408 4966
rect 6368 4684 6420 4690
rect 6368 4626 6420 4632
rect 6148 4380 6456 4389
rect 6148 4378 6154 4380
rect 6210 4378 6234 4380
rect 6290 4378 6314 4380
rect 6370 4378 6394 4380
rect 6450 4378 6456 4380
rect 6210 4326 6212 4378
rect 6392 4326 6394 4378
rect 6148 4324 6154 4326
rect 6210 4324 6234 4326
rect 6290 4324 6314 4326
rect 6370 4324 6394 4326
rect 6450 4324 6456 4326
rect 6148 4315 6456 4324
rect 6184 4276 6236 4282
rect 6184 4218 6236 4224
rect 5908 4072 5960 4078
rect 5908 4014 5960 4020
rect 5998 3904 6054 3913
rect 5998 3839 6054 3848
rect 5816 3732 5868 3738
rect 5816 3674 5868 3680
rect 5908 3732 5960 3738
rect 5908 3674 5960 3680
rect 5920 3194 5948 3674
rect 5908 3188 5960 3194
rect 5908 3130 5960 3136
rect 5814 2952 5870 2961
rect 5814 2887 5816 2896
rect 5868 2887 5870 2896
rect 5816 2858 5868 2864
rect 5816 2304 5868 2310
rect 5816 2246 5868 2252
rect 5828 1562 5856 2246
rect 5816 1556 5868 1562
rect 5816 1498 5868 1504
rect 6012 1306 6040 3839
rect 6196 3466 6224 4218
rect 6184 3460 6236 3466
rect 6184 3402 6236 3408
rect 6148 3292 6456 3301
rect 6148 3290 6154 3292
rect 6210 3290 6234 3292
rect 6290 3290 6314 3292
rect 6370 3290 6394 3292
rect 6450 3290 6456 3292
rect 6210 3238 6212 3290
rect 6392 3238 6394 3290
rect 6148 3236 6154 3238
rect 6210 3236 6234 3238
rect 6290 3236 6314 3238
rect 6370 3236 6394 3238
rect 6450 3236 6456 3238
rect 6148 3227 6456 3236
rect 6148 2204 6456 2213
rect 6148 2202 6154 2204
rect 6210 2202 6234 2204
rect 6290 2202 6314 2204
rect 6370 2202 6394 2204
rect 6450 2202 6456 2204
rect 6210 2150 6212 2202
rect 6392 2150 6394 2202
rect 6148 2148 6154 2150
rect 6210 2148 6234 2150
rect 6290 2148 6314 2150
rect 6370 2148 6394 2150
rect 6450 2148 6456 2150
rect 6148 2139 6456 2148
rect 6460 2100 6512 2106
rect 6460 2042 6512 2048
rect 6012 1278 6132 1306
rect 6104 800 6132 1278
rect 6472 800 6500 2042
rect 2516 734 2728 762
rect 2778 0 2834 800
rect 3146 0 3202 800
rect 3514 0 3570 800
rect 3882 0 3938 800
rect 4250 0 4306 800
rect 4618 0 4674 800
rect 4986 0 5042 800
rect 5354 0 5410 800
rect 5722 0 5778 800
rect 6090 0 6146 800
rect 6458 0 6514 800
rect 6564 762 6592 6151
rect 6656 6066 6684 8486
rect 6736 6656 6788 6662
rect 6736 6598 6788 6604
rect 6748 6458 6776 6598
rect 6736 6452 6788 6458
rect 6736 6394 6788 6400
rect 6840 6361 6868 9862
rect 7208 9450 7236 12838
rect 7668 12646 7696 12922
rect 7656 12640 7708 12646
rect 7656 12582 7708 12588
rect 7470 12336 7526 12345
rect 7470 12271 7472 12280
rect 7524 12271 7526 12280
rect 7472 12242 7524 12248
rect 7668 12170 7696 12582
rect 7656 12164 7708 12170
rect 7656 12106 7708 12112
rect 7380 12096 7432 12102
rect 7380 12038 7432 12044
rect 7392 11898 7420 12038
rect 7760 11898 7788 15438
rect 7840 14544 7892 14550
rect 7840 14486 7892 14492
rect 7852 12986 7880 14486
rect 8392 14408 8444 14414
rect 8392 14350 8444 14356
rect 8208 14340 8260 14346
rect 8208 14282 8260 14288
rect 8220 14074 8248 14282
rect 8208 14068 8260 14074
rect 8208 14010 8260 14016
rect 8300 13388 8352 13394
rect 8220 13348 8300 13376
rect 7932 13184 7984 13190
rect 7932 13126 7984 13132
rect 7840 12980 7892 12986
rect 7840 12922 7892 12928
rect 7944 12850 7972 13126
rect 7932 12844 7984 12850
rect 7932 12786 7984 12792
rect 7944 12434 7972 12786
rect 8024 12776 8076 12782
rect 8024 12718 8076 12724
rect 8036 12442 8064 12718
rect 8116 12640 8168 12646
rect 8116 12582 8168 12588
rect 7852 12406 7972 12434
rect 8024 12436 8076 12442
rect 7380 11892 7432 11898
rect 7380 11834 7432 11840
rect 7748 11892 7800 11898
rect 7748 11834 7800 11840
rect 7380 11552 7432 11558
rect 7380 11494 7432 11500
rect 7392 10470 7420 11494
rect 7746 11248 7802 11257
rect 7746 11183 7802 11192
rect 7472 11076 7524 11082
rect 7472 11018 7524 11024
rect 7484 10810 7512 11018
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 7484 10266 7512 10746
rect 7760 10305 7788 11183
rect 7746 10296 7802 10305
rect 7472 10260 7524 10266
rect 7746 10231 7802 10240
rect 7472 10202 7524 10208
rect 7760 10198 7788 10231
rect 7748 10192 7800 10198
rect 7748 10134 7800 10140
rect 7852 10062 7880 12406
rect 8024 12378 8076 12384
rect 8024 12300 8076 12306
rect 8024 12242 8076 12248
rect 7932 11552 7984 11558
rect 7932 11494 7984 11500
rect 7944 11286 7972 11494
rect 7932 11280 7984 11286
rect 7932 11222 7984 11228
rect 8036 10577 8064 12242
rect 8128 12238 8156 12582
rect 8220 12306 8248 13348
rect 8300 13330 8352 13336
rect 8404 12434 8432 14350
rect 8484 14272 8536 14278
rect 8484 14214 8536 14220
rect 8496 13734 8524 14214
rect 8484 13728 8536 13734
rect 8484 13670 8536 13676
rect 8588 12442 8616 16526
rect 9140 16454 9168 19314
rect 9404 17672 9456 17678
rect 9404 17614 9456 17620
rect 9128 16448 9180 16454
rect 9128 16390 9180 16396
rect 8747 15804 9055 15813
rect 8747 15802 8753 15804
rect 8809 15802 8833 15804
rect 8889 15802 8913 15804
rect 8969 15802 8993 15804
rect 9049 15802 9055 15804
rect 8809 15750 8811 15802
rect 8991 15750 8993 15802
rect 8747 15748 8753 15750
rect 8809 15748 8833 15750
rect 8889 15748 8913 15750
rect 8969 15748 8993 15750
rect 9049 15748 9055 15750
rect 8747 15739 9055 15748
rect 9312 15360 9364 15366
rect 9312 15302 9364 15308
rect 8747 14716 9055 14725
rect 8747 14714 8753 14716
rect 8809 14714 8833 14716
rect 8889 14714 8913 14716
rect 8969 14714 8993 14716
rect 9049 14714 9055 14716
rect 8809 14662 8811 14714
rect 8991 14662 8993 14714
rect 8747 14660 8753 14662
rect 8809 14660 8833 14662
rect 8889 14660 8913 14662
rect 8969 14660 8993 14662
rect 9049 14660 9055 14662
rect 8747 14651 9055 14660
rect 9324 14618 9352 15302
rect 9312 14612 9364 14618
rect 9312 14554 9364 14560
rect 9416 14074 9444 17614
rect 10324 14408 10376 14414
rect 10324 14350 10376 14356
rect 9680 14272 9732 14278
rect 9680 14214 9732 14220
rect 9404 14068 9456 14074
rect 9404 14010 9456 14016
rect 9036 13864 9088 13870
rect 9034 13832 9036 13841
rect 9088 13832 9090 13841
rect 9034 13767 9090 13776
rect 8747 13628 9055 13637
rect 8747 13626 8753 13628
rect 8809 13626 8833 13628
rect 8889 13626 8913 13628
rect 8969 13626 8993 13628
rect 9049 13626 9055 13628
rect 8809 13574 8811 13626
rect 8991 13574 8993 13626
rect 8747 13572 8753 13574
rect 8809 13572 8833 13574
rect 8889 13572 8913 13574
rect 8969 13572 8993 13574
rect 9049 13572 9055 13574
rect 8747 13563 9055 13572
rect 9692 12986 9720 14214
rect 9772 13932 9824 13938
rect 9772 13874 9824 13880
rect 9784 13394 9812 13874
rect 9956 13796 10008 13802
rect 9956 13738 10008 13744
rect 10140 13796 10192 13802
rect 10140 13738 10192 13744
rect 9772 13388 9824 13394
rect 9772 13330 9824 13336
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 9128 12844 9180 12850
rect 9128 12786 9180 12792
rect 9140 12646 9168 12786
rect 9128 12640 9180 12646
rect 9128 12582 9180 12588
rect 8747 12540 9055 12549
rect 8747 12538 8753 12540
rect 8809 12538 8833 12540
rect 8889 12538 8913 12540
rect 8969 12538 8993 12540
rect 9049 12538 9055 12540
rect 8809 12486 8811 12538
rect 8991 12486 8993 12538
rect 8747 12484 8753 12486
rect 8809 12484 8833 12486
rect 8889 12484 8913 12486
rect 8969 12484 8993 12486
rect 9049 12484 9055 12486
rect 8747 12475 9055 12484
rect 8576 12436 8628 12442
rect 8404 12406 8524 12434
rect 8300 12368 8352 12374
rect 8300 12310 8352 12316
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 8116 12232 8168 12238
rect 8116 12174 8168 12180
rect 8022 10568 8078 10577
rect 8022 10503 8078 10512
rect 7932 10464 7984 10470
rect 7932 10406 7984 10412
rect 7840 10056 7892 10062
rect 7840 9998 7892 10004
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 7852 9654 7880 9862
rect 7840 9648 7892 9654
rect 7840 9590 7892 9596
rect 7196 9444 7248 9450
rect 7196 9386 7248 9392
rect 7654 9072 7710 9081
rect 7654 9007 7710 9016
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 7012 8900 7064 8906
rect 7012 8842 7064 8848
rect 7024 7426 7052 8842
rect 7380 8832 7432 8838
rect 7380 8774 7432 8780
rect 7196 8356 7248 8362
rect 7196 8298 7248 8304
rect 7102 8256 7158 8265
rect 7102 8191 7158 8200
rect 7116 7546 7144 8191
rect 7104 7540 7156 7546
rect 7104 7482 7156 7488
rect 7024 7398 7144 7426
rect 6920 7336 6972 7342
rect 6920 7278 6972 7284
rect 6826 6352 6882 6361
rect 6826 6287 6882 6296
rect 6656 6038 6868 6066
rect 6644 5568 6696 5574
rect 6644 5510 6696 5516
rect 6656 5302 6684 5510
rect 6644 5296 6696 5302
rect 6644 5238 6696 5244
rect 6736 5092 6788 5098
rect 6736 5034 6788 5040
rect 6644 4072 6696 4078
rect 6644 4014 6696 4020
rect 6656 2650 6684 4014
rect 6748 3602 6776 5034
rect 6840 4570 6868 6038
rect 6932 5846 6960 7278
rect 7012 6112 7064 6118
rect 7012 6054 7064 6060
rect 6920 5840 6972 5846
rect 6920 5782 6972 5788
rect 6932 5574 6960 5782
rect 6920 5568 6972 5574
rect 6920 5510 6972 5516
rect 7024 5370 7052 6054
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 7024 5001 7052 5170
rect 7010 4992 7066 5001
rect 7010 4927 7066 4936
rect 7116 4690 7144 7398
rect 7104 4684 7156 4690
rect 7104 4626 7156 4632
rect 7012 4616 7064 4622
rect 6840 4542 6960 4570
rect 7064 4564 7144 4570
rect 7012 4558 7144 4564
rect 7024 4542 7144 4558
rect 6828 4480 6880 4486
rect 6828 4422 6880 4428
rect 6840 4146 6868 4422
rect 6932 4214 6960 4542
rect 7012 4480 7064 4486
rect 7012 4422 7064 4428
rect 6920 4208 6972 4214
rect 6920 4150 6972 4156
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 6920 3392 6972 3398
rect 6920 3334 6972 3340
rect 6932 3194 6960 3334
rect 7024 3194 7052 4422
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 7116 2990 7144 4542
rect 6920 2984 6972 2990
rect 6920 2926 6972 2932
rect 7104 2984 7156 2990
rect 7104 2926 7156 2932
rect 6644 2644 6696 2650
rect 6644 2586 6696 2592
rect 6736 2576 6788 2582
rect 6932 2553 6960 2926
rect 6736 2518 6788 2524
rect 6918 2544 6974 2553
rect 6748 1766 6776 2518
rect 6918 2479 6974 2488
rect 7208 2446 7236 8298
rect 7392 7546 7420 8774
rect 7380 7540 7432 7546
rect 7380 7482 7432 7488
rect 7484 6882 7512 8910
rect 7668 8430 7696 9007
rect 7564 8424 7616 8430
rect 7564 8366 7616 8372
rect 7656 8424 7708 8430
rect 7656 8366 7708 8372
rect 7576 8090 7604 8366
rect 7748 8356 7800 8362
rect 7748 8298 7800 8304
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 7484 6854 7696 6882
rect 7472 6724 7524 6730
rect 7472 6666 7524 6672
rect 7288 6248 7340 6254
rect 7288 6190 7340 6196
rect 7300 5710 7328 6190
rect 7288 5704 7340 5710
rect 7288 5646 7340 5652
rect 7380 5160 7432 5166
rect 7380 5102 7432 5108
rect 7286 4720 7342 4729
rect 7286 4655 7288 4664
rect 7340 4655 7342 4664
rect 7288 4626 7340 4632
rect 7288 4548 7340 4554
rect 7288 4490 7340 4496
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 7300 2106 7328 4490
rect 7392 2922 7420 5102
rect 7484 3670 7512 6666
rect 7668 5710 7696 6854
rect 7760 6798 7788 8298
rect 7838 7984 7894 7993
rect 7838 7919 7840 7928
rect 7892 7919 7894 7928
rect 7840 7890 7892 7896
rect 7838 7576 7894 7585
rect 7838 7511 7894 7520
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 7656 5704 7708 5710
rect 7656 5646 7708 5652
rect 7472 3664 7524 3670
rect 7472 3606 7524 3612
rect 7470 3496 7526 3505
rect 7576 3466 7604 5646
rect 7668 5370 7696 5646
rect 7656 5364 7708 5370
rect 7656 5306 7708 5312
rect 7656 3664 7708 3670
rect 7656 3606 7708 3612
rect 7470 3431 7472 3440
rect 7524 3431 7526 3440
rect 7564 3460 7616 3466
rect 7472 3402 7524 3408
rect 7564 3402 7616 3408
rect 7380 2916 7432 2922
rect 7380 2858 7432 2864
rect 7668 2774 7696 3606
rect 7748 3596 7800 3602
rect 7748 3538 7800 3544
rect 7760 3369 7788 3538
rect 7746 3360 7802 3369
rect 7746 3295 7802 3304
rect 7484 2746 7696 2774
rect 7852 2774 7880 7511
rect 7944 3194 7972 10406
rect 8024 10192 8076 10198
rect 8022 10160 8024 10169
rect 8076 10160 8078 10169
rect 8022 10095 8078 10104
rect 8024 7744 8076 7750
rect 8024 7686 8076 7692
rect 8036 4282 8064 7686
rect 8024 4276 8076 4282
rect 8024 4218 8076 4224
rect 8024 4072 8076 4078
rect 8024 4014 8076 4020
rect 7932 3188 7984 3194
rect 7932 3130 7984 3136
rect 8036 3058 8064 4014
rect 8024 3052 8076 3058
rect 8024 2994 8076 3000
rect 7852 2746 7972 2774
rect 7288 2100 7340 2106
rect 7288 2042 7340 2048
rect 6736 1760 6788 1766
rect 6736 1702 6788 1708
rect 6748 870 6868 898
rect 6748 762 6776 870
rect 6840 800 6868 870
rect 7208 870 7328 898
rect 7208 800 7236 870
rect 6564 734 6776 762
rect 6826 0 6882 800
rect 7194 0 7250 800
rect 7300 762 7328 870
rect 7484 762 7512 2746
rect 7564 1420 7616 1426
rect 7564 1362 7616 1368
rect 7576 800 7604 1362
rect 7944 800 7972 2746
rect 8128 1426 8156 12174
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 8220 11354 8248 12038
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 8208 10736 8260 10742
rect 8208 10678 8260 10684
rect 8220 7818 8248 10678
rect 8312 10266 8340 12310
rect 8392 11824 8444 11830
rect 8392 11766 8444 11772
rect 8404 11354 8432 11766
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 8390 11248 8446 11257
rect 8390 11183 8392 11192
rect 8444 11183 8446 11192
rect 8392 11154 8444 11160
rect 8392 11076 8444 11082
rect 8392 11018 8444 11024
rect 8404 10538 8432 11018
rect 8392 10532 8444 10538
rect 8392 10474 8444 10480
rect 8300 10260 8352 10266
rect 8300 10202 8352 10208
rect 8298 10024 8354 10033
rect 8298 9959 8354 9968
rect 8312 8906 8340 9959
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 8300 8900 8352 8906
rect 8300 8842 8352 8848
rect 8298 8120 8354 8129
rect 8404 8090 8432 9318
rect 8298 8055 8354 8064
rect 8392 8084 8444 8090
rect 8208 7812 8260 7818
rect 8208 7754 8260 7760
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 8220 2514 8248 7278
rect 8312 5930 8340 8055
rect 8392 8026 8444 8032
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 8404 6458 8432 6938
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 8312 5902 8432 5930
rect 8300 5772 8352 5778
rect 8300 5714 8352 5720
rect 8312 4185 8340 5714
rect 8404 4690 8432 5902
rect 8392 4684 8444 4690
rect 8392 4626 8444 4632
rect 8298 4176 8354 4185
rect 8298 4111 8354 4120
rect 8390 3496 8446 3505
rect 8300 3460 8352 3466
rect 8390 3431 8446 3440
rect 8300 3402 8352 3408
rect 8312 2582 8340 3402
rect 8300 2576 8352 2582
rect 8300 2518 8352 2524
rect 8208 2508 8260 2514
rect 8208 2450 8260 2456
rect 8208 2372 8260 2378
rect 8208 2314 8260 2320
rect 8220 1970 8248 2314
rect 8208 1964 8260 1970
rect 8208 1906 8260 1912
rect 8116 1420 8168 1426
rect 8116 1362 8168 1368
rect 8404 1034 8432 3431
rect 8496 2774 8524 12406
rect 8576 12378 8628 12384
rect 8576 12300 8628 12306
rect 8576 12242 8628 12248
rect 8588 10742 8616 12242
rect 9140 11762 9168 12582
rect 9968 12442 9996 13738
rect 10152 13433 10180 13738
rect 10138 13424 10194 13433
rect 10138 13359 10194 13368
rect 10232 12776 10284 12782
rect 10232 12718 10284 12724
rect 9956 12436 10008 12442
rect 9956 12378 10008 12384
rect 9588 12300 9640 12306
rect 9588 12242 9640 12248
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 9128 11756 9180 11762
rect 9128 11698 9180 11704
rect 8680 11218 8708 11698
rect 9140 11558 9168 11698
rect 9312 11688 9364 11694
rect 9312 11630 9364 11636
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 8747 11452 9055 11461
rect 8747 11450 8753 11452
rect 8809 11450 8833 11452
rect 8889 11450 8913 11452
rect 8969 11450 8993 11452
rect 9049 11450 9055 11452
rect 8809 11398 8811 11450
rect 8991 11398 8993 11450
rect 8747 11396 8753 11398
rect 8809 11396 8833 11398
rect 8889 11396 8913 11398
rect 8969 11396 8993 11398
rect 9049 11396 9055 11398
rect 8747 11387 9055 11396
rect 8668 11212 8720 11218
rect 8668 11154 8720 11160
rect 9324 11082 9352 11630
rect 9312 11076 9364 11082
rect 9312 11018 9364 11024
rect 8576 10736 8628 10742
rect 8576 10678 8628 10684
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 8956 10452 8984 10610
rect 8680 10424 8984 10452
rect 8576 8424 8628 8430
rect 8576 8366 8628 8372
rect 8588 7886 8616 8366
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 8576 7404 8628 7410
rect 8576 7346 8628 7352
rect 8588 7002 8616 7346
rect 8576 6996 8628 7002
rect 8576 6938 8628 6944
rect 8680 6254 8708 10424
rect 8747 10364 9055 10373
rect 8747 10362 8753 10364
rect 8809 10362 8833 10364
rect 8889 10362 8913 10364
rect 8969 10362 8993 10364
rect 9049 10362 9055 10364
rect 8809 10310 8811 10362
rect 8991 10310 8993 10362
rect 8747 10308 8753 10310
rect 8809 10308 8833 10310
rect 8889 10308 8913 10310
rect 8969 10308 8993 10310
rect 9049 10308 9055 10310
rect 8747 10299 9055 10308
rect 9128 9920 9180 9926
rect 9128 9862 9180 9868
rect 8747 9276 9055 9285
rect 8747 9274 8753 9276
rect 8809 9274 8833 9276
rect 8889 9274 8913 9276
rect 8969 9274 8993 9276
rect 9049 9274 9055 9276
rect 8809 9222 8811 9274
rect 8991 9222 8993 9274
rect 8747 9220 8753 9222
rect 8809 9220 8833 9222
rect 8889 9220 8913 9222
rect 8969 9220 8993 9222
rect 9049 9220 9055 9222
rect 8747 9211 9055 9220
rect 9140 8974 9168 9862
rect 9220 9376 9272 9382
rect 9220 9318 9272 9324
rect 9128 8968 9180 8974
rect 9128 8910 9180 8916
rect 8747 8188 9055 8197
rect 8747 8186 8753 8188
rect 8809 8186 8833 8188
rect 8889 8186 8913 8188
rect 8969 8186 8993 8188
rect 9049 8186 9055 8188
rect 8809 8134 8811 8186
rect 8991 8134 8993 8186
rect 8747 8132 8753 8134
rect 8809 8132 8833 8134
rect 8889 8132 8913 8134
rect 8969 8132 8993 8134
rect 9049 8132 9055 8134
rect 8747 8123 9055 8132
rect 8747 7100 9055 7109
rect 8747 7098 8753 7100
rect 8809 7098 8833 7100
rect 8889 7098 8913 7100
rect 8969 7098 8993 7100
rect 9049 7098 9055 7100
rect 8809 7046 8811 7098
rect 8991 7046 8993 7098
rect 8747 7044 8753 7046
rect 8809 7044 8833 7046
rect 8889 7044 8913 7046
rect 8969 7044 8993 7046
rect 9049 7044 9055 7046
rect 8747 7035 9055 7044
rect 9128 6860 9180 6866
rect 9128 6802 9180 6808
rect 9036 6656 9088 6662
rect 9036 6598 9088 6604
rect 9048 6458 9076 6598
rect 9140 6458 9168 6802
rect 9036 6452 9088 6458
rect 9036 6394 9088 6400
rect 9128 6452 9180 6458
rect 9128 6394 9180 6400
rect 8668 6248 8720 6254
rect 8668 6190 8720 6196
rect 8680 6118 8708 6190
rect 8668 6112 8720 6118
rect 8668 6054 8720 6060
rect 8747 6012 9055 6021
rect 8747 6010 8753 6012
rect 8809 6010 8833 6012
rect 8889 6010 8913 6012
rect 8969 6010 8993 6012
rect 9049 6010 9055 6012
rect 8809 5958 8811 6010
rect 8991 5958 8993 6010
rect 8747 5956 8753 5958
rect 8809 5956 8833 5958
rect 8889 5956 8913 5958
rect 8969 5956 8993 5958
rect 9049 5956 9055 5958
rect 8747 5947 9055 5956
rect 8666 5672 8722 5681
rect 8666 5607 8722 5616
rect 8576 5568 8628 5574
rect 8576 5510 8628 5516
rect 8588 5370 8616 5510
rect 8576 5364 8628 5370
rect 8576 5306 8628 5312
rect 8576 5024 8628 5030
rect 8576 4966 8628 4972
rect 8588 3534 8616 4966
rect 8576 3528 8628 3534
rect 8576 3470 8628 3476
rect 8680 3398 8708 5607
rect 8944 5568 8996 5574
rect 8944 5510 8996 5516
rect 8956 5234 8984 5510
rect 8944 5228 8996 5234
rect 8944 5170 8996 5176
rect 9128 5024 9180 5030
rect 9128 4966 9180 4972
rect 8747 4924 9055 4933
rect 8747 4922 8753 4924
rect 8809 4922 8833 4924
rect 8889 4922 8913 4924
rect 8969 4922 8993 4924
rect 9049 4922 9055 4924
rect 8809 4870 8811 4922
rect 8991 4870 8993 4922
rect 8747 4868 8753 4870
rect 8809 4868 8833 4870
rect 8889 4868 8913 4870
rect 8969 4868 8993 4870
rect 9049 4868 9055 4870
rect 8747 4859 9055 4868
rect 9140 4622 9168 4966
rect 9128 4616 9180 4622
rect 9128 4558 9180 4564
rect 9128 4480 9180 4486
rect 9128 4422 9180 4428
rect 9140 4282 9168 4422
rect 9128 4276 9180 4282
rect 9128 4218 9180 4224
rect 9128 4004 9180 4010
rect 9128 3946 9180 3952
rect 8747 3836 9055 3845
rect 8747 3834 8753 3836
rect 8809 3834 8833 3836
rect 8889 3834 8913 3836
rect 8969 3834 8993 3836
rect 9049 3834 9055 3836
rect 8809 3782 8811 3834
rect 8991 3782 8993 3834
rect 8747 3780 8753 3782
rect 8809 3780 8833 3782
rect 8889 3780 8913 3782
rect 8969 3780 8993 3782
rect 9049 3780 9055 3782
rect 8747 3771 9055 3780
rect 9140 3738 9168 3946
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 9126 3632 9182 3641
rect 9126 3567 9182 3576
rect 8668 3392 8720 3398
rect 8668 3334 8720 3340
rect 8758 3224 8814 3233
rect 8758 3159 8814 3168
rect 9036 3188 9088 3194
rect 8772 3058 8800 3159
rect 9036 3130 9088 3136
rect 9048 3058 9076 3130
rect 8760 3052 8812 3058
rect 8760 2994 8812 3000
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 8496 2746 8708 2774
rect 8312 1006 8432 1034
rect 8312 800 8340 1006
rect 8680 800 8708 2746
rect 8747 2748 9055 2757
rect 8747 2746 8753 2748
rect 8809 2746 8833 2748
rect 8889 2746 8913 2748
rect 8969 2746 8993 2748
rect 9049 2746 9055 2748
rect 8809 2694 8811 2746
rect 8991 2694 8993 2746
rect 8747 2692 8753 2694
rect 8809 2692 8833 2694
rect 8889 2692 8913 2694
rect 8969 2692 8993 2694
rect 9049 2692 9055 2694
rect 8747 2683 9055 2692
rect 9036 2508 9088 2514
rect 9036 2450 9088 2456
rect 9048 2378 9076 2450
rect 9036 2372 9088 2378
rect 9036 2314 9088 2320
rect 9048 2281 9076 2314
rect 9034 2272 9090 2281
rect 9034 2207 9090 2216
rect 9048 1630 9076 2207
rect 9036 1624 9088 1630
rect 9036 1566 9088 1572
rect 9140 1034 9168 3567
rect 9232 3233 9260 9318
rect 9324 7585 9352 11018
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 9404 9920 9456 9926
rect 9404 9862 9456 9868
rect 9416 8673 9444 9862
rect 9508 8922 9536 10066
rect 9600 10033 9628 12242
rect 10048 12232 10100 12238
rect 10048 12174 10100 12180
rect 10140 12232 10192 12238
rect 10140 12174 10192 12180
rect 9956 11620 10008 11626
rect 9956 11562 10008 11568
rect 9968 10538 9996 11562
rect 10060 11150 10088 12174
rect 10048 11144 10100 11150
rect 10048 11086 10100 11092
rect 10060 10810 10088 11086
rect 10152 11082 10180 12174
rect 10140 11076 10192 11082
rect 10140 11018 10192 11024
rect 10048 10804 10100 10810
rect 10048 10746 10100 10752
rect 9864 10532 9916 10538
rect 9864 10474 9916 10480
rect 9956 10532 10008 10538
rect 9956 10474 10008 10480
rect 9680 10124 9732 10130
rect 9680 10066 9732 10072
rect 9586 10024 9642 10033
rect 9586 9959 9642 9968
rect 9692 9722 9720 10066
rect 9680 9716 9732 9722
rect 9680 9658 9732 9664
rect 9508 8894 9628 8922
rect 9496 8832 9548 8838
rect 9496 8774 9548 8780
rect 9402 8664 9458 8673
rect 9508 8634 9536 8774
rect 9402 8599 9458 8608
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9404 8288 9456 8294
rect 9404 8230 9456 8236
rect 9310 7576 9366 7585
rect 9310 7511 9366 7520
rect 9312 6248 9364 6254
rect 9312 6190 9364 6196
rect 9324 5710 9352 6190
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 9416 5030 9444 8230
rect 9600 7274 9628 8894
rect 9588 7268 9640 7274
rect 9588 7210 9640 7216
rect 9588 6860 9640 6866
rect 9588 6802 9640 6808
rect 9600 5914 9628 6802
rect 9588 5908 9640 5914
rect 9588 5850 9640 5856
rect 9588 5772 9640 5778
rect 9588 5714 9640 5720
rect 9600 5302 9628 5714
rect 9588 5296 9640 5302
rect 9588 5238 9640 5244
rect 9404 5024 9456 5030
rect 9404 4966 9456 4972
rect 9312 4548 9364 4554
rect 9364 4508 9536 4536
rect 9312 4490 9364 4496
rect 9218 3224 9274 3233
rect 9218 3159 9274 3168
rect 9508 2582 9536 4508
rect 9588 4072 9640 4078
rect 9588 4014 9640 4020
rect 9600 3738 9628 4014
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 9586 3632 9642 3641
rect 9692 3602 9720 9658
rect 9876 9654 9904 10474
rect 9864 9648 9916 9654
rect 9864 9590 9916 9596
rect 9772 9036 9824 9042
rect 9772 8978 9824 8984
rect 9784 8838 9812 8978
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 9586 3567 9642 3576
rect 9680 3596 9732 3602
rect 9600 3398 9628 3567
rect 9680 3538 9732 3544
rect 9680 3460 9732 3466
rect 9680 3402 9732 3408
rect 9588 3392 9640 3398
rect 9588 3334 9640 3340
rect 9588 2984 9640 2990
rect 9588 2926 9640 2932
rect 9600 2666 9628 2926
rect 9692 2854 9720 3402
rect 9784 3058 9812 8774
rect 9864 8424 9916 8430
rect 9864 8366 9916 8372
rect 9876 8090 9904 8366
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9876 3194 9904 7142
rect 10048 6316 10100 6322
rect 10048 6258 10100 6264
rect 9956 5568 10008 5574
rect 9956 5510 10008 5516
rect 9968 4214 9996 5510
rect 10060 5098 10088 6258
rect 10048 5092 10100 5098
rect 10048 5034 10100 5040
rect 9956 4208 10008 4214
rect 9956 4150 10008 4156
rect 10048 4140 10100 4146
rect 10048 4082 10100 4088
rect 10060 3942 10088 4082
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 9956 3664 10008 3670
rect 9956 3606 10008 3612
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 9772 3052 9824 3058
rect 9772 2994 9824 3000
rect 9680 2848 9732 2854
rect 9968 2825 9996 3606
rect 9680 2790 9732 2796
rect 9954 2816 10010 2825
rect 9954 2751 10010 2760
rect 9678 2680 9734 2689
rect 9600 2638 9678 2666
rect 9678 2615 9734 2624
rect 9496 2576 9548 2582
rect 9496 2518 9548 2524
rect 9956 2576 10008 2582
rect 9956 2518 10008 2524
rect 9220 2304 9272 2310
rect 9218 2272 9220 2281
rect 9496 2304 9548 2310
rect 9272 2272 9274 2281
rect 9218 2207 9274 2216
rect 9494 2272 9496 2281
rect 9548 2272 9550 2281
rect 9494 2207 9550 2216
rect 9402 2136 9458 2145
rect 9968 2106 9996 2518
rect 9402 2071 9458 2080
rect 9956 2100 10008 2106
rect 9048 1006 9168 1034
rect 9048 800 9076 1006
rect 9416 800 9444 2071
rect 9956 2042 10008 2048
rect 9772 944 9824 950
rect 9772 886 9824 892
rect 9784 800 9812 886
rect 10152 800 10180 11018
rect 10244 4486 10272 12718
rect 10336 8974 10364 14350
rect 10428 14074 10456 19790
rect 11346 19612 11654 19621
rect 11346 19610 11352 19612
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11648 19610 11654 19612
rect 11408 19558 11410 19610
rect 11590 19558 11592 19610
rect 11346 19556 11352 19558
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11648 19556 11654 19558
rect 11346 19547 11654 19556
rect 16544 19612 16852 19621
rect 16544 19610 16550 19612
rect 16606 19610 16630 19612
rect 16686 19610 16710 19612
rect 16766 19610 16790 19612
rect 16846 19610 16852 19612
rect 16606 19558 16608 19610
rect 16788 19558 16790 19610
rect 16544 19556 16550 19558
rect 16606 19556 16630 19558
rect 16686 19556 16710 19558
rect 16766 19556 16790 19558
rect 16846 19556 16852 19558
rect 16544 19547 16852 19556
rect 21742 19612 22050 19621
rect 21742 19610 21748 19612
rect 21804 19610 21828 19612
rect 21884 19610 21908 19612
rect 21964 19610 21988 19612
rect 22044 19610 22050 19612
rect 21804 19558 21806 19610
rect 21986 19558 21988 19610
rect 21742 19556 21748 19558
rect 21804 19556 21828 19558
rect 21884 19556 21908 19558
rect 21964 19556 21988 19558
rect 22044 19556 22050 19558
rect 21742 19547 22050 19556
rect 13945 19068 14253 19077
rect 13945 19066 13951 19068
rect 14007 19066 14031 19068
rect 14087 19066 14111 19068
rect 14167 19066 14191 19068
rect 14247 19066 14253 19068
rect 14007 19014 14009 19066
rect 14189 19014 14191 19066
rect 13945 19012 13951 19014
rect 14007 19012 14031 19014
rect 14087 19012 14111 19014
rect 14167 19012 14191 19014
rect 14247 19012 14253 19014
rect 13945 19003 14253 19012
rect 19143 19068 19451 19077
rect 19143 19066 19149 19068
rect 19205 19066 19229 19068
rect 19285 19066 19309 19068
rect 19365 19066 19389 19068
rect 19445 19066 19451 19068
rect 19205 19014 19207 19066
rect 19387 19014 19389 19066
rect 19143 19012 19149 19014
rect 19205 19012 19229 19014
rect 19285 19012 19309 19014
rect 19365 19012 19389 19014
rect 19445 19012 19451 19014
rect 19143 19003 19451 19012
rect 11346 18524 11654 18533
rect 11346 18522 11352 18524
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11648 18522 11654 18524
rect 11408 18470 11410 18522
rect 11590 18470 11592 18522
rect 11346 18468 11352 18470
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11648 18468 11654 18470
rect 11346 18459 11654 18468
rect 16544 18524 16852 18533
rect 16544 18522 16550 18524
rect 16606 18522 16630 18524
rect 16686 18522 16710 18524
rect 16766 18522 16790 18524
rect 16846 18522 16852 18524
rect 16606 18470 16608 18522
rect 16788 18470 16790 18522
rect 16544 18468 16550 18470
rect 16606 18468 16630 18470
rect 16686 18468 16710 18470
rect 16766 18468 16790 18470
rect 16846 18468 16852 18470
rect 16544 18459 16852 18468
rect 21742 18524 22050 18533
rect 21742 18522 21748 18524
rect 21804 18522 21828 18524
rect 21884 18522 21908 18524
rect 21964 18522 21988 18524
rect 22044 18522 22050 18524
rect 21804 18470 21806 18522
rect 21986 18470 21988 18522
rect 21742 18468 21748 18470
rect 21804 18468 21828 18470
rect 21884 18468 21908 18470
rect 21964 18468 21988 18470
rect 22044 18468 22050 18470
rect 21742 18459 22050 18468
rect 13945 17980 14253 17989
rect 13945 17978 13951 17980
rect 14007 17978 14031 17980
rect 14087 17978 14111 17980
rect 14167 17978 14191 17980
rect 14247 17978 14253 17980
rect 14007 17926 14009 17978
rect 14189 17926 14191 17978
rect 13945 17924 13951 17926
rect 14007 17924 14031 17926
rect 14087 17924 14111 17926
rect 14167 17924 14191 17926
rect 14247 17924 14253 17926
rect 13945 17915 14253 17924
rect 19143 17980 19451 17989
rect 19143 17978 19149 17980
rect 19205 17978 19229 17980
rect 19285 17978 19309 17980
rect 19365 17978 19389 17980
rect 19445 17978 19451 17980
rect 19205 17926 19207 17978
rect 19387 17926 19389 17978
rect 19143 17924 19149 17926
rect 19205 17924 19229 17926
rect 19285 17924 19309 17926
rect 19365 17924 19389 17926
rect 19445 17924 19451 17926
rect 19143 17915 19451 17924
rect 11346 17436 11654 17445
rect 11346 17434 11352 17436
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11648 17434 11654 17436
rect 11408 17382 11410 17434
rect 11590 17382 11592 17434
rect 11346 17380 11352 17382
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11648 17380 11654 17382
rect 11346 17371 11654 17380
rect 16544 17436 16852 17445
rect 16544 17434 16550 17436
rect 16606 17434 16630 17436
rect 16686 17434 16710 17436
rect 16766 17434 16790 17436
rect 16846 17434 16852 17436
rect 16606 17382 16608 17434
rect 16788 17382 16790 17434
rect 16544 17380 16550 17382
rect 16606 17380 16630 17382
rect 16686 17380 16710 17382
rect 16766 17380 16790 17382
rect 16846 17380 16852 17382
rect 16544 17371 16852 17380
rect 21742 17436 22050 17445
rect 21742 17434 21748 17436
rect 21804 17434 21828 17436
rect 21884 17434 21908 17436
rect 21964 17434 21988 17436
rect 22044 17434 22050 17436
rect 21804 17382 21806 17434
rect 21986 17382 21988 17434
rect 21742 17380 21748 17382
rect 21804 17380 21828 17382
rect 21884 17380 21908 17382
rect 21964 17380 21988 17382
rect 22044 17380 22050 17382
rect 21742 17371 22050 17380
rect 21454 17232 21510 17241
rect 12164 17196 12216 17202
rect 21454 17167 21510 17176
rect 12164 17138 12216 17144
rect 10876 16720 10928 16726
rect 10876 16662 10928 16668
rect 10600 14476 10652 14482
rect 10600 14418 10652 14424
rect 10416 14068 10468 14074
rect 10416 14010 10468 14016
rect 10508 13252 10560 13258
rect 10508 13194 10560 13200
rect 10416 12300 10468 12306
rect 10416 12242 10468 12248
rect 10428 12102 10456 12242
rect 10416 12096 10468 12102
rect 10416 12038 10468 12044
rect 10324 8968 10376 8974
rect 10324 8910 10376 8916
rect 10324 6656 10376 6662
rect 10324 6598 10376 6604
rect 10336 6390 10364 6598
rect 10324 6384 10376 6390
rect 10324 6326 10376 6332
rect 10232 4480 10284 4486
rect 10232 4422 10284 4428
rect 10414 4040 10470 4049
rect 10414 3975 10470 3984
rect 10428 3534 10456 3975
rect 10416 3528 10468 3534
rect 10416 3470 10468 3476
rect 10324 2644 10376 2650
rect 10324 2586 10376 2592
rect 10336 2446 10364 2586
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 10520 800 10548 13194
rect 10612 11257 10640 14418
rect 10784 14272 10836 14278
rect 10784 14214 10836 14220
rect 10796 14074 10824 14214
rect 10784 14068 10836 14074
rect 10784 14010 10836 14016
rect 10888 13530 10916 16662
rect 11346 16348 11654 16357
rect 11346 16346 11352 16348
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11648 16346 11654 16348
rect 11408 16294 11410 16346
rect 11590 16294 11592 16346
rect 11346 16292 11352 16294
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11648 16292 11654 16294
rect 11346 16283 11654 16292
rect 11796 15564 11848 15570
rect 11796 15506 11848 15512
rect 11346 15260 11654 15269
rect 11346 15258 11352 15260
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11648 15258 11654 15260
rect 11408 15206 11410 15258
rect 11590 15206 11592 15258
rect 11346 15204 11352 15206
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11648 15204 11654 15206
rect 11346 15195 11654 15204
rect 11152 14408 11204 14414
rect 11152 14350 11204 14356
rect 10876 13524 10928 13530
rect 10876 13466 10928 13472
rect 10876 13388 10928 13394
rect 10876 13330 10928 13336
rect 10692 13320 10744 13326
rect 10692 13262 10744 13268
rect 10704 13190 10732 13262
rect 10692 13184 10744 13190
rect 10692 13126 10744 13132
rect 10598 11248 10654 11257
rect 10598 11183 10654 11192
rect 10612 11082 10640 11183
rect 10600 11076 10652 11082
rect 10600 11018 10652 11024
rect 10598 2680 10654 2689
rect 10598 2615 10654 2624
rect 10612 2446 10640 2615
rect 10600 2440 10652 2446
rect 10600 2382 10652 2388
rect 10704 950 10732 13126
rect 10888 12434 10916 13330
rect 10796 12406 10916 12434
rect 11164 12434 11192 14350
rect 11346 14172 11654 14181
rect 11346 14170 11352 14172
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11648 14170 11654 14172
rect 11408 14118 11410 14170
rect 11590 14118 11592 14170
rect 11346 14116 11352 14118
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11648 14116 11654 14118
rect 11346 14107 11654 14116
rect 11704 13320 11756 13326
rect 11704 13262 11756 13268
rect 11346 13084 11654 13093
rect 11346 13082 11352 13084
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11648 13082 11654 13084
rect 11408 13030 11410 13082
rect 11590 13030 11592 13082
rect 11346 13028 11352 13030
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11648 13028 11654 13030
rect 11346 13019 11654 13028
rect 11716 12986 11744 13262
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 11808 12434 11836 15506
rect 11888 14544 11940 14550
rect 11888 14486 11940 14492
rect 11900 14278 11928 14486
rect 11888 14272 11940 14278
rect 11888 14214 11940 14220
rect 11900 14006 11928 14214
rect 11888 14000 11940 14006
rect 11888 13942 11940 13948
rect 11980 13864 12032 13870
rect 11980 13806 12032 13812
rect 11992 13258 12020 13806
rect 11980 13252 12032 13258
rect 11980 13194 12032 13200
rect 12072 13184 12124 13190
rect 12072 13126 12124 13132
rect 11980 12912 12032 12918
rect 11980 12854 12032 12860
rect 11164 12406 11284 12434
rect 11808 12406 11928 12434
rect 10796 11830 10824 12406
rect 10876 12300 10928 12306
rect 10876 12242 10928 12248
rect 10784 11824 10836 11830
rect 10784 11766 10836 11772
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 10796 11150 10824 11494
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 10784 10804 10836 10810
rect 10784 10746 10836 10752
rect 10796 9586 10824 10746
rect 10888 10062 10916 12242
rect 10966 11112 11022 11121
rect 10966 11047 11022 11056
rect 10876 10056 10928 10062
rect 10876 9998 10928 10004
rect 10980 9586 11008 11047
rect 11060 11008 11112 11014
rect 11060 10950 11112 10956
rect 11072 9994 11100 10950
rect 11060 9988 11112 9994
rect 11060 9930 11112 9936
rect 10784 9580 10836 9586
rect 10784 9522 10836 9528
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 11060 9512 11112 9518
rect 11060 9454 11112 9460
rect 10876 8968 10928 8974
rect 10876 8910 10928 8916
rect 10888 8838 10916 8910
rect 10876 8832 10928 8838
rect 10876 8774 10928 8780
rect 10966 7712 11022 7721
rect 10966 7647 11022 7656
rect 10980 7478 11008 7647
rect 10968 7472 11020 7478
rect 10968 7414 11020 7420
rect 10874 5808 10930 5817
rect 10874 5743 10930 5752
rect 10888 5234 10916 5743
rect 10876 5228 10928 5234
rect 10876 5170 10928 5176
rect 10888 4826 10916 5170
rect 10876 4820 10928 4826
rect 10876 4762 10928 4768
rect 11072 4554 11100 9454
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 11164 8634 11192 8910
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 11150 7848 11206 7857
rect 11150 7783 11206 7792
rect 11164 7546 11192 7783
rect 11152 7540 11204 7546
rect 11152 7482 11204 7488
rect 11152 6724 11204 6730
rect 11152 6666 11204 6672
rect 11164 5846 11192 6666
rect 11152 5840 11204 5846
rect 11152 5782 11204 5788
rect 11152 5568 11204 5574
rect 11152 5510 11204 5516
rect 11164 5234 11192 5510
rect 11152 5228 11204 5234
rect 11152 5170 11204 5176
rect 11164 4690 11192 5170
rect 11152 4684 11204 4690
rect 11152 4626 11204 4632
rect 11060 4548 11112 4554
rect 11060 4490 11112 4496
rect 10876 4480 10928 4486
rect 10876 4422 10928 4428
rect 10692 944 10744 950
rect 10692 886 10744 892
rect 10888 800 10916 4422
rect 11072 2582 11100 4490
rect 11164 4282 11192 4626
rect 11152 4276 11204 4282
rect 11152 4218 11204 4224
rect 11164 3602 11192 4218
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 11164 3058 11192 3538
rect 11152 3052 11204 3058
rect 11152 2994 11204 3000
rect 11164 2650 11192 2994
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 11060 2576 11112 2582
rect 11060 2518 11112 2524
rect 11256 800 11284 12406
rect 11796 12232 11848 12238
rect 11796 12174 11848 12180
rect 11704 12164 11756 12170
rect 11704 12106 11756 12112
rect 11346 11996 11654 12005
rect 11346 11994 11352 11996
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11648 11994 11654 11996
rect 11408 11942 11410 11994
rect 11590 11942 11592 11994
rect 11346 11940 11352 11942
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11648 11940 11654 11942
rect 11346 11931 11654 11940
rect 11716 11898 11744 12106
rect 11704 11892 11756 11898
rect 11704 11834 11756 11840
rect 11336 11824 11388 11830
rect 11336 11766 11388 11772
rect 11348 11558 11376 11766
rect 11704 11756 11756 11762
rect 11704 11698 11756 11704
rect 11336 11552 11388 11558
rect 11336 11494 11388 11500
rect 11346 10908 11654 10917
rect 11346 10906 11352 10908
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11648 10906 11654 10908
rect 11408 10854 11410 10906
rect 11590 10854 11592 10906
rect 11346 10852 11352 10854
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11648 10852 11654 10854
rect 11346 10843 11654 10852
rect 11346 9820 11654 9829
rect 11346 9818 11352 9820
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11648 9818 11654 9820
rect 11408 9766 11410 9818
rect 11590 9766 11592 9818
rect 11346 9764 11352 9766
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11648 9764 11654 9766
rect 11346 9755 11654 9764
rect 11716 9722 11744 11698
rect 11808 11694 11836 12174
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 11900 11354 11928 12406
rect 11888 11348 11940 11354
rect 11888 11290 11940 11296
rect 11794 10160 11850 10169
rect 11794 10095 11850 10104
rect 11704 9716 11756 9722
rect 11704 9658 11756 9664
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 11346 8732 11654 8741
rect 11346 8730 11352 8732
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11648 8730 11654 8732
rect 11408 8678 11410 8730
rect 11590 8678 11592 8730
rect 11346 8676 11352 8678
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11648 8676 11654 8678
rect 11346 8667 11654 8676
rect 11336 8084 11388 8090
rect 11336 8026 11388 8032
rect 11348 7818 11376 8026
rect 11336 7812 11388 7818
rect 11336 7754 11388 7760
rect 11346 7644 11654 7653
rect 11346 7642 11352 7644
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11648 7642 11654 7644
rect 11408 7590 11410 7642
rect 11590 7590 11592 7642
rect 11346 7588 11352 7590
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11648 7588 11654 7590
rect 11346 7579 11654 7588
rect 11346 6556 11654 6565
rect 11346 6554 11352 6556
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11648 6554 11654 6556
rect 11408 6502 11410 6554
rect 11590 6502 11592 6554
rect 11346 6500 11352 6502
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11648 6500 11654 6502
rect 11346 6491 11654 6500
rect 11346 5468 11654 5477
rect 11346 5466 11352 5468
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11648 5466 11654 5468
rect 11408 5414 11410 5466
rect 11590 5414 11592 5466
rect 11346 5412 11352 5414
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11648 5412 11654 5414
rect 11346 5403 11654 5412
rect 11612 5024 11664 5030
rect 11612 4966 11664 4972
rect 11716 4978 11744 9522
rect 11808 6254 11836 10095
rect 11888 9988 11940 9994
rect 11888 9930 11940 9936
rect 11796 6248 11848 6254
rect 11796 6190 11848 6196
rect 11808 5098 11836 6190
rect 11900 6118 11928 9930
rect 11992 8906 12020 12854
rect 11980 8900 12032 8906
rect 11980 8842 12032 8848
rect 11992 8362 12020 8842
rect 11980 8356 12032 8362
rect 11980 8298 12032 8304
rect 11888 6112 11940 6118
rect 11888 6054 11940 6060
rect 11796 5092 11848 5098
rect 11796 5034 11848 5040
rect 11624 4826 11652 4966
rect 11716 4950 11836 4978
rect 11612 4820 11664 4826
rect 11612 4762 11664 4768
rect 11702 4584 11758 4593
rect 11702 4519 11758 4528
rect 11346 4380 11654 4389
rect 11346 4378 11352 4380
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11648 4378 11654 4380
rect 11408 4326 11410 4378
rect 11590 4326 11592 4378
rect 11346 4324 11352 4326
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11648 4324 11654 4326
rect 11346 4315 11654 4324
rect 11716 4146 11744 4519
rect 11704 4140 11756 4146
rect 11704 4082 11756 4088
rect 11716 3618 11744 4082
rect 11624 3602 11744 3618
rect 11612 3596 11744 3602
rect 11664 3590 11744 3596
rect 11612 3538 11664 3544
rect 11346 3292 11654 3301
rect 11346 3290 11352 3292
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11648 3290 11654 3292
rect 11408 3238 11410 3290
rect 11590 3238 11592 3290
rect 11346 3236 11352 3238
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11648 3236 11654 3238
rect 11346 3227 11654 3236
rect 11428 3188 11480 3194
rect 11428 3130 11480 3136
rect 11440 2990 11468 3130
rect 11428 2984 11480 2990
rect 11428 2926 11480 2932
rect 11808 2774 11836 4950
rect 11808 2746 12020 2774
rect 11704 2304 11756 2310
rect 11704 2246 11756 2252
rect 11346 2204 11654 2213
rect 11346 2202 11352 2204
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11648 2202 11654 2204
rect 11408 2150 11410 2202
rect 11590 2150 11592 2202
rect 11346 2148 11352 2150
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11648 2148 11654 2150
rect 11346 2139 11654 2148
rect 11716 1902 11744 2246
rect 11704 1896 11756 1902
rect 11704 1838 11756 1844
rect 11992 1290 12020 2746
rect 11980 1284 12032 1290
rect 11980 1226 12032 1232
rect 12084 1170 12112 13126
rect 12176 12986 12204 17138
rect 13945 16892 14253 16901
rect 13945 16890 13951 16892
rect 14007 16890 14031 16892
rect 14087 16890 14111 16892
rect 14167 16890 14191 16892
rect 14247 16890 14253 16892
rect 14007 16838 14009 16890
rect 14189 16838 14191 16890
rect 13945 16836 13951 16838
rect 14007 16836 14031 16838
rect 14087 16836 14111 16838
rect 14167 16836 14191 16838
rect 14247 16836 14253 16838
rect 13945 16827 14253 16836
rect 19143 16892 19451 16901
rect 19143 16890 19149 16892
rect 19205 16890 19229 16892
rect 19285 16890 19309 16892
rect 19365 16890 19389 16892
rect 19445 16890 19451 16892
rect 19205 16838 19207 16890
rect 19387 16838 19389 16890
rect 19143 16836 19149 16838
rect 19205 16836 19229 16838
rect 19285 16836 19309 16838
rect 19365 16836 19389 16838
rect 19445 16836 19451 16838
rect 19143 16827 19451 16836
rect 21468 16658 21496 17167
rect 21456 16652 21508 16658
rect 21456 16594 21508 16600
rect 16544 16348 16852 16357
rect 16544 16346 16550 16348
rect 16606 16346 16630 16348
rect 16686 16346 16710 16348
rect 16766 16346 16790 16348
rect 16846 16346 16852 16348
rect 16606 16294 16608 16346
rect 16788 16294 16790 16346
rect 16544 16292 16550 16294
rect 16606 16292 16630 16294
rect 16686 16292 16710 16294
rect 16766 16292 16790 16294
rect 16846 16292 16852 16294
rect 16544 16283 16852 16292
rect 13945 15804 14253 15813
rect 13945 15802 13951 15804
rect 14007 15802 14031 15804
rect 14087 15802 14111 15804
rect 14167 15802 14191 15804
rect 14247 15802 14253 15804
rect 14007 15750 14009 15802
rect 14189 15750 14191 15802
rect 13945 15748 13951 15750
rect 14007 15748 14031 15750
rect 14087 15748 14111 15750
rect 14167 15748 14191 15750
rect 14247 15748 14253 15750
rect 13945 15739 14253 15748
rect 19143 15804 19451 15813
rect 19143 15802 19149 15804
rect 19205 15802 19229 15804
rect 19285 15802 19309 15804
rect 19365 15802 19389 15804
rect 19445 15802 19451 15804
rect 19205 15750 19207 15802
rect 19387 15750 19389 15802
rect 19143 15748 19149 15750
rect 19205 15748 19229 15750
rect 19285 15748 19309 15750
rect 19365 15748 19389 15750
rect 19445 15748 19451 15750
rect 19143 15739 19451 15748
rect 16544 15260 16852 15269
rect 16544 15258 16550 15260
rect 16606 15258 16630 15260
rect 16686 15258 16710 15260
rect 16766 15258 16790 15260
rect 16846 15258 16852 15260
rect 16606 15206 16608 15258
rect 16788 15206 16790 15258
rect 16544 15204 16550 15206
rect 16606 15204 16630 15206
rect 16686 15204 16710 15206
rect 16766 15204 16790 15206
rect 16846 15204 16852 15206
rect 16544 15195 16852 15204
rect 15568 14952 15620 14958
rect 15568 14894 15620 14900
rect 13945 14716 14253 14725
rect 13945 14714 13951 14716
rect 14007 14714 14031 14716
rect 14087 14714 14111 14716
rect 14167 14714 14191 14716
rect 14247 14714 14253 14716
rect 14007 14662 14009 14714
rect 14189 14662 14191 14714
rect 13945 14660 13951 14662
rect 14007 14660 14031 14662
rect 14087 14660 14111 14662
rect 14167 14660 14191 14662
rect 14247 14660 14253 14662
rect 13945 14651 14253 14660
rect 12348 14408 12400 14414
rect 12348 14350 12400 14356
rect 12360 14006 12388 14350
rect 12900 14272 12952 14278
rect 12900 14214 12952 14220
rect 12912 14074 12940 14214
rect 12900 14068 12952 14074
rect 12900 14010 12952 14016
rect 12348 14000 12400 14006
rect 12348 13942 12400 13948
rect 13084 13728 13136 13734
rect 13084 13670 13136 13676
rect 12164 12980 12216 12986
rect 12164 12922 12216 12928
rect 12716 12640 12768 12646
rect 12716 12582 12768 12588
rect 12348 12164 12400 12170
rect 12348 12106 12400 12112
rect 12254 11792 12310 11801
rect 12360 11762 12388 12106
rect 12254 11727 12310 11736
rect 12348 11756 12400 11762
rect 12268 11014 12296 11727
rect 12348 11698 12400 11704
rect 12256 11008 12308 11014
rect 12256 10950 12308 10956
rect 12268 10010 12296 10950
rect 12624 10532 12676 10538
rect 12624 10474 12676 10480
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12452 10266 12480 10406
rect 12440 10260 12492 10266
rect 12440 10202 12492 10208
rect 12268 9982 12388 10010
rect 12256 9920 12308 9926
rect 12256 9862 12308 9868
rect 12268 8498 12296 9862
rect 12256 8492 12308 8498
rect 12256 8434 12308 8440
rect 12360 7410 12388 9982
rect 12636 9654 12664 10474
rect 12728 9994 12756 12582
rect 13096 10470 13124 13670
rect 13945 13628 14253 13637
rect 13945 13626 13951 13628
rect 14007 13626 14031 13628
rect 14087 13626 14111 13628
rect 14167 13626 14191 13628
rect 14247 13626 14253 13628
rect 14007 13574 14009 13626
rect 14189 13574 14191 13626
rect 13945 13572 13951 13574
rect 14007 13572 14031 13574
rect 14087 13572 14111 13574
rect 14167 13572 14191 13574
rect 14247 13572 14253 13574
rect 13945 13563 14253 13572
rect 13945 12540 14253 12549
rect 13945 12538 13951 12540
rect 14007 12538 14031 12540
rect 14087 12538 14111 12540
rect 14167 12538 14191 12540
rect 14247 12538 14253 12540
rect 14007 12486 14009 12538
rect 14189 12486 14191 12538
rect 13945 12484 13951 12486
rect 14007 12484 14031 12486
rect 14087 12484 14111 12486
rect 14167 12484 14191 12486
rect 14247 12484 14253 12486
rect 13945 12475 14253 12484
rect 13176 12436 13228 12442
rect 13176 12378 13228 12384
rect 13188 12102 13216 12378
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 13728 12096 13780 12102
rect 13728 12038 13780 12044
rect 13188 11898 13216 12038
rect 13176 11892 13228 11898
rect 13176 11834 13228 11840
rect 13740 11762 13768 12038
rect 15580 11898 15608 14894
rect 19143 14716 19451 14725
rect 19143 14714 19149 14716
rect 19205 14714 19229 14716
rect 19285 14714 19309 14716
rect 19365 14714 19389 14716
rect 19445 14714 19451 14716
rect 19205 14662 19207 14714
rect 19387 14662 19389 14714
rect 19143 14660 19149 14662
rect 19205 14660 19229 14662
rect 19285 14660 19309 14662
rect 19365 14660 19389 14662
rect 19445 14660 19451 14662
rect 19143 14651 19451 14660
rect 16544 14172 16852 14181
rect 16544 14170 16550 14172
rect 16606 14170 16630 14172
rect 16686 14170 16710 14172
rect 16766 14170 16790 14172
rect 16846 14170 16852 14172
rect 16606 14118 16608 14170
rect 16788 14118 16790 14170
rect 16544 14116 16550 14118
rect 16606 14116 16630 14118
rect 16686 14116 16710 14118
rect 16766 14116 16790 14118
rect 16846 14116 16852 14118
rect 16544 14107 16852 14116
rect 19984 13796 20036 13802
rect 19984 13738 20036 13744
rect 15660 13728 15712 13734
rect 15660 13670 15712 13676
rect 15672 12102 15700 13670
rect 19143 13628 19451 13637
rect 19143 13626 19149 13628
rect 19205 13626 19229 13628
rect 19285 13626 19309 13628
rect 19365 13626 19389 13628
rect 19445 13626 19451 13628
rect 19205 13574 19207 13626
rect 19387 13574 19389 13626
rect 19143 13572 19149 13574
rect 19205 13572 19229 13574
rect 19285 13572 19309 13574
rect 19365 13572 19389 13574
rect 19445 13572 19451 13574
rect 19143 13563 19451 13572
rect 19522 13424 19578 13433
rect 17960 13388 18012 13394
rect 19522 13359 19578 13368
rect 17960 13330 18012 13336
rect 16544 13084 16852 13093
rect 16544 13082 16550 13084
rect 16606 13082 16630 13084
rect 16686 13082 16710 13084
rect 16766 13082 16790 13084
rect 16846 13082 16852 13084
rect 16606 13030 16608 13082
rect 16788 13030 16790 13082
rect 16544 13028 16550 13030
rect 16606 13028 16630 13030
rect 16686 13028 16710 13030
rect 16766 13028 16790 13030
rect 16846 13028 16852 13030
rect 16544 13019 16852 13028
rect 17132 12776 17184 12782
rect 17132 12718 17184 12724
rect 17144 12170 17172 12718
rect 17132 12164 17184 12170
rect 17132 12106 17184 12112
rect 15660 12096 15712 12102
rect 15660 12038 15712 12044
rect 17040 12096 17092 12102
rect 17040 12038 17092 12044
rect 15568 11892 15620 11898
rect 15568 11834 15620 11840
rect 13728 11756 13780 11762
rect 13728 11698 13780 11704
rect 13450 11656 13506 11665
rect 13450 11591 13506 11600
rect 13464 11558 13492 11591
rect 13740 11558 13768 11698
rect 13452 11552 13504 11558
rect 13452 11494 13504 11500
rect 13728 11552 13780 11558
rect 13728 11494 13780 11500
rect 13360 11076 13412 11082
rect 13360 11018 13412 11024
rect 13084 10464 13136 10470
rect 13084 10406 13136 10412
rect 12716 9988 12768 9994
rect 12716 9930 12768 9936
rect 12532 9648 12584 9654
rect 12532 9590 12584 9596
rect 12624 9648 12676 9654
rect 12624 9590 12676 9596
rect 12544 7818 12572 9590
rect 12992 9104 13044 9110
rect 12992 9046 13044 9052
rect 12900 9036 12952 9042
rect 12900 8978 12952 8984
rect 12912 8566 12940 8978
rect 13004 8838 13032 9046
rect 12992 8832 13044 8838
rect 12992 8774 13044 8780
rect 13096 8566 13124 10406
rect 13268 10260 13320 10266
rect 13268 10202 13320 10208
rect 13280 9654 13308 10202
rect 13268 9648 13320 9654
rect 13268 9590 13320 9596
rect 13280 9382 13308 9590
rect 13268 9376 13320 9382
rect 13268 9318 13320 9324
rect 13280 8838 13308 9318
rect 13268 8832 13320 8838
rect 13268 8774 13320 8780
rect 12900 8560 12952 8566
rect 12900 8502 12952 8508
rect 13084 8560 13136 8566
rect 13084 8502 13136 8508
rect 13280 8430 13308 8774
rect 13372 8634 13400 11018
rect 13464 8974 13492 11494
rect 13740 11150 13768 11494
rect 13945 11452 14253 11461
rect 13945 11450 13951 11452
rect 14007 11450 14031 11452
rect 14087 11450 14111 11452
rect 14167 11450 14191 11452
rect 14247 11450 14253 11452
rect 14007 11398 14009 11450
rect 14189 11398 14191 11450
rect 13945 11396 13951 11398
rect 14007 11396 14031 11398
rect 14087 11396 14111 11398
rect 14167 11396 14191 11398
rect 14247 11396 14253 11398
rect 13945 11387 14253 11396
rect 13820 11348 13872 11354
rect 13820 11290 13872 11296
rect 15476 11348 15528 11354
rect 15476 11290 15528 11296
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13452 8968 13504 8974
rect 13452 8910 13504 8916
rect 13360 8628 13412 8634
rect 13360 8570 13412 8576
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 13280 7886 13308 8366
rect 13268 7880 13320 7886
rect 13268 7822 13320 7828
rect 13728 7880 13780 7886
rect 13728 7822 13780 7828
rect 12532 7812 12584 7818
rect 12532 7754 12584 7760
rect 12348 7404 12400 7410
rect 12348 7346 12400 7352
rect 12440 6724 12492 6730
rect 12440 6666 12492 6672
rect 12348 6656 12400 6662
rect 12348 6598 12400 6604
rect 12360 6338 12388 6598
rect 12452 6338 12480 6666
rect 12360 6310 12480 6338
rect 12256 5704 12308 5710
rect 12256 5646 12308 5652
rect 12268 4468 12296 5646
rect 12440 5296 12492 5302
rect 12440 5238 12492 5244
rect 12452 4758 12480 5238
rect 12544 4826 12572 7754
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 12636 5302 12664 7482
rect 13360 7472 13412 7478
rect 13360 7414 13412 7420
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 13188 7002 13216 7142
rect 13372 7002 13400 7414
rect 13740 7410 13768 7822
rect 13832 7818 13860 11290
rect 14464 11280 14516 11286
rect 14462 11248 14464 11257
rect 14516 11248 14518 11257
rect 14462 11183 14518 11192
rect 14464 11008 14516 11014
rect 14464 10950 14516 10956
rect 14476 10606 14504 10950
rect 15488 10674 15516 11290
rect 15580 11082 15608 11834
rect 15568 11076 15620 11082
rect 15568 11018 15620 11024
rect 15672 10742 15700 12038
rect 16544 11996 16852 12005
rect 16544 11994 16550 11996
rect 16606 11994 16630 11996
rect 16686 11994 16710 11996
rect 16766 11994 16790 11996
rect 16846 11994 16852 11996
rect 16606 11942 16608 11994
rect 16788 11942 16790 11994
rect 16544 11940 16550 11942
rect 16606 11940 16630 11942
rect 16686 11940 16710 11942
rect 16766 11940 16790 11942
rect 16846 11940 16852 11942
rect 16544 11931 16852 11940
rect 16488 11824 16540 11830
rect 16488 11766 16540 11772
rect 16120 11756 16172 11762
rect 16120 11698 16172 11704
rect 16132 11150 16160 11698
rect 16500 11354 16528 11766
rect 16488 11348 16540 11354
rect 16488 11290 16540 11296
rect 16120 11144 16172 11150
rect 16120 11086 16172 11092
rect 15660 10736 15712 10742
rect 15660 10678 15712 10684
rect 15476 10668 15528 10674
rect 15476 10610 15528 10616
rect 15568 10668 15620 10674
rect 15568 10610 15620 10616
rect 14464 10600 14516 10606
rect 14464 10542 14516 10548
rect 13945 10364 14253 10373
rect 13945 10362 13951 10364
rect 14007 10362 14031 10364
rect 14087 10362 14111 10364
rect 14167 10362 14191 10364
rect 14247 10362 14253 10364
rect 14007 10310 14009 10362
rect 14189 10310 14191 10362
rect 13945 10308 13951 10310
rect 14007 10308 14031 10310
rect 14087 10308 14111 10310
rect 14167 10308 14191 10310
rect 14247 10308 14253 10310
rect 13945 10299 14253 10308
rect 14476 10266 14504 10542
rect 14464 10260 14516 10266
rect 14464 10202 14516 10208
rect 14462 9480 14518 9489
rect 14462 9415 14518 9424
rect 13945 9276 14253 9285
rect 13945 9274 13951 9276
rect 14007 9274 14031 9276
rect 14087 9274 14111 9276
rect 14167 9274 14191 9276
rect 14247 9274 14253 9276
rect 14007 9222 14009 9274
rect 14189 9222 14191 9274
rect 13945 9220 13951 9222
rect 14007 9220 14031 9222
rect 14087 9220 14111 9222
rect 14167 9220 14191 9222
rect 14247 9220 14253 9222
rect 13945 9211 14253 9220
rect 14370 8936 14426 8945
rect 14370 8871 14426 8880
rect 14384 8838 14412 8871
rect 14372 8832 14424 8838
rect 14372 8774 14424 8780
rect 14188 8492 14240 8498
rect 14240 8452 14320 8480
rect 14188 8434 14240 8440
rect 13945 8188 14253 8197
rect 13945 8186 13951 8188
rect 14007 8186 14031 8188
rect 14087 8186 14111 8188
rect 14167 8186 14191 8188
rect 14247 8186 14253 8188
rect 14007 8134 14009 8186
rect 14189 8134 14191 8186
rect 13945 8132 13951 8134
rect 14007 8132 14031 8134
rect 14087 8132 14111 8134
rect 14167 8132 14191 8134
rect 14247 8132 14253 8134
rect 13945 8123 14253 8132
rect 13820 7812 13872 7818
rect 13820 7754 13872 7760
rect 13728 7404 13780 7410
rect 13728 7346 13780 7352
rect 13740 7002 13768 7346
rect 13945 7100 14253 7109
rect 13945 7098 13951 7100
rect 14007 7098 14031 7100
rect 14087 7098 14111 7100
rect 14167 7098 14191 7100
rect 14247 7098 14253 7100
rect 14007 7046 14009 7098
rect 14189 7046 14191 7098
rect 13945 7044 13951 7046
rect 14007 7044 14031 7046
rect 14087 7044 14111 7046
rect 14167 7044 14191 7046
rect 14247 7044 14253 7046
rect 13945 7035 14253 7044
rect 13176 6996 13228 7002
rect 13176 6938 13228 6944
rect 13360 6996 13412 7002
rect 13360 6938 13412 6944
rect 13728 6996 13780 7002
rect 13728 6938 13780 6944
rect 13740 6798 13768 6938
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 13740 6322 13768 6734
rect 14292 6662 14320 8452
rect 14280 6656 14332 6662
rect 14280 6598 14332 6604
rect 14292 6322 14320 6598
rect 13728 6316 13780 6322
rect 13728 6258 13780 6264
rect 14280 6316 14332 6322
rect 14280 6258 14332 6264
rect 13740 5914 13768 6258
rect 13945 6012 14253 6021
rect 13945 6010 13951 6012
rect 14007 6010 14031 6012
rect 14087 6010 14111 6012
rect 14167 6010 14191 6012
rect 14247 6010 14253 6012
rect 14007 5958 14009 6010
rect 14189 5958 14191 6010
rect 13945 5956 13951 5958
rect 14007 5956 14031 5958
rect 14087 5956 14111 5958
rect 14167 5956 14191 5958
rect 14247 5956 14253 5958
rect 13945 5947 14253 5956
rect 13452 5908 13504 5914
rect 13452 5850 13504 5856
rect 13728 5908 13780 5914
rect 13728 5850 13780 5856
rect 13464 5778 13492 5850
rect 13452 5772 13504 5778
rect 13452 5714 13504 5720
rect 13464 5370 13492 5714
rect 14384 5642 14412 8774
rect 14476 8498 14504 9415
rect 14556 9104 14608 9110
rect 14556 9046 14608 9052
rect 14568 8838 14596 9046
rect 14556 8832 14608 8838
rect 14556 8774 14608 8780
rect 14464 8492 14516 8498
rect 14464 8434 14516 8440
rect 14476 7546 14504 8434
rect 15476 8084 15528 8090
rect 15580 8072 15608 10610
rect 16132 10606 16160 11086
rect 16304 11008 16356 11014
rect 16304 10950 16356 10956
rect 16316 10810 16344 10950
rect 16544 10908 16852 10917
rect 16544 10906 16550 10908
rect 16606 10906 16630 10908
rect 16686 10906 16710 10908
rect 16766 10906 16790 10908
rect 16846 10906 16852 10908
rect 16606 10854 16608 10906
rect 16788 10854 16790 10906
rect 16544 10852 16550 10854
rect 16606 10852 16630 10854
rect 16686 10852 16710 10854
rect 16766 10852 16790 10854
rect 16846 10852 16852 10854
rect 16544 10843 16852 10852
rect 16304 10804 16356 10810
rect 16304 10746 16356 10752
rect 16948 10668 17000 10674
rect 16948 10610 17000 10616
rect 16120 10600 16172 10606
rect 16120 10542 16172 10548
rect 16132 10266 16160 10542
rect 16120 10260 16172 10266
rect 16120 10202 16172 10208
rect 16544 9820 16852 9829
rect 16544 9818 16550 9820
rect 16606 9818 16630 9820
rect 16686 9818 16710 9820
rect 16766 9818 16790 9820
rect 16846 9818 16852 9820
rect 16606 9766 16608 9818
rect 16788 9766 16790 9818
rect 16544 9764 16550 9766
rect 16606 9764 16630 9766
rect 16686 9764 16710 9766
rect 16766 9764 16790 9766
rect 16846 9764 16852 9766
rect 16544 9755 16852 9764
rect 16960 9178 16988 10610
rect 17052 9450 17080 12038
rect 17144 10266 17172 12106
rect 17132 10260 17184 10266
rect 17132 10202 17184 10208
rect 17040 9444 17092 9450
rect 17040 9386 17092 9392
rect 16948 9172 17000 9178
rect 16948 9114 17000 9120
rect 15752 8968 15804 8974
rect 15752 8910 15804 8916
rect 15764 8634 15792 8910
rect 16948 8900 17000 8906
rect 16948 8842 17000 8848
rect 16544 8732 16852 8741
rect 16544 8730 16550 8732
rect 16606 8730 16630 8732
rect 16686 8730 16710 8732
rect 16766 8730 16790 8732
rect 16846 8730 16852 8732
rect 16606 8678 16608 8730
rect 16788 8678 16790 8730
rect 16544 8676 16550 8678
rect 16606 8676 16630 8678
rect 16686 8676 16710 8678
rect 16766 8676 16790 8678
rect 16846 8676 16852 8678
rect 16544 8667 16852 8676
rect 15752 8628 15804 8634
rect 15752 8570 15804 8576
rect 15658 8392 15714 8401
rect 15658 8327 15714 8336
rect 15672 8090 15700 8327
rect 15528 8044 15608 8072
rect 15660 8084 15712 8090
rect 15476 8026 15528 8032
rect 15660 8026 15712 8032
rect 15764 7954 15792 8570
rect 16960 8090 16988 8842
rect 17972 8634 18000 13330
rect 19143 12540 19451 12549
rect 19143 12538 19149 12540
rect 19205 12538 19229 12540
rect 19285 12538 19309 12540
rect 19365 12538 19389 12540
rect 19445 12538 19451 12540
rect 19205 12486 19207 12538
rect 19387 12486 19389 12538
rect 19143 12484 19149 12486
rect 19205 12484 19229 12486
rect 19285 12484 19309 12486
rect 19365 12484 19389 12486
rect 19445 12484 19451 12486
rect 19143 12475 19451 12484
rect 18602 12336 18658 12345
rect 18602 12271 18658 12280
rect 18328 12096 18380 12102
rect 18328 12038 18380 12044
rect 18340 11694 18368 12038
rect 18616 11830 18644 12271
rect 18604 11824 18656 11830
rect 18604 11766 18656 11772
rect 18328 11688 18380 11694
rect 18328 11630 18380 11636
rect 18052 11552 18104 11558
rect 18052 11494 18104 11500
rect 18064 9654 18092 11494
rect 18340 11014 18368 11630
rect 18328 11008 18380 11014
rect 18328 10950 18380 10956
rect 18616 10810 18644 11766
rect 19143 11452 19451 11461
rect 19143 11450 19149 11452
rect 19205 11450 19229 11452
rect 19285 11450 19309 11452
rect 19365 11450 19389 11452
rect 19445 11450 19451 11452
rect 19205 11398 19207 11450
rect 19387 11398 19389 11450
rect 19143 11396 19149 11398
rect 19205 11396 19229 11398
rect 19285 11396 19309 11398
rect 19365 11396 19389 11398
rect 19445 11396 19451 11398
rect 19143 11387 19451 11396
rect 19536 11354 19564 13359
rect 19996 11898 20024 13738
rect 21364 12096 21416 12102
rect 21364 12038 21416 12044
rect 19984 11892 20036 11898
rect 19984 11834 20036 11840
rect 19524 11348 19576 11354
rect 19524 11290 19576 11296
rect 19996 11150 20024 11834
rect 21376 11762 21404 12038
rect 21088 11756 21140 11762
rect 21088 11698 21140 11704
rect 21364 11756 21416 11762
rect 21364 11698 21416 11704
rect 20628 11552 20680 11558
rect 20628 11494 20680 11500
rect 19984 11144 20036 11150
rect 19984 11086 20036 11092
rect 19800 11008 19852 11014
rect 19800 10950 19852 10956
rect 18604 10804 18656 10810
rect 18604 10746 18656 10752
rect 19812 10742 19840 10950
rect 19800 10736 19852 10742
rect 19800 10678 19852 10684
rect 19432 10668 19484 10674
rect 19432 10610 19484 10616
rect 19444 10554 19472 10610
rect 19444 10526 19564 10554
rect 19143 10364 19451 10373
rect 19143 10362 19149 10364
rect 19205 10362 19229 10364
rect 19285 10362 19309 10364
rect 19365 10362 19389 10364
rect 19445 10362 19451 10364
rect 19205 10310 19207 10362
rect 19387 10310 19389 10362
rect 19143 10308 19149 10310
rect 19205 10308 19229 10310
rect 19285 10308 19309 10310
rect 19365 10308 19389 10310
rect 19445 10308 19451 10310
rect 19143 10299 19451 10308
rect 19340 10056 19392 10062
rect 19340 9998 19392 10004
rect 18420 9988 18472 9994
rect 18420 9930 18472 9936
rect 18052 9648 18104 9654
rect 18052 9590 18104 9596
rect 18432 9178 18460 9930
rect 19352 9586 19380 9998
rect 19432 9988 19484 9994
rect 19432 9930 19484 9936
rect 19444 9722 19472 9930
rect 19432 9716 19484 9722
rect 19432 9658 19484 9664
rect 19340 9580 19392 9586
rect 19340 9522 19392 9528
rect 19143 9276 19451 9285
rect 19143 9274 19149 9276
rect 19205 9274 19229 9276
rect 19285 9274 19309 9276
rect 19365 9274 19389 9276
rect 19445 9274 19451 9276
rect 19205 9222 19207 9274
rect 19387 9222 19389 9274
rect 19143 9220 19149 9222
rect 19205 9220 19229 9222
rect 19285 9220 19309 9222
rect 19365 9220 19389 9222
rect 19445 9220 19451 9222
rect 19143 9211 19451 9220
rect 18420 9172 18472 9178
rect 18420 9114 18472 9120
rect 18328 8968 18380 8974
rect 18328 8910 18380 8916
rect 18052 8900 18104 8906
rect 18052 8842 18104 8848
rect 17960 8628 18012 8634
rect 17960 8570 18012 8576
rect 16948 8084 17000 8090
rect 16948 8026 17000 8032
rect 15752 7948 15804 7954
rect 15752 7890 15804 7896
rect 15764 7546 15792 7890
rect 16212 7812 16264 7818
rect 16212 7754 16264 7760
rect 14464 7540 14516 7546
rect 14464 7482 14516 7488
rect 15752 7540 15804 7546
rect 15752 7482 15804 7488
rect 15764 7002 15792 7482
rect 15752 6996 15804 7002
rect 15752 6938 15804 6944
rect 15476 6792 15528 6798
rect 15474 6760 15476 6769
rect 15528 6760 15530 6769
rect 15474 6695 15530 6704
rect 15384 6656 15436 6662
rect 15384 6598 15436 6604
rect 14740 6112 14792 6118
rect 14740 6054 14792 6060
rect 14752 5710 14780 6054
rect 14740 5704 14792 5710
rect 14740 5646 14792 5652
rect 14372 5636 14424 5642
rect 14372 5578 14424 5584
rect 14096 5568 14148 5574
rect 14096 5510 14148 5516
rect 13452 5364 13504 5370
rect 13452 5306 13504 5312
rect 14108 5302 14136 5510
rect 12624 5296 12676 5302
rect 12624 5238 12676 5244
rect 14096 5296 14148 5302
rect 14096 5238 14148 5244
rect 12992 5228 13044 5234
rect 12992 5170 13044 5176
rect 13004 4826 13032 5170
rect 15200 5024 15252 5030
rect 15200 4966 15252 4972
rect 13945 4924 14253 4933
rect 13945 4922 13951 4924
rect 14007 4922 14031 4924
rect 14087 4922 14111 4924
rect 14167 4922 14191 4924
rect 14247 4922 14253 4924
rect 14007 4870 14009 4922
rect 14189 4870 14191 4922
rect 13945 4868 13951 4870
rect 14007 4868 14031 4870
rect 14087 4868 14111 4870
rect 14167 4868 14191 4870
rect 14247 4868 14253 4870
rect 13945 4859 14253 4868
rect 12532 4820 12584 4826
rect 12532 4762 12584 4768
rect 12992 4820 13044 4826
rect 12992 4762 13044 4768
rect 13636 4820 13688 4826
rect 13636 4762 13688 4768
rect 12440 4752 12492 4758
rect 12440 4694 12492 4700
rect 12440 4480 12492 4486
rect 12268 4440 12440 4468
rect 12360 3466 12388 4440
rect 12440 4422 12492 4428
rect 12808 4072 12860 4078
rect 12808 4014 12860 4020
rect 12624 3936 12676 3942
rect 12624 3878 12676 3884
rect 12348 3460 12400 3466
rect 12348 3402 12400 3408
rect 12346 2816 12402 2825
rect 12346 2751 12402 2760
rect 11900 1142 12112 1170
rect 11624 870 11744 898
rect 11624 800 11652 870
rect 7300 734 7512 762
rect 7562 0 7618 800
rect 7930 0 7986 800
rect 8298 0 8354 800
rect 8666 0 8722 800
rect 9034 0 9090 800
rect 9402 0 9458 800
rect 9770 0 9826 800
rect 10138 0 10194 800
rect 10506 0 10562 800
rect 10874 0 10930 800
rect 11242 0 11298 800
rect 11610 0 11666 800
rect 11716 762 11744 870
rect 11900 762 11928 1142
rect 11980 1080 12032 1086
rect 11980 1022 12032 1028
rect 11992 800 12020 1022
rect 12360 800 12388 2751
rect 12636 2378 12664 3878
rect 12716 3732 12768 3738
rect 12716 3674 12768 3680
rect 12728 3466 12756 3674
rect 12820 3534 12848 4014
rect 13004 3738 13032 4762
rect 13648 4214 13676 4762
rect 15108 4752 15160 4758
rect 15108 4694 15160 4700
rect 15120 4486 15148 4694
rect 15108 4480 15160 4486
rect 15108 4422 15160 4428
rect 13636 4208 13688 4214
rect 13636 4150 13688 4156
rect 13176 4140 13228 4146
rect 13176 4082 13228 4088
rect 12992 3732 13044 3738
rect 12992 3674 13044 3680
rect 12808 3528 12860 3534
rect 12808 3470 12860 3476
rect 12716 3460 12768 3466
rect 12716 3402 12768 3408
rect 12808 3188 12860 3194
rect 12808 3130 12860 3136
rect 12820 3097 12848 3130
rect 12806 3088 12862 3097
rect 12806 3023 12862 3032
rect 13004 2774 13032 3674
rect 13188 3194 13216 4082
rect 14278 4040 14334 4049
rect 14278 3975 14280 3984
rect 14332 3975 14334 3984
rect 14280 3946 14332 3952
rect 13728 3936 13780 3942
rect 13728 3878 13780 3884
rect 13452 3392 13504 3398
rect 13452 3334 13504 3340
rect 13176 3188 13228 3194
rect 13176 3130 13228 3136
rect 13084 3120 13136 3126
rect 13082 3088 13084 3097
rect 13136 3088 13138 3097
rect 13082 3023 13138 3032
rect 13176 3052 13228 3058
rect 13176 2994 13228 3000
rect 12912 2746 13032 2774
rect 12912 2514 12940 2746
rect 12900 2508 12952 2514
rect 12900 2450 12952 2456
rect 12624 2372 12676 2378
rect 12624 2314 12676 2320
rect 13084 2304 13136 2310
rect 13084 2246 13136 2252
rect 12716 1692 12768 1698
rect 12716 1634 12768 1640
rect 12728 800 12756 1634
rect 13096 800 13124 2246
rect 13188 1970 13216 2994
rect 13176 1964 13228 1970
rect 13176 1906 13228 1912
rect 13464 800 13492 3334
rect 13740 3058 13768 3878
rect 13945 3836 14253 3845
rect 13945 3834 13951 3836
rect 14007 3834 14031 3836
rect 14087 3834 14111 3836
rect 14167 3834 14191 3836
rect 14247 3834 14253 3836
rect 14007 3782 14009 3834
rect 14189 3782 14191 3834
rect 13945 3780 13951 3782
rect 14007 3780 14031 3782
rect 14087 3780 14111 3782
rect 14167 3780 14191 3782
rect 14247 3780 14253 3782
rect 13945 3771 14253 3780
rect 15212 3534 15240 4966
rect 15396 4146 15424 6598
rect 15764 6458 15792 6938
rect 15752 6452 15804 6458
rect 15752 6394 15804 6400
rect 15764 6322 15792 6394
rect 15752 6316 15804 6322
rect 15752 6258 15804 6264
rect 15764 5914 15792 6258
rect 15752 5908 15804 5914
rect 15752 5850 15804 5856
rect 15764 5778 15792 5850
rect 15752 5772 15804 5778
rect 15752 5714 15804 5720
rect 15764 5370 15792 5714
rect 15752 5364 15804 5370
rect 15752 5306 15804 5312
rect 16224 4758 16252 7754
rect 16544 7644 16852 7653
rect 16544 7642 16550 7644
rect 16606 7642 16630 7644
rect 16686 7642 16710 7644
rect 16766 7642 16790 7644
rect 16846 7642 16852 7644
rect 16606 7590 16608 7642
rect 16788 7590 16790 7642
rect 16544 7588 16550 7590
rect 16606 7588 16630 7590
rect 16686 7588 16710 7590
rect 16766 7588 16790 7590
rect 16846 7588 16852 7590
rect 16544 7579 16852 7588
rect 16960 6662 16988 8026
rect 17408 7744 17460 7750
rect 17408 7686 17460 7692
rect 17420 7546 17448 7686
rect 18064 7546 18092 8842
rect 18340 8498 18368 8910
rect 18972 8832 19024 8838
rect 18972 8774 19024 8780
rect 18510 8528 18566 8537
rect 18328 8492 18380 8498
rect 18328 8434 18380 8440
rect 18420 8492 18472 8498
rect 18510 8463 18566 8472
rect 18420 8434 18472 8440
rect 18340 8090 18368 8434
rect 18328 8084 18380 8090
rect 18328 8026 18380 8032
rect 17408 7540 17460 7546
rect 17408 7482 17460 7488
rect 18052 7540 18104 7546
rect 18052 7482 18104 7488
rect 18064 7449 18092 7482
rect 18340 7478 18368 8026
rect 18432 8022 18460 8434
rect 18524 8294 18552 8463
rect 18512 8288 18564 8294
rect 18512 8230 18564 8236
rect 18420 8016 18472 8022
rect 18420 7958 18472 7964
rect 18328 7472 18380 7478
rect 18050 7440 18106 7449
rect 18328 7414 18380 7420
rect 18050 7375 18106 7384
rect 17038 7304 17094 7313
rect 17038 7239 17094 7248
rect 16948 6656 17000 6662
rect 16948 6598 17000 6604
rect 16544 6556 16852 6565
rect 16544 6554 16550 6556
rect 16606 6554 16630 6556
rect 16686 6554 16710 6556
rect 16766 6554 16790 6556
rect 16846 6554 16852 6556
rect 16606 6502 16608 6554
rect 16788 6502 16790 6554
rect 16544 6500 16550 6502
rect 16606 6500 16630 6502
rect 16686 6500 16710 6502
rect 16766 6500 16790 6502
rect 16846 6500 16852 6502
rect 16544 6491 16852 6500
rect 16396 5636 16448 5642
rect 16396 5578 16448 5584
rect 16212 4752 16264 4758
rect 16212 4694 16264 4700
rect 16120 4684 16172 4690
rect 16120 4626 16172 4632
rect 16132 4282 16160 4626
rect 16120 4276 16172 4282
rect 16120 4218 16172 4224
rect 15384 4140 15436 4146
rect 15384 4082 15436 4088
rect 16132 3738 16160 4218
rect 16408 4196 16436 5578
rect 16544 5468 16852 5477
rect 16544 5466 16550 5468
rect 16606 5466 16630 5468
rect 16686 5466 16710 5468
rect 16766 5466 16790 5468
rect 16846 5466 16852 5468
rect 16606 5414 16608 5466
rect 16788 5414 16790 5466
rect 16544 5412 16550 5414
rect 16606 5412 16630 5414
rect 16686 5412 16710 5414
rect 16766 5412 16790 5414
rect 16846 5412 16852 5414
rect 16544 5403 16852 5412
rect 17052 5302 17080 7239
rect 18340 7002 18368 7414
rect 18524 7410 18552 8230
rect 18512 7404 18564 7410
rect 18512 7346 18564 7352
rect 18328 6996 18380 7002
rect 18328 6938 18380 6944
rect 18236 6792 18288 6798
rect 18236 6734 18288 6740
rect 17776 6724 17828 6730
rect 17776 6666 17828 6672
rect 17788 5642 17816 6666
rect 17776 5636 17828 5642
rect 17776 5578 17828 5584
rect 17040 5296 17092 5302
rect 17040 5238 17092 5244
rect 16488 5228 16540 5234
rect 16488 5170 16540 5176
rect 16948 5228 17000 5234
rect 16948 5170 17000 5176
rect 16500 4826 16528 5170
rect 16488 4820 16540 4826
rect 16488 4762 16540 4768
rect 16544 4380 16852 4389
rect 16544 4378 16550 4380
rect 16606 4378 16630 4380
rect 16686 4378 16710 4380
rect 16766 4378 16790 4380
rect 16846 4378 16852 4380
rect 16606 4326 16608 4378
rect 16788 4326 16790 4378
rect 16544 4324 16550 4326
rect 16606 4324 16630 4326
rect 16686 4324 16710 4326
rect 16766 4324 16790 4326
rect 16846 4324 16852 4326
rect 16544 4315 16852 4324
rect 16408 4168 16528 4196
rect 16120 3732 16172 3738
rect 16120 3674 16172 3680
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 15200 3528 15252 3534
rect 15200 3470 15252 3476
rect 13728 3052 13780 3058
rect 13728 2994 13780 3000
rect 13820 2916 13872 2922
rect 13820 2858 13872 2864
rect 13832 800 13860 2858
rect 13945 2748 14253 2757
rect 13945 2746 13951 2748
rect 14007 2746 14031 2748
rect 14087 2746 14111 2748
rect 14167 2746 14191 2748
rect 14247 2746 14253 2748
rect 14007 2694 14009 2746
rect 14189 2694 14191 2746
rect 13945 2692 13951 2694
rect 14007 2692 14031 2694
rect 14087 2692 14111 2694
rect 14167 2692 14191 2694
rect 14247 2692 14253 2694
rect 13945 2683 14253 2692
rect 14292 1442 14320 3470
rect 16500 3398 16528 4168
rect 16764 4140 16816 4146
rect 16764 4082 16816 4088
rect 16776 3641 16804 4082
rect 16960 3942 16988 5170
rect 17788 4729 17816 5578
rect 18144 5024 18196 5030
rect 18144 4966 18196 4972
rect 17774 4720 17830 4729
rect 17774 4655 17830 4664
rect 17040 4480 17092 4486
rect 17040 4422 17092 4428
rect 18052 4480 18104 4486
rect 18052 4422 18104 4428
rect 16948 3936 17000 3942
rect 16948 3878 17000 3884
rect 17052 3738 17080 4422
rect 18064 4185 18092 4422
rect 18050 4176 18106 4185
rect 18050 4111 18106 4120
rect 17960 4004 18012 4010
rect 17960 3946 18012 3952
rect 17040 3732 17092 3738
rect 17040 3674 17092 3680
rect 16762 3632 16818 3641
rect 16762 3567 16818 3576
rect 14648 3392 14700 3398
rect 14648 3334 14700 3340
rect 16396 3392 16448 3398
rect 16396 3334 16448 3340
rect 16488 3392 16540 3398
rect 16488 3334 16540 3340
rect 14660 3194 14688 3334
rect 14648 3188 14700 3194
rect 14648 3130 14700 3136
rect 15752 3120 15804 3126
rect 15566 3088 15622 3097
rect 14660 3058 15240 3074
rect 14648 3052 15240 3058
rect 14700 3046 15240 3052
rect 14648 2994 14700 3000
rect 15212 2774 15240 3046
rect 15752 3062 15804 3068
rect 15566 3023 15568 3032
rect 15620 3023 15622 3032
rect 15568 2994 15620 3000
rect 15658 2952 15714 2961
rect 15658 2887 15714 2896
rect 15212 2746 15332 2774
rect 14924 1760 14976 1766
rect 14924 1702 14976 1708
rect 14556 1556 14608 1562
rect 14556 1498 14608 1504
rect 14200 1414 14320 1442
rect 14200 800 14228 1414
rect 14568 800 14596 1498
rect 14936 800 14964 1702
rect 15304 800 15332 2746
rect 15672 800 15700 2887
rect 15764 1630 15792 3062
rect 16028 1896 16080 1902
rect 16028 1838 16080 1844
rect 15752 1624 15804 1630
rect 15752 1566 15804 1572
rect 16040 800 16068 1838
rect 16408 800 16436 3334
rect 16544 3292 16852 3301
rect 16544 3290 16550 3292
rect 16606 3290 16630 3292
rect 16686 3290 16710 3292
rect 16766 3290 16790 3292
rect 16846 3290 16852 3292
rect 16606 3238 16608 3290
rect 16788 3238 16790 3290
rect 16544 3236 16550 3238
rect 16606 3236 16630 3238
rect 16686 3236 16710 3238
rect 16766 3236 16790 3238
rect 16846 3236 16852 3238
rect 16544 3227 16852 3236
rect 17132 3188 17184 3194
rect 17132 3130 17184 3136
rect 17040 2916 17092 2922
rect 17040 2858 17092 2864
rect 16948 2848 17000 2854
rect 16948 2790 17000 2796
rect 16544 2204 16852 2213
rect 16544 2202 16550 2204
rect 16606 2202 16630 2204
rect 16686 2202 16710 2204
rect 16766 2202 16790 2204
rect 16846 2202 16852 2204
rect 16606 2150 16608 2202
rect 16788 2150 16790 2202
rect 16544 2148 16550 2150
rect 16606 2148 16630 2150
rect 16686 2148 16710 2150
rect 16766 2148 16790 2150
rect 16846 2148 16852 2150
rect 16544 2139 16852 2148
rect 16960 1442 16988 2790
rect 16776 1414 16988 1442
rect 17052 1442 17080 2858
rect 17144 2650 17172 3130
rect 17972 3126 18000 3946
rect 18064 3534 18092 4111
rect 18052 3528 18104 3534
rect 18156 3505 18184 4966
rect 18248 4010 18276 6734
rect 18340 6458 18368 6938
rect 18328 6452 18380 6458
rect 18328 6394 18380 6400
rect 18340 5914 18368 6394
rect 18328 5908 18380 5914
rect 18328 5850 18380 5856
rect 18340 5370 18368 5850
rect 18328 5364 18380 5370
rect 18328 5306 18380 5312
rect 18604 5296 18656 5302
rect 18604 5238 18656 5244
rect 18236 4004 18288 4010
rect 18236 3946 18288 3952
rect 18328 3596 18380 3602
rect 18328 3538 18380 3544
rect 18052 3470 18104 3476
rect 18142 3496 18198 3505
rect 18142 3431 18198 3440
rect 17960 3120 18012 3126
rect 17960 3062 18012 3068
rect 17776 3052 17828 3058
rect 17776 2994 17828 3000
rect 17788 2650 17816 2994
rect 17132 2644 17184 2650
rect 17132 2586 17184 2592
rect 17776 2644 17828 2650
rect 17776 2586 17828 2592
rect 18156 2378 18184 3431
rect 18340 3194 18368 3538
rect 18328 3188 18380 3194
rect 18328 3130 18380 3136
rect 18340 3058 18368 3130
rect 18328 3052 18380 3058
rect 18328 2994 18380 3000
rect 18234 2408 18290 2417
rect 18144 2372 18196 2378
rect 18234 2343 18290 2352
rect 18144 2314 18196 2320
rect 17500 2304 17552 2310
rect 17500 2246 17552 2252
rect 17052 1414 17172 1442
rect 16776 800 16804 1414
rect 17144 800 17172 1414
rect 17512 800 17540 2246
rect 17866 1864 17922 1873
rect 17866 1799 17922 1808
rect 17880 800 17908 1799
rect 18248 800 18276 2343
rect 18616 800 18644 5238
rect 18788 4276 18840 4282
rect 18788 4218 18840 4224
rect 18800 3058 18828 4218
rect 18788 3052 18840 3058
rect 18788 2994 18840 3000
rect 18800 2106 18828 2994
rect 18788 2100 18840 2106
rect 18788 2042 18840 2048
rect 18984 800 19012 8774
rect 19143 8188 19451 8197
rect 19143 8186 19149 8188
rect 19205 8186 19229 8188
rect 19285 8186 19309 8188
rect 19365 8186 19389 8188
rect 19445 8186 19451 8188
rect 19205 8134 19207 8186
rect 19387 8134 19389 8186
rect 19143 8132 19149 8134
rect 19205 8132 19229 8134
rect 19285 8132 19309 8134
rect 19365 8132 19389 8134
rect 19445 8132 19451 8134
rect 19143 8123 19451 8132
rect 19062 7984 19118 7993
rect 19062 7919 19118 7928
rect 19076 6440 19104 7919
rect 19536 7834 19564 10526
rect 19812 10062 19840 10678
rect 20640 10674 20668 11494
rect 20720 11348 20772 11354
rect 20720 11290 20772 11296
rect 20628 10668 20680 10674
rect 20628 10610 20680 10616
rect 19982 10568 20038 10577
rect 19982 10503 19984 10512
rect 20036 10503 20038 10512
rect 19984 10474 20036 10480
rect 19800 10056 19852 10062
rect 19800 9998 19852 10004
rect 19996 9654 20024 10474
rect 20626 10024 20682 10033
rect 20626 9959 20682 9968
rect 20640 9926 20668 9959
rect 20628 9920 20680 9926
rect 20628 9862 20680 9868
rect 19984 9648 20036 9654
rect 19984 9590 20036 9596
rect 19798 9072 19854 9081
rect 19798 9007 19854 9016
rect 19444 7806 19564 7834
rect 19616 7812 19668 7818
rect 19444 7750 19472 7806
rect 19616 7754 19668 7760
rect 19432 7744 19484 7750
rect 19432 7686 19484 7692
rect 19524 7200 19576 7206
rect 19524 7142 19576 7148
rect 19143 7100 19451 7109
rect 19143 7098 19149 7100
rect 19205 7098 19229 7100
rect 19285 7098 19309 7100
rect 19365 7098 19389 7100
rect 19445 7098 19451 7100
rect 19205 7046 19207 7098
rect 19387 7046 19389 7098
rect 19143 7044 19149 7046
rect 19205 7044 19229 7046
rect 19285 7044 19309 7046
rect 19365 7044 19389 7046
rect 19445 7044 19451 7046
rect 19143 7035 19451 7044
rect 19536 7002 19564 7142
rect 19524 6996 19576 7002
rect 19524 6938 19576 6944
rect 19628 6882 19656 7754
rect 19536 6854 19656 6882
rect 19156 6452 19208 6458
rect 19076 6412 19156 6440
rect 19076 5710 19104 6412
rect 19156 6394 19208 6400
rect 19536 6322 19564 6854
rect 19812 6798 19840 9007
rect 19984 8968 20036 8974
rect 19984 8910 20036 8916
rect 19996 8498 20024 8910
rect 20732 8906 20760 11290
rect 21100 9926 21128 11698
rect 21376 11354 21404 11698
rect 21364 11348 21416 11354
rect 21364 11290 21416 11296
rect 21376 10674 21404 11290
rect 21364 10668 21416 10674
rect 21364 10610 21416 10616
rect 21376 10266 21404 10610
rect 21364 10260 21416 10266
rect 21364 10202 21416 10208
rect 21088 9920 21140 9926
rect 21088 9862 21140 9868
rect 21376 9722 21404 10202
rect 21364 9716 21416 9722
rect 21364 9658 21416 9664
rect 21376 9042 21404 9658
rect 21364 9036 21416 9042
rect 21364 8978 21416 8984
rect 20720 8900 20772 8906
rect 20720 8842 20772 8848
rect 21468 8634 21496 16594
rect 21742 16348 22050 16357
rect 21742 16346 21748 16348
rect 21804 16346 21828 16348
rect 21884 16346 21908 16348
rect 21964 16346 21988 16348
rect 22044 16346 22050 16348
rect 21804 16294 21806 16346
rect 21986 16294 21988 16346
rect 21742 16292 21748 16294
rect 21804 16292 21828 16294
rect 21884 16292 21908 16294
rect 21964 16292 21988 16294
rect 22044 16292 22050 16294
rect 21742 16283 22050 16292
rect 21742 15260 22050 15269
rect 21742 15258 21748 15260
rect 21804 15258 21828 15260
rect 21884 15258 21908 15260
rect 21964 15258 21988 15260
rect 22044 15258 22050 15260
rect 21804 15206 21806 15258
rect 21986 15206 21988 15258
rect 21742 15204 21748 15206
rect 21804 15204 21828 15206
rect 21884 15204 21908 15206
rect 21964 15204 21988 15206
rect 22044 15204 22050 15206
rect 21742 15195 22050 15204
rect 21742 14172 22050 14181
rect 21742 14170 21748 14172
rect 21804 14170 21828 14172
rect 21884 14170 21908 14172
rect 21964 14170 21988 14172
rect 22044 14170 22050 14172
rect 21804 14118 21806 14170
rect 21986 14118 21988 14170
rect 21742 14116 21748 14118
rect 21804 14116 21828 14118
rect 21884 14116 21908 14118
rect 21964 14116 21988 14118
rect 22044 14116 22050 14118
rect 21742 14107 22050 14116
rect 21742 13084 22050 13093
rect 21742 13082 21748 13084
rect 21804 13082 21828 13084
rect 21884 13082 21908 13084
rect 21964 13082 21988 13084
rect 22044 13082 22050 13084
rect 21804 13030 21806 13082
rect 21986 13030 21988 13082
rect 21742 13028 21748 13030
rect 21804 13028 21828 13030
rect 21884 13028 21908 13030
rect 21964 13028 21988 13030
rect 22044 13028 22050 13030
rect 21742 13019 22050 13028
rect 21742 11996 22050 12005
rect 21742 11994 21748 11996
rect 21804 11994 21828 11996
rect 21884 11994 21908 11996
rect 21964 11994 21988 11996
rect 22044 11994 22050 11996
rect 21804 11942 21806 11994
rect 21986 11942 21988 11994
rect 21742 11940 21748 11942
rect 21804 11940 21828 11942
rect 21884 11940 21908 11942
rect 21964 11940 21988 11942
rect 22044 11940 22050 11942
rect 21742 11931 22050 11940
rect 21742 10908 22050 10917
rect 21742 10906 21748 10908
rect 21804 10906 21828 10908
rect 21884 10906 21908 10908
rect 21964 10906 21988 10908
rect 22044 10906 22050 10908
rect 21804 10854 21806 10906
rect 21986 10854 21988 10906
rect 21742 10852 21748 10854
rect 21804 10852 21828 10854
rect 21884 10852 21908 10854
rect 21964 10852 21988 10854
rect 22044 10852 22050 10854
rect 21742 10843 22050 10852
rect 21742 9820 22050 9829
rect 21742 9818 21748 9820
rect 21804 9818 21828 9820
rect 21884 9818 21908 9820
rect 21964 9818 21988 9820
rect 22044 9818 22050 9820
rect 21804 9766 21806 9818
rect 21986 9766 21988 9818
rect 21742 9764 21748 9766
rect 21804 9764 21828 9766
rect 21884 9764 21908 9766
rect 21964 9764 21988 9766
rect 22044 9764 22050 9766
rect 21742 9755 22050 9764
rect 21742 8732 22050 8741
rect 21742 8730 21748 8732
rect 21804 8730 21828 8732
rect 21884 8730 21908 8732
rect 21964 8730 21988 8732
rect 22044 8730 22050 8732
rect 21804 8678 21806 8730
rect 21986 8678 21988 8730
rect 21742 8676 21748 8678
rect 21804 8676 21828 8678
rect 21884 8676 21908 8678
rect 21964 8676 21988 8678
rect 22044 8676 22050 8678
rect 21742 8667 22050 8676
rect 21456 8628 21508 8634
rect 21456 8570 21508 8576
rect 19984 8492 20036 8498
rect 19984 8434 20036 8440
rect 19996 8090 20024 8434
rect 20720 8288 20772 8294
rect 20720 8230 20772 8236
rect 19984 8084 20036 8090
rect 19984 8026 20036 8032
rect 20628 7744 20680 7750
rect 20628 7686 20680 7692
rect 20640 6905 20668 7686
rect 20732 7546 20760 8230
rect 21088 8084 21140 8090
rect 21088 8026 21140 8032
rect 21100 7546 21128 8026
rect 21742 7644 22050 7653
rect 21742 7642 21748 7644
rect 21804 7642 21828 7644
rect 21884 7642 21908 7644
rect 21964 7642 21988 7644
rect 22044 7642 22050 7644
rect 21804 7590 21806 7642
rect 21986 7590 21988 7642
rect 21742 7588 21748 7590
rect 21804 7588 21828 7590
rect 21884 7588 21908 7590
rect 21964 7588 21988 7590
rect 22044 7588 22050 7590
rect 21742 7579 22050 7588
rect 20720 7540 20772 7546
rect 20720 7482 20772 7488
rect 21088 7540 21140 7546
rect 21088 7482 21140 7488
rect 21100 7002 21128 7482
rect 21088 6996 21140 7002
rect 21088 6938 21140 6944
rect 20626 6896 20682 6905
rect 20682 6854 20852 6882
rect 20626 6831 20682 6840
rect 19800 6792 19852 6798
rect 19800 6734 19852 6740
rect 19708 6656 19760 6662
rect 19708 6598 19760 6604
rect 19720 6322 19748 6598
rect 19524 6316 19576 6322
rect 19524 6258 19576 6264
rect 19708 6316 19760 6322
rect 19708 6258 19760 6264
rect 19143 6012 19451 6021
rect 19143 6010 19149 6012
rect 19205 6010 19229 6012
rect 19285 6010 19309 6012
rect 19365 6010 19389 6012
rect 19445 6010 19451 6012
rect 19205 5958 19207 6010
rect 19387 5958 19389 6010
rect 19143 5956 19149 5958
rect 19205 5956 19229 5958
rect 19285 5956 19309 5958
rect 19365 5956 19389 5958
rect 19445 5956 19451 5958
rect 19143 5947 19451 5956
rect 19812 5914 19840 6734
rect 19800 5908 19852 5914
rect 19800 5850 19852 5856
rect 19708 5840 19760 5846
rect 19760 5788 19840 5794
rect 19708 5782 19840 5788
rect 19720 5766 19840 5782
rect 19064 5704 19116 5710
rect 19064 5646 19116 5652
rect 19708 5636 19760 5642
rect 19708 5578 19760 5584
rect 19720 5370 19748 5578
rect 19708 5364 19760 5370
rect 19708 5306 19760 5312
rect 19143 4924 19451 4933
rect 19143 4922 19149 4924
rect 19205 4922 19229 4924
rect 19285 4922 19309 4924
rect 19365 4922 19389 4924
rect 19445 4922 19451 4924
rect 19205 4870 19207 4922
rect 19387 4870 19389 4922
rect 19143 4868 19149 4870
rect 19205 4868 19229 4870
rect 19285 4868 19309 4870
rect 19365 4868 19389 4870
rect 19445 4868 19451 4870
rect 19143 4859 19451 4868
rect 19616 4684 19668 4690
rect 19616 4626 19668 4632
rect 19524 4548 19576 4554
rect 19524 4490 19576 4496
rect 19064 4140 19116 4146
rect 19064 4082 19116 4088
rect 19076 3126 19104 4082
rect 19143 3836 19451 3845
rect 19143 3834 19149 3836
rect 19205 3834 19229 3836
rect 19285 3834 19309 3836
rect 19365 3834 19389 3836
rect 19445 3834 19451 3836
rect 19205 3782 19207 3834
rect 19387 3782 19389 3834
rect 19143 3780 19149 3782
rect 19205 3780 19229 3782
rect 19285 3780 19309 3782
rect 19365 3780 19389 3782
rect 19445 3780 19451 3782
rect 19143 3771 19451 3780
rect 19536 3466 19564 4490
rect 19628 4146 19656 4626
rect 19616 4140 19668 4146
rect 19616 4082 19668 4088
rect 19628 3738 19656 4082
rect 19616 3732 19668 3738
rect 19616 3674 19668 3680
rect 19812 3534 19840 5766
rect 20720 5296 20772 5302
rect 20720 5238 20772 5244
rect 19984 4616 20036 4622
rect 19984 4558 20036 4564
rect 19996 4282 20024 4558
rect 19984 4276 20036 4282
rect 19984 4218 20036 4224
rect 20628 3596 20680 3602
rect 20628 3538 20680 3544
rect 19800 3528 19852 3534
rect 19800 3470 19852 3476
rect 19524 3460 19576 3466
rect 19524 3402 19576 3408
rect 19064 3120 19116 3126
rect 19064 3062 19116 3068
rect 20352 3052 20404 3058
rect 20352 2994 20404 3000
rect 19800 2848 19852 2854
rect 19800 2790 19852 2796
rect 19143 2748 19451 2757
rect 19143 2746 19149 2748
rect 19205 2746 19229 2748
rect 19285 2746 19309 2748
rect 19365 2746 19389 2748
rect 19445 2746 19451 2748
rect 19205 2694 19207 2746
rect 19387 2694 19389 2746
rect 19143 2692 19149 2694
rect 19205 2692 19229 2694
rect 19285 2692 19309 2694
rect 19365 2692 19389 2694
rect 19445 2692 19451 2694
rect 19143 2683 19451 2692
rect 19340 2440 19392 2446
rect 19340 2382 19392 2388
rect 19352 2038 19380 2382
rect 19812 2122 19840 2790
rect 20364 2650 20392 2994
rect 20640 2990 20668 3538
rect 20628 2984 20680 2990
rect 20628 2926 20680 2932
rect 20640 2650 20668 2926
rect 20352 2644 20404 2650
rect 20352 2586 20404 2592
rect 20628 2644 20680 2650
rect 20628 2586 20680 2592
rect 20640 2446 20668 2586
rect 20732 2582 20760 5238
rect 20824 4146 20852 6854
rect 21100 6458 21128 6938
rect 21742 6556 22050 6565
rect 21742 6554 21748 6556
rect 21804 6554 21828 6556
rect 21884 6554 21908 6556
rect 21964 6554 21988 6556
rect 22044 6554 22050 6556
rect 21804 6502 21806 6554
rect 21986 6502 21988 6554
rect 21742 6500 21748 6502
rect 21804 6500 21828 6502
rect 21884 6500 21908 6502
rect 21964 6500 21988 6502
rect 22044 6500 22050 6502
rect 21742 6491 22050 6500
rect 21088 6452 21140 6458
rect 21088 6394 21140 6400
rect 21100 5914 21128 6394
rect 21088 5908 21140 5914
rect 21088 5850 21140 5856
rect 21100 5234 21128 5850
rect 21742 5468 22050 5477
rect 21742 5466 21748 5468
rect 21804 5466 21828 5468
rect 21884 5466 21908 5468
rect 21964 5466 21988 5468
rect 22044 5466 22050 5468
rect 21804 5414 21806 5466
rect 21986 5414 21988 5466
rect 21742 5412 21748 5414
rect 21804 5412 21828 5414
rect 21884 5412 21908 5414
rect 21964 5412 21988 5414
rect 22044 5412 22050 5414
rect 21742 5403 22050 5412
rect 21088 5228 21140 5234
rect 21088 5170 21140 5176
rect 21100 4826 21128 5170
rect 21088 4820 21140 4826
rect 21088 4762 21140 4768
rect 21742 4380 22050 4389
rect 21742 4378 21748 4380
rect 21804 4378 21828 4380
rect 21884 4378 21908 4380
rect 21964 4378 21988 4380
rect 22044 4378 22050 4380
rect 21804 4326 21806 4378
rect 21986 4326 21988 4378
rect 21742 4324 21748 4326
rect 21804 4324 21828 4326
rect 21884 4324 21908 4326
rect 21964 4324 21988 4326
rect 22044 4324 22050 4326
rect 21742 4315 22050 4324
rect 20812 4140 20864 4146
rect 20812 4082 20864 4088
rect 21742 3292 22050 3301
rect 21742 3290 21748 3292
rect 21804 3290 21828 3292
rect 21884 3290 21908 3292
rect 21964 3290 21988 3292
rect 22044 3290 22050 3292
rect 21804 3238 21806 3290
rect 21986 3238 21988 3290
rect 21742 3236 21748 3238
rect 21804 3236 21828 3238
rect 21884 3236 21908 3238
rect 21964 3236 21988 3238
rect 22044 3236 22050 3238
rect 21742 3227 22050 3236
rect 20812 3052 20864 3058
rect 20812 2994 20864 3000
rect 20720 2576 20772 2582
rect 20718 2544 20720 2553
rect 20772 2544 20774 2553
rect 20718 2479 20774 2488
rect 20628 2440 20680 2446
rect 20628 2382 20680 2388
rect 20444 2304 20496 2310
rect 20444 2246 20496 2252
rect 19720 2094 19840 2122
rect 19340 2032 19392 2038
rect 19340 1974 19392 1980
rect 19338 1728 19394 1737
rect 19338 1663 19394 1672
rect 19352 800 19380 1663
rect 19720 800 19748 2094
rect 20076 2032 20128 2038
rect 20076 1974 20128 1980
rect 20088 800 20116 1974
rect 20456 800 20484 2246
rect 20824 800 20852 2994
rect 21742 2204 22050 2213
rect 21742 2202 21748 2204
rect 21804 2202 21828 2204
rect 21884 2202 21908 2204
rect 21964 2202 21988 2204
rect 22044 2202 22050 2204
rect 21804 2150 21806 2202
rect 21986 2150 21988 2202
rect 21742 2148 21748 2150
rect 21804 2148 21828 2150
rect 21884 2148 21908 2150
rect 21964 2148 21988 2150
rect 22044 2148 22050 2150
rect 21742 2139 22050 2148
rect 11716 734 11928 762
rect 11978 0 12034 800
rect 12346 0 12402 800
rect 12714 0 12770 800
rect 13082 0 13138 800
rect 13450 0 13506 800
rect 13818 0 13874 800
rect 14186 0 14242 800
rect 14554 0 14610 800
rect 14922 0 14978 800
rect 15290 0 15346 800
rect 15658 0 15714 800
rect 16026 0 16082 800
rect 16394 0 16450 800
rect 16762 0 16818 800
rect 17130 0 17186 800
rect 17498 0 17554 800
rect 17866 0 17922 800
rect 18234 0 18290 800
rect 18602 0 18658 800
rect 18970 0 19026 800
rect 19338 0 19394 800
rect 19706 0 19762 800
rect 20074 0 20130 800
rect 20442 0 20498 800
rect 20810 0 20866 800
<< via2 >>
rect 2962 21256 3018 21312
rect 3882 20848 3938 20904
rect 4066 20440 4122 20496
rect 3555 20154 3611 20156
rect 3635 20154 3691 20156
rect 3715 20154 3771 20156
rect 3795 20154 3851 20156
rect 3555 20102 3601 20154
rect 3601 20102 3611 20154
rect 3635 20102 3665 20154
rect 3665 20102 3677 20154
rect 3677 20102 3691 20154
rect 3715 20102 3729 20154
rect 3729 20102 3741 20154
rect 3741 20102 3771 20154
rect 3795 20102 3805 20154
rect 3805 20102 3851 20154
rect 3555 20100 3611 20102
rect 3635 20100 3691 20102
rect 3715 20100 3771 20102
rect 3795 20100 3851 20102
rect 3238 20032 3294 20088
rect 4158 19624 4214 19680
rect 4066 19216 4122 19272
rect 3555 19066 3611 19068
rect 3635 19066 3691 19068
rect 3715 19066 3771 19068
rect 3795 19066 3851 19068
rect 3555 19014 3601 19066
rect 3601 19014 3611 19066
rect 3635 19014 3665 19066
rect 3665 19014 3677 19066
rect 3677 19014 3691 19066
rect 3715 19014 3729 19066
rect 3729 19014 3741 19066
rect 3741 19014 3771 19066
rect 3795 19014 3805 19066
rect 3805 19014 3851 19066
rect 3555 19012 3611 19014
rect 3635 19012 3691 19014
rect 3715 19012 3771 19014
rect 3795 19012 3851 19014
rect 3974 18400 4030 18456
rect 4158 18808 4214 18864
rect 1950 17992 2006 18048
rect 3555 17978 3611 17980
rect 3635 17978 3691 17980
rect 3715 17978 3771 17980
rect 3795 17978 3851 17980
rect 3555 17926 3601 17978
rect 3601 17926 3611 17978
rect 3635 17926 3665 17978
rect 3665 17926 3677 17978
rect 3677 17926 3691 17978
rect 3715 17926 3729 17978
rect 3729 17926 3741 17978
rect 3741 17926 3771 17978
rect 3795 17926 3805 17978
rect 3805 17926 3851 17978
rect 3555 17924 3611 17926
rect 3635 17924 3691 17926
rect 3715 17924 3771 17926
rect 3795 17924 3851 17926
rect 3698 17584 3754 17640
rect 1582 17176 1638 17232
rect 3555 16890 3611 16892
rect 3635 16890 3691 16892
rect 3715 16890 3771 16892
rect 3795 16890 3851 16892
rect 3555 16838 3601 16890
rect 3601 16838 3611 16890
rect 3635 16838 3665 16890
rect 3665 16838 3677 16890
rect 3677 16838 3691 16890
rect 3715 16838 3729 16890
rect 3729 16838 3741 16890
rect 3741 16838 3771 16890
rect 3795 16838 3805 16890
rect 3805 16838 3851 16890
rect 3555 16836 3611 16838
rect 3635 16836 3691 16838
rect 3715 16836 3771 16838
rect 3795 16836 3851 16838
rect 1950 16768 2006 16824
rect 1674 16360 1730 16416
rect 2778 15952 2834 16008
rect 3555 15802 3611 15804
rect 3635 15802 3691 15804
rect 3715 15802 3771 15804
rect 3795 15802 3851 15804
rect 3555 15750 3601 15802
rect 3601 15750 3611 15802
rect 3635 15750 3665 15802
rect 3665 15750 3677 15802
rect 3677 15750 3691 15802
rect 3715 15750 3729 15802
rect 3729 15750 3741 15802
rect 3741 15750 3771 15802
rect 3795 15750 3805 15802
rect 3805 15750 3851 15802
rect 3555 15748 3611 15750
rect 3635 15748 3691 15750
rect 3715 15748 3771 15750
rect 3795 15748 3851 15750
rect 2226 15580 2228 15600
rect 2228 15580 2280 15600
rect 2280 15580 2282 15600
rect 2226 15544 2282 15580
rect 1490 15136 1546 15192
rect 1950 14764 1952 14784
rect 1952 14764 2004 14784
rect 2004 14764 2006 14784
rect 1950 14728 2006 14764
rect 3555 14714 3611 14716
rect 3635 14714 3691 14716
rect 3715 14714 3771 14716
rect 3795 14714 3851 14716
rect 3555 14662 3601 14714
rect 3601 14662 3611 14714
rect 3635 14662 3665 14714
rect 3665 14662 3677 14714
rect 3677 14662 3691 14714
rect 3715 14662 3729 14714
rect 3729 14662 3741 14714
rect 3741 14662 3771 14714
rect 3795 14662 3805 14714
rect 3805 14662 3851 14714
rect 3555 14660 3611 14662
rect 3635 14660 3691 14662
rect 3715 14660 3771 14662
rect 3795 14660 3851 14662
rect 1950 14320 2006 14376
rect 2778 13912 2834 13968
rect 1490 4936 1546 4992
rect 1398 4528 1454 4584
rect 1674 13096 1730 13152
rect 2778 13504 2834 13560
rect 1950 11872 2006 11928
rect 1674 6604 1676 6624
rect 1676 6604 1728 6624
rect 1728 6604 1730 6624
rect 1674 6568 1730 6604
rect 1674 5752 1730 5808
rect 1582 3712 1638 3768
rect 1398 2896 1454 2952
rect 1214 1672 1270 1728
rect 1858 4528 1914 4584
rect 2042 7268 2098 7304
rect 2042 7248 2044 7268
rect 2044 7248 2096 7268
rect 2096 7248 2098 7268
rect 2778 12688 2834 12744
rect 2686 11736 2742 11792
rect 2962 12280 3018 12336
rect 2410 7928 2466 7984
rect 2318 3984 2374 4040
rect 2226 2488 2282 2544
rect 2134 2352 2190 2408
rect 2042 1672 2098 1728
rect 3555 13626 3611 13628
rect 3635 13626 3691 13628
rect 3715 13626 3771 13628
rect 3795 13626 3851 13628
rect 3555 13574 3601 13626
rect 3601 13574 3611 13626
rect 3635 13574 3665 13626
rect 3665 13574 3677 13626
rect 3677 13574 3691 13626
rect 3715 13574 3729 13626
rect 3729 13574 3741 13626
rect 3741 13574 3771 13626
rect 3795 13574 3805 13626
rect 3805 13574 3851 13626
rect 3555 13572 3611 13574
rect 3635 13572 3691 13574
rect 3715 13572 3771 13574
rect 3795 13572 3851 13574
rect 3555 12538 3611 12540
rect 3635 12538 3691 12540
rect 3715 12538 3771 12540
rect 3795 12538 3851 12540
rect 3555 12486 3601 12538
rect 3601 12486 3611 12538
rect 3635 12486 3665 12538
rect 3665 12486 3677 12538
rect 3677 12486 3691 12538
rect 3715 12486 3729 12538
rect 3729 12486 3741 12538
rect 3741 12486 3771 12538
rect 3795 12486 3805 12538
rect 3805 12486 3851 12538
rect 3555 12484 3611 12486
rect 3635 12484 3691 12486
rect 3715 12484 3771 12486
rect 3795 12484 3851 12486
rect 3422 11464 3478 11520
rect 3555 11450 3611 11452
rect 3635 11450 3691 11452
rect 3715 11450 3771 11452
rect 3795 11450 3851 11452
rect 3555 11398 3601 11450
rect 3601 11398 3611 11450
rect 3635 11398 3665 11450
rect 3665 11398 3677 11450
rect 3677 11398 3691 11450
rect 3715 11398 3729 11450
rect 3729 11398 3741 11450
rect 3741 11398 3771 11450
rect 3795 11398 3805 11450
rect 3805 11398 3851 11450
rect 3555 11396 3611 11398
rect 3635 11396 3691 11398
rect 3715 11396 3771 11398
rect 3795 11396 3851 11398
rect 6154 20698 6210 20700
rect 6234 20698 6290 20700
rect 6314 20698 6370 20700
rect 6394 20698 6450 20700
rect 6154 20646 6200 20698
rect 6200 20646 6210 20698
rect 6234 20646 6264 20698
rect 6264 20646 6276 20698
rect 6276 20646 6290 20698
rect 6314 20646 6328 20698
rect 6328 20646 6340 20698
rect 6340 20646 6370 20698
rect 6394 20646 6404 20698
rect 6404 20646 6450 20698
rect 6154 20644 6210 20646
rect 6234 20644 6290 20646
rect 6314 20644 6370 20646
rect 6394 20644 6450 20646
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11398 20698
rect 11398 20646 11408 20698
rect 11432 20646 11462 20698
rect 11462 20646 11474 20698
rect 11474 20646 11488 20698
rect 11512 20646 11526 20698
rect 11526 20646 11538 20698
rect 11538 20646 11568 20698
rect 11592 20646 11602 20698
rect 11602 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 16550 20698 16606 20700
rect 16630 20698 16686 20700
rect 16710 20698 16766 20700
rect 16790 20698 16846 20700
rect 16550 20646 16596 20698
rect 16596 20646 16606 20698
rect 16630 20646 16660 20698
rect 16660 20646 16672 20698
rect 16672 20646 16686 20698
rect 16710 20646 16724 20698
rect 16724 20646 16736 20698
rect 16736 20646 16766 20698
rect 16790 20646 16800 20698
rect 16800 20646 16846 20698
rect 16550 20644 16606 20646
rect 16630 20644 16686 20646
rect 16710 20644 16766 20646
rect 16790 20644 16846 20646
rect 21748 20698 21804 20700
rect 21828 20698 21884 20700
rect 21908 20698 21964 20700
rect 21988 20698 22044 20700
rect 21748 20646 21794 20698
rect 21794 20646 21804 20698
rect 21828 20646 21858 20698
rect 21858 20646 21870 20698
rect 21870 20646 21884 20698
rect 21908 20646 21922 20698
rect 21922 20646 21934 20698
rect 21934 20646 21964 20698
rect 21988 20646 21998 20698
rect 21998 20646 22044 20698
rect 21748 20644 21804 20646
rect 21828 20644 21884 20646
rect 21908 20644 21964 20646
rect 21988 20644 22044 20646
rect 8753 20154 8809 20156
rect 8833 20154 8889 20156
rect 8913 20154 8969 20156
rect 8993 20154 9049 20156
rect 8753 20102 8799 20154
rect 8799 20102 8809 20154
rect 8833 20102 8863 20154
rect 8863 20102 8875 20154
rect 8875 20102 8889 20154
rect 8913 20102 8927 20154
rect 8927 20102 8939 20154
rect 8939 20102 8969 20154
rect 8993 20102 9003 20154
rect 9003 20102 9049 20154
rect 8753 20100 8809 20102
rect 8833 20100 8889 20102
rect 8913 20100 8969 20102
rect 8993 20100 9049 20102
rect 13951 20154 14007 20156
rect 14031 20154 14087 20156
rect 14111 20154 14167 20156
rect 14191 20154 14247 20156
rect 13951 20102 13997 20154
rect 13997 20102 14007 20154
rect 14031 20102 14061 20154
rect 14061 20102 14073 20154
rect 14073 20102 14087 20154
rect 14111 20102 14125 20154
rect 14125 20102 14137 20154
rect 14137 20102 14167 20154
rect 14191 20102 14201 20154
rect 14201 20102 14247 20154
rect 13951 20100 14007 20102
rect 14031 20100 14087 20102
rect 14111 20100 14167 20102
rect 14191 20100 14247 20102
rect 19149 20154 19205 20156
rect 19229 20154 19285 20156
rect 19309 20154 19365 20156
rect 19389 20154 19445 20156
rect 19149 20102 19195 20154
rect 19195 20102 19205 20154
rect 19229 20102 19259 20154
rect 19259 20102 19271 20154
rect 19271 20102 19285 20154
rect 19309 20102 19323 20154
rect 19323 20102 19335 20154
rect 19335 20102 19365 20154
rect 19389 20102 19399 20154
rect 19399 20102 19445 20154
rect 19149 20100 19205 20102
rect 19229 20100 19285 20102
rect 19309 20100 19365 20102
rect 19389 20100 19445 20102
rect 6154 19610 6210 19612
rect 6234 19610 6290 19612
rect 6314 19610 6370 19612
rect 6394 19610 6450 19612
rect 6154 19558 6200 19610
rect 6200 19558 6210 19610
rect 6234 19558 6264 19610
rect 6264 19558 6276 19610
rect 6276 19558 6290 19610
rect 6314 19558 6328 19610
rect 6328 19558 6340 19610
rect 6340 19558 6370 19610
rect 6394 19558 6404 19610
rect 6404 19558 6450 19610
rect 6154 19556 6210 19558
rect 6234 19556 6290 19558
rect 6314 19556 6370 19558
rect 6394 19556 6450 19558
rect 8753 19066 8809 19068
rect 8833 19066 8889 19068
rect 8913 19066 8969 19068
rect 8993 19066 9049 19068
rect 8753 19014 8799 19066
rect 8799 19014 8809 19066
rect 8833 19014 8863 19066
rect 8863 19014 8875 19066
rect 8875 19014 8889 19066
rect 8913 19014 8927 19066
rect 8927 19014 8939 19066
rect 8939 19014 8969 19066
rect 8993 19014 9003 19066
rect 9003 19014 9049 19066
rect 8753 19012 8809 19014
rect 8833 19012 8889 19014
rect 8913 19012 8969 19014
rect 8993 19012 9049 19014
rect 6154 18522 6210 18524
rect 6234 18522 6290 18524
rect 6314 18522 6370 18524
rect 6394 18522 6450 18524
rect 6154 18470 6200 18522
rect 6200 18470 6210 18522
rect 6234 18470 6264 18522
rect 6264 18470 6276 18522
rect 6276 18470 6290 18522
rect 6314 18470 6328 18522
rect 6328 18470 6340 18522
rect 6340 18470 6370 18522
rect 6394 18470 6404 18522
rect 6404 18470 6450 18522
rect 6154 18468 6210 18470
rect 6234 18468 6290 18470
rect 6314 18468 6370 18470
rect 6394 18468 6450 18470
rect 6154 17434 6210 17436
rect 6234 17434 6290 17436
rect 6314 17434 6370 17436
rect 6394 17434 6450 17436
rect 6154 17382 6200 17434
rect 6200 17382 6210 17434
rect 6234 17382 6264 17434
rect 6264 17382 6276 17434
rect 6276 17382 6290 17434
rect 6314 17382 6328 17434
rect 6328 17382 6340 17434
rect 6340 17382 6370 17434
rect 6394 17382 6404 17434
rect 6404 17382 6450 17434
rect 6154 17380 6210 17382
rect 6234 17380 6290 17382
rect 6314 17380 6370 17382
rect 6394 17380 6450 17382
rect 6154 16346 6210 16348
rect 6234 16346 6290 16348
rect 6314 16346 6370 16348
rect 6394 16346 6450 16348
rect 6154 16294 6200 16346
rect 6200 16294 6210 16346
rect 6234 16294 6264 16346
rect 6264 16294 6276 16346
rect 6276 16294 6290 16346
rect 6314 16294 6328 16346
rect 6328 16294 6340 16346
rect 6340 16294 6370 16346
rect 6394 16294 6404 16346
rect 6404 16294 6450 16346
rect 6154 16292 6210 16294
rect 6234 16292 6290 16294
rect 6314 16292 6370 16294
rect 6394 16292 6450 16294
rect 8753 17978 8809 17980
rect 8833 17978 8889 17980
rect 8913 17978 8969 17980
rect 8993 17978 9049 17980
rect 8753 17926 8799 17978
rect 8799 17926 8809 17978
rect 8833 17926 8863 17978
rect 8863 17926 8875 17978
rect 8875 17926 8889 17978
rect 8913 17926 8927 17978
rect 8927 17926 8939 17978
rect 8939 17926 8969 17978
rect 8993 17926 9003 17978
rect 9003 17926 9049 17978
rect 8753 17924 8809 17926
rect 8833 17924 8889 17926
rect 8913 17924 8969 17926
rect 8993 17924 9049 17926
rect 8753 16890 8809 16892
rect 8833 16890 8889 16892
rect 8913 16890 8969 16892
rect 8993 16890 9049 16892
rect 8753 16838 8799 16890
rect 8799 16838 8809 16890
rect 8833 16838 8863 16890
rect 8863 16838 8875 16890
rect 8875 16838 8889 16890
rect 8913 16838 8927 16890
rect 8927 16838 8939 16890
rect 8939 16838 8969 16890
rect 8993 16838 9003 16890
rect 9003 16838 9049 16890
rect 8753 16836 8809 16838
rect 8833 16836 8889 16838
rect 8913 16836 8969 16838
rect 8993 16836 9049 16838
rect 4986 12588 4988 12608
rect 4988 12588 5040 12608
rect 5040 12588 5042 12608
rect 4986 12552 5042 12588
rect 3422 10648 3478 10704
rect 3330 10240 3386 10296
rect 3555 10362 3611 10364
rect 3635 10362 3691 10364
rect 3715 10362 3771 10364
rect 3795 10362 3851 10364
rect 3555 10310 3601 10362
rect 3601 10310 3611 10362
rect 3635 10310 3665 10362
rect 3665 10310 3677 10362
rect 3677 10310 3691 10362
rect 3715 10310 3729 10362
rect 3729 10310 3741 10362
rect 3741 10310 3771 10362
rect 3795 10310 3805 10362
rect 3805 10310 3851 10362
rect 3555 10308 3611 10310
rect 3635 10308 3691 10310
rect 3715 10308 3771 10310
rect 3795 10308 3851 10310
rect 3054 6976 3110 7032
rect 2870 5616 2926 5672
rect 2778 4120 2834 4176
rect 3882 9832 3938 9888
rect 3790 9444 3846 9480
rect 3790 9424 3792 9444
rect 3792 9424 3844 9444
rect 3844 9424 3846 9444
rect 3555 9274 3611 9276
rect 3635 9274 3691 9276
rect 3715 9274 3771 9276
rect 3795 9274 3851 9276
rect 3555 9222 3601 9274
rect 3601 9222 3611 9274
rect 3635 9222 3665 9274
rect 3665 9222 3677 9274
rect 3677 9222 3691 9274
rect 3715 9222 3729 9274
rect 3729 9222 3741 9274
rect 3741 9222 3771 9274
rect 3795 9222 3805 9274
rect 3805 9222 3851 9274
rect 3555 9220 3611 9222
rect 3635 9220 3691 9222
rect 3715 9220 3771 9222
rect 3795 9220 3851 9222
rect 3330 8200 3386 8256
rect 3555 8186 3611 8188
rect 3635 8186 3691 8188
rect 3715 8186 3771 8188
rect 3795 8186 3851 8188
rect 3555 8134 3601 8186
rect 3601 8134 3611 8186
rect 3635 8134 3665 8186
rect 3665 8134 3677 8186
rect 3677 8134 3691 8186
rect 3715 8134 3729 8186
rect 3729 8134 3741 8186
rect 3741 8134 3771 8186
rect 3795 8134 3805 8186
rect 3805 8134 3851 8186
rect 3555 8132 3611 8134
rect 3635 8132 3691 8134
rect 3715 8132 3771 8134
rect 3795 8132 3851 8134
rect 4066 11092 4068 11112
rect 4068 11092 4120 11112
rect 4120 11092 4122 11112
rect 4066 11056 4122 11092
rect 4066 9968 4122 10024
rect 4066 9460 4068 9480
rect 4068 9460 4120 9480
rect 4120 9460 4122 9480
rect 4066 9424 4122 9460
rect 4066 9016 4122 9072
rect 3974 8200 4030 8256
rect 3974 7792 4030 7848
rect 3422 7384 3478 7440
rect 3555 7098 3611 7100
rect 3635 7098 3691 7100
rect 3715 7098 3771 7100
rect 3795 7098 3851 7100
rect 3555 7046 3601 7098
rect 3601 7046 3611 7098
rect 3635 7046 3665 7098
rect 3665 7046 3677 7098
rect 3677 7046 3691 7098
rect 3715 7046 3729 7098
rect 3729 7046 3741 7098
rect 3741 7046 3771 7098
rect 3795 7046 3805 7098
rect 3805 7046 3851 7098
rect 3555 7044 3611 7046
rect 3635 7044 3691 7046
rect 3715 7044 3771 7046
rect 3795 7044 3851 7046
rect 3555 6010 3611 6012
rect 3635 6010 3691 6012
rect 3715 6010 3771 6012
rect 3795 6010 3851 6012
rect 3555 5958 3601 6010
rect 3601 5958 3611 6010
rect 3635 5958 3665 6010
rect 3665 5958 3677 6010
rect 3677 5958 3691 6010
rect 3715 5958 3729 6010
rect 3729 5958 3741 6010
rect 3741 5958 3771 6010
rect 3795 5958 3805 6010
rect 3805 5958 3851 6010
rect 3555 5956 3611 5958
rect 3635 5956 3691 5958
rect 3715 5956 3771 5958
rect 3795 5956 3851 5958
rect 4158 6160 4214 6216
rect 3330 5616 3386 5672
rect 2594 1808 2650 1864
rect 4066 5344 4122 5400
rect 3555 4922 3611 4924
rect 3635 4922 3691 4924
rect 3715 4922 3771 4924
rect 3795 4922 3851 4924
rect 3555 4870 3601 4922
rect 3601 4870 3611 4922
rect 3635 4870 3665 4922
rect 3665 4870 3677 4922
rect 3677 4870 3691 4922
rect 3715 4870 3729 4922
rect 3729 4870 3741 4922
rect 3741 4870 3771 4922
rect 3795 4870 3805 4922
rect 3805 4870 3851 4922
rect 3555 4868 3611 4870
rect 3635 4868 3691 4870
rect 3715 4868 3771 4870
rect 3795 4868 3851 4870
rect 3330 3304 3386 3360
rect 3555 3834 3611 3836
rect 3635 3834 3691 3836
rect 3715 3834 3771 3836
rect 3795 3834 3851 3836
rect 3555 3782 3601 3834
rect 3601 3782 3611 3834
rect 3635 3782 3665 3834
rect 3665 3782 3677 3834
rect 3677 3782 3691 3834
rect 3715 3782 3729 3834
rect 3729 3782 3741 3834
rect 3741 3782 3771 3834
rect 3795 3782 3805 3834
rect 3805 3782 3851 3834
rect 3555 3780 3611 3782
rect 3635 3780 3691 3782
rect 3715 3780 3771 3782
rect 3795 3780 3851 3782
rect 3555 2746 3611 2748
rect 3635 2746 3691 2748
rect 3715 2746 3771 2748
rect 3795 2746 3851 2748
rect 3555 2694 3601 2746
rect 3601 2694 3611 2746
rect 3635 2694 3665 2746
rect 3665 2694 3677 2746
rect 3677 2694 3691 2746
rect 3715 2694 3729 2746
rect 3729 2694 3741 2746
rect 3741 2694 3771 2746
rect 3795 2694 3805 2746
rect 3805 2694 3851 2746
rect 3555 2692 3611 2694
rect 3635 2692 3691 2694
rect 3715 2692 3771 2694
rect 3795 2692 3851 2694
rect 4250 5616 4306 5672
rect 3974 2080 4030 2136
rect 5170 9016 5226 9072
rect 4986 7792 5042 7848
rect 4802 7384 4858 7440
rect 4802 3440 4858 3496
rect 6154 15258 6210 15260
rect 6234 15258 6290 15260
rect 6314 15258 6370 15260
rect 6394 15258 6450 15260
rect 6154 15206 6200 15258
rect 6200 15206 6210 15258
rect 6234 15206 6264 15258
rect 6264 15206 6276 15258
rect 6276 15206 6290 15258
rect 6314 15206 6328 15258
rect 6328 15206 6340 15258
rect 6340 15206 6370 15258
rect 6394 15206 6404 15258
rect 6404 15206 6450 15258
rect 6154 15204 6210 15206
rect 6234 15204 6290 15206
rect 6314 15204 6370 15206
rect 6394 15204 6450 15206
rect 6154 14170 6210 14172
rect 6234 14170 6290 14172
rect 6314 14170 6370 14172
rect 6394 14170 6450 14172
rect 6154 14118 6200 14170
rect 6200 14118 6210 14170
rect 6234 14118 6264 14170
rect 6264 14118 6276 14170
rect 6276 14118 6290 14170
rect 6314 14118 6328 14170
rect 6328 14118 6340 14170
rect 6340 14118 6370 14170
rect 6394 14118 6404 14170
rect 6404 14118 6450 14170
rect 6154 14116 6210 14118
rect 6234 14116 6290 14118
rect 6314 14116 6370 14118
rect 6394 14116 6450 14118
rect 6550 13912 6606 13968
rect 6154 13082 6210 13084
rect 6234 13082 6290 13084
rect 6314 13082 6370 13084
rect 6394 13082 6450 13084
rect 6154 13030 6200 13082
rect 6200 13030 6210 13082
rect 6234 13030 6264 13082
rect 6264 13030 6276 13082
rect 6276 13030 6290 13082
rect 6314 13030 6328 13082
rect 6328 13030 6340 13082
rect 6340 13030 6370 13082
rect 6394 13030 6404 13082
rect 6404 13030 6450 13082
rect 6154 13028 6210 13030
rect 6234 13028 6290 13030
rect 6314 13028 6370 13030
rect 6394 13028 6450 13030
rect 6154 11994 6210 11996
rect 6234 11994 6290 11996
rect 6314 11994 6370 11996
rect 6394 11994 6450 11996
rect 6154 11942 6200 11994
rect 6200 11942 6210 11994
rect 6234 11942 6264 11994
rect 6264 11942 6276 11994
rect 6276 11942 6290 11994
rect 6314 11942 6328 11994
rect 6328 11942 6340 11994
rect 6340 11942 6370 11994
rect 6394 11942 6404 11994
rect 6404 11942 6450 11994
rect 6154 11940 6210 11942
rect 6234 11940 6290 11942
rect 6314 11940 6370 11942
rect 6394 11940 6450 11942
rect 5630 11636 5632 11656
rect 5632 11636 5684 11656
rect 5684 11636 5686 11656
rect 5630 11600 5686 11636
rect 5538 8608 5594 8664
rect 5446 8472 5502 8528
rect 5538 8064 5594 8120
rect 5538 6704 5594 6760
rect 6642 11056 6698 11112
rect 6154 10906 6210 10908
rect 6234 10906 6290 10908
rect 6314 10906 6370 10908
rect 6394 10906 6450 10908
rect 6154 10854 6200 10906
rect 6200 10854 6210 10906
rect 6234 10854 6264 10906
rect 6264 10854 6276 10906
rect 6276 10854 6290 10906
rect 6314 10854 6328 10906
rect 6328 10854 6340 10906
rect 6340 10854 6370 10906
rect 6394 10854 6404 10906
rect 6404 10854 6450 10906
rect 6154 10852 6210 10854
rect 6234 10852 6290 10854
rect 6314 10852 6370 10854
rect 6394 10852 6450 10854
rect 6154 9818 6210 9820
rect 6234 9818 6290 9820
rect 6314 9818 6370 9820
rect 6394 9818 6450 9820
rect 6154 9766 6200 9818
rect 6200 9766 6210 9818
rect 6234 9766 6264 9818
rect 6264 9766 6276 9818
rect 6276 9766 6290 9818
rect 6314 9766 6328 9818
rect 6328 9766 6340 9818
rect 6340 9766 6370 9818
rect 6394 9766 6404 9818
rect 6404 9766 6450 9818
rect 6154 9764 6210 9766
rect 6234 9764 6290 9766
rect 6314 9764 6370 9766
rect 6394 9764 6450 9766
rect 6154 8730 6210 8732
rect 6234 8730 6290 8732
rect 6314 8730 6370 8732
rect 6394 8730 6450 8732
rect 6154 8678 6200 8730
rect 6200 8678 6210 8730
rect 6234 8678 6264 8730
rect 6264 8678 6276 8730
rect 6276 8678 6290 8730
rect 6314 8678 6328 8730
rect 6328 8678 6340 8730
rect 6340 8678 6370 8730
rect 6394 8678 6404 8730
rect 6404 8678 6450 8730
rect 6154 8676 6210 8678
rect 6234 8676 6290 8678
rect 6314 8676 6370 8678
rect 6394 8676 6450 8678
rect 5906 8336 5962 8392
rect 6154 7642 6210 7644
rect 6234 7642 6290 7644
rect 6314 7642 6370 7644
rect 6394 7642 6450 7644
rect 6154 7590 6200 7642
rect 6200 7590 6210 7642
rect 6234 7590 6264 7642
rect 6264 7590 6276 7642
rect 6276 7590 6290 7642
rect 6314 7590 6328 7642
rect 6328 7590 6340 7642
rect 6340 7590 6370 7642
rect 6394 7590 6404 7642
rect 6404 7590 6450 7642
rect 6154 7588 6210 7590
rect 6234 7588 6290 7590
rect 6314 7588 6370 7590
rect 6394 7588 6450 7590
rect 5906 6840 5962 6896
rect 6154 6554 6210 6556
rect 6234 6554 6290 6556
rect 6314 6554 6370 6556
rect 6394 6554 6450 6556
rect 6154 6502 6200 6554
rect 6200 6502 6210 6554
rect 6234 6502 6264 6554
rect 6264 6502 6276 6554
rect 6276 6502 6290 6554
rect 6314 6502 6328 6554
rect 6328 6502 6340 6554
rect 6340 6502 6370 6554
rect 6394 6502 6404 6554
rect 6404 6502 6450 6554
rect 6154 6500 6210 6502
rect 6234 6500 6290 6502
rect 6314 6500 6370 6502
rect 6394 6500 6450 6502
rect 6550 6160 6606 6216
rect 6154 5466 6210 5468
rect 6234 5466 6290 5468
rect 6314 5466 6370 5468
rect 6394 5466 6450 5468
rect 6154 5414 6200 5466
rect 6200 5414 6210 5466
rect 6234 5414 6264 5466
rect 6264 5414 6276 5466
rect 6276 5414 6290 5466
rect 6314 5414 6328 5466
rect 6328 5414 6340 5466
rect 6340 5414 6370 5466
rect 6394 5414 6404 5466
rect 6404 5414 6450 5466
rect 6154 5412 6210 5414
rect 6234 5412 6290 5414
rect 6314 5412 6370 5414
rect 6394 5412 6450 5414
rect 6154 4378 6210 4380
rect 6234 4378 6290 4380
rect 6314 4378 6370 4380
rect 6394 4378 6450 4380
rect 6154 4326 6200 4378
rect 6200 4326 6210 4378
rect 6234 4326 6264 4378
rect 6264 4326 6276 4378
rect 6276 4326 6290 4378
rect 6314 4326 6328 4378
rect 6328 4326 6340 4378
rect 6340 4326 6370 4378
rect 6394 4326 6404 4378
rect 6404 4326 6450 4378
rect 6154 4324 6210 4326
rect 6234 4324 6290 4326
rect 6314 4324 6370 4326
rect 6394 4324 6450 4326
rect 5998 3848 6054 3904
rect 5814 2916 5870 2952
rect 5814 2896 5816 2916
rect 5816 2896 5868 2916
rect 5868 2896 5870 2916
rect 6154 3290 6210 3292
rect 6234 3290 6290 3292
rect 6314 3290 6370 3292
rect 6394 3290 6450 3292
rect 6154 3238 6200 3290
rect 6200 3238 6210 3290
rect 6234 3238 6264 3290
rect 6264 3238 6276 3290
rect 6276 3238 6290 3290
rect 6314 3238 6328 3290
rect 6328 3238 6340 3290
rect 6340 3238 6370 3290
rect 6394 3238 6404 3290
rect 6404 3238 6450 3290
rect 6154 3236 6210 3238
rect 6234 3236 6290 3238
rect 6314 3236 6370 3238
rect 6394 3236 6450 3238
rect 6154 2202 6210 2204
rect 6234 2202 6290 2204
rect 6314 2202 6370 2204
rect 6394 2202 6450 2204
rect 6154 2150 6200 2202
rect 6200 2150 6210 2202
rect 6234 2150 6264 2202
rect 6264 2150 6276 2202
rect 6276 2150 6290 2202
rect 6314 2150 6328 2202
rect 6328 2150 6340 2202
rect 6340 2150 6370 2202
rect 6394 2150 6404 2202
rect 6404 2150 6450 2202
rect 6154 2148 6210 2150
rect 6234 2148 6290 2150
rect 6314 2148 6370 2150
rect 6394 2148 6450 2150
rect 7470 12300 7526 12336
rect 7470 12280 7472 12300
rect 7472 12280 7524 12300
rect 7524 12280 7526 12300
rect 7746 11192 7802 11248
rect 7746 10240 7802 10296
rect 8753 15802 8809 15804
rect 8833 15802 8889 15804
rect 8913 15802 8969 15804
rect 8993 15802 9049 15804
rect 8753 15750 8799 15802
rect 8799 15750 8809 15802
rect 8833 15750 8863 15802
rect 8863 15750 8875 15802
rect 8875 15750 8889 15802
rect 8913 15750 8927 15802
rect 8927 15750 8939 15802
rect 8939 15750 8969 15802
rect 8993 15750 9003 15802
rect 9003 15750 9049 15802
rect 8753 15748 8809 15750
rect 8833 15748 8889 15750
rect 8913 15748 8969 15750
rect 8993 15748 9049 15750
rect 8753 14714 8809 14716
rect 8833 14714 8889 14716
rect 8913 14714 8969 14716
rect 8993 14714 9049 14716
rect 8753 14662 8799 14714
rect 8799 14662 8809 14714
rect 8833 14662 8863 14714
rect 8863 14662 8875 14714
rect 8875 14662 8889 14714
rect 8913 14662 8927 14714
rect 8927 14662 8939 14714
rect 8939 14662 8969 14714
rect 8993 14662 9003 14714
rect 9003 14662 9049 14714
rect 8753 14660 8809 14662
rect 8833 14660 8889 14662
rect 8913 14660 8969 14662
rect 8993 14660 9049 14662
rect 9034 13812 9036 13832
rect 9036 13812 9088 13832
rect 9088 13812 9090 13832
rect 9034 13776 9090 13812
rect 8753 13626 8809 13628
rect 8833 13626 8889 13628
rect 8913 13626 8969 13628
rect 8993 13626 9049 13628
rect 8753 13574 8799 13626
rect 8799 13574 8809 13626
rect 8833 13574 8863 13626
rect 8863 13574 8875 13626
rect 8875 13574 8889 13626
rect 8913 13574 8927 13626
rect 8927 13574 8939 13626
rect 8939 13574 8969 13626
rect 8993 13574 9003 13626
rect 9003 13574 9049 13626
rect 8753 13572 8809 13574
rect 8833 13572 8889 13574
rect 8913 13572 8969 13574
rect 8993 13572 9049 13574
rect 8753 12538 8809 12540
rect 8833 12538 8889 12540
rect 8913 12538 8969 12540
rect 8993 12538 9049 12540
rect 8753 12486 8799 12538
rect 8799 12486 8809 12538
rect 8833 12486 8863 12538
rect 8863 12486 8875 12538
rect 8875 12486 8889 12538
rect 8913 12486 8927 12538
rect 8927 12486 8939 12538
rect 8939 12486 8969 12538
rect 8993 12486 9003 12538
rect 9003 12486 9049 12538
rect 8753 12484 8809 12486
rect 8833 12484 8889 12486
rect 8913 12484 8969 12486
rect 8993 12484 9049 12486
rect 8022 10512 8078 10568
rect 7654 9016 7710 9072
rect 7102 8200 7158 8256
rect 6826 6296 6882 6352
rect 7010 4936 7066 4992
rect 6918 2488 6974 2544
rect 7286 4684 7342 4720
rect 7286 4664 7288 4684
rect 7288 4664 7340 4684
rect 7340 4664 7342 4684
rect 7838 7948 7894 7984
rect 7838 7928 7840 7948
rect 7840 7928 7892 7948
rect 7892 7928 7894 7948
rect 7838 7520 7894 7576
rect 7470 3460 7526 3496
rect 7470 3440 7472 3460
rect 7472 3440 7524 3460
rect 7524 3440 7526 3460
rect 7746 3304 7802 3360
rect 8022 10140 8024 10160
rect 8024 10140 8076 10160
rect 8076 10140 8078 10160
rect 8022 10104 8078 10140
rect 8390 11212 8446 11248
rect 8390 11192 8392 11212
rect 8392 11192 8444 11212
rect 8444 11192 8446 11212
rect 8298 9968 8354 10024
rect 8298 8064 8354 8120
rect 8298 4120 8354 4176
rect 8390 3440 8446 3496
rect 10138 13368 10194 13424
rect 8753 11450 8809 11452
rect 8833 11450 8889 11452
rect 8913 11450 8969 11452
rect 8993 11450 9049 11452
rect 8753 11398 8799 11450
rect 8799 11398 8809 11450
rect 8833 11398 8863 11450
rect 8863 11398 8875 11450
rect 8875 11398 8889 11450
rect 8913 11398 8927 11450
rect 8927 11398 8939 11450
rect 8939 11398 8969 11450
rect 8993 11398 9003 11450
rect 9003 11398 9049 11450
rect 8753 11396 8809 11398
rect 8833 11396 8889 11398
rect 8913 11396 8969 11398
rect 8993 11396 9049 11398
rect 8753 10362 8809 10364
rect 8833 10362 8889 10364
rect 8913 10362 8969 10364
rect 8993 10362 9049 10364
rect 8753 10310 8799 10362
rect 8799 10310 8809 10362
rect 8833 10310 8863 10362
rect 8863 10310 8875 10362
rect 8875 10310 8889 10362
rect 8913 10310 8927 10362
rect 8927 10310 8939 10362
rect 8939 10310 8969 10362
rect 8993 10310 9003 10362
rect 9003 10310 9049 10362
rect 8753 10308 8809 10310
rect 8833 10308 8889 10310
rect 8913 10308 8969 10310
rect 8993 10308 9049 10310
rect 8753 9274 8809 9276
rect 8833 9274 8889 9276
rect 8913 9274 8969 9276
rect 8993 9274 9049 9276
rect 8753 9222 8799 9274
rect 8799 9222 8809 9274
rect 8833 9222 8863 9274
rect 8863 9222 8875 9274
rect 8875 9222 8889 9274
rect 8913 9222 8927 9274
rect 8927 9222 8939 9274
rect 8939 9222 8969 9274
rect 8993 9222 9003 9274
rect 9003 9222 9049 9274
rect 8753 9220 8809 9222
rect 8833 9220 8889 9222
rect 8913 9220 8969 9222
rect 8993 9220 9049 9222
rect 8753 8186 8809 8188
rect 8833 8186 8889 8188
rect 8913 8186 8969 8188
rect 8993 8186 9049 8188
rect 8753 8134 8799 8186
rect 8799 8134 8809 8186
rect 8833 8134 8863 8186
rect 8863 8134 8875 8186
rect 8875 8134 8889 8186
rect 8913 8134 8927 8186
rect 8927 8134 8939 8186
rect 8939 8134 8969 8186
rect 8993 8134 9003 8186
rect 9003 8134 9049 8186
rect 8753 8132 8809 8134
rect 8833 8132 8889 8134
rect 8913 8132 8969 8134
rect 8993 8132 9049 8134
rect 8753 7098 8809 7100
rect 8833 7098 8889 7100
rect 8913 7098 8969 7100
rect 8993 7098 9049 7100
rect 8753 7046 8799 7098
rect 8799 7046 8809 7098
rect 8833 7046 8863 7098
rect 8863 7046 8875 7098
rect 8875 7046 8889 7098
rect 8913 7046 8927 7098
rect 8927 7046 8939 7098
rect 8939 7046 8969 7098
rect 8993 7046 9003 7098
rect 9003 7046 9049 7098
rect 8753 7044 8809 7046
rect 8833 7044 8889 7046
rect 8913 7044 8969 7046
rect 8993 7044 9049 7046
rect 8753 6010 8809 6012
rect 8833 6010 8889 6012
rect 8913 6010 8969 6012
rect 8993 6010 9049 6012
rect 8753 5958 8799 6010
rect 8799 5958 8809 6010
rect 8833 5958 8863 6010
rect 8863 5958 8875 6010
rect 8875 5958 8889 6010
rect 8913 5958 8927 6010
rect 8927 5958 8939 6010
rect 8939 5958 8969 6010
rect 8993 5958 9003 6010
rect 9003 5958 9049 6010
rect 8753 5956 8809 5958
rect 8833 5956 8889 5958
rect 8913 5956 8969 5958
rect 8993 5956 9049 5958
rect 8666 5616 8722 5672
rect 8753 4922 8809 4924
rect 8833 4922 8889 4924
rect 8913 4922 8969 4924
rect 8993 4922 9049 4924
rect 8753 4870 8799 4922
rect 8799 4870 8809 4922
rect 8833 4870 8863 4922
rect 8863 4870 8875 4922
rect 8875 4870 8889 4922
rect 8913 4870 8927 4922
rect 8927 4870 8939 4922
rect 8939 4870 8969 4922
rect 8993 4870 9003 4922
rect 9003 4870 9049 4922
rect 8753 4868 8809 4870
rect 8833 4868 8889 4870
rect 8913 4868 8969 4870
rect 8993 4868 9049 4870
rect 8753 3834 8809 3836
rect 8833 3834 8889 3836
rect 8913 3834 8969 3836
rect 8993 3834 9049 3836
rect 8753 3782 8799 3834
rect 8799 3782 8809 3834
rect 8833 3782 8863 3834
rect 8863 3782 8875 3834
rect 8875 3782 8889 3834
rect 8913 3782 8927 3834
rect 8927 3782 8939 3834
rect 8939 3782 8969 3834
rect 8993 3782 9003 3834
rect 9003 3782 9049 3834
rect 8753 3780 8809 3782
rect 8833 3780 8889 3782
rect 8913 3780 8969 3782
rect 8993 3780 9049 3782
rect 9126 3576 9182 3632
rect 8758 3168 8814 3224
rect 8753 2746 8809 2748
rect 8833 2746 8889 2748
rect 8913 2746 8969 2748
rect 8993 2746 9049 2748
rect 8753 2694 8799 2746
rect 8799 2694 8809 2746
rect 8833 2694 8863 2746
rect 8863 2694 8875 2746
rect 8875 2694 8889 2746
rect 8913 2694 8927 2746
rect 8927 2694 8939 2746
rect 8939 2694 8969 2746
rect 8993 2694 9003 2746
rect 9003 2694 9049 2746
rect 8753 2692 8809 2694
rect 8833 2692 8889 2694
rect 8913 2692 8969 2694
rect 8993 2692 9049 2694
rect 9034 2216 9090 2272
rect 9586 9968 9642 10024
rect 9402 8608 9458 8664
rect 9310 7520 9366 7576
rect 9218 3168 9274 3224
rect 9586 3576 9642 3632
rect 9954 2760 10010 2816
rect 9678 2624 9734 2680
rect 9218 2252 9220 2272
rect 9220 2252 9272 2272
rect 9272 2252 9274 2272
rect 9218 2216 9274 2252
rect 9494 2252 9496 2272
rect 9496 2252 9548 2272
rect 9548 2252 9550 2272
rect 9494 2216 9550 2252
rect 9402 2080 9458 2136
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11398 19610
rect 11398 19558 11408 19610
rect 11432 19558 11462 19610
rect 11462 19558 11474 19610
rect 11474 19558 11488 19610
rect 11512 19558 11526 19610
rect 11526 19558 11538 19610
rect 11538 19558 11568 19610
rect 11592 19558 11602 19610
rect 11602 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 16550 19610 16606 19612
rect 16630 19610 16686 19612
rect 16710 19610 16766 19612
rect 16790 19610 16846 19612
rect 16550 19558 16596 19610
rect 16596 19558 16606 19610
rect 16630 19558 16660 19610
rect 16660 19558 16672 19610
rect 16672 19558 16686 19610
rect 16710 19558 16724 19610
rect 16724 19558 16736 19610
rect 16736 19558 16766 19610
rect 16790 19558 16800 19610
rect 16800 19558 16846 19610
rect 16550 19556 16606 19558
rect 16630 19556 16686 19558
rect 16710 19556 16766 19558
rect 16790 19556 16846 19558
rect 21748 19610 21804 19612
rect 21828 19610 21884 19612
rect 21908 19610 21964 19612
rect 21988 19610 22044 19612
rect 21748 19558 21794 19610
rect 21794 19558 21804 19610
rect 21828 19558 21858 19610
rect 21858 19558 21870 19610
rect 21870 19558 21884 19610
rect 21908 19558 21922 19610
rect 21922 19558 21934 19610
rect 21934 19558 21964 19610
rect 21988 19558 21998 19610
rect 21998 19558 22044 19610
rect 21748 19556 21804 19558
rect 21828 19556 21884 19558
rect 21908 19556 21964 19558
rect 21988 19556 22044 19558
rect 13951 19066 14007 19068
rect 14031 19066 14087 19068
rect 14111 19066 14167 19068
rect 14191 19066 14247 19068
rect 13951 19014 13997 19066
rect 13997 19014 14007 19066
rect 14031 19014 14061 19066
rect 14061 19014 14073 19066
rect 14073 19014 14087 19066
rect 14111 19014 14125 19066
rect 14125 19014 14137 19066
rect 14137 19014 14167 19066
rect 14191 19014 14201 19066
rect 14201 19014 14247 19066
rect 13951 19012 14007 19014
rect 14031 19012 14087 19014
rect 14111 19012 14167 19014
rect 14191 19012 14247 19014
rect 19149 19066 19205 19068
rect 19229 19066 19285 19068
rect 19309 19066 19365 19068
rect 19389 19066 19445 19068
rect 19149 19014 19195 19066
rect 19195 19014 19205 19066
rect 19229 19014 19259 19066
rect 19259 19014 19271 19066
rect 19271 19014 19285 19066
rect 19309 19014 19323 19066
rect 19323 19014 19335 19066
rect 19335 19014 19365 19066
rect 19389 19014 19399 19066
rect 19399 19014 19445 19066
rect 19149 19012 19205 19014
rect 19229 19012 19285 19014
rect 19309 19012 19365 19014
rect 19389 19012 19445 19014
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11398 18522
rect 11398 18470 11408 18522
rect 11432 18470 11462 18522
rect 11462 18470 11474 18522
rect 11474 18470 11488 18522
rect 11512 18470 11526 18522
rect 11526 18470 11538 18522
rect 11538 18470 11568 18522
rect 11592 18470 11602 18522
rect 11602 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 16550 18522 16606 18524
rect 16630 18522 16686 18524
rect 16710 18522 16766 18524
rect 16790 18522 16846 18524
rect 16550 18470 16596 18522
rect 16596 18470 16606 18522
rect 16630 18470 16660 18522
rect 16660 18470 16672 18522
rect 16672 18470 16686 18522
rect 16710 18470 16724 18522
rect 16724 18470 16736 18522
rect 16736 18470 16766 18522
rect 16790 18470 16800 18522
rect 16800 18470 16846 18522
rect 16550 18468 16606 18470
rect 16630 18468 16686 18470
rect 16710 18468 16766 18470
rect 16790 18468 16846 18470
rect 21748 18522 21804 18524
rect 21828 18522 21884 18524
rect 21908 18522 21964 18524
rect 21988 18522 22044 18524
rect 21748 18470 21794 18522
rect 21794 18470 21804 18522
rect 21828 18470 21858 18522
rect 21858 18470 21870 18522
rect 21870 18470 21884 18522
rect 21908 18470 21922 18522
rect 21922 18470 21934 18522
rect 21934 18470 21964 18522
rect 21988 18470 21998 18522
rect 21998 18470 22044 18522
rect 21748 18468 21804 18470
rect 21828 18468 21884 18470
rect 21908 18468 21964 18470
rect 21988 18468 22044 18470
rect 13951 17978 14007 17980
rect 14031 17978 14087 17980
rect 14111 17978 14167 17980
rect 14191 17978 14247 17980
rect 13951 17926 13997 17978
rect 13997 17926 14007 17978
rect 14031 17926 14061 17978
rect 14061 17926 14073 17978
rect 14073 17926 14087 17978
rect 14111 17926 14125 17978
rect 14125 17926 14137 17978
rect 14137 17926 14167 17978
rect 14191 17926 14201 17978
rect 14201 17926 14247 17978
rect 13951 17924 14007 17926
rect 14031 17924 14087 17926
rect 14111 17924 14167 17926
rect 14191 17924 14247 17926
rect 19149 17978 19205 17980
rect 19229 17978 19285 17980
rect 19309 17978 19365 17980
rect 19389 17978 19445 17980
rect 19149 17926 19195 17978
rect 19195 17926 19205 17978
rect 19229 17926 19259 17978
rect 19259 17926 19271 17978
rect 19271 17926 19285 17978
rect 19309 17926 19323 17978
rect 19323 17926 19335 17978
rect 19335 17926 19365 17978
rect 19389 17926 19399 17978
rect 19399 17926 19445 17978
rect 19149 17924 19205 17926
rect 19229 17924 19285 17926
rect 19309 17924 19365 17926
rect 19389 17924 19445 17926
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11398 17434
rect 11398 17382 11408 17434
rect 11432 17382 11462 17434
rect 11462 17382 11474 17434
rect 11474 17382 11488 17434
rect 11512 17382 11526 17434
rect 11526 17382 11538 17434
rect 11538 17382 11568 17434
rect 11592 17382 11602 17434
rect 11602 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 16550 17434 16606 17436
rect 16630 17434 16686 17436
rect 16710 17434 16766 17436
rect 16790 17434 16846 17436
rect 16550 17382 16596 17434
rect 16596 17382 16606 17434
rect 16630 17382 16660 17434
rect 16660 17382 16672 17434
rect 16672 17382 16686 17434
rect 16710 17382 16724 17434
rect 16724 17382 16736 17434
rect 16736 17382 16766 17434
rect 16790 17382 16800 17434
rect 16800 17382 16846 17434
rect 16550 17380 16606 17382
rect 16630 17380 16686 17382
rect 16710 17380 16766 17382
rect 16790 17380 16846 17382
rect 21748 17434 21804 17436
rect 21828 17434 21884 17436
rect 21908 17434 21964 17436
rect 21988 17434 22044 17436
rect 21748 17382 21794 17434
rect 21794 17382 21804 17434
rect 21828 17382 21858 17434
rect 21858 17382 21870 17434
rect 21870 17382 21884 17434
rect 21908 17382 21922 17434
rect 21922 17382 21934 17434
rect 21934 17382 21964 17434
rect 21988 17382 21998 17434
rect 21998 17382 22044 17434
rect 21748 17380 21804 17382
rect 21828 17380 21884 17382
rect 21908 17380 21964 17382
rect 21988 17380 22044 17382
rect 21454 17176 21510 17232
rect 10414 3984 10470 4040
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11398 16346
rect 11398 16294 11408 16346
rect 11432 16294 11462 16346
rect 11462 16294 11474 16346
rect 11474 16294 11488 16346
rect 11512 16294 11526 16346
rect 11526 16294 11538 16346
rect 11538 16294 11568 16346
rect 11592 16294 11602 16346
rect 11602 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11398 15258
rect 11398 15206 11408 15258
rect 11432 15206 11462 15258
rect 11462 15206 11474 15258
rect 11474 15206 11488 15258
rect 11512 15206 11526 15258
rect 11526 15206 11538 15258
rect 11538 15206 11568 15258
rect 11592 15206 11602 15258
rect 11602 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 10598 11192 10654 11248
rect 10598 2624 10654 2680
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11398 14170
rect 11398 14118 11408 14170
rect 11432 14118 11462 14170
rect 11462 14118 11474 14170
rect 11474 14118 11488 14170
rect 11512 14118 11526 14170
rect 11526 14118 11538 14170
rect 11538 14118 11568 14170
rect 11592 14118 11602 14170
rect 11602 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11398 13082
rect 11398 13030 11408 13082
rect 11432 13030 11462 13082
rect 11462 13030 11474 13082
rect 11474 13030 11488 13082
rect 11512 13030 11526 13082
rect 11526 13030 11538 13082
rect 11538 13030 11568 13082
rect 11592 13030 11602 13082
rect 11602 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 10966 11056 11022 11112
rect 10966 7656 11022 7712
rect 10874 5752 10930 5808
rect 11150 7792 11206 7848
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11398 11994
rect 11398 11942 11408 11994
rect 11432 11942 11462 11994
rect 11462 11942 11474 11994
rect 11474 11942 11488 11994
rect 11512 11942 11526 11994
rect 11526 11942 11538 11994
rect 11538 11942 11568 11994
rect 11592 11942 11602 11994
rect 11602 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11398 10906
rect 11398 10854 11408 10906
rect 11432 10854 11462 10906
rect 11462 10854 11474 10906
rect 11474 10854 11488 10906
rect 11512 10854 11526 10906
rect 11526 10854 11538 10906
rect 11538 10854 11568 10906
rect 11592 10854 11602 10906
rect 11602 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11398 9818
rect 11398 9766 11408 9818
rect 11432 9766 11462 9818
rect 11462 9766 11474 9818
rect 11474 9766 11488 9818
rect 11512 9766 11526 9818
rect 11526 9766 11538 9818
rect 11538 9766 11568 9818
rect 11592 9766 11602 9818
rect 11602 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11794 10104 11850 10160
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11398 8730
rect 11398 8678 11408 8730
rect 11432 8678 11462 8730
rect 11462 8678 11474 8730
rect 11474 8678 11488 8730
rect 11512 8678 11526 8730
rect 11526 8678 11538 8730
rect 11538 8678 11568 8730
rect 11592 8678 11602 8730
rect 11602 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11398 7642
rect 11398 7590 11408 7642
rect 11432 7590 11462 7642
rect 11462 7590 11474 7642
rect 11474 7590 11488 7642
rect 11512 7590 11526 7642
rect 11526 7590 11538 7642
rect 11538 7590 11568 7642
rect 11592 7590 11602 7642
rect 11602 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11398 6554
rect 11398 6502 11408 6554
rect 11432 6502 11462 6554
rect 11462 6502 11474 6554
rect 11474 6502 11488 6554
rect 11512 6502 11526 6554
rect 11526 6502 11538 6554
rect 11538 6502 11568 6554
rect 11592 6502 11602 6554
rect 11602 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11398 5466
rect 11398 5414 11408 5466
rect 11432 5414 11462 5466
rect 11462 5414 11474 5466
rect 11474 5414 11488 5466
rect 11512 5414 11526 5466
rect 11526 5414 11538 5466
rect 11538 5414 11568 5466
rect 11592 5414 11602 5466
rect 11602 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 11702 4528 11758 4584
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11398 4378
rect 11398 4326 11408 4378
rect 11432 4326 11462 4378
rect 11462 4326 11474 4378
rect 11474 4326 11488 4378
rect 11512 4326 11526 4378
rect 11526 4326 11538 4378
rect 11538 4326 11568 4378
rect 11592 4326 11602 4378
rect 11602 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11398 3290
rect 11398 3238 11408 3290
rect 11432 3238 11462 3290
rect 11462 3238 11474 3290
rect 11474 3238 11488 3290
rect 11512 3238 11526 3290
rect 11526 3238 11538 3290
rect 11538 3238 11568 3290
rect 11592 3238 11602 3290
rect 11602 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11398 2202
rect 11398 2150 11408 2202
rect 11432 2150 11462 2202
rect 11462 2150 11474 2202
rect 11474 2150 11488 2202
rect 11512 2150 11526 2202
rect 11526 2150 11538 2202
rect 11538 2150 11568 2202
rect 11592 2150 11602 2202
rect 11602 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 13951 16890 14007 16892
rect 14031 16890 14087 16892
rect 14111 16890 14167 16892
rect 14191 16890 14247 16892
rect 13951 16838 13997 16890
rect 13997 16838 14007 16890
rect 14031 16838 14061 16890
rect 14061 16838 14073 16890
rect 14073 16838 14087 16890
rect 14111 16838 14125 16890
rect 14125 16838 14137 16890
rect 14137 16838 14167 16890
rect 14191 16838 14201 16890
rect 14201 16838 14247 16890
rect 13951 16836 14007 16838
rect 14031 16836 14087 16838
rect 14111 16836 14167 16838
rect 14191 16836 14247 16838
rect 19149 16890 19205 16892
rect 19229 16890 19285 16892
rect 19309 16890 19365 16892
rect 19389 16890 19445 16892
rect 19149 16838 19195 16890
rect 19195 16838 19205 16890
rect 19229 16838 19259 16890
rect 19259 16838 19271 16890
rect 19271 16838 19285 16890
rect 19309 16838 19323 16890
rect 19323 16838 19335 16890
rect 19335 16838 19365 16890
rect 19389 16838 19399 16890
rect 19399 16838 19445 16890
rect 19149 16836 19205 16838
rect 19229 16836 19285 16838
rect 19309 16836 19365 16838
rect 19389 16836 19445 16838
rect 16550 16346 16606 16348
rect 16630 16346 16686 16348
rect 16710 16346 16766 16348
rect 16790 16346 16846 16348
rect 16550 16294 16596 16346
rect 16596 16294 16606 16346
rect 16630 16294 16660 16346
rect 16660 16294 16672 16346
rect 16672 16294 16686 16346
rect 16710 16294 16724 16346
rect 16724 16294 16736 16346
rect 16736 16294 16766 16346
rect 16790 16294 16800 16346
rect 16800 16294 16846 16346
rect 16550 16292 16606 16294
rect 16630 16292 16686 16294
rect 16710 16292 16766 16294
rect 16790 16292 16846 16294
rect 13951 15802 14007 15804
rect 14031 15802 14087 15804
rect 14111 15802 14167 15804
rect 14191 15802 14247 15804
rect 13951 15750 13997 15802
rect 13997 15750 14007 15802
rect 14031 15750 14061 15802
rect 14061 15750 14073 15802
rect 14073 15750 14087 15802
rect 14111 15750 14125 15802
rect 14125 15750 14137 15802
rect 14137 15750 14167 15802
rect 14191 15750 14201 15802
rect 14201 15750 14247 15802
rect 13951 15748 14007 15750
rect 14031 15748 14087 15750
rect 14111 15748 14167 15750
rect 14191 15748 14247 15750
rect 19149 15802 19205 15804
rect 19229 15802 19285 15804
rect 19309 15802 19365 15804
rect 19389 15802 19445 15804
rect 19149 15750 19195 15802
rect 19195 15750 19205 15802
rect 19229 15750 19259 15802
rect 19259 15750 19271 15802
rect 19271 15750 19285 15802
rect 19309 15750 19323 15802
rect 19323 15750 19335 15802
rect 19335 15750 19365 15802
rect 19389 15750 19399 15802
rect 19399 15750 19445 15802
rect 19149 15748 19205 15750
rect 19229 15748 19285 15750
rect 19309 15748 19365 15750
rect 19389 15748 19445 15750
rect 16550 15258 16606 15260
rect 16630 15258 16686 15260
rect 16710 15258 16766 15260
rect 16790 15258 16846 15260
rect 16550 15206 16596 15258
rect 16596 15206 16606 15258
rect 16630 15206 16660 15258
rect 16660 15206 16672 15258
rect 16672 15206 16686 15258
rect 16710 15206 16724 15258
rect 16724 15206 16736 15258
rect 16736 15206 16766 15258
rect 16790 15206 16800 15258
rect 16800 15206 16846 15258
rect 16550 15204 16606 15206
rect 16630 15204 16686 15206
rect 16710 15204 16766 15206
rect 16790 15204 16846 15206
rect 13951 14714 14007 14716
rect 14031 14714 14087 14716
rect 14111 14714 14167 14716
rect 14191 14714 14247 14716
rect 13951 14662 13997 14714
rect 13997 14662 14007 14714
rect 14031 14662 14061 14714
rect 14061 14662 14073 14714
rect 14073 14662 14087 14714
rect 14111 14662 14125 14714
rect 14125 14662 14137 14714
rect 14137 14662 14167 14714
rect 14191 14662 14201 14714
rect 14201 14662 14247 14714
rect 13951 14660 14007 14662
rect 14031 14660 14087 14662
rect 14111 14660 14167 14662
rect 14191 14660 14247 14662
rect 12254 11736 12310 11792
rect 13951 13626 14007 13628
rect 14031 13626 14087 13628
rect 14111 13626 14167 13628
rect 14191 13626 14247 13628
rect 13951 13574 13997 13626
rect 13997 13574 14007 13626
rect 14031 13574 14061 13626
rect 14061 13574 14073 13626
rect 14073 13574 14087 13626
rect 14111 13574 14125 13626
rect 14125 13574 14137 13626
rect 14137 13574 14167 13626
rect 14191 13574 14201 13626
rect 14201 13574 14247 13626
rect 13951 13572 14007 13574
rect 14031 13572 14087 13574
rect 14111 13572 14167 13574
rect 14191 13572 14247 13574
rect 13951 12538 14007 12540
rect 14031 12538 14087 12540
rect 14111 12538 14167 12540
rect 14191 12538 14247 12540
rect 13951 12486 13997 12538
rect 13997 12486 14007 12538
rect 14031 12486 14061 12538
rect 14061 12486 14073 12538
rect 14073 12486 14087 12538
rect 14111 12486 14125 12538
rect 14125 12486 14137 12538
rect 14137 12486 14167 12538
rect 14191 12486 14201 12538
rect 14201 12486 14247 12538
rect 13951 12484 14007 12486
rect 14031 12484 14087 12486
rect 14111 12484 14167 12486
rect 14191 12484 14247 12486
rect 19149 14714 19205 14716
rect 19229 14714 19285 14716
rect 19309 14714 19365 14716
rect 19389 14714 19445 14716
rect 19149 14662 19195 14714
rect 19195 14662 19205 14714
rect 19229 14662 19259 14714
rect 19259 14662 19271 14714
rect 19271 14662 19285 14714
rect 19309 14662 19323 14714
rect 19323 14662 19335 14714
rect 19335 14662 19365 14714
rect 19389 14662 19399 14714
rect 19399 14662 19445 14714
rect 19149 14660 19205 14662
rect 19229 14660 19285 14662
rect 19309 14660 19365 14662
rect 19389 14660 19445 14662
rect 16550 14170 16606 14172
rect 16630 14170 16686 14172
rect 16710 14170 16766 14172
rect 16790 14170 16846 14172
rect 16550 14118 16596 14170
rect 16596 14118 16606 14170
rect 16630 14118 16660 14170
rect 16660 14118 16672 14170
rect 16672 14118 16686 14170
rect 16710 14118 16724 14170
rect 16724 14118 16736 14170
rect 16736 14118 16766 14170
rect 16790 14118 16800 14170
rect 16800 14118 16846 14170
rect 16550 14116 16606 14118
rect 16630 14116 16686 14118
rect 16710 14116 16766 14118
rect 16790 14116 16846 14118
rect 19149 13626 19205 13628
rect 19229 13626 19285 13628
rect 19309 13626 19365 13628
rect 19389 13626 19445 13628
rect 19149 13574 19195 13626
rect 19195 13574 19205 13626
rect 19229 13574 19259 13626
rect 19259 13574 19271 13626
rect 19271 13574 19285 13626
rect 19309 13574 19323 13626
rect 19323 13574 19335 13626
rect 19335 13574 19365 13626
rect 19389 13574 19399 13626
rect 19399 13574 19445 13626
rect 19149 13572 19205 13574
rect 19229 13572 19285 13574
rect 19309 13572 19365 13574
rect 19389 13572 19445 13574
rect 19522 13368 19578 13424
rect 16550 13082 16606 13084
rect 16630 13082 16686 13084
rect 16710 13082 16766 13084
rect 16790 13082 16846 13084
rect 16550 13030 16596 13082
rect 16596 13030 16606 13082
rect 16630 13030 16660 13082
rect 16660 13030 16672 13082
rect 16672 13030 16686 13082
rect 16710 13030 16724 13082
rect 16724 13030 16736 13082
rect 16736 13030 16766 13082
rect 16790 13030 16800 13082
rect 16800 13030 16846 13082
rect 16550 13028 16606 13030
rect 16630 13028 16686 13030
rect 16710 13028 16766 13030
rect 16790 13028 16846 13030
rect 13450 11600 13506 11656
rect 13951 11450 14007 11452
rect 14031 11450 14087 11452
rect 14111 11450 14167 11452
rect 14191 11450 14247 11452
rect 13951 11398 13997 11450
rect 13997 11398 14007 11450
rect 14031 11398 14061 11450
rect 14061 11398 14073 11450
rect 14073 11398 14087 11450
rect 14111 11398 14125 11450
rect 14125 11398 14137 11450
rect 14137 11398 14167 11450
rect 14191 11398 14201 11450
rect 14201 11398 14247 11450
rect 13951 11396 14007 11398
rect 14031 11396 14087 11398
rect 14111 11396 14167 11398
rect 14191 11396 14247 11398
rect 14462 11228 14464 11248
rect 14464 11228 14516 11248
rect 14516 11228 14518 11248
rect 14462 11192 14518 11228
rect 16550 11994 16606 11996
rect 16630 11994 16686 11996
rect 16710 11994 16766 11996
rect 16790 11994 16846 11996
rect 16550 11942 16596 11994
rect 16596 11942 16606 11994
rect 16630 11942 16660 11994
rect 16660 11942 16672 11994
rect 16672 11942 16686 11994
rect 16710 11942 16724 11994
rect 16724 11942 16736 11994
rect 16736 11942 16766 11994
rect 16790 11942 16800 11994
rect 16800 11942 16846 11994
rect 16550 11940 16606 11942
rect 16630 11940 16686 11942
rect 16710 11940 16766 11942
rect 16790 11940 16846 11942
rect 13951 10362 14007 10364
rect 14031 10362 14087 10364
rect 14111 10362 14167 10364
rect 14191 10362 14247 10364
rect 13951 10310 13997 10362
rect 13997 10310 14007 10362
rect 14031 10310 14061 10362
rect 14061 10310 14073 10362
rect 14073 10310 14087 10362
rect 14111 10310 14125 10362
rect 14125 10310 14137 10362
rect 14137 10310 14167 10362
rect 14191 10310 14201 10362
rect 14201 10310 14247 10362
rect 13951 10308 14007 10310
rect 14031 10308 14087 10310
rect 14111 10308 14167 10310
rect 14191 10308 14247 10310
rect 14462 9424 14518 9480
rect 13951 9274 14007 9276
rect 14031 9274 14087 9276
rect 14111 9274 14167 9276
rect 14191 9274 14247 9276
rect 13951 9222 13997 9274
rect 13997 9222 14007 9274
rect 14031 9222 14061 9274
rect 14061 9222 14073 9274
rect 14073 9222 14087 9274
rect 14111 9222 14125 9274
rect 14125 9222 14137 9274
rect 14137 9222 14167 9274
rect 14191 9222 14201 9274
rect 14201 9222 14247 9274
rect 13951 9220 14007 9222
rect 14031 9220 14087 9222
rect 14111 9220 14167 9222
rect 14191 9220 14247 9222
rect 14370 8880 14426 8936
rect 13951 8186 14007 8188
rect 14031 8186 14087 8188
rect 14111 8186 14167 8188
rect 14191 8186 14247 8188
rect 13951 8134 13997 8186
rect 13997 8134 14007 8186
rect 14031 8134 14061 8186
rect 14061 8134 14073 8186
rect 14073 8134 14087 8186
rect 14111 8134 14125 8186
rect 14125 8134 14137 8186
rect 14137 8134 14167 8186
rect 14191 8134 14201 8186
rect 14201 8134 14247 8186
rect 13951 8132 14007 8134
rect 14031 8132 14087 8134
rect 14111 8132 14167 8134
rect 14191 8132 14247 8134
rect 13951 7098 14007 7100
rect 14031 7098 14087 7100
rect 14111 7098 14167 7100
rect 14191 7098 14247 7100
rect 13951 7046 13997 7098
rect 13997 7046 14007 7098
rect 14031 7046 14061 7098
rect 14061 7046 14073 7098
rect 14073 7046 14087 7098
rect 14111 7046 14125 7098
rect 14125 7046 14137 7098
rect 14137 7046 14167 7098
rect 14191 7046 14201 7098
rect 14201 7046 14247 7098
rect 13951 7044 14007 7046
rect 14031 7044 14087 7046
rect 14111 7044 14167 7046
rect 14191 7044 14247 7046
rect 13951 6010 14007 6012
rect 14031 6010 14087 6012
rect 14111 6010 14167 6012
rect 14191 6010 14247 6012
rect 13951 5958 13997 6010
rect 13997 5958 14007 6010
rect 14031 5958 14061 6010
rect 14061 5958 14073 6010
rect 14073 5958 14087 6010
rect 14111 5958 14125 6010
rect 14125 5958 14137 6010
rect 14137 5958 14167 6010
rect 14191 5958 14201 6010
rect 14201 5958 14247 6010
rect 13951 5956 14007 5958
rect 14031 5956 14087 5958
rect 14111 5956 14167 5958
rect 14191 5956 14247 5958
rect 16550 10906 16606 10908
rect 16630 10906 16686 10908
rect 16710 10906 16766 10908
rect 16790 10906 16846 10908
rect 16550 10854 16596 10906
rect 16596 10854 16606 10906
rect 16630 10854 16660 10906
rect 16660 10854 16672 10906
rect 16672 10854 16686 10906
rect 16710 10854 16724 10906
rect 16724 10854 16736 10906
rect 16736 10854 16766 10906
rect 16790 10854 16800 10906
rect 16800 10854 16846 10906
rect 16550 10852 16606 10854
rect 16630 10852 16686 10854
rect 16710 10852 16766 10854
rect 16790 10852 16846 10854
rect 16550 9818 16606 9820
rect 16630 9818 16686 9820
rect 16710 9818 16766 9820
rect 16790 9818 16846 9820
rect 16550 9766 16596 9818
rect 16596 9766 16606 9818
rect 16630 9766 16660 9818
rect 16660 9766 16672 9818
rect 16672 9766 16686 9818
rect 16710 9766 16724 9818
rect 16724 9766 16736 9818
rect 16736 9766 16766 9818
rect 16790 9766 16800 9818
rect 16800 9766 16846 9818
rect 16550 9764 16606 9766
rect 16630 9764 16686 9766
rect 16710 9764 16766 9766
rect 16790 9764 16846 9766
rect 16550 8730 16606 8732
rect 16630 8730 16686 8732
rect 16710 8730 16766 8732
rect 16790 8730 16846 8732
rect 16550 8678 16596 8730
rect 16596 8678 16606 8730
rect 16630 8678 16660 8730
rect 16660 8678 16672 8730
rect 16672 8678 16686 8730
rect 16710 8678 16724 8730
rect 16724 8678 16736 8730
rect 16736 8678 16766 8730
rect 16790 8678 16800 8730
rect 16800 8678 16846 8730
rect 16550 8676 16606 8678
rect 16630 8676 16686 8678
rect 16710 8676 16766 8678
rect 16790 8676 16846 8678
rect 15658 8336 15714 8392
rect 19149 12538 19205 12540
rect 19229 12538 19285 12540
rect 19309 12538 19365 12540
rect 19389 12538 19445 12540
rect 19149 12486 19195 12538
rect 19195 12486 19205 12538
rect 19229 12486 19259 12538
rect 19259 12486 19271 12538
rect 19271 12486 19285 12538
rect 19309 12486 19323 12538
rect 19323 12486 19335 12538
rect 19335 12486 19365 12538
rect 19389 12486 19399 12538
rect 19399 12486 19445 12538
rect 19149 12484 19205 12486
rect 19229 12484 19285 12486
rect 19309 12484 19365 12486
rect 19389 12484 19445 12486
rect 18602 12280 18658 12336
rect 19149 11450 19205 11452
rect 19229 11450 19285 11452
rect 19309 11450 19365 11452
rect 19389 11450 19445 11452
rect 19149 11398 19195 11450
rect 19195 11398 19205 11450
rect 19229 11398 19259 11450
rect 19259 11398 19271 11450
rect 19271 11398 19285 11450
rect 19309 11398 19323 11450
rect 19323 11398 19335 11450
rect 19335 11398 19365 11450
rect 19389 11398 19399 11450
rect 19399 11398 19445 11450
rect 19149 11396 19205 11398
rect 19229 11396 19285 11398
rect 19309 11396 19365 11398
rect 19389 11396 19445 11398
rect 19149 10362 19205 10364
rect 19229 10362 19285 10364
rect 19309 10362 19365 10364
rect 19389 10362 19445 10364
rect 19149 10310 19195 10362
rect 19195 10310 19205 10362
rect 19229 10310 19259 10362
rect 19259 10310 19271 10362
rect 19271 10310 19285 10362
rect 19309 10310 19323 10362
rect 19323 10310 19335 10362
rect 19335 10310 19365 10362
rect 19389 10310 19399 10362
rect 19399 10310 19445 10362
rect 19149 10308 19205 10310
rect 19229 10308 19285 10310
rect 19309 10308 19365 10310
rect 19389 10308 19445 10310
rect 19149 9274 19205 9276
rect 19229 9274 19285 9276
rect 19309 9274 19365 9276
rect 19389 9274 19445 9276
rect 19149 9222 19195 9274
rect 19195 9222 19205 9274
rect 19229 9222 19259 9274
rect 19259 9222 19271 9274
rect 19271 9222 19285 9274
rect 19309 9222 19323 9274
rect 19323 9222 19335 9274
rect 19335 9222 19365 9274
rect 19389 9222 19399 9274
rect 19399 9222 19445 9274
rect 19149 9220 19205 9222
rect 19229 9220 19285 9222
rect 19309 9220 19365 9222
rect 19389 9220 19445 9222
rect 15474 6740 15476 6760
rect 15476 6740 15528 6760
rect 15528 6740 15530 6760
rect 15474 6704 15530 6740
rect 13951 4922 14007 4924
rect 14031 4922 14087 4924
rect 14111 4922 14167 4924
rect 14191 4922 14247 4924
rect 13951 4870 13997 4922
rect 13997 4870 14007 4922
rect 14031 4870 14061 4922
rect 14061 4870 14073 4922
rect 14073 4870 14087 4922
rect 14111 4870 14125 4922
rect 14125 4870 14137 4922
rect 14137 4870 14167 4922
rect 14191 4870 14201 4922
rect 14201 4870 14247 4922
rect 13951 4868 14007 4870
rect 14031 4868 14087 4870
rect 14111 4868 14167 4870
rect 14191 4868 14247 4870
rect 12346 2760 12402 2816
rect 12806 3032 12862 3088
rect 14278 4004 14334 4040
rect 14278 3984 14280 4004
rect 14280 3984 14332 4004
rect 14332 3984 14334 4004
rect 13082 3068 13084 3088
rect 13084 3068 13136 3088
rect 13136 3068 13138 3088
rect 13082 3032 13138 3068
rect 13951 3834 14007 3836
rect 14031 3834 14087 3836
rect 14111 3834 14167 3836
rect 14191 3834 14247 3836
rect 13951 3782 13997 3834
rect 13997 3782 14007 3834
rect 14031 3782 14061 3834
rect 14061 3782 14073 3834
rect 14073 3782 14087 3834
rect 14111 3782 14125 3834
rect 14125 3782 14137 3834
rect 14137 3782 14167 3834
rect 14191 3782 14201 3834
rect 14201 3782 14247 3834
rect 13951 3780 14007 3782
rect 14031 3780 14087 3782
rect 14111 3780 14167 3782
rect 14191 3780 14247 3782
rect 16550 7642 16606 7644
rect 16630 7642 16686 7644
rect 16710 7642 16766 7644
rect 16790 7642 16846 7644
rect 16550 7590 16596 7642
rect 16596 7590 16606 7642
rect 16630 7590 16660 7642
rect 16660 7590 16672 7642
rect 16672 7590 16686 7642
rect 16710 7590 16724 7642
rect 16724 7590 16736 7642
rect 16736 7590 16766 7642
rect 16790 7590 16800 7642
rect 16800 7590 16846 7642
rect 16550 7588 16606 7590
rect 16630 7588 16686 7590
rect 16710 7588 16766 7590
rect 16790 7588 16846 7590
rect 18510 8472 18566 8528
rect 18050 7384 18106 7440
rect 17038 7248 17094 7304
rect 16550 6554 16606 6556
rect 16630 6554 16686 6556
rect 16710 6554 16766 6556
rect 16790 6554 16846 6556
rect 16550 6502 16596 6554
rect 16596 6502 16606 6554
rect 16630 6502 16660 6554
rect 16660 6502 16672 6554
rect 16672 6502 16686 6554
rect 16710 6502 16724 6554
rect 16724 6502 16736 6554
rect 16736 6502 16766 6554
rect 16790 6502 16800 6554
rect 16800 6502 16846 6554
rect 16550 6500 16606 6502
rect 16630 6500 16686 6502
rect 16710 6500 16766 6502
rect 16790 6500 16846 6502
rect 16550 5466 16606 5468
rect 16630 5466 16686 5468
rect 16710 5466 16766 5468
rect 16790 5466 16846 5468
rect 16550 5414 16596 5466
rect 16596 5414 16606 5466
rect 16630 5414 16660 5466
rect 16660 5414 16672 5466
rect 16672 5414 16686 5466
rect 16710 5414 16724 5466
rect 16724 5414 16736 5466
rect 16736 5414 16766 5466
rect 16790 5414 16800 5466
rect 16800 5414 16846 5466
rect 16550 5412 16606 5414
rect 16630 5412 16686 5414
rect 16710 5412 16766 5414
rect 16790 5412 16846 5414
rect 16550 4378 16606 4380
rect 16630 4378 16686 4380
rect 16710 4378 16766 4380
rect 16790 4378 16846 4380
rect 16550 4326 16596 4378
rect 16596 4326 16606 4378
rect 16630 4326 16660 4378
rect 16660 4326 16672 4378
rect 16672 4326 16686 4378
rect 16710 4326 16724 4378
rect 16724 4326 16736 4378
rect 16736 4326 16766 4378
rect 16790 4326 16800 4378
rect 16800 4326 16846 4378
rect 16550 4324 16606 4326
rect 16630 4324 16686 4326
rect 16710 4324 16766 4326
rect 16790 4324 16846 4326
rect 13951 2746 14007 2748
rect 14031 2746 14087 2748
rect 14111 2746 14167 2748
rect 14191 2746 14247 2748
rect 13951 2694 13997 2746
rect 13997 2694 14007 2746
rect 14031 2694 14061 2746
rect 14061 2694 14073 2746
rect 14073 2694 14087 2746
rect 14111 2694 14125 2746
rect 14125 2694 14137 2746
rect 14137 2694 14167 2746
rect 14191 2694 14201 2746
rect 14201 2694 14247 2746
rect 13951 2692 14007 2694
rect 14031 2692 14087 2694
rect 14111 2692 14167 2694
rect 14191 2692 14247 2694
rect 17774 4664 17830 4720
rect 18050 4120 18106 4176
rect 16762 3576 16818 3632
rect 15566 3052 15622 3088
rect 15566 3032 15568 3052
rect 15568 3032 15620 3052
rect 15620 3032 15622 3052
rect 15658 2896 15714 2952
rect 16550 3290 16606 3292
rect 16630 3290 16686 3292
rect 16710 3290 16766 3292
rect 16790 3290 16846 3292
rect 16550 3238 16596 3290
rect 16596 3238 16606 3290
rect 16630 3238 16660 3290
rect 16660 3238 16672 3290
rect 16672 3238 16686 3290
rect 16710 3238 16724 3290
rect 16724 3238 16736 3290
rect 16736 3238 16766 3290
rect 16790 3238 16800 3290
rect 16800 3238 16846 3290
rect 16550 3236 16606 3238
rect 16630 3236 16686 3238
rect 16710 3236 16766 3238
rect 16790 3236 16846 3238
rect 16550 2202 16606 2204
rect 16630 2202 16686 2204
rect 16710 2202 16766 2204
rect 16790 2202 16846 2204
rect 16550 2150 16596 2202
rect 16596 2150 16606 2202
rect 16630 2150 16660 2202
rect 16660 2150 16672 2202
rect 16672 2150 16686 2202
rect 16710 2150 16724 2202
rect 16724 2150 16736 2202
rect 16736 2150 16766 2202
rect 16790 2150 16800 2202
rect 16800 2150 16846 2202
rect 16550 2148 16606 2150
rect 16630 2148 16686 2150
rect 16710 2148 16766 2150
rect 16790 2148 16846 2150
rect 18142 3440 18198 3496
rect 18234 2352 18290 2408
rect 17866 1808 17922 1864
rect 19149 8186 19205 8188
rect 19229 8186 19285 8188
rect 19309 8186 19365 8188
rect 19389 8186 19445 8188
rect 19149 8134 19195 8186
rect 19195 8134 19205 8186
rect 19229 8134 19259 8186
rect 19259 8134 19271 8186
rect 19271 8134 19285 8186
rect 19309 8134 19323 8186
rect 19323 8134 19335 8186
rect 19335 8134 19365 8186
rect 19389 8134 19399 8186
rect 19399 8134 19445 8186
rect 19149 8132 19205 8134
rect 19229 8132 19285 8134
rect 19309 8132 19365 8134
rect 19389 8132 19445 8134
rect 19062 7928 19118 7984
rect 19982 10532 20038 10568
rect 19982 10512 19984 10532
rect 19984 10512 20036 10532
rect 20036 10512 20038 10532
rect 20626 9968 20682 10024
rect 19798 9016 19854 9072
rect 19149 7098 19205 7100
rect 19229 7098 19285 7100
rect 19309 7098 19365 7100
rect 19389 7098 19445 7100
rect 19149 7046 19195 7098
rect 19195 7046 19205 7098
rect 19229 7046 19259 7098
rect 19259 7046 19271 7098
rect 19271 7046 19285 7098
rect 19309 7046 19323 7098
rect 19323 7046 19335 7098
rect 19335 7046 19365 7098
rect 19389 7046 19399 7098
rect 19399 7046 19445 7098
rect 19149 7044 19205 7046
rect 19229 7044 19285 7046
rect 19309 7044 19365 7046
rect 19389 7044 19445 7046
rect 21748 16346 21804 16348
rect 21828 16346 21884 16348
rect 21908 16346 21964 16348
rect 21988 16346 22044 16348
rect 21748 16294 21794 16346
rect 21794 16294 21804 16346
rect 21828 16294 21858 16346
rect 21858 16294 21870 16346
rect 21870 16294 21884 16346
rect 21908 16294 21922 16346
rect 21922 16294 21934 16346
rect 21934 16294 21964 16346
rect 21988 16294 21998 16346
rect 21998 16294 22044 16346
rect 21748 16292 21804 16294
rect 21828 16292 21884 16294
rect 21908 16292 21964 16294
rect 21988 16292 22044 16294
rect 21748 15258 21804 15260
rect 21828 15258 21884 15260
rect 21908 15258 21964 15260
rect 21988 15258 22044 15260
rect 21748 15206 21794 15258
rect 21794 15206 21804 15258
rect 21828 15206 21858 15258
rect 21858 15206 21870 15258
rect 21870 15206 21884 15258
rect 21908 15206 21922 15258
rect 21922 15206 21934 15258
rect 21934 15206 21964 15258
rect 21988 15206 21998 15258
rect 21998 15206 22044 15258
rect 21748 15204 21804 15206
rect 21828 15204 21884 15206
rect 21908 15204 21964 15206
rect 21988 15204 22044 15206
rect 21748 14170 21804 14172
rect 21828 14170 21884 14172
rect 21908 14170 21964 14172
rect 21988 14170 22044 14172
rect 21748 14118 21794 14170
rect 21794 14118 21804 14170
rect 21828 14118 21858 14170
rect 21858 14118 21870 14170
rect 21870 14118 21884 14170
rect 21908 14118 21922 14170
rect 21922 14118 21934 14170
rect 21934 14118 21964 14170
rect 21988 14118 21998 14170
rect 21998 14118 22044 14170
rect 21748 14116 21804 14118
rect 21828 14116 21884 14118
rect 21908 14116 21964 14118
rect 21988 14116 22044 14118
rect 21748 13082 21804 13084
rect 21828 13082 21884 13084
rect 21908 13082 21964 13084
rect 21988 13082 22044 13084
rect 21748 13030 21794 13082
rect 21794 13030 21804 13082
rect 21828 13030 21858 13082
rect 21858 13030 21870 13082
rect 21870 13030 21884 13082
rect 21908 13030 21922 13082
rect 21922 13030 21934 13082
rect 21934 13030 21964 13082
rect 21988 13030 21998 13082
rect 21998 13030 22044 13082
rect 21748 13028 21804 13030
rect 21828 13028 21884 13030
rect 21908 13028 21964 13030
rect 21988 13028 22044 13030
rect 21748 11994 21804 11996
rect 21828 11994 21884 11996
rect 21908 11994 21964 11996
rect 21988 11994 22044 11996
rect 21748 11942 21794 11994
rect 21794 11942 21804 11994
rect 21828 11942 21858 11994
rect 21858 11942 21870 11994
rect 21870 11942 21884 11994
rect 21908 11942 21922 11994
rect 21922 11942 21934 11994
rect 21934 11942 21964 11994
rect 21988 11942 21998 11994
rect 21998 11942 22044 11994
rect 21748 11940 21804 11942
rect 21828 11940 21884 11942
rect 21908 11940 21964 11942
rect 21988 11940 22044 11942
rect 21748 10906 21804 10908
rect 21828 10906 21884 10908
rect 21908 10906 21964 10908
rect 21988 10906 22044 10908
rect 21748 10854 21794 10906
rect 21794 10854 21804 10906
rect 21828 10854 21858 10906
rect 21858 10854 21870 10906
rect 21870 10854 21884 10906
rect 21908 10854 21922 10906
rect 21922 10854 21934 10906
rect 21934 10854 21964 10906
rect 21988 10854 21998 10906
rect 21998 10854 22044 10906
rect 21748 10852 21804 10854
rect 21828 10852 21884 10854
rect 21908 10852 21964 10854
rect 21988 10852 22044 10854
rect 21748 9818 21804 9820
rect 21828 9818 21884 9820
rect 21908 9818 21964 9820
rect 21988 9818 22044 9820
rect 21748 9766 21794 9818
rect 21794 9766 21804 9818
rect 21828 9766 21858 9818
rect 21858 9766 21870 9818
rect 21870 9766 21884 9818
rect 21908 9766 21922 9818
rect 21922 9766 21934 9818
rect 21934 9766 21964 9818
rect 21988 9766 21998 9818
rect 21998 9766 22044 9818
rect 21748 9764 21804 9766
rect 21828 9764 21884 9766
rect 21908 9764 21964 9766
rect 21988 9764 22044 9766
rect 21748 8730 21804 8732
rect 21828 8730 21884 8732
rect 21908 8730 21964 8732
rect 21988 8730 22044 8732
rect 21748 8678 21794 8730
rect 21794 8678 21804 8730
rect 21828 8678 21858 8730
rect 21858 8678 21870 8730
rect 21870 8678 21884 8730
rect 21908 8678 21922 8730
rect 21922 8678 21934 8730
rect 21934 8678 21964 8730
rect 21988 8678 21998 8730
rect 21998 8678 22044 8730
rect 21748 8676 21804 8678
rect 21828 8676 21884 8678
rect 21908 8676 21964 8678
rect 21988 8676 22044 8678
rect 21748 7642 21804 7644
rect 21828 7642 21884 7644
rect 21908 7642 21964 7644
rect 21988 7642 22044 7644
rect 21748 7590 21794 7642
rect 21794 7590 21804 7642
rect 21828 7590 21858 7642
rect 21858 7590 21870 7642
rect 21870 7590 21884 7642
rect 21908 7590 21922 7642
rect 21922 7590 21934 7642
rect 21934 7590 21964 7642
rect 21988 7590 21998 7642
rect 21998 7590 22044 7642
rect 21748 7588 21804 7590
rect 21828 7588 21884 7590
rect 21908 7588 21964 7590
rect 21988 7588 22044 7590
rect 20626 6840 20682 6896
rect 19149 6010 19205 6012
rect 19229 6010 19285 6012
rect 19309 6010 19365 6012
rect 19389 6010 19445 6012
rect 19149 5958 19195 6010
rect 19195 5958 19205 6010
rect 19229 5958 19259 6010
rect 19259 5958 19271 6010
rect 19271 5958 19285 6010
rect 19309 5958 19323 6010
rect 19323 5958 19335 6010
rect 19335 5958 19365 6010
rect 19389 5958 19399 6010
rect 19399 5958 19445 6010
rect 19149 5956 19205 5958
rect 19229 5956 19285 5958
rect 19309 5956 19365 5958
rect 19389 5956 19445 5958
rect 19149 4922 19205 4924
rect 19229 4922 19285 4924
rect 19309 4922 19365 4924
rect 19389 4922 19445 4924
rect 19149 4870 19195 4922
rect 19195 4870 19205 4922
rect 19229 4870 19259 4922
rect 19259 4870 19271 4922
rect 19271 4870 19285 4922
rect 19309 4870 19323 4922
rect 19323 4870 19335 4922
rect 19335 4870 19365 4922
rect 19389 4870 19399 4922
rect 19399 4870 19445 4922
rect 19149 4868 19205 4870
rect 19229 4868 19285 4870
rect 19309 4868 19365 4870
rect 19389 4868 19445 4870
rect 19149 3834 19205 3836
rect 19229 3834 19285 3836
rect 19309 3834 19365 3836
rect 19389 3834 19445 3836
rect 19149 3782 19195 3834
rect 19195 3782 19205 3834
rect 19229 3782 19259 3834
rect 19259 3782 19271 3834
rect 19271 3782 19285 3834
rect 19309 3782 19323 3834
rect 19323 3782 19335 3834
rect 19335 3782 19365 3834
rect 19389 3782 19399 3834
rect 19399 3782 19445 3834
rect 19149 3780 19205 3782
rect 19229 3780 19285 3782
rect 19309 3780 19365 3782
rect 19389 3780 19445 3782
rect 19149 2746 19205 2748
rect 19229 2746 19285 2748
rect 19309 2746 19365 2748
rect 19389 2746 19445 2748
rect 19149 2694 19195 2746
rect 19195 2694 19205 2746
rect 19229 2694 19259 2746
rect 19259 2694 19271 2746
rect 19271 2694 19285 2746
rect 19309 2694 19323 2746
rect 19323 2694 19335 2746
rect 19335 2694 19365 2746
rect 19389 2694 19399 2746
rect 19399 2694 19445 2746
rect 19149 2692 19205 2694
rect 19229 2692 19285 2694
rect 19309 2692 19365 2694
rect 19389 2692 19445 2694
rect 21748 6554 21804 6556
rect 21828 6554 21884 6556
rect 21908 6554 21964 6556
rect 21988 6554 22044 6556
rect 21748 6502 21794 6554
rect 21794 6502 21804 6554
rect 21828 6502 21858 6554
rect 21858 6502 21870 6554
rect 21870 6502 21884 6554
rect 21908 6502 21922 6554
rect 21922 6502 21934 6554
rect 21934 6502 21964 6554
rect 21988 6502 21998 6554
rect 21998 6502 22044 6554
rect 21748 6500 21804 6502
rect 21828 6500 21884 6502
rect 21908 6500 21964 6502
rect 21988 6500 22044 6502
rect 21748 5466 21804 5468
rect 21828 5466 21884 5468
rect 21908 5466 21964 5468
rect 21988 5466 22044 5468
rect 21748 5414 21794 5466
rect 21794 5414 21804 5466
rect 21828 5414 21858 5466
rect 21858 5414 21870 5466
rect 21870 5414 21884 5466
rect 21908 5414 21922 5466
rect 21922 5414 21934 5466
rect 21934 5414 21964 5466
rect 21988 5414 21998 5466
rect 21998 5414 22044 5466
rect 21748 5412 21804 5414
rect 21828 5412 21884 5414
rect 21908 5412 21964 5414
rect 21988 5412 22044 5414
rect 21748 4378 21804 4380
rect 21828 4378 21884 4380
rect 21908 4378 21964 4380
rect 21988 4378 22044 4380
rect 21748 4326 21794 4378
rect 21794 4326 21804 4378
rect 21828 4326 21858 4378
rect 21858 4326 21870 4378
rect 21870 4326 21884 4378
rect 21908 4326 21922 4378
rect 21922 4326 21934 4378
rect 21934 4326 21964 4378
rect 21988 4326 21998 4378
rect 21998 4326 22044 4378
rect 21748 4324 21804 4326
rect 21828 4324 21884 4326
rect 21908 4324 21964 4326
rect 21988 4324 22044 4326
rect 21748 3290 21804 3292
rect 21828 3290 21884 3292
rect 21908 3290 21964 3292
rect 21988 3290 22044 3292
rect 21748 3238 21794 3290
rect 21794 3238 21804 3290
rect 21828 3238 21858 3290
rect 21858 3238 21870 3290
rect 21870 3238 21884 3290
rect 21908 3238 21922 3290
rect 21922 3238 21934 3290
rect 21934 3238 21964 3290
rect 21988 3238 21998 3290
rect 21998 3238 22044 3290
rect 21748 3236 21804 3238
rect 21828 3236 21884 3238
rect 21908 3236 21964 3238
rect 21988 3236 22044 3238
rect 20718 2524 20720 2544
rect 20720 2524 20772 2544
rect 20772 2524 20774 2544
rect 20718 2488 20774 2524
rect 19338 1672 19394 1728
rect 21748 2202 21804 2204
rect 21828 2202 21884 2204
rect 21908 2202 21964 2204
rect 21988 2202 22044 2204
rect 21748 2150 21794 2202
rect 21794 2150 21804 2202
rect 21828 2150 21858 2202
rect 21858 2150 21870 2202
rect 21870 2150 21884 2202
rect 21908 2150 21922 2202
rect 21922 2150 21934 2202
rect 21934 2150 21964 2202
rect 21988 2150 21998 2202
rect 21998 2150 22044 2202
rect 21748 2148 21804 2150
rect 21828 2148 21884 2150
rect 21908 2148 21964 2150
rect 21988 2148 22044 2150
<< metal3 >>
rect 0 21314 800 21344
rect 2957 21314 3023 21317
rect 0 21312 3023 21314
rect 0 21256 2962 21312
rect 3018 21256 3023 21312
rect 0 21254 3023 21256
rect 0 21224 800 21254
rect 2957 21251 3023 21254
rect 0 20906 800 20936
rect 3877 20906 3943 20909
rect 0 20904 3943 20906
rect 0 20848 3882 20904
rect 3938 20848 3943 20904
rect 0 20846 3943 20848
rect 0 20816 800 20846
rect 3877 20843 3943 20846
rect 6144 20704 6460 20705
rect 6144 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6460 20704
rect 6144 20639 6460 20640
rect 11342 20704 11658 20705
rect 11342 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11658 20704
rect 11342 20639 11658 20640
rect 16540 20704 16856 20705
rect 16540 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16856 20704
rect 16540 20639 16856 20640
rect 21738 20704 22054 20705
rect 21738 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22054 20704
rect 21738 20639 22054 20640
rect 0 20498 800 20528
rect 4061 20498 4127 20501
rect 0 20496 4127 20498
rect 0 20440 4066 20496
rect 4122 20440 4127 20496
rect 0 20438 4127 20440
rect 0 20408 800 20438
rect 4061 20435 4127 20438
rect 3545 20160 3861 20161
rect 0 20090 800 20120
rect 3545 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3861 20160
rect 3545 20095 3861 20096
rect 8743 20160 9059 20161
rect 8743 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9059 20160
rect 8743 20095 9059 20096
rect 13941 20160 14257 20161
rect 13941 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14257 20160
rect 13941 20095 14257 20096
rect 19139 20160 19455 20161
rect 19139 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19455 20160
rect 19139 20095 19455 20096
rect 3233 20090 3299 20093
rect 0 20088 3299 20090
rect 0 20032 3238 20088
rect 3294 20032 3299 20088
rect 0 20030 3299 20032
rect 0 20000 800 20030
rect 3233 20027 3299 20030
rect 0 19682 800 19712
rect 4153 19682 4219 19685
rect 0 19680 4219 19682
rect 0 19624 4158 19680
rect 4214 19624 4219 19680
rect 0 19622 4219 19624
rect 0 19592 800 19622
rect 4153 19619 4219 19622
rect 6144 19616 6460 19617
rect 6144 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6460 19616
rect 6144 19551 6460 19552
rect 11342 19616 11658 19617
rect 11342 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11658 19616
rect 11342 19551 11658 19552
rect 16540 19616 16856 19617
rect 16540 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16856 19616
rect 16540 19551 16856 19552
rect 21738 19616 22054 19617
rect 21738 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22054 19616
rect 21738 19551 22054 19552
rect 0 19274 800 19304
rect 4061 19274 4127 19277
rect 0 19272 4127 19274
rect 0 19216 4066 19272
rect 4122 19216 4127 19272
rect 0 19214 4127 19216
rect 0 19184 800 19214
rect 4061 19211 4127 19214
rect 3545 19072 3861 19073
rect 3545 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3861 19072
rect 3545 19007 3861 19008
rect 8743 19072 9059 19073
rect 8743 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9059 19072
rect 8743 19007 9059 19008
rect 13941 19072 14257 19073
rect 13941 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14257 19072
rect 13941 19007 14257 19008
rect 19139 19072 19455 19073
rect 19139 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19455 19072
rect 19139 19007 19455 19008
rect 0 18866 800 18896
rect 4153 18866 4219 18869
rect 0 18864 4219 18866
rect 0 18808 4158 18864
rect 4214 18808 4219 18864
rect 0 18806 4219 18808
rect 0 18776 800 18806
rect 4153 18803 4219 18806
rect 6144 18528 6460 18529
rect 0 18458 800 18488
rect 6144 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6460 18528
rect 6144 18463 6460 18464
rect 11342 18528 11658 18529
rect 11342 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11658 18528
rect 11342 18463 11658 18464
rect 16540 18528 16856 18529
rect 16540 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16856 18528
rect 16540 18463 16856 18464
rect 21738 18528 22054 18529
rect 21738 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22054 18528
rect 21738 18463 22054 18464
rect 3969 18458 4035 18461
rect 0 18456 4035 18458
rect 0 18400 3974 18456
rect 4030 18400 4035 18456
rect 0 18398 4035 18400
rect 0 18368 800 18398
rect 3969 18395 4035 18398
rect 0 18050 800 18080
rect 1945 18050 2011 18053
rect 0 18048 2011 18050
rect 0 17992 1950 18048
rect 2006 17992 2011 18048
rect 0 17990 2011 17992
rect 0 17960 800 17990
rect 1945 17987 2011 17990
rect 3545 17984 3861 17985
rect 3545 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3861 17984
rect 3545 17919 3861 17920
rect 8743 17984 9059 17985
rect 8743 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9059 17984
rect 8743 17919 9059 17920
rect 13941 17984 14257 17985
rect 13941 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14257 17984
rect 13941 17919 14257 17920
rect 19139 17984 19455 17985
rect 19139 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19455 17984
rect 19139 17919 19455 17920
rect 0 17642 800 17672
rect 3693 17642 3759 17645
rect 0 17640 3759 17642
rect 0 17584 3698 17640
rect 3754 17584 3759 17640
rect 0 17582 3759 17584
rect 0 17552 800 17582
rect 3693 17579 3759 17582
rect 6144 17440 6460 17441
rect 6144 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6460 17440
rect 6144 17375 6460 17376
rect 11342 17440 11658 17441
rect 11342 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11658 17440
rect 11342 17375 11658 17376
rect 16540 17440 16856 17441
rect 16540 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16856 17440
rect 16540 17375 16856 17376
rect 21738 17440 22054 17441
rect 21738 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22054 17440
rect 21738 17375 22054 17376
rect 0 17234 800 17264
rect 1577 17234 1643 17237
rect 0 17232 1643 17234
rect 0 17176 1582 17232
rect 1638 17176 1643 17232
rect 0 17174 1643 17176
rect 0 17144 800 17174
rect 1577 17171 1643 17174
rect 21449 17234 21515 17237
rect 22200 17234 23000 17264
rect 21449 17232 23000 17234
rect 21449 17176 21454 17232
rect 21510 17176 23000 17232
rect 21449 17174 23000 17176
rect 21449 17171 21515 17174
rect 22200 17144 23000 17174
rect 3545 16896 3861 16897
rect 0 16826 800 16856
rect 3545 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3861 16896
rect 3545 16831 3861 16832
rect 8743 16896 9059 16897
rect 8743 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9059 16896
rect 8743 16831 9059 16832
rect 13941 16896 14257 16897
rect 13941 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14257 16896
rect 13941 16831 14257 16832
rect 19139 16896 19455 16897
rect 19139 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19455 16896
rect 19139 16831 19455 16832
rect 1945 16826 2011 16829
rect 0 16824 2011 16826
rect 0 16768 1950 16824
rect 2006 16768 2011 16824
rect 0 16766 2011 16768
rect 0 16736 800 16766
rect 1945 16763 2011 16766
rect 0 16418 800 16448
rect 1669 16418 1735 16421
rect 0 16416 1735 16418
rect 0 16360 1674 16416
rect 1730 16360 1735 16416
rect 0 16358 1735 16360
rect 0 16328 800 16358
rect 1669 16355 1735 16358
rect 6144 16352 6460 16353
rect 6144 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6460 16352
rect 6144 16287 6460 16288
rect 11342 16352 11658 16353
rect 11342 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11658 16352
rect 11342 16287 11658 16288
rect 16540 16352 16856 16353
rect 16540 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16856 16352
rect 16540 16287 16856 16288
rect 21738 16352 22054 16353
rect 21738 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22054 16352
rect 21738 16287 22054 16288
rect 0 16010 800 16040
rect 2773 16010 2839 16013
rect 0 16008 2839 16010
rect 0 15952 2778 16008
rect 2834 15952 2839 16008
rect 0 15950 2839 15952
rect 0 15920 800 15950
rect 2773 15947 2839 15950
rect 3545 15808 3861 15809
rect 3545 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3861 15808
rect 3545 15743 3861 15744
rect 8743 15808 9059 15809
rect 8743 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9059 15808
rect 8743 15743 9059 15744
rect 13941 15808 14257 15809
rect 13941 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14257 15808
rect 13941 15743 14257 15744
rect 19139 15808 19455 15809
rect 19139 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19455 15808
rect 19139 15743 19455 15744
rect 0 15602 800 15632
rect 2221 15602 2287 15605
rect 0 15600 2287 15602
rect 0 15544 2226 15600
rect 2282 15544 2287 15600
rect 0 15542 2287 15544
rect 0 15512 800 15542
rect 2221 15539 2287 15542
rect 6144 15264 6460 15265
rect 0 15194 800 15224
rect 6144 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6460 15264
rect 6144 15199 6460 15200
rect 11342 15264 11658 15265
rect 11342 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11658 15264
rect 11342 15199 11658 15200
rect 16540 15264 16856 15265
rect 16540 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16856 15264
rect 16540 15199 16856 15200
rect 21738 15264 22054 15265
rect 21738 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22054 15264
rect 21738 15199 22054 15200
rect 1485 15194 1551 15197
rect 0 15192 1551 15194
rect 0 15136 1490 15192
rect 1546 15136 1551 15192
rect 0 15134 1551 15136
rect 0 15104 800 15134
rect 1485 15131 1551 15134
rect 0 14786 800 14816
rect 1945 14786 2011 14789
rect 0 14784 2011 14786
rect 0 14728 1950 14784
rect 2006 14728 2011 14784
rect 0 14726 2011 14728
rect 0 14696 800 14726
rect 1945 14723 2011 14726
rect 3545 14720 3861 14721
rect 3545 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3861 14720
rect 3545 14655 3861 14656
rect 8743 14720 9059 14721
rect 8743 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9059 14720
rect 8743 14655 9059 14656
rect 13941 14720 14257 14721
rect 13941 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14257 14720
rect 13941 14655 14257 14656
rect 19139 14720 19455 14721
rect 19139 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19455 14720
rect 19139 14655 19455 14656
rect 0 14378 800 14408
rect 1945 14378 2011 14381
rect 0 14376 2011 14378
rect 0 14320 1950 14376
rect 2006 14320 2011 14376
rect 0 14318 2011 14320
rect 0 14288 800 14318
rect 1945 14315 2011 14318
rect 6144 14176 6460 14177
rect 6144 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6460 14176
rect 6144 14111 6460 14112
rect 11342 14176 11658 14177
rect 11342 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11658 14176
rect 11342 14111 11658 14112
rect 16540 14176 16856 14177
rect 16540 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16856 14176
rect 16540 14111 16856 14112
rect 21738 14176 22054 14177
rect 21738 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22054 14176
rect 21738 14111 22054 14112
rect 0 13970 800 14000
rect 2773 13970 2839 13973
rect 0 13968 2839 13970
rect 0 13912 2778 13968
rect 2834 13912 2839 13968
rect 0 13910 2839 13912
rect 0 13880 800 13910
rect 2773 13907 2839 13910
rect 6545 13970 6611 13973
rect 8334 13970 8340 13972
rect 6545 13968 8340 13970
rect 6545 13912 6550 13968
rect 6606 13912 8340 13968
rect 6545 13910 8340 13912
rect 6545 13907 6611 13910
rect 8334 13908 8340 13910
rect 8404 13908 8410 13972
rect 9029 13834 9095 13837
rect 9254 13834 9260 13836
rect 9029 13832 9260 13834
rect 9029 13776 9034 13832
rect 9090 13776 9260 13832
rect 9029 13774 9260 13776
rect 9029 13771 9095 13774
rect 9254 13772 9260 13774
rect 9324 13772 9330 13836
rect 3545 13632 3861 13633
rect 0 13562 800 13592
rect 3545 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3861 13632
rect 3545 13567 3861 13568
rect 8743 13632 9059 13633
rect 8743 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9059 13632
rect 8743 13567 9059 13568
rect 13941 13632 14257 13633
rect 13941 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14257 13632
rect 13941 13567 14257 13568
rect 19139 13632 19455 13633
rect 19139 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19455 13632
rect 19139 13567 19455 13568
rect 2773 13562 2839 13565
rect 0 13560 2839 13562
rect 0 13504 2778 13560
rect 2834 13504 2839 13560
rect 0 13502 2839 13504
rect 0 13472 800 13502
rect 2773 13499 2839 13502
rect 10133 13426 10199 13429
rect 19517 13426 19583 13429
rect 10133 13424 19583 13426
rect 10133 13368 10138 13424
rect 10194 13368 19522 13424
rect 19578 13368 19583 13424
rect 10133 13366 19583 13368
rect 10133 13363 10199 13366
rect 19517 13363 19583 13366
rect 0 13154 800 13184
rect 1669 13154 1735 13157
rect 0 13152 1735 13154
rect 0 13096 1674 13152
rect 1730 13096 1735 13152
rect 0 13094 1735 13096
rect 0 13064 800 13094
rect 1669 13091 1735 13094
rect 6144 13088 6460 13089
rect 6144 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6460 13088
rect 6144 13023 6460 13024
rect 11342 13088 11658 13089
rect 11342 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11658 13088
rect 11342 13023 11658 13024
rect 16540 13088 16856 13089
rect 16540 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16856 13088
rect 16540 13023 16856 13024
rect 21738 13088 22054 13089
rect 21738 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22054 13088
rect 21738 13023 22054 13024
rect 0 12746 800 12776
rect 2773 12746 2839 12749
rect 0 12744 2839 12746
rect 0 12688 2778 12744
rect 2834 12688 2839 12744
rect 0 12686 2839 12688
rect 0 12656 800 12686
rect 2773 12683 2839 12686
rect 4981 12610 5047 12613
rect 5574 12610 5580 12612
rect 4981 12608 5580 12610
rect 4981 12552 4986 12608
rect 5042 12552 5580 12608
rect 4981 12550 5580 12552
rect 4981 12547 5047 12550
rect 5574 12548 5580 12550
rect 5644 12548 5650 12612
rect 3545 12544 3861 12545
rect 3545 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3861 12544
rect 3545 12479 3861 12480
rect 8743 12544 9059 12545
rect 8743 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9059 12544
rect 8743 12479 9059 12480
rect 13941 12544 14257 12545
rect 13941 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14257 12544
rect 13941 12479 14257 12480
rect 19139 12544 19455 12545
rect 19139 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19455 12544
rect 19139 12479 19455 12480
rect 0 12338 800 12368
rect 2957 12338 3023 12341
rect 0 12336 3023 12338
rect 0 12280 2962 12336
rect 3018 12280 3023 12336
rect 0 12278 3023 12280
rect 0 12248 800 12278
rect 2957 12275 3023 12278
rect 7465 12338 7531 12341
rect 18597 12338 18663 12341
rect 7465 12336 18663 12338
rect 7465 12280 7470 12336
rect 7526 12280 18602 12336
rect 18658 12280 18663 12336
rect 7465 12278 18663 12280
rect 7465 12275 7531 12278
rect 18597 12275 18663 12278
rect 6144 12000 6460 12001
rect 0 11930 800 11960
rect 6144 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6460 12000
rect 6144 11935 6460 11936
rect 11342 12000 11658 12001
rect 11342 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11658 12000
rect 11342 11935 11658 11936
rect 16540 12000 16856 12001
rect 16540 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16856 12000
rect 16540 11935 16856 11936
rect 21738 12000 22054 12001
rect 21738 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22054 12000
rect 21738 11935 22054 11936
rect 1945 11930 2011 11933
rect 0 11928 2011 11930
rect 0 11872 1950 11928
rect 2006 11872 2011 11928
rect 0 11870 2011 11872
rect 0 11840 800 11870
rect 1945 11867 2011 11870
rect 2681 11794 2747 11797
rect 12249 11794 12315 11797
rect 2681 11792 12315 11794
rect 2681 11736 2686 11792
rect 2742 11736 12254 11792
rect 12310 11736 12315 11792
rect 2681 11734 12315 11736
rect 2681 11731 2747 11734
rect 12249 11731 12315 11734
rect 5625 11658 5691 11661
rect 13445 11658 13511 11661
rect 5625 11656 13511 11658
rect 5625 11600 5630 11656
rect 5686 11600 13450 11656
rect 13506 11600 13511 11656
rect 5625 11598 13511 11600
rect 5625 11595 5691 11598
rect 13445 11595 13511 11598
rect 0 11522 800 11552
rect 3417 11522 3483 11525
rect 0 11520 3483 11522
rect 0 11464 3422 11520
rect 3478 11464 3483 11520
rect 0 11462 3483 11464
rect 0 11432 800 11462
rect 3417 11459 3483 11462
rect 3545 11456 3861 11457
rect 3545 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3861 11456
rect 3545 11391 3861 11392
rect 8743 11456 9059 11457
rect 8743 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9059 11456
rect 8743 11391 9059 11392
rect 13941 11456 14257 11457
rect 13941 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14257 11456
rect 13941 11391 14257 11392
rect 19139 11456 19455 11457
rect 19139 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19455 11456
rect 19139 11391 19455 11392
rect 7741 11250 7807 11253
rect 8385 11250 8451 11253
rect 7741 11248 8451 11250
rect 7741 11192 7746 11248
rect 7802 11192 8390 11248
rect 8446 11192 8451 11248
rect 7741 11190 8451 11192
rect 7741 11187 7807 11190
rect 8385 11187 8451 11190
rect 10593 11250 10659 11253
rect 14457 11250 14523 11253
rect 10593 11248 14523 11250
rect 10593 11192 10598 11248
rect 10654 11192 14462 11248
rect 14518 11192 14523 11248
rect 10593 11190 14523 11192
rect 10593 11187 10659 11190
rect 14457 11187 14523 11190
rect 0 11114 800 11144
rect 4061 11114 4127 11117
rect 0 11112 4127 11114
rect 0 11056 4066 11112
rect 4122 11056 4127 11112
rect 0 11054 4127 11056
rect 0 11024 800 11054
rect 4061 11051 4127 11054
rect 6637 11114 6703 11117
rect 10961 11114 11027 11117
rect 6637 11112 11027 11114
rect 6637 11056 6642 11112
rect 6698 11056 10966 11112
rect 11022 11056 11027 11112
rect 6637 11054 11027 11056
rect 6637 11051 6703 11054
rect 10961 11051 11027 11054
rect 6144 10912 6460 10913
rect 6144 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6460 10912
rect 6144 10847 6460 10848
rect 11342 10912 11658 10913
rect 11342 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11658 10912
rect 11342 10847 11658 10848
rect 16540 10912 16856 10913
rect 16540 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16856 10912
rect 16540 10847 16856 10848
rect 21738 10912 22054 10913
rect 21738 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22054 10912
rect 21738 10847 22054 10848
rect 0 10706 800 10736
rect 3417 10706 3483 10709
rect 0 10704 3483 10706
rect 0 10648 3422 10704
rect 3478 10648 3483 10704
rect 0 10646 3483 10648
rect 0 10616 800 10646
rect 3417 10643 3483 10646
rect 8017 10570 8083 10573
rect 19977 10570 20043 10573
rect 8017 10568 20043 10570
rect 8017 10512 8022 10568
rect 8078 10512 19982 10568
rect 20038 10512 20043 10568
rect 8017 10510 20043 10512
rect 8017 10507 8083 10510
rect 19977 10507 20043 10510
rect 3545 10368 3861 10369
rect 0 10298 800 10328
rect 3545 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3861 10368
rect 3545 10303 3861 10304
rect 8743 10368 9059 10369
rect 8743 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9059 10368
rect 8743 10303 9059 10304
rect 13941 10368 14257 10369
rect 13941 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14257 10368
rect 13941 10303 14257 10304
rect 19139 10368 19455 10369
rect 19139 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19455 10368
rect 19139 10303 19455 10304
rect 3325 10298 3391 10301
rect 0 10296 3391 10298
rect 0 10240 3330 10296
rect 3386 10240 3391 10296
rect 0 10238 3391 10240
rect 0 10208 800 10238
rect 3325 10235 3391 10238
rect 7741 10298 7807 10301
rect 7741 10296 8356 10298
rect 7741 10240 7746 10296
rect 7802 10240 8356 10296
rect 7741 10238 8356 10240
rect 7741 10235 7807 10238
rect 8017 10162 8083 10165
rect 8150 10162 8156 10164
rect 8017 10160 8156 10162
rect 8017 10104 8022 10160
rect 8078 10104 8156 10160
rect 8017 10102 8156 10104
rect 8017 10099 8083 10102
rect 8150 10100 8156 10102
rect 8220 10100 8226 10164
rect 8296 10162 8356 10238
rect 11789 10162 11855 10165
rect 8296 10160 11855 10162
rect 8296 10104 11794 10160
rect 11850 10104 11855 10160
rect 8296 10102 11855 10104
rect 11789 10099 11855 10102
rect 4061 10026 4127 10029
rect 8293 10026 8359 10029
rect 4061 10024 8359 10026
rect 4061 9968 4066 10024
rect 4122 9968 8298 10024
rect 8354 9968 8359 10024
rect 4061 9966 8359 9968
rect 4061 9963 4127 9966
rect 8293 9963 8359 9966
rect 9581 10026 9647 10029
rect 20621 10026 20687 10029
rect 9581 10024 20687 10026
rect 9581 9968 9586 10024
rect 9642 9968 20626 10024
rect 20682 9968 20687 10024
rect 9581 9966 20687 9968
rect 9581 9963 9647 9966
rect 20621 9963 20687 9966
rect 0 9890 800 9920
rect 3877 9890 3943 9893
rect 0 9888 3943 9890
rect 0 9832 3882 9888
rect 3938 9832 3943 9888
rect 0 9830 3943 9832
rect 0 9800 800 9830
rect 3877 9827 3943 9830
rect 6144 9824 6460 9825
rect 6144 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6460 9824
rect 6144 9759 6460 9760
rect 11342 9824 11658 9825
rect 11342 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11658 9824
rect 11342 9759 11658 9760
rect 16540 9824 16856 9825
rect 16540 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16856 9824
rect 16540 9759 16856 9760
rect 21738 9824 22054 9825
rect 21738 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22054 9824
rect 21738 9759 22054 9760
rect 0 9482 800 9512
rect 3785 9482 3851 9485
rect 0 9480 3851 9482
rect 0 9424 3790 9480
rect 3846 9424 3851 9480
rect 0 9422 3851 9424
rect 0 9392 800 9422
rect 3785 9419 3851 9422
rect 4061 9482 4127 9485
rect 14457 9482 14523 9485
rect 4061 9480 14523 9482
rect 4061 9424 4066 9480
rect 4122 9424 14462 9480
rect 14518 9424 14523 9480
rect 4061 9422 14523 9424
rect 4061 9419 4127 9422
rect 14457 9419 14523 9422
rect 3545 9280 3861 9281
rect 3545 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3861 9280
rect 3545 9215 3861 9216
rect 8743 9280 9059 9281
rect 8743 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9059 9280
rect 8743 9215 9059 9216
rect 13941 9280 14257 9281
rect 13941 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14257 9280
rect 13941 9215 14257 9216
rect 19139 9280 19455 9281
rect 19139 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19455 9280
rect 19139 9215 19455 9216
rect 0 9074 800 9104
rect 4061 9074 4127 9077
rect 0 9072 4127 9074
rect 0 9016 4066 9072
rect 4122 9016 4127 9072
rect 0 9014 4127 9016
rect 0 8984 800 9014
rect 4061 9011 4127 9014
rect 5165 9074 5231 9077
rect 7649 9074 7715 9077
rect 19793 9074 19859 9077
rect 5165 9072 5274 9074
rect 5165 9016 5170 9072
rect 5226 9016 5274 9072
rect 5165 9011 5274 9016
rect 7649 9072 19859 9074
rect 7649 9016 7654 9072
rect 7710 9016 19798 9072
rect 19854 9016 19859 9072
rect 7649 9014 19859 9016
rect 7649 9011 7715 9014
rect 19793 9011 19859 9014
rect 5214 8938 5274 9011
rect 14365 8938 14431 8941
rect 5214 8936 14431 8938
rect 5214 8880 14370 8936
rect 14426 8880 14431 8936
rect 5214 8878 14431 8880
rect 14365 8875 14431 8878
rect 6144 8736 6460 8737
rect 0 8666 800 8696
rect 6144 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6460 8736
rect 6144 8671 6460 8672
rect 11342 8736 11658 8737
rect 11342 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11658 8736
rect 11342 8671 11658 8672
rect 16540 8736 16856 8737
rect 16540 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16856 8736
rect 16540 8671 16856 8672
rect 21738 8736 22054 8737
rect 21738 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22054 8736
rect 21738 8671 22054 8672
rect 5533 8666 5599 8669
rect 0 8664 5599 8666
rect 0 8608 5538 8664
rect 5594 8608 5599 8664
rect 0 8606 5599 8608
rect 0 8576 800 8606
rect 5533 8603 5599 8606
rect 9397 8668 9463 8669
rect 9397 8664 9444 8668
rect 9508 8666 9514 8668
rect 9397 8608 9402 8664
rect 9397 8604 9444 8608
rect 9508 8606 9554 8666
rect 9508 8604 9514 8606
rect 9397 8603 9463 8604
rect 5441 8530 5507 8533
rect 18505 8530 18571 8533
rect 5441 8528 18571 8530
rect 5441 8472 5446 8528
rect 5502 8472 18510 8528
rect 18566 8472 18571 8528
rect 5441 8470 18571 8472
rect 5441 8467 5507 8470
rect 18505 8467 18571 8470
rect 5901 8394 5967 8397
rect 15653 8394 15719 8397
rect 5901 8392 15719 8394
rect 5901 8336 5906 8392
rect 5962 8336 15658 8392
rect 15714 8336 15719 8392
rect 5901 8334 15719 8336
rect 5901 8331 5967 8334
rect 15653 8331 15719 8334
rect 0 8258 800 8288
rect 3325 8258 3391 8261
rect 0 8256 3391 8258
rect 0 8200 3330 8256
rect 3386 8200 3391 8256
rect 0 8198 3391 8200
rect 0 8168 800 8198
rect 3325 8195 3391 8198
rect 3969 8258 4035 8261
rect 7097 8258 7163 8261
rect 3969 8256 7163 8258
rect 3969 8200 3974 8256
rect 4030 8200 7102 8256
rect 7158 8200 7163 8256
rect 3969 8198 7163 8200
rect 3969 8195 4035 8198
rect 7097 8195 7163 8198
rect 3545 8192 3861 8193
rect 3545 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3861 8192
rect 3545 8127 3861 8128
rect 8743 8192 9059 8193
rect 8743 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9059 8192
rect 8743 8127 9059 8128
rect 13941 8192 14257 8193
rect 13941 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14257 8192
rect 13941 8127 14257 8128
rect 19139 8192 19455 8193
rect 19139 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19455 8192
rect 19139 8127 19455 8128
rect 5533 8122 5599 8125
rect 8293 8122 8359 8125
rect 5533 8120 8359 8122
rect 5533 8064 5538 8120
rect 5594 8064 8298 8120
rect 8354 8064 8359 8120
rect 5533 8062 8359 8064
rect 5533 8059 5599 8062
rect 8293 8059 8359 8062
rect 2405 7986 2471 7989
rect 7833 7986 7899 7989
rect 19057 7986 19123 7989
rect 2405 7984 7666 7986
rect 2405 7928 2410 7984
rect 2466 7928 7666 7984
rect 2405 7926 7666 7928
rect 2405 7923 2471 7926
rect 0 7850 800 7880
rect 3969 7850 4035 7853
rect 0 7848 4035 7850
rect 0 7792 3974 7848
rect 4030 7792 4035 7848
rect 0 7790 4035 7792
rect 0 7760 800 7790
rect 3969 7787 4035 7790
rect 4981 7850 5047 7853
rect 7606 7850 7666 7926
rect 7833 7984 19123 7986
rect 7833 7928 7838 7984
rect 7894 7928 19062 7984
rect 19118 7928 19123 7984
rect 7833 7926 19123 7928
rect 7833 7923 7899 7926
rect 19057 7923 19123 7926
rect 11145 7850 11211 7853
rect 4981 7848 6746 7850
rect 4981 7792 4986 7848
rect 5042 7792 6746 7848
rect 4981 7790 6746 7792
rect 7606 7848 11211 7850
rect 7606 7792 11150 7848
rect 11206 7792 11211 7848
rect 7606 7790 11211 7792
rect 4981 7787 5047 7790
rect 6686 7714 6746 7790
rect 11145 7787 11211 7790
rect 10961 7714 11027 7717
rect 6686 7712 11027 7714
rect 6686 7656 10966 7712
rect 11022 7656 11027 7712
rect 6686 7654 11027 7656
rect 10961 7651 11027 7654
rect 6144 7648 6460 7649
rect 6144 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6460 7648
rect 6144 7583 6460 7584
rect 11342 7648 11658 7649
rect 11342 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11658 7648
rect 11342 7583 11658 7584
rect 16540 7648 16856 7649
rect 16540 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16856 7648
rect 16540 7583 16856 7584
rect 21738 7648 22054 7649
rect 21738 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22054 7648
rect 21738 7583 22054 7584
rect 7833 7578 7899 7581
rect 9305 7578 9371 7581
rect 7833 7576 9371 7578
rect 7833 7520 7838 7576
rect 7894 7520 9310 7576
rect 9366 7520 9371 7576
rect 7833 7518 9371 7520
rect 7833 7515 7899 7518
rect 9305 7515 9371 7518
rect 0 7442 800 7472
rect 3417 7442 3483 7445
rect 0 7440 3483 7442
rect 0 7384 3422 7440
rect 3478 7384 3483 7440
rect 0 7382 3483 7384
rect 0 7352 800 7382
rect 3417 7379 3483 7382
rect 4797 7442 4863 7445
rect 18045 7442 18111 7445
rect 4797 7440 18111 7442
rect 4797 7384 4802 7440
rect 4858 7384 18050 7440
rect 18106 7384 18111 7440
rect 4797 7382 18111 7384
rect 4797 7379 4863 7382
rect 18045 7379 18111 7382
rect 2037 7306 2103 7309
rect 17033 7306 17099 7309
rect 2037 7304 17099 7306
rect 2037 7248 2042 7304
rect 2098 7248 17038 7304
rect 17094 7248 17099 7304
rect 2037 7246 17099 7248
rect 2037 7243 2103 7246
rect 17033 7243 17099 7246
rect 3545 7104 3861 7105
rect 0 7034 800 7064
rect 3545 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3861 7104
rect 3545 7039 3861 7040
rect 8743 7104 9059 7105
rect 8743 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9059 7104
rect 8743 7039 9059 7040
rect 13941 7104 14257 7105
rect 13941 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14257 7104
rect 13941 7039 14257 7040
rect 19139 7104 19455 7105
rect 19139 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19455 7104
rect 19139 7039 19455 7040
rect 3049 7034 3115 7037
rect 0 7032 3115 7034
rect 0 6976 3054 7032
rect 3110 6976 3115 7032
rect 0 6974 3115 6976
rect 0 6944 800 6974
rect 3049 6971 3115 6974
rect 5901 6898 5967 6901
rect 20621 6898 20687 6901
rect 5901 6896 20687 6898
rect 5901 6840 5906 6896
rect 5962 6840 20626 6896
rect 20682 6840 20687 6896
rect 5901 6838 20687 6840
rect 5901 6835 5967 6838
rect 20621 6835 20687 6838
rect 5533 6762 5599 6765
rect 15469 6762 15535 6765
rect 5533 6760 15535 6762
rect 5533 6704 5538 6760
rect 5594 6704 15474 6760
rect 15530 6704 15535 6760
rect 5533 6702 15535 6704
rect 5533 6699 5599 6702
rect 15469 6699 15535 6702
rect 0 6626 800 6656
rect 1669 6626 1735 6629
rect 0 6624 1735 6626
rect 0 6568 1674 6624
rect 1730 6568 1735 6624
rect 0 6566 1735 6568
rect 0 6536 800 6566
rect 1669 6563 1735 6566
rect 6144 6560 6460 6561
rect 6144 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6460 6560
rect 6144 6495 6460 6496
rect 11342 6560 11658 6561
rect 11342 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11658 6560
rect 11342 6495 11658 6496
rect 16540 6560 16856 6561
rect 16540 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16856 6560
rect 16540 6495 16856 6496
rect 21738 6560 22054 6561
rect 21738 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22054 6560
rect 21738 6495 22054 6496
rect 6821 6354 6887 6357
rect 6686 6352 6887 6354
rect 6686 6296 6826 6352
rect 6882 6296 6887 6352
rect 6686 6294 6887 6296
rect 0 6218 800 6248
rect 4153 6218 4219 6221
rect 0 6216 4219 6218
rect 0 6160 4158 6216
rect 4214 6160 4219 6216
rect 0 6158 4219 6160
rect 0 6128 800 6158
rect 4153 6155 4219 6158
rect 6545 6218 6611 6221
rect 6686 6218 6746 6294
rect 6821 6291 6887 6294
rect 6545 6216 6746 6218
rect 6545 6160 6550 6216
rect 6606 6160 6746 6216
rect 6545 6158 6746 6160
rect 6545 6155 6611 6158
rect 3545 6016 3861 6017
rect 3545 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3861 6016
rect 3545 5951 3861 5952
rect 8743 6016 9059 6017
rect 8743 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9059 6016
rect 8743 5951 9059 5952
rect 13941 6016 14257 6017
rect 13941 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14257 6016
rect 13941 5951 14257 5952
rect 19139 6016 19455 6017
rect 19139 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19455 6016
rect 19139 5951 19455 5952
rect 0 5810 800 5840
rect 1669 5810 1735 5813
rect 0 5808 1735 5810
rect 0 5752 1674 5808
rect 1730 5752 1735 5808
rect 0 5750 1735 5752
rect 0 5720 800 5750
rect 1669 5747 1735 5750
rect 10869 5810 10935 5813
rect 22200 5810 23000 5840
rect 10869 5808 23000 5810
rect 10869 5752 10874 5808
rect 10930 5752 23000 5808
rect 10869 5750 23000 5752
rect 10869 5747 10935 5750
rect 22200 5720 23000 5750
rect 2865 5674 2931 5677
rect 3325 5674 3391 5677
rect 2865 5672 3391 5674
rect 2865 5616 2870 5672
rect 2926 5616 3330 5672
rect 3386 5616 3391 5672
rect 2865 5614 3391 5616
rect 2865 5611 2931 5614
rect 3325 5611 3391 5614
rect 4245 5674 4311 5677
rect 8661 5674 8727 5677
rect 4245 5672 8727 5674
rect 4245 5616 4250 5672
rect 4306 5616 8666 5672
rect 8722 5616 8727 5672
rect 4245 5614 8727 5616
rect 4245 5611 4311 5614
rect 8661 5611 8727 5614
rect 6144 5472 6460 5473
rect 0 5402 800 5432
rect 6144 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6460 5472
rect 6144 5407 6460 5408
rect 11342 5472 11658 5473
rect 11342 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11658 5472
rect 11342 5407 11658 5408
rect 16540 5472 16856 5473
rect 16540 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16856 5472
rect 16540 5407 16856 5408
rect 21738 5472 22054 5473
rect 21738 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22054 5472
rect 21738 5407 22054 5408
rect 4061 5402 4127 5405
rect 0 5400 4127 5402
rect 0 5344 4066 5400
rect 4122 5344 4127 5400
rect 0 5342 4127 5344
rect 0 5312 800 5342
rect 4061 5339 4127 5342
rect 0 4994 800 5024
rect 1485 4994 1551 4997
rect 7005 4996 7071 4997
rect 7005 4994 7052 4996
rect 0 4992 1551 4994
rect 0 4936 1490 4992
rect 1546 4936 1551 4992
rect 0 4934 1551 4936
rect 6960 4992 7052 4994
rect 6960 4936 7010 4992
rect 6960 4934 7052 4936
rect 0 4904 800 4934
rect 1485 4931 1551 4934
rect 7005 4932 7052 4934
rect 7116 4932 7122 4996
rect 7005 4931 7071 4932
rect 3545 4928 3861 4929
rect 3545 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3861 4928
rect 3545 4863 3861 4864
rect 8743 4928 9059 4929
rect 8743 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9059 4928
rect 8743 4863 9059 4864
rect 13941 4928 14257 4929
rect 13941 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14257 4928
rect 13941 4863 14257 4864
rect 19139 4928 19455 4929
rect 19139 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19455 4928
rect 19139 4863 19455 4864
rect 7281 4722 7347 4725
rect 17769 4722 17835 4725
rect 7281 4720 17835 4722
rect 7281 4664 7286 4720
rect 7342 4664 17774 4720
rect 17830 4664 17835 4720
rect 7281 4662 17835 4664
rect 7281 4659 7347 4662
rect 17769 4659 17835 4662
rect 0 4586 800 4616
rect 1393 4586 1459 4589
rect 0 4584 1459 4586
rect 0 4528 1398 4584
rect 1454 4528 1459 4584
rect 0 4526 1459 4528
rect 0 4496 800 4526
rect 1393 4523 1459 4526
rect 1853 4586 1919 4589
rect 11697 4586 11763 4589
rect 1853 4584 11763 4586
rect 1853 4528 1858 4584
rect 1914 4528 11702 4584
rect 11758 4528 11763 4584
rect 1853 4526 11763 4528
rect 1853 4523 1919 4526
rect 11697 4523 11763 4526
rect 6144 4384 6460 4385
rect 6144 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6460 4384
rect 6144 4319 6460 4320
rect 11342 4384 11658 4385
rect 11342 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11658 4384
rect 11342 4319 11658 4320
rect 16540 4384 16856 4385
rect 16540 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16856 4384
rect 16540 4319 16856 4320
rect 21738 4384 22054 4385
rect 21738 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22054 4384
rect 21738 4319 22054 4320
rect 0 4178 800 4208
rect 2773 4178 2839 4181
rect 0 4176 2839 4178
rect 0 4120 2778 4176
rect 2834 4120 2839 4176
rect 0 4118 2839 4120
rect 0 4088 800 4118
rect 2773 4115 2839 4118
rect 8293 4178 8359 4181
rect 18045 4178 18111 4181
rect 8293 4176 18111 4178
rect 8293 4120 8298 4176
rect 8354 4120 18050 4176
rect 18106 4120 18111 4176
rect 8293 4118 18111 4120
rect 8293 4115 8359 4118
rect 18045 4115 18111 4118
rect 2313 4042 2379 4045
rect 10409 4042 10475 4045
rect 14273 4042 14339 4045
rect 2313 4040 14339 4042
rect 2313 3984 2318 4040
rect 2374 3984 10414 4040
rect 10470 3984 14278 4040
rect 14334 3984 14339 4040
rect 2313 3982 14339 3984
rect 2313 3979 2379 3982
rect 10409 3979 10475 3982
rect 14273 3979 14339 3982
rect 5574 3844 5580 3908
rect 5644 3906 5650 3908
rect 5993 3906 6059 3909
rect 5644 3904 6059 3906
rect 5644 3848 5998 3904
rect 6054 3848 6059 3904
rect 5644 3846 6059 3848
rect 5644 3844 5650 3846
rect 5993 3843 6059 3846
rect 3545 3840 3861 3841
rect 0 3770 800 3800
rect 3545 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3861 3840
rect 3545 3775 3861 3776
rect 8743 3840 9059 3841
rect 8743 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9059 3840
rect 8743 3775 9059 3776
rect 13941 3840 14257 3841
rect 13941 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14257 3840
rect 13941 3775 14257 3776
rect 19139 3840 19455 3841
rect 19139 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19455 3840
rect 19139 3775 19455 3776
rect 1577 3770 1643 3773
rect 0 3768 1643 3770
rect 0 3712 1582 3768
rect 1638 3712 1643 3768
rect 0 3710 1643 3712
rect 0 3680 800 3710
rect 1577 3707 1643 3710
rect 8334 3572 8340 3636
rect 8404 3634 8410 3636
rect 9121 3634 9187 3637
rect 8404 3632 9187 3634
rect 8404 3576 9126 3632
rect 9182 3576 9187 3632
rect 8404 3574 9187 3576
rect 8404 3572 8410 3574
rect 9121 3571 9187 3574
rect 9581 3634 9647 3637
rect 16757 3634 16823 3637
rect 9581 3632 16823 3634
rect 9581 3576 9586 3632
rect 9642 3576 16762 3632
rect 16818 3576 16823 3632
rect 9581 3574 16823 3576
rect 9581 3571 9647 3574
rect 16757 3571 16823 3574
rect 4797 3498 4863 3501
rect 7465 3498 7531 3501
rect 4797 3496 7531 3498
rect 4797 3440 4802 3496
rect 4858 3440 7470 3496
rect 7526 3440 7531 3496
rect 4797 3438 7531 3440
rect 4797 3435 4863 3438
rect 7465 3435 7531 3438
rect 8385 3498 8451 3501
rect 9254 3498 9260 3500
rect 8385 3496 9260 3498
rect 8385 3440 8390 3496
rect 8446 3440 9260 3496
rect 8385 3438 9260 3440
rect 8385 3435 8451 3438
rect 9254 3436 9260 3438
rect 9324 3436 9330 3500
rect 18137 3498 18203 3501
rect 9446 3496 18203 3498
rect 9446 3440 18142 3496
rect 18198 3440 18203 3496
rect 9446 3438 18203 3440
rect 0 3362 800 3392
rect 3325 3362 3391 3365
rect 0 3360 3391 3362
rect 0 3304 3330 3360
rect 3386 3304 3391 3360
rect 0 3302 3391 3304
rect 0 3272 800 3302
rect 3325 3299 3391 3302
rect 7741 3362 7807 3365
rect 9446 3362 9506 3438
rect 18137 3435 18203 3438
rect 7741 3360 9506 3362
rect 7741 3304 7746 3360
rect 7802 3304 9506 3360
rect 7741 3302 9506 3304
rect 7741 3299 7807 3302
rect 6144 3296 6460 3297
rect 6144 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6460 3296
rect 6144 3231 6460 3232
rect 11342 3296 11658 3297
rect 11342 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11658 3296
rect 11342 3231 11658 3232
rect 16540 3296 16856 3297
rect 16540 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16856 3296
rect 16540 3231 16856 3232
rect 21738 3296 22054 3297
rect 21738 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22054 3296
rect 21738 3231 22054 3232
rect 8753 3226 8819 3229
rect 9213 3226 9279 3229
rect 8753 3224 9279 3226
rect 8753 3168 8758 3224
rect 8814 3168 9218 3224
rect 9274 3168 9279 3224
rect 8753 3166 9279 3168
rect 8753 3163 8819 3166
rect 9213 3163 9279 3166
rect 8150 3028 8156 3092
rect 8220 3090 8226 3092
rect 12801 3090 12867 3093
rect 8220 3088 12867 3090
rect 8220 3032 12806 3088
rect 12862 3032 12867 3088
rect 8220 3030 12867 3032
rect 8220 3028 8226 3030
rect 12801 3027 12867 3030
rect 13077 3090 13143 3093
rect 15561 3090 15627 3093
rect 13077 3088 15627 3090
rect 13077 3032 13082 3088
rect 13138 3032 15566 3088
rect 15622 3032 15627 3088
rect 13077 3030 15627 3032
rect 13077 3027 13143 3030
rect 15561 3027 15627 3030
rect 0 2954 800 2984
rect 1393 2954 1459 2957
rect 0 2952 1459 2954
rect 0 2896 1398 2952
rect 1454 2896 1459 2952
rect 0 2894 1459 2896
rect 0 2864 800 2894
rect 1393 2891 1459 2894
rect 5809 2954 5875 2957
rect 15653 2954 15719 2957
rect 5809 2952 15719 2954
rect 5809 2896 5814 2952
rect 5870 2896 15658 2952
rect 15714 2896 15719 2952
rect 5809 2894 15719 2896
rect 5809 2891 5875 2894
rect 15653 2891 15719 2894
rect 9949 2818 10015 2821
rect 12341 2818 12407 2821
rect 9949 2816 12407 2818
rect 9949 2760 9954 2816
rect 10010 2760 12346 2816
rect 12402 2760 12407 2816
rect 9949 2758 12407 2760
rect 9949 2755 10015 2758
rect 12341 2755 12407 2758
rect 3545 2752 3861 2753
rect 3545 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3861 2752
rect 3545 2687 3861 2688
rect 8743 2752 9059 2753
rect 8743 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9059 2752
rect 8743 2687 9059 2688
rect 13941 2752 14257 2753
rect 13941 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14257 2752
rect 13941 2687 14257 2688
rect 19139 2752 19455 2753
rect 19139 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19455 2752
rect 19139 2687 19455 2688
rect 9673 2682 9739 2685
rect 10593 2682 10659 2685
rect 9673 2680 10659 2682
rect 9673 2624 9678 2680
rect 9734 2624 10598 2680
rect 10654 2624 10659 2680
rect 9673 2622 10659 2624
rect 9673 2619 9739 2622
rect 10593 2619 10659 2622
rect 0 2546 800 2576
rect 2221 2546 2287 2549
rect 0 2544 2287 2546
rect 0 2488 2226 2544
rect 2282 2488 2287 2544
rect 0 2486 2287 2488
rect 0 2456 800 2486
rect 2221 2483 2287 2486
rect 6913 2546 6979 2549
rect 20713 2546 20779 2549
rect 6913 2544 20779 2546
rect 6913 2488 6918 2544
rect 6974 2488 20718 2544
rect 20774 2488 20779 2544
rect 6913 2486 20779 2488
rect 6913 2483 6979 2486
rect 20713 2483 20779 2486
rect 2129 2410 2195 2413
rect 18229 2410 18295 2413
rect 2129 2408 18295 2410
rect 2129 2352 2134 2408
rect 2190 2352 18234 2408
rect 18290 2352 18295 2408
rect 2129 2350 18295 2352
rect 2129 2347 2195 2350
rect 18229 2347 18295 2350
rect 7046 2212 7052 2276
rect 7116 2274 7122 2276
rect 9029 2274 9095 2277
rect 7116 2272 9095 2274
rect 7116 2216 9034 2272
rect 9090 2216 9095 2272
rect 7116 2214 9095 2216
rect 7116 2212 7122 2214
rect 9029 2211 9095 2214
rect 9213 2274 9279 2277
rect 9489 2274 9555 2277
rect 9213 2272 9555 2274
rect 9213 2216 9218 2272
rect 9274 2216 9494 2272
rect 9550 2216 9555 2272
rect 9213 2214 9555 2216
rect 9213 2211 9279 2214
rect 9489 2211 9555 2214
rect 6144 2208 6460 2209
rect 0 2138 800 2168
rect 6144 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6460 2208
rect 6144 2143 6460 2144
rect 11342 2208 11658 2209
rect 11342 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11658 2208
rect 11342 2143 11658 2144
rect 16540 2208 16856 2209
rect 16540 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16856 2208
rect 16540 2143 16856 2144
rect 21738 2208 22054 2209
rect 21738 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22054 2208
rect 21738 2143 22054 2144
rect 3969 2138 4035 2141
rect 9397 2140 9463 2141
rect 9397 2138 9444 2140
rect 0 2136 4035 2138
rect 0 2080 3974 2136
rect 4030 2080 4035 2136
rect 0 2078 4035 2080
rect 9352 2136 9444 2138
rect 9352 2080 9402 2136
rect 9352 2078 9444 2080
rect 0 2048 800 2078
rect 3969 2075 4035 2078
rect 9397 2076 9444 2078
rect 9508 2076 9514 2140
rect 9397 2075 9463 2076
rect 2589 1866 2655 1869
rect 17861 1866 17927 1869
rect 2589 1864 17927 1866
rect 2589 1808 2594 1864
rect 2650 1808 17866 1864
rect 17922 1808 17927 1864
rect 2589 1806 17927 1808
rect 2589 1803 2655 1806
rect 17861 1803 17927 1806
rect 0 1730 800 1760
rect 1209 1730 1275 1733
rect 0 1728 1275 1730
rect 0 1672 1214 1728
rect 1270 1672 1275 1728
rect 0 1670 1275 1672
rect 0 1640 800 1670
rect 1209 1667 1275 1670
rect 2037 1730 2103 1733
rect 19333 1730 19399 1733
rect 2037 1728 19399 1730
rect 2037 1672 2042 1728
rect 2098 1672 19338 1728
rect 19394 1672 19399 1728
rect 2037 1670 19399 1672
rect 2037 1667 2103 1670
rect 19333 1667 19399 1670
<< via3 >>
rect 6150 20700 6214 20704
rect 6150 20644 6154 20700
rect 6154 20644 6210 20700
rect 6210 20644 6214 20700
rect 6150 20640 6214 20644
rect 6230 20700 6294 20704
rect 6230 20644 6234 20700
rect 6234 20644 6290 20700
rect 6290 20644 6294 20700
rect 6230 20640 6294 20644
rect 6310 20700 6374 20704
rect 6310 20644 6314 20700
rect 6314 20644 6370 20700
rect 6370 20644 6374 20700
rect 6310 20640 6374 20644
rect 6390 20700 6454 20704
rect 6390 20644 6394 20700
rect 6394 20644 6450 20700
rect 6450 20644 6454 20700
rect 6390 20640 6454 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 16546 20700 16610 20704
rect 16546 20644 16550 20700
rect 16550 20644 16606 20700
rect 16606 20644 16610 20700
rect 16546 20640 16610 20644
rect 16626 20700 16690 20704
rect 16626 20644 16630 20700
rect 16630 20644 16686 20700
rect 16686 20644 16690 20700
rect 16626 20640 16690 20644
rect 16706 20700 16770 20704
rect 16706 20644 16710 20700
rect 16710 20644 16766 20700
rect 16766 20644 16770 20700
rect 16706 20640 16770 20644
rect 16786 20700 16850 20704
rect 16786 20644 16790 20700
rect 16790 20644 16846 20700
rect 16846 20644 16850 20700
rect 16786 20640 16850 20644
rect 21744 20700 21808 20704
rect 21744 20644 21748 20700
rect 21748 20644 21804 20700
rect 21804 20644 21808 20700
rect 21744 20640 21808 20644
rect 21824 20700 21888 20704
rect 21824 20644 21828 20700
rect 21828 20644 21884 20700
rect 21884 20644 21888 20700
rect 21824 20640 21888 20644
rect 21904 20700 21968 20704
rect 21904 20644 21908 20700
rect 21908 20644 21964 20700
rect 21964 20644 21968 20700
rect 21904 20640 21968 20644
rect 21984 20700 22048 20704
rect 21984 20644 21988 20700
rect 21988 20644 22044 20700
rect 22044 20644 22048 20700
rect 21984 20640 22048 20644
rect 3551 20156 3615 20160
rect 3551 20100 3555 20156
rect 3555 20100 3611 20156
rect 3611 20100 3615 20156
rect 3551 20096 3615 20100
rect 3631 20156 3695 20160
rect 3631 20100 3635 20156
rect 3635 20100 3691 20156
rect 3691 20100 3695 20156
rect 3631 20096 3695 20100
rect 3711 20156 3775 20160
rect 3711 20100 3715 20156
rect 3715 20100 3771 20156
rect 3771 20100 3775 20156
rect 3711 20096 3775 20100
rect 3791 20156 3855 20160
rect 3791 20100 3795 20156
rect 3795 20100 3851 20156
rect 3851 20100 3855 20156
rect 3791 20096 3855 20100
rect 8749 20156 8813 20160
rect 8749 20100 8753 20156
rect 8753 20100 8809 20156
rect 8809 20100 8813 20156
rect 8749 20096 8813 20100
rect 8829 20156 8893 20160
rect 8829 20100 8833 20156
rect 8833 20100 8889 20156
rect 8889 20100 8893 20156
rect 8829 20096 8893 20100
rect 8909 20156 8973 20160
rect 8909 20100 8913 20156
rect 8913 20100 8969 20156
rect 8969 20100 8973 20156
rect 8909 20096 8973 20100
rect 8989 20156 9053 20160
rect 8989 20100 8993 20156
rect 8993 20100 9049 20156
rect 9049 20100 9053 20156
rect 8989 20096 9053 20100
rect 13947 20156 14011 20160
rect 13947 20100 13951 20156
rect 13951 20100 14007 20156
rect 14007 20100 14011 20156
rect 13947 20096 14011 20100
rect 14027 20156 14091 20160
rect 14027 20100 14031 20156
rect 14031 20100 14087 20156
rect 14087 20100 14091 20156
rect 14027 20096 14091 20100
rect 14107 20156 14171 20160
rect 14107 20100 14111 20156
rect 14111 20100 14167 20156
rect 14167 20100 14171 20156
rect 14107 20096 14171 20100
rect 14187 20156 14251 20160
rect 14187 20100 14191 20156
rect 14191 20100 14247 20156
rect 14247 20100 14251 20156
rect 14187 20096 14251 20100
rect 19145 20156 19209 20160
rect 19145 20100 19149 20156
rect 19149 20100 19205 20156
rect 19205 20100 19209 20156
rect 19145 20096 19209 20100
rect 19225 20156 19289 20160
rect 19225 20100 19229 20156
rect 19229 20100 19285 20156
rect 19285 20100 19289 20156
rect 19225 20096 19289 20100
rect 19305 20156 19369 20160
rect 19305 20100 19309 20156
rect 19309 20100 19365 20156
rect 19365 20100 19369 20156
rect 19305 20096 19369 20100
rect 19385 20156 19449 20160
rect 19385 20100 19389 20156
rect 19389 20100 19445 20156
rect 19445 20100 19449 20156
rect 19385 20096 19449 20100
rect 6150 19612 6214 19616
rect 6150 19556 6154 19612
rect 6154 19556 6210 19612
rect 6210 19556 6214 19612
rect 6150 19552 6214 19556
rect 6230 19612 6294 19616
rect 6230 19556 6234 19612
rect 6234 19556 6290 19612
rect 6290 19556 6294 19612
rect 6230 19552 6294 19556
rect 6310 19612 6374 19616
rect 6310 19556 6314 19612
rect 6314 19556 6370 19612
rect 6370 19556 6374 19612
rect 6310 19552 6374 19556
rect 6390 19612 6454 19616
rect 6390 19556 6394 19612
rect 6394 19556 6450 19612
rect 6450 19556 6454 19612
rect 6390 19552 6454 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 16546 19612 16610 19616
rect 16546 19556 16550 19612
rect 16550 19556 16606 19612
rect 16606 19556 16610 19612
rect 16546 19552 16610 19556
rect 16626 19612 16690 19616
rect 16626 19556 16630 19612
rect 16630 19556 16686 19612
rect 16686 19556 16690 19612
rect 16626 19552 16690 19556
rect 16706 19612 16770 19616
rect 16706 19556 16710 19612
rect 16710 19556 16766 19612
rect 16766 19556 16770 19612
rect 16706 19552 16770 19556
rect 16786 19612 16850 19616
rect 16786 19556 16790 19612
rect 16790 19556 16846 19612
rect 16846 19556 16850 19612
rect 16786 19552 16850 19556
rect 21744 19612 21808 19616
rect 21744 19556 21748 19612
rect 21748 19556 21804 19612
rect 21804 19556 21808 19612
rect 21744 19552 21808 19556
rect 21824 19612 21888 19616
rect 21824 19556 21828 19612
rect 21828 19556 21884 19612
rect 21884 19556 21888 19612
rect 21824 19552 21888 19556
rect 21904 19612 21968 19616
rect 21904 19556 21908 19612
rect 21908 19556 21964 19612
rect 21964 19556 21968 19612
rect 21904 19552 21968 19556
rect 21984 19612 22048 19616
rect 21984 19556 21988 19612
rect 21988 19556 22044 19612
rect 22044 19556 22048 19612
rect 21984 19552 22048 19556
rect 3551 19068 3615 19072
rect 3551 19012 3555 19068
rect 3555 19012 3611 19068
rect 3611 19012 3615 19068
rect 3551 19008 3615 19012
rect 3631 19068 3695 19072
rect 3631 19012 3635 19068
rect 3635 19012 3691 19068
rect 3691 19012 3695 19068
rect 3631 19008 3695 19012
rect 3711 19068 3775 19072
rect 3711 19012 3715 19068
rect 3715 19012 3771 19068
rect 3771 19012 3775 19068
rect 3711 19008 3775 19012
rect 3791 19068 3855 19072
rect 3791 19012 3795 19068
rect 3795 19012 3851 19068
rect 3851 19012 3855 19068
rect 3791 19008 3855 19012
rect 8749 19068 8813 19072
rect 8749 19012 8753 19068
rect 8753 19012 8809 19068
rect 8809 19012 8813 19068
rect 8749 19008 8813 19012
rect 8829 19068 8893 19072
rect 8829 19012 8833 19068
rect 8833 19012 8889 19068
rect 8889 19012 8893 19068
rect 8829 19008 8893 19012
rect 8909 19068 8973 19072
rect 8909 19012 8913 19068
rect 8913 19012 8969 19068
rect 8969 19012 8973 19068
rect 8909 19008 8973 19012
rect 8989 19068 9053 19072
rect 8989 19012 8993 19068
rect 8993 19012 9049 19068
rect 9049 19012 9053 19068
rect 8989 19008 9053 19012
rect 13947 19068 14011 19072
rect 13947 19012 13951 19068
rect 13951 19012 14007 19068
rect 14007 19012 14011 19068
rect 13947 19008 14011 19012
rect 14027 19068 14091 19072
rect 14027 19012 14031 19068
rect 14031 19012 14087 19068
rect 14087 19012 14091 19068
rect 14027 19008 14091 19012
rect 14107 19068 14171 19072
rect 14107 19012 14111 19068
rect 14111 19012 14167 19068
rect 14167 19012 14171 19068
rect 14107 19008 14171 19012
rect 14187 19068 14251 19072
rect 14187 19012 14191 19068
rect 14191 19012 14247 19068
rect 14247 19012 14251 19068
rect 14187 19008 14251 19012
rect 19145 19068 19209 19072
rect 19145 19012 19149 19068
rect 19149 19012 19205 19068
rect 19205 19012 19209 19068
rect 19145 19008 19209 19012
rect 19225 19068 19289 19072
rect 19225 19012 19229 19068
rect 19229 19012 19285 19068
rect 19285 19012 19289 19068
rect 19225 19008 19289 19012
rect 19305 19068 19369 19072
rect 19305 19012 19309 19068
rect 19309 19012 19365 19068
rect 19365 19012 19369 19068
rect 19305 19008 19369 19012
rect 19385 19068 19449 19072
rect 19385 19012 19389 19068
rect 19389 19012 19445 19068
rect 19445 19012 19449 19068
rect 19385 19008 19449 19012
rect 6150 18524 6214 18528
rect 6150 18468 6154 18524
rect 6154 18468 6210 18524
rect 6210 18468 6214 18524
rect 6150 18464 6214 18468
rect 6230 18524 6294 18528
rect 6230 18468 6234 18524
rect 6234 18468 6290 18524
rect 6290 18468 6294 18524
rect 6230 18464 6294 18468
rect 6310 18524 6374 18528
rect 6310 18468 6314 18524
rect 6314 18468 6370 18524
rect 6370 18468 6374 18524
rect 6310 18464 6374 18468
rect 6390 18524 6454 18528
rect 6390 18468 6394 18524
rect 6394 18468 6450 18524
rect 6450 18468 6454 18524
rect 6390 18464 6454 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 16546 18524 16610 18528
rect 16546 18468 16550 18524
rect 16550 18468 16606 18524
rect 16606 18468 16610 18524
rect 16546 18464 16610 18468
rect 16626 18524 16690 18528
rect 16626 18468 16630 18524
rect 16630 18468 16686 18524
rect 16686 18468 16690 18524
rect 16626 18464 16690 18468
rect 16706 18524 16770 18528
rect 16706 18468 16710 18524
rect 16710 18468 16766 18524
rect 16766 18468 16770 18524
rect 16706 18464 16770 18468
rect 16786 18524 16850 18528
rect 16786 18468 16790 18524
rect 16790 18468 16846 18524
rect 16846 18468 16850 18524
rect 16786 18464 16850 18468
rect 21744 18524 21808 18528
rect 21744 18468 21748 18524
rect 21748 18468 21804 18524
rect 21804 18468 21808 18524
rect 21744 18464 21808 18468
rect 21824 18524 21888 18528
rect 21824 18468 21828 18524
rect 21828 18468 21884 18524
rect 21884 18468 21888 18524
rect 21824 18464 21888 18468
rect 21904 18524 21968 18528
rect 21904 18468 21908 18524
rect 21908 18468 21964 18524
rect 21964 18468 21968 18524
rect 21904 18464 21968 18468
rect 21984 18524 22048 18528
rect 21984 18468 21988 18524
rect 21988 18468 22044 18524
rect 22044 18468 22048 18524
rect 21984 18464 22048 18468
rect 3551 17980 3615 17984
rect 3551 17924 3555 17980
rect 3555 17924 3611 17980
rect 3611 17924 3615 17980
rect 3551 17920 3615 17924
rect 3631 17980 3695 17984
rect 3631 17924 3635 17980
rect 3635 17924 3691 17980
rect 3691 17924 3695 17980
rect 3631 17920 3695 17924
rect 3711 17980 3775 17984
rect 3711 17924 3715 17980
rect 3715 17924 3771 17980
rect 3771 17924 3775 17980
rect 3711 17920 3775 17924
rect 3791 17980 3855 17984
rect 3791 17924 3795 17980
rect 3795 17924 3851 17980
rect 3851 17924 3855 17980
rect 3791 17920 3855 17924
rect 8749 17980 8813 17984
rect 8749 17924 8753 17980
rect 8753 17924 8809 17980
rect 8809 17924 8813 17980
rect 8749 17920 8813 17924
rect 8829 17980 8893 17984
rect 8829 17924 8833 17980
rect 8833 17924 8889 17980
rect 8889 17924 8893 17980
rect 8829 17920 8893 17924
rect 8909 17980 8973 17984
rect 8909 17924 8913 17980
rect 8913 17924 8969 17980
rect 8969 17924 8973 17980
rect 8909 17920 8973 17924
rect 8989 17980 9053 17984
rect 8989 17924 8993 17980
rect 8993 17924 9049 17980
rect 9049 17924 9053 17980
rect 8989 17920 9053 17924
rect 13947 17980 14011 17984
rect 13947 17924 13951 17980
rect 13951 17924 14007 17980
rect 14007 17924 14011 17980
rect 13947 17920 14011 17924
rect 14027 17980 14091 17984
rect 14027 17924 14031 17980
rect 14031 17924 14087 17980
rect 14087 17924 14091 17980
rect 14027 17920 14091 17924
rect 14107 17980 14171 17984
rect 14107 17924 14111 17980
rect 14111 17924 14167 17980
rect 14167 17924 14171 17980
rect 14107 17920 14171 17924
rect 14187 17980 14251 17984
rect 14187 17924 14191 17980
rect 14191 17924 14247 17980
rect 14247 17924 14251 17980
rect 14187 17920 14251 17924
rect 19145 17980 19209 17984
rect 19145 17924 19149 17980
rect 19149 17924 19205 17980
rect 19205 17924 19209 17980
rect 19145 17920 19209 17924
rect 19225 17980 19289 17984
rect 19225 17924 19229 17980
rect 19229 17924 19285 17980
rect 19285 17924 19289 17980
rect 19225 17920 19289 17924
rect 19305 17980 19369 17984
rect 19305 17924 19309 17980
rect 19309 17924 19365 17980
rect 19365 17924 19369 17980
rect 19305 17920 19369 17924
rect 19385 17980 19449 17984
rect 19385 17924 19389 17980
rect 19389 17924 19445 17980
rect 19445 17924 19449 17980
rect 19385 17920 19449 17924
rect 6150 17436 6214 17440
rect 6150 17380 6154 17436
rect 6154 17380 6210 17436
rect 6210 17380 6214 17436
rect 6150 17376 6214 17380
rect 6230 17436 6294 17440
rect 6230 17380 6234 17436
rect 6234 17380 6290 17436
rect 6290 17380 6294 17436
rect 6230 17376 6294 17380
rect 6310 17436 6374 17440
rect 6310 17380 6314 17436
rect 6314 17380 6370 17436
rect 6370 17380 6374 17436
rect 6310 17376 6374 17380
rect 6390 17436 6454 17440
rect 6390 17380 6394 17436
rect 6394 17380 6450 17436
rect 6450 17380 6454 17436
rect 6390 17376 6454 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 16546 17436 16610 17440
rect 16546 17380 16550 17436
rect 16550 17380 16606 17436
rect 16606 17380 16610 17436
rect 16546 17376 16610 17380
rect 16626 17436 16690 17440
rect 16626 17380 16630 17436
rect 16630 17380 16686 17436
rect 16686 17380 16690 17436
rect 16626 17376 16690 17380
rect 16706 17436 16770 17440
rect 16706 17380 16710 17436
rect 16710 17380 16766 17436
rect 16766 17380 16770 17436
rect 16706 17376 16770 17380
rect 16786 17436 16850 17440
rect 16786 17380 16790 17436
rect 16790 17380 16846 17436
rect 16846 17380 16850 17436
rect 16786 17376 16850 17380
rect 21744 17436 21808 17440
rect 21744 17380 21748 17436
rect 21748 17380 21804 17436
rect 21804 17380 21808 17436
rect 21744 17376 21808 17380
rect 21824 17436 21888 17440
rect 21824 17380 21828 17436
rect 21828 17380 21884 17436
rect 21884 17380 21888 17436
rect 21824 17376 21888 17380
rect 21904 17436 21968 17440
rect 21904 17380 21908 17436
rect 21908 17380 21964 17436
rect 21964 17380 21968 17436
rect 21904 17376 21968 17380
rect 21984 17436 22048 17440
rect 21984 17380 21988 17436
rect 21988 17380 22044 17436
rect 22044 17380 22048 17436
rect 21984 17376 22048 17380
rect 3551 16892 3615 16896
rect 3551 16836 3555 16892
rect 3555 16836 3611 16892
rect 3611 16836 3615 16892
rect 3551 16832 3615 16836
rect 3631 16892 3695 16896
rect 3631 16836 3635 16892
rect 3635 16836 3691 16892
rect 3691 16836 3695 16892
rect 3631 16832 3695 16836
rect 3711 16892 3775 16896
rect 3711 16836 3715 16892
rect 3715 16836 3771 16892
rect 3771 16836 3775 16892
rect 3711 16832 3775 16836
rect 3791 16892 3855 16896
rect 3791 16836 3795 16892
rect 3795 16836 3851 16892
rect 3851 16836 3855 16892
rect 3791 16832 3855 16836
rect 8749 16892 8813 16896
rect 8749 16836 8753 16892
rect 8753 16836 8809 16892
rect 8809 16836 8813 16892
rect 8749 16832 8813 16836
rect 8829 16892 8893 16896
rect 8829 16836 8833 16892
rect 8833 16836 8889 16892
rect 8889 16836 8893 16892
rect 8829 16832 8893 16836
rect 8909 16892 8973 16896
rect 8909 16836 8913 16892
rect 8913 16836 8969 16892
rect 8969 16836 8973 16892
rect 8909 16832 8973 16836
rect 8989 16892 9053 16896
rect 8989 16836 8993 16892
rect 8993 16836 9049 16892
rect 9049 16836 9053 16892
rect 8989 16832 9053 16836
rect 13947 16892 14011 16896
rect 13947 16836 13951 16892
rect 13951 16836 14007 16892
rect 14007 16836 14011 16892
rect 13947 16832 14011 16836
rect 14027 16892 14091 16896
rect 14027 16836 14031 16892
rect 14031 16836 14087 16892
rect 14087 16836 14091 16892
rect 14027 16832 14091 16836
rect 14107 16892 14171 16896
rect 14107 16836 14111 16892
rect 14111 16836 14167 16892
rect 14167 16836 14171 16892
rect 14107 16832 14171 16836
rect 14187 16892 14251 16896
rect 14187 16836 14191 16892
rect 14191 16836 14247 16892
rect 14247 16836 14251 16892
rect 14187 16832 14251 16836
rect 19145 16892 19209 16896
rect 19145 16836 19149 16892
rect 19149 16836 19205 16892
rect 19205 16836 19209 16892
rect 19145 16832 19209 16836
rect 19225 16892 19289 16896
rect 19225 16836 19229 16892
rect 19229 16836 19285 16892
rect 19285 16836 19289 16892
rect 19225 16832 19289 16836
rect 19305 16892 19369 16896
rect 19305 16836 19309 16892
rect 19309 16836 19365 16892
rect 19365 16836 19369 16892
rect 19305 16832 19369 16836
rect 19385 16892 19449 16896
rect 19385 16836 19389 16892
rect 19389 16836 19445 16892
rect 19445 16836 19449 16892
rect 19385 16832 19449 16836
rect 6150 16348 6214 16352
rect 6150 16292 6154 16348
rect 6154 16292 6210 16348
rect 6210 16292 6214 16348
rect 6150 16288 6214 16292
rect 6230 16348 6294 16352
rect 6230 16292 6234 16348
rect 6234 16292 6290 16348
rect 6290 16292 6294 16348
rect 6230 16288 6294 16292
rect 6310 16348 6374 16352
rect 6310 16292 6314 16348
rect 6314 16292 6370 16348
rect 6370 16292 6374 16348
rect 6310 16288 6374 16292
rect 6390 16348 6454 16352
rect 6390 16292 6394 16348
rect 6394 16292 6450 16348
rect 6450 16292 6454 16348
rect 6390 16288 6454 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 16546 16348 16610 16352
rect 16546 16292 16550 16348
rect 16550 16292 16606 16348
rect 16606 16292 16610 16348
rect 16546 16288 16610 16292
rect 16626 16348 16690 16352
rect 16626 16292 16630 16348
rect 16630 16292 16686 16348
rect 16686 16292 16690 16348
rect 16626 16288 16690 16292
rect 16706 16348 16770 16352
rect 16706 16292 16710 16348
rect 16710 16292 16766 16348
rect 16766 16292 16770 16348
rect 16706 16288 16770 16292
rect 16786 16348 16850 16352
rect 16786 16292 16790 16348
rect 16790 16292 16846 16348
rect 16846 16292 16850 16348
rect 16786 16288 16850 16292
rect 21744 16348 21808 16352
rect 21744 16292 21748 16348
rect 21748 16292 21804 16348
rect 21804 16292 21808 16348
rect 21744 16288 21808 16292
rect 21824 16348 21888 16352
rect 21824 16292 21828 16348
rect 21828 16292 21884 16348
rect 21884 16292 21888 16348
rect 21824 16288 21888 16292
rect 21904 16348 21968 16352
rect 21904 16292 21908 16348
rect 21908 16292 21964 16348
rect 21964 16292 21968 16348
rect 21904 16288 21968 16292
rect 21984 16348 22048 16352
rect 21984 16292 21988 16348
rect 21988 16292 22044 16348
rect 22044 16292 22048 16348
rect 21984 16288 22048 16292
rect 3551 15804 3615 15808
rect 3551 15748 3555 15804
rect 3555 15748 3611 15804
rect 3611 15748 3615 15804
rect 3551 15744 3615 15748
rect 3631 15804 3695 15808
rect 3631 15748 3635 15804
rect 3635 15748 3691 15804
rect 3691 15748 3695 15804
rect 3631 15744 3695 15748
rect 3711 15804 3775 15808
rect 3711 15748 3715 15804
rect 3715 15748 3771 15804
rect 3771 15748 3775 15804
rect 3711 15744 3775 15748
rect 3791 15804 3855 15808
rect 3791 15748 3795 15804
rect 3795 15748 3851 15804
rect 3851 15748 3855 15804
rect 3791 15744 3855 15748
rect 8749 15804 8813 15808
rect 8749 15748 8753 15804
rect 8753 15748 8809 15804
rect 8809 15748 8813 15804
rect 8749 15744 8813 15748
rect 8829 15804 8893 15808
rect 8829 15748 8833 15804
rect 8833 15748 8889 15804
rect 8889 15748 8893 15804
rect 8829 15744 8893 15748
rect 8909 15804 8973 15808
rect 8909 15748 8913 15804
rect 8913 15748 8969 15804
rect 8969 15748 8973 15804
rect 8909 15744 8973 15748
rect 8989 15804 9053 15808
rect 8989 15748 8993 15804
rect 8993 15748 9049 15804
rect 9049 15748 9053 15804
rect 8989 15744 9053 15748
rect 13947 15804 14011 15808
rect 13947 15748 13951 15804
rect 13951 15748 14007 15804
rect 14007 15748 14011 15804
rect 13947 15744 14011 15748
rect 14027 15804 14091 15808
rect 14027 15748 14031 15804
rect 14031 15748 14087 15804
rect 14087 15748 14091 15804
rect 14027 15744 14091 15748
rect 14107 15804 14171 15808
rect 14107 15748 14111 15804
rect 14111 15748 14167 15804
rect 14167 15748 14171 15804
rect 14107 15744 14171 15748
rect 14187 15804 14251 15808
rect 14187 15748 14191 15804
rect 14191 15748 14247 15804
rect 14247 15748 14251 15804
rect 14187 15744 14251 15748
rect 19145 15804 19209 15808
rect 19145 15748 19149 15804
rect 19149 15748 19205 15804
rect 19205 15748 19209 15804
rect 19145 15744 19209 15748
rect 19225 15804 19289 15808
rect 19225 15748 19229 15804
rect 19229 15748 19285 15804
rect 19285 15748 19289 15804
rect 19225 15744 19289 15748
rect 19305 15804 19369 15808
rect 19305 15748 19309 15804
rect 19309 15748 19365 15804
rect 19365 15748 19369 15804
rect 19305 15744 19369 15748
rect 19385 15804 19449 15808
rect 19385 15748 19389 15804
rect 19389 15748 19445 15804
rect 19445 15748 19449 15804
rect 19385 15744 19449 15748
rect 6150 15260 6214 15264
rect 6150 15204 6154 15260
rect 6154 15204 6210 15260
rect 6210 15204 6214 15260
rect 6150 15200 6214 15204
rect 6230 15260 6294 15264
rect 6230 15204 6234 15260
rect 6234 15204 6290 15260
rect 6290 15204 6294 15260
rect 6230 15200 6294 15204
rect 6310 15260 6374 15264
rect 6310 15204 6314 15260
rect 6314 15204 6370 15260
rect 6370 15204 6374 15260
rect 6310 15200 6374 15204
rect 6390 15260 6454 15264
rect 6390 15204 6394 15260
rect 6394 15204 6450 15260
rect 6450 15204 6454 15260
rect 6390 15200 6454 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 16546 15260 16610 15264
rect 16546 15204 16550 15260
rect 16550 15204 16606 15260
rect 16606 15204 16610 15260
rect 16546 15200 16610 15204
rect 16626 15260 16690 15264
rect 16626 15204 16630 15260
rect 16630 15204 16686 15260
rect 16686 15204 16690 15260
rect 16626 15200 16690 15204
rect 16706 15260 16770 15264
rect 16706 15204 16710 15260
rect 16710 15204 16766 15260
rect 16766 15204 16770 15260
rect 16706 15200 16770 15204
rect 16786 15260 16850 15264
rect 16786 15204 16790 15260
rect 16790 15204 16846 15260
rect 16846 15204 16850 15260
rect 16786 15200 16850 15204
rect 21744 15260 21808 15264
rect 21744 15204 21748 15260
rect 21748 15204 21804 15260
rect 21804 15204 21808 15260
rect 21744 15200 21808 15204
rect 21824 15260 21888 15264
rect 21824 15204 21828 15260
rect 21828 15204 21884 15260
rect 21884 15204 21888 15260
rect 21824 15200 21888 15204
rect 21904 15260 21968 15264
rect 21904 15204 21908 15260
rect 21908 15204 21964 15260
rect 21964 15204 21968 15260
rect 21904 15200 21968 15204
rect 21984 15260 22048 15264
rect 21984 15204 21988 15260
rect 21988 15204 22044 15260
rect 22044 15204 22048 15260
rect 21984 15200 22048 15204
rect 3551 14716 3615 14720
rect 3551 14660 3555 14716
rect 3555 14660 3611 14716
rect 3611 14660 3615 14716
rect 3551 14656 3615 14660
rect 3631 14716 3695 14720
rect 3631 14660 3635 14716
rect 3635 14660 3691 14716
rect 3691 14660 3695 14716
rect 3631 14656 3695 14660
rect 3711 14716 3775 14720
rect 3711 14660 3715 14716
rect 3715 14660 3771 14716
rect 3771 14660 3775 14716
rect 3711 14656 3775 14660
rect 3791 14716 3855 14720
rect 3791 14660 3795 14716
rect 3795 14660 3851 14716
rect 3851 14660 3855 14716
rect 3791 14656 3855 14660
rect 8749 14716 8813 14720
rect 8749 14660 8753 14716
rect 8753 14660 8809 14716
rect 8809 14660 8813 14716
rect 8749 14656 8813 14660
rect 8829 14716 8893 14720
rect 8829 14660 8833 14716
rect 8833 14660 8889 14716
rect 8889 14660 8893 14716
rect 8829 14656 8893 14660
rect 8909 14716 8973 14720
rect 8909 14660 8913 14716
rect 8913 14660 8969 14716
rect 8969 14660 8973 14716
rect 8909 14656 8973 14660
rect 8989 14716 9053 14720
rect 8989 14660 8993 14716
rect 8993 14660 9049 14716
rect 9049 14660 9053 14716
rect 8989 14656 9053 14660
rect 13947 14716 14011 14720
rect 13947 14660 13951 14716
rect 13951 14660 14007 14716
rect 14007 14660 14011 14716
rect 13947 14656 14011 14660
rect 14027 14716 14091 14720
rect 14027 14660 14031 14716
rect 14031 14660 14087 14716
rect 14087 14660 14091 14716
rect 14027 14656 14091 14660
rect 14107 14716 14171 14720
rect 14107 14660 14111 14716
rect 14111 14660 14167 14716
rect 14167 14660 14171 14716
rect 14107 14656 14171 14660
rect 14187 14716 14251 14720
rect 14187 14660 14191 14716
rect 14191 14660 14247 14716
rect 14247 14660 14251 14716
rect 14187 14656 14251 14660
rect 19145 14716 19209 14720
rect 19145 14660 19149 14716
rect 19149 14660 19205 14716
rect 19205 14660 19209 14716
rect 19145 14656 19209 14660
rect 19225 14716 19289 14720
rect 19225 14660 19229 14716
rect 19229 14660 19285 14716
rect 19285 14660 19289 14716
rect 19225 14656 19289 14660
rect 19305 14716 19369 14720
rect 19305 14660 19309 14716
rect 19309 14660 19365 14716
rect 19365 14660 19369 14716
rect 19305 14656 19369 14660
rect 19385 14716 19449 14720
rect 19385 14660 19389 14716
rect 19389 14660 19445 14716
rect 19445 14660 19449 14716
rect 19385 14656 19449 14660
rect 6150 14172 6214 14176
rect 6150 14116 6154 14172
rect 6154 14116 6210 14172
rect 6210 14116 6214 14172
rect 6150 14112 6214 14116
rect 6230 14172 6294 14176
rect 6230 14116 6234 14172
rect 6234 14116 6290 14172
rect 6290 14116 6294 14172
rect 6230 14112 6294 14116
rect 6310 14172 6374 14176
rect 6310 14116 6314 14172
rect 6314 14116 6370 14172
rect 6370 14116 6374 14172
rect 6310 14112 6374 14116
rect 6390 14172 6454 14176
rect 6390 14116 6394 14172
rect 6394 14116 6450 14172
rect 6450 14116 6454 14172
rect 6390 14112 6454 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 16546 14172 16610 14176
rect 16546 14116 16550 14172
rect 16550 14116 16606 14172
rect 16606 14116 16610 14172
rect 16546 14112 16610 14116
rect 16626 14172 16690 14176
rect 16626 14116 16630 14172
rect 16630 14116 16686 14172
rect 16686 14116 16690 14172
rect 16626 14112 16690 14116
rect 16706 14172 16770 14176
rect 16706 14116 16710 14172
rect 16710 14116 16766 14172
rect 16766 14116 16770 14172
rect 16706 14112 16770 14116
rect 16786 14172 16850 14176
rect 16786 14116 16790 14172
rect 16790 14116 16846 14172
rect 16846 14116 16850 14172
rect 16786 14112 16850 14116
rect 21744 14172 21808 14176
rect 21744 14116 21748 14172
rect 21748 14116 21804 14172
rect 21804 14116 21808 14172
rect 21744 14112 21808 14116
rect 21824 14172 21888 14176
rect 21824 14116 21828 14172
rect 21828 14116 21884 14172
rect 21884 14116 21888 14172
rect 21824 14112 21888 14116
rect 21904 14172 21968 14176
rect 21904 14116 21908 14172
rect 21908 14116 21964 14172
rect 21964 14116 21968 14172
rect 21904 14112 21968 14116
rect 21984 14172 22048 14176
rect 21984 14116 21988 14172
rect 21988 14116 22044 14172
rect 22044 14116 22048 14172
rect 21984 14112 22048 14116
rect 8340 13908 8404 13972
rect 9260 13772 9324 13836
rect 3551 13628 3615 13632
rect 3551 13572 3555 13628
rect 3555 13572 3611 13628
rect 3611 13572 3615 13628
rect 3551 13568 3615 13572
rect 3631 13628 3695 13632
rect 3631 13572 3635 13628
rect 3635 13572 3691 13628
rect 3691 13572 3695 13628
rect 3631 13568 3695 13572
rect 3711 13628 3775 13632
rect 3711 13572 3715 13628
rect 3715 13572 3771 13628
rect 3771 13572 3775 13628
rect 3711 13568 3775 13572
rect 3791 13628 3855 13632
rect 3791 13572 3795 13628
rect 3795 13572 3851 13628
rect 3851 13572 3855 13628
rect 3791 13568 3855 13572
rect 8749 13628 8813 13632
rect 8749 13572 8753 13628
rect 8753 13572 8809 13628
rect 8809 13572 8813 13628
rect 8749 13568 8813 13572
rect 8829 13628 8893 13632
rect 8829 13572 8833 13628
rect 8833 13572 8889 13628
rect 8889 13572 8893 13628
rect 8829 13568 8893 13572
rect 8909 13628 8973 13632
rect 8909 13572 8913 13628
rect 8913 13572 8969 13628
rect 8969 13572 8973 13628
rect 8909 13568 8973 13572
rect 8989 13628 9053 13632
rect 8989 13572 8993 13628
rect 8993 13572 9049 13628
rect 9049 13572 9053 13628
rect 8989 13568 9053 13572
rect 13947 13628 14011 13632
rect 13947 13572 13951 13628
rect 13951 13572 14007 13628
rect 14007 13572 14011 13628
rect 13947 13568 14011 13572
rect 14027 13628 14091 13632
rect 14027 13572 14031 13628
rect 14031 13572 14087 13628
rect 14087 13572 14091 13628
rect 14027 13568 14091 13572
rect 14107 13628 14171 13632
rect 14107 13572 14111 13628
rect 14111 13572 14167 13628
rect 14167 13572 14171 13628
rect 14107 13568 14171 13572
rect 14187 13628 14251 13632
rect 14187 13572 14191 13628
rect 14191 13572 14247 13628
rect 14247 13572 14251 13628
rect 14187 13568 14251 13572
rect 19145 13628 19209 13632
rect 19145 13572 19149 13628
rect 19149 13572 19205 13628
rect 19205 13572 19209 13628
rect 19145 13568 19209 13572
rect 19225 13628 19289 13632
rect 19225 13572 19229 13628
rect 19229 13572 19285 13628
rect 19285 13572 19289 13628
rect 19225 13568 19289 13572
rect 19305 13628 19369 13632
rect 19305 13572 19309 13628
rect 19309 13572 19365 13628
rect 19365 13572 19369 13628
rect 19305 13568 19369 13572
rect 19385 13628 19449 13632
rect 19385 13572 19389 13628
rect 19389 13572 19445 13628
rect 19445 13572 19449 13628
rect 19385 13568 19449 13572
rect 6150 13084 6214 13088
rect 6150 13028 6154 13084
rect 6154 13028 6210 13084
rect 6210 13028 6214 13084
rect 6150 13024 6214 13028
rect 6230 13084 6294 13088
rect 6230 13028 6234 13084
rect 6234 13028 6290 13084
rect 6290 13028 6294 13084
rect 6230 13024 6294 13028
rect 6310 13084 6374 13088
rect 6310 13028 6314 13084
rect 6314 13028 6370 13084
rect 6370 13028 6374 13084
rect 6310 13024 6374 13028
rect 6390 13084 6454 13088
rect 6390 13028 6394 13084
rect 6394 13028 6450 13084
rect 6450 13028 6454 13084
rect 6390 13024 6454 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 16546 13084 16610 13088
rect 16546 13028 16550 13084
rect 16550 13028 16606 13084
rect 16606 13028 16610 13084
rect 16546 13024 16610 13028
rect 16626 13084 16690 13088
rect 16626 13028 16630 13084
rect 16630 13028 16686 13084
rect 16686 13028 16690 13084
rect 16626 13024 16690 13028
rect 16706 13084 16770 13088
rect 16706 13028 16710 13084
rect 16710 13028 16766 13084
rect 16766 13028 16770 13084
rect 16706 13024 16770 13028
rect 16786 13084 16850 13088
rect 16786 13028 16790 13084
rect 16790 13028 16846 13084
rect 16846 13028 16850 13084
rect 16786 13024 16850 13028
rect 21744 13084 21808 13088
rect 21744 13028 21748 13084
rect 21748 13028 21804 13084
rect 21804 13028 21808 13084
rect 21744 13024 21808 13028
rect 21824 13084 21888 13088
rect 21824 13028 21828 13084
rect 21828 13028 21884 13084
rect 21884 13028 21888 13084
rect 21824 13024 21888 13028
rect 21904 13084 21968 13088
rect 21904 13028 21908 13084
rect 21908 13028 21964 13084
rect 21964 13028 21968 13084
rect 21904 13024 21968 13028
rect 21984 13084 22048 13088
rect 21984 13028 21988 13084
rect 21988 13028 22044 13084
rect 22044 13028 22048 13084
rect 21984 13024 22048 13028
rect 5580 12548 5644 12612
rect 3551 12540 3615 12544
rect 3551 12484 3555 12540
rect 3555 12484 3611 12540
rect 3611 12484 3615 12540
rect 3551 12480 3615 12484
rect 3631 12540 3695 12544
rect 3631 12484 3635 12540
rect 3635 12484 3691 12540
rect 3691 12484 3695 12540
rect 3631 12480 3695 12484
rect 3711 12540 3775 12544
rect 3711 12484 3715 12540
rect 3715 12484 3771 12540
rect 3771 12484 3775 12540
rect 3711 12480 3775 12484
rect 3791 12540 3855 12544
rect 3791 12484 3795 12540
rect 3795 12484 3851 12540
rect 3851 12484 3855 12540
rect 3791 12480 3855 12484
rect 8749 12540 8813 12544
rect 8749 12484 8753 12540
rect 8753 12484 8809 12540
rect 8809 12484 8813 12540
rect 8749 12480 8813 12484
rect 8829 12540 8893 12544
rect 8829 12484 8833 12540
rect 8833 12484 8889 12540
rect 8889 12484 8893 12540
rect 8829 12480 8893 12484
rect 8909 12540 8973 12544
rect 8909 12484 8913 12540
rect 8913 12484 8969 12540
rect 8969 12484 8973 12540
rect 8909 12480 8973 12484
rect 8989 12540 9053 12544
rect 8989 12484 8993 12540
rect 8993 12484 9049 12540
rect 9049 12484 9053 12540
rect 8989 12480 9053 12484
rect 13947 12540 14011 12544
rect 13947 12484 13951 12540
rect 13951 12484 14007 12540
rect 14007 12484 14011 12540
rect 13947 12480 14011 12484
rect 14027 12540 14091 12544
rect 14027 12484 14031 12540
rect 14031 12484 14087 12540
rect 14087 12484 14091 12540
rect 14027 12480 14091 12484
rect 14107 12540 14171 12544
rect 14107 12484 14111 12540
rect 14111 12484 14167 12540
rect 14167 12484 14171 12540
rect 14107 12480 14171 12484
rect 14187 12540 14251 12544
rect 14187 12484 14191 12540
rect 14191 12484 14247 12540
rect 14247 12484 14251 12540
rect 14187 12480 14251 12484
rect 19145 12540 19209 12544
rect 19145 12484 19149 12540
rect 19149 12484 19205 12540
rect 19205 12484 19209 12540
rect 19145 12480 19209 12484
rect 19225 12540 19289 12544
rect 19225 12484 19229 12540
rect 19229 12484 19285 12540
rect 19285 12484 19289 12540
rect 19225 12480 19289 12484
rect 19305 12540 19369 12544
rect 19305 12484 19309 12540
rect 19309 12484 19365 12540
rect 19365 12484 19369 12540
rect 19305 12480 19369 12484
rect 19385 12540 19449 12544
rect 19385 12484 19389 12540
rect 19389 12484 19445 12540
rect 19445 12484 19449 12540
rect 19385 12480 19449 12484
rect 6150 11996 6214 12000
rect 6150 11940 6154 11996
rect 6154 11940 6210 11996
rect 6210 11940 6214 11996
rect 6150 11936 6214 11940
rect 6230 11996 6294 12000
rect 6230 11940 6234 11996
rect 6234 11940 6290 11996
rect 6290 11940 6294 11996
rect 6230 11936 6294 11940
rect 6310 11996 6374 12000
rect 6310 11940 6314 11996
rect 6314 11940 6370 11996
rect 6370 11940 6374 11996
rect 6310 11936 6374 11940
rect 6390 11996 6454 12000
rect 6390 11940 6394 11996
rect 6394 11940 6450 11996
rect 6450 11940 6454 11996
rect 6390 11936 6454 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 16546 11996 16610 12000
rect 16546 11940 16550 11996
rect 16550 11940 16606 11996
rect 16606 11940 16610 11996
rect 16546 11936 16610 11940
rect 16626 11996 16690 12000
rect 16626 11940 16630 11996
rect 16630 11940 16686 11996
rect 16686 11940 16690 11996
rect 16626 11936 16690 11940
rect 16706 11996 16770 12000
rect 16706 11940 16710 11996
rect 16710 11940 16766 11996
rect 16766 11940 16770 11996
rect 16706 11936 16770 11940
rect 16786 11996 16850 12000
rect 16786 11940 16790 11996
rect 16790 11940 16846 11996
rect 16846 11940 16850 11996
rect 16786 11936 16850 11940
rect 21744 11996 21808 12000
rect 21744 11940 21748 11996
rect 21748 11940 21804 11996
rect 21804 11940 21808 11996
rect 21744 11936 21808 11940
rect 21824 11996 21888 12000
rect 21824 11940 21828 11996
rect 21828 11940 21884 11996
rect 21884 11940 21888 11996
rect 21824 11936 21888 11940
rect 21904 11996 21968 12000
rect 21904 11940 21908 11996
rect 21908 11940 21964 11996
rect 21964 11940 21968 11996
rect 21904 11936 21968 11940
rect 21984 11996 22048 12000
rect 21984 11940 21988 11996
rect 21988 11940 22044 11996
rect 22044 11940 22048 11996
rect 21984 11936 22048 11940
rect 3551 11452 3615 11456
rect 3551 11396 3555 11452
rect 3555 11396 3611 11452
rect 3611 11396 3615 11452
rect 3551 11392 3615 11396
rect 3631 11452 3695 11456
rect 3631 11396 3635 11452
rect 3635 11396 3691 11452
rect 3691 11396 3695 11452
rect 3631 11392 3695 11396
rect 3711 11452 3775 11456
rect 3711 11396 3715 11452
rect 3715 11396 3771 11452
rect 3771 11396 3775 11452
rect 3711 11392 3775 11396
rect 3791 11452 3855 11456
rect 3791 11396 3795 11452
rect 3795 11396 3851 11452
rect 3851 11396 3855 11452
rect 3791 11392 3855 11396
rect 8749 11452 8813 11456
rect 8749 11396 8753 11452
rect 8753 11396 8809 11452
rect 8809 11396 8813 11452
rect 8749 11392 8813 11396
rect 8829 11452 8893 11456
rect 8829 11396 8833 11452
rect 8833 11396 8889 11452
rect 8889 11396 8893 11452
rect 8829 11392 8893 11396
rect 8909 11452 8973 11456
rect 8909 11396 8913 11452
rect 8913 11396 8969 11452
rect 8969 11396 8973 11452
rect 8909 11392 8973 11396
rect 8989 11452 9053 11456
rect 8989 11396 8993 11452
rect 8993 11396 9049 11452
rect 9049 11396 9053 11452
rect 8989 11392 9053 11396
rect 13947 11452 14011 11456
rect 13947 11396 13951 11452
rect 13951 11396 14007 11452
rect 14007 11396 14011 11452
rect 13947 11392 14011 11396
rect 14027 11452 14091 11456
rect 14027 11396 14031 11452
rect 14031 11396 14087 11452
rect 14087 11396 14091 11452
rect 14027 11392 14091 11396
rect 14107 11452 14171 11456
rect 14107 11396 14111 11452
rect 14111 11396 14167 11452
rect 14167 11396 14171 11452
rect 14107 11392 14171 11396
rect 14187 11452 14251 11456
rect 14187 11396 14191 11452
rect 14191 11396 14247 11452
rect 14247 11396 14251 11452
rect 14187 11392 14251 11396
rect 19145 11452 19209 11456
rect 19145 11396 19149 11452
rect 19149 11396 19205 11452
rect 19205 11396 19209 11452
rect 19145 11392 19209 11396
rect 19225 11452 19289 11456
rect 19225 11396 19229 11452
rect 19229 11396 19285 11452
rect 19285 11396 19289 11452
rect 19225 11392 19289 11396
rect 19305 11452 19369 11456
rect 19305 11396 19309 11452
rect 19309 11396 19365 11452
rect 19365 11396 19369 11452
rect 19305 11392 19369 11396
rect 19385 11452 19449 11456
rect 19385 11396 19389 11452
rect 19389 11396 19445 11452
rect 19445 11396 19449 11452
rect 19385 11392 19449 11396
rect 6150 10908 6214 10912
rect 6150 10852 6154 10908
rect 6154 10852 6210 10908
rect 6210 10852 6214 10908
rect 6150 10848 6214 10852
rect 6230 10908 6294 10912
rect 6230 10852 6234 10908
rect 6234 10852 6290 10908
rect 6290 10852 6294 10908
rect 6230 10848 6294 10852
rect 6310 10908 6374 10912
rect 6310 10852 6314 10908
rect 6314 10852 6370 10908
rect 6370 10852 6374 10908
rect 6310 10848 6374 10852
rect 6390 10908 6454 10912
rect 6390 10852 6394 10908
rect 6394 10852 6450 10908
rect 6450 10852 6454 10908
rect 6390 10848 6454 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 16546 10908 16610 10912
rect 16546 10852 16550 10908
rect 16550 10852 16606 10908
rect 16606 10852 16610 10908
rect 16546 10848 16610 10852
rect 16626 10908 16690 10912
rect 16626 10852 16630 10908
rect 16630 10852 16686 10908
rect 16686 10852 16690 10908
rect 16626 10848 16690 10852
rect 16706 10908 16770 10912
rect 16706 10852 16710 10908
rect 16710 10852 16766 10908
rect 16766 10852 16770 10908
rect 16706 10848 16770 10852
rect 16786 10908 16850 10912
rect 16786 10852 16790 10908
rect 16790 10852 16846 10908
rect 16846 10852 16850 10908
rect 16786 10848 16850 10852
rect 21744 10908 21808 10912
rect 21744 10852 21748 10908
rect 21748 10852 21804 10908
rect 21804 10852 21808 10908
rect 21744 10848 21808 10852
rect 21824 10908 21888 10912
rect 21824 10852 21828 10908
rect 21828 10852 21884 10908
rect 21884 10852 21888 10908
rect 21824 10848 21888 10852
rect 21904 10908 21968 10912
rect 21904 10852 21908 10908
rect 21908 10852 21964 10908
rect 21964 10852 21968 10908
rect 21904 10848 21968 10852
rect 21984 10908 22048 10912
rect 21984 10852 21988 10908
rect 21988 10852 22044 10908
rect 22044 10852 22048 10908
rect 21984 10848 22048 10852
rect 3551 10364 3615 10368
rect 3551 10308 3555 10364
rect 3555 10308 3611 10364
rect 3611 10308 3615 10364
rect 3551 10304 3615 10308
rect 3631 10364 3695 10368
rect 3631 10308 3635 10364
rect 3635 10308 3691 10364
rect 3691 10308 3695 10364
rect 3631 10304 3695 10308
rect 3711 10364 3775 10368
rect 3711 10308 3715 10364
rect 3715 10308 3771 10364
rect 3771 10308 3775 10364
rect 3711 10304 3775 10308
rect 3791 10364 3855 10368
rect 3791 10308 3795 10364
rect 3795 10308 3851 10364
rect 3851 10308 3855 10364
rect 3791 10304 3855 10308
rect 8749 10364 8813 10368
rect 8749 10308 8753 10364
rect 8753 10308 8809 10364
rect 8809 10308 8813 10364
rect 8749 10304 8813 10308
rect 8829 10364 8893 10368
rect 8829 10308 8833 10364
rect 8833 10308 8889 10364
rect 8889 10308 8893 10364
rect 8829 10304 8893 10308
rect 8909 10364 8973 10368
rect 8909 10308 8913 10364
rect 8913 10308 8969 10364
rect 8969 10308 8973 10364
rect 8909 10304 8973 10308
rect 8989 10364 9053 10368
rect 8989 10308 8993 10364
rect 8993 10308 9049 10364
rect 9049 10308 9053 10364
rect 8989 10304 9053 10308
rect 13947 10364 14011 10368
rect 13947 10308 13951 10364
rect 13951 10308 14007 10364
rect 14007 10308 14011 10364
rect 13947 10304 14011 10308
rect 14027 10364 14091 10368
rect 14027 10308 14031 10364
rect 14031 10308 14087 10364
rect 14087 10308 14091 10364
rect 14027 10304 14091 10308
rect 14107 10364 14171 10368
rect 14107 10308 14111 10364
rect 14111 10308 14167 10364
rect 14167 10308 14171 10364
rect 14107 10304 14171 10308
rect 14187 10364 14251 10368
rect 14187 10308 14191 10364
rect 14191 10308 14247 10364
rect 14247 10308 14251 10364
rect 14187 10304 14251 10308
rect 19145 10364 19209 10368
rect 19145 10308 19149 10364
rect 19149 10308 19205 10364
rect 19205 10308 19209 10364
rect 19145 10304 19209 10308
rect 19225 10364 19289 10368
rect 19225 10308 19229 10364
rect 19229 10308 19285 10364
rect 19285 10308 19289 10364
rect 19225 10304 19289 10308
rect 19305 10364 19369 10368
rect 19305 10308 19309 10364
rect 19309 10308 19365 10364
rect 19365 10308 19369 10364
rect 19305 10304 19369 10308
rect 19385 10364 19449 10368
rect 19385 10308 19389 10364
rect 19389 10308 19445 10364
rect 19445 10308 19449 10364
rect 19385 10304 19449 10308
rect 8156 10100 8220 10164
rect 6150 9820 6214 9824
rect 6150 9764 6154 9820
rect 6154 9764 6210 9820
rect 6210 9764 6214 9820
rect 6150 9760 6214 9764
rect 6230 9820 6294 9824
rect 6230 9764 6234 9820
rect 6234 9764 6290 9820
rect 6290 9764 6294 9820
rect 6230 9760 6294 9764
rect 6310 9820 6374 9824
rect 6310 9764 6314 9820
rect 6314 9764 6370 9820
rect 6370 9764 6374 9820
rect 6310 9760 6374 9764
rect 6390 9820 6454 9824
rect 6390 9764 6394 9820
rect 6394 9764 6450 9820
rect 6450 9764 6454 9820
rect 6390 9760 6454 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 16546 9820 16610 9824
rect 16546 9764 16550 9820
rect 16550 9764 16606 9820
rect 16606 9764 16610 9820
rect 16546 9760 16610 9764
rect 16626 9820 16690 9824
rect 16626 9764 16630 9820
rect 16630 9764 16686 9820
rect 16686 9764 16690 9820
rect 16626 9760 16690 9764
rect 16706 9820 16770 9824
rect 16706 9764 16710 9820
rect 16710 9764 16766 9820
rect 16766 9764 16770 9820
rect 16706 9760 16770 9764
rect 16786 9820 16850 9824
rect 16786 9764 16790 9820
rect 16790 9764 16846 9820
rect 16846 9764 16850 9820
rect 16786 9760 16850 9764
rect 21744 9820 21808 9824
rect 21744 9764 21748 9820
rect 21748 9764 21804 9820
rect 21804 9764 21808 9820
rect 21744 9760 21808 9764
rect 21824 9820 21888 9824
rect 21824 9764 21828 9820
rect 21828 9764 21884 9820
rect 21884 9764 21888 9820
rect 21824 9760 21888 9764
rect 21904 9820 21968 9824
rect 21904 9764 21908 9820
rect 21908 9764 21964 9820
rect 21964 9764 21968 9820
rect 21904 9760 21968 9764
rect 21984 9820 22048 9824
rect 21984 9764 21988 9820
rect 21988 9764 22044 9820
rect 22044 9764 22048 9820
rect 21984 9760 22048 9764
rect 3551 9276 3615 9280
rect 3551 9220 3555 9276
rect 3555 9220 3611 9276
rect 3611 9220 3615 9276
rect 3551 9216 3615 9220
rect 3631 9276 3695 9280
rect 3631 9220 3635 9276
rect 3635 9220 3691 9276
rect 3691 9220 3695 9276
rect 3631 9216 3695 9220
rect 3711 9276 3775 9280
rect 3711 9220 3715 9276
rect 3715 9220 3771 9276
rect 3771 9220 3775 9276
rect 3711 9216 3775 9220
rect 3791 9276 3855 9280
rect 3791 9220 3795 9276
rect 3795 9220 3851 9276
rect 3851 9220 3855 9276
rect 3791 9216 3855 9220
rect 8749 9276 8813 9280
rect 8749 9220 8753 9276
rect 8753 9220 8809 9276
rect 8809 9220 8813 9276
rect 8749 9216 8813 9220
rect 8829 9276 8893 9280
rect 8829 9220 8833 9276
rect 8833 9220 8889 9276
rect 8889 9220 8893 9276
rect 8829 9216 8893 9220
rect 8909 9276 8973 9280
rect 8909 9220 8913 9276
rect 8913 9220 8969 9276
rect 8969 9220 8973 9276
rect 8909 9216 8973 9220
rect 8989 9276 9053 9280
rect 8989 9220 8993 9276
rect 8993 9220 9049 9276
rect 9049 9220 9053 9276
rect 8989 9216 9053 9220
rect 13947 9276 14011 9280
rect 13947 9220 13951 9276
rect 13951 9220 14007 9276
rect 14007 9220 14011 9276
rect 13947 9216 14011 9220
rect 14027 9276 14091 9280
rect 14027 9220 14031 9276
rect 14031 9220 14087 9276
rect 14087 9220 14091 9276
rect 14027 9216 14091 9220
rect 14107 9276 14171 9280
rect 14107 9220 14111 9276
rect 14111 9220 14167 9276
rect 14167 9220 14171 9276
rect 14107 9216 14171 9220
rect 14187 9276 14251 9280
rect 14187 9220 14191 9276
rect 14191 9220 14247 9276
rect 14247 9220 14251 9276
rect 14187 9216 14251 9220
rect 19145 9276 19209 9280
rect 19145 9220 19149 9276
rect 19149 9220 19205 9276
rect 19205 9220 19209 9276
rect 19145 9216 19209 9220
rect 19225 9276 19289 9280
rect 19225 9220 19229 9276
rect 19229 9220 19285 9276
rect 19285 9220 19289 9276
rect 19225 9216 19289 9220
rect 19305 9276 19369 9280
rect 19305 9220 19309 9276
rect 19309 9220 19365 9276
rect 19365 9220 19369 9276
rect 19305 9216 19369 9220
rect 19385 9276 19449 9280
rect 19385 9220 19389 9276
rect 19389 9220 19445 9276
rect 19445 9220 19449 9276
rect 19385 9216 19449 9220
rect 6150 8732 6214 8736
rect 6150 8676 6154 8732
rect 6154 8676 6210 8732
rect 6210 8676 6214 8732
rect 6150 8672 6214 8676
rect 6230 8732 6294 8736
rect 6230 8676 6234 8732
rect 6234 8676 6290 8732
rect 6290 8676 6294 8732
rect 6230 8672 6294 8676
rect 6310 8732 6374 8736
rect 6310 8676 6314 8732
rect 6314 8676 6370 8732
rect 6370 8676 6374 8732
rect 6310 8672 6374 8676
rect 6390 8732 6454 8736
rect 6390 8676 6394 8732
rect 6394 8676 6450 8732
rect 6450 8676 6454 8732
rect 6390 8672 6454 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 16546 8732 16610 8736
rect 16546 8676 16550 8732
rect 16550 8676 16606 8732
rect 16606 8676 16610 8732
rect 16546 8672 16610 8676
rect 16626 8732 16690 8736
rect 16626 8676 16630 8732
rect 16630 8676 16686 8732
rect 16686 8676 16690 8732
rect 16626 8672 16690 8676
rect 16706 8732 16770 8736
rect 16706 8676 16710 8732
rect 16710 8676 16766 8732
rect 16766 8676 16770 8732
rect 16706 8672 16770 8676
rect 16786 8732 16850 8736
rect 16786 8676 16790 8732
rect 16790 8676 16846 8732
rect 16846 8676 16850 8732
rect 16786 8672 16850 8676
rect 21744 8732 21808 8736
rect 21744 8676 21748 8732
rect 21748 8676 21804 8732
rect 21804 8676 21808 8732
rect 21744 8672 21808 8676
rect 21824 8732 21888 8736
rect 21824 8676 21828 8732
rect 21828 8676 21884 8732
rect 21884 8676 21888 8732
rect 21824 8672 21888 8676
rect 21904 8732 21968 8736
rect 21904 8676 21908 8732
rect 21908 8676 21964 8732
rect 21964 8676 21968 8732
rect 21904 8672 21968 8676
rect 21984 8732 22048 8736
rect 21984 8676 21988 8732
rect 21988 8676 22044 8732
rect 22044 8676 22048 8732
rect 21984 8672 22048 8676
rect 9444 8664 9508 8668
rect 9444 8608 9458 8664
rect 9458 8608 9508 8664
rect 9444 8604 9508 8608
rect 3551 8188 3615 8192
rect 3551 8132 3555 8188
rect 3555 8132 3611 8188
rect 3611 8132 3615 8188
rect 3551 8128 3615 8132
rect 3631 8188 3695 8192
rect 3631 8132 3635 8188
rect 3635 8132 3691 8188
rect 3691 8132 3695 8188
rect 3631 8128 3695 8132
rect 3711 8188 3775 8192
rect 3711 8132 3715 8188
rect 3715 8132 3771 8188
rect 3771 8132 3775 8188
rect 3711 8128 3775 8132
rect 3791 8188 3855 8192
rect 3791 8132 3795 8188
rect 3795 8132 3851 8188
rect 3851 8132 3855 8188
rect 3791 8128 3855 8132
rect 8749 8188 8813 8192
rect 8749 8132 8753 8188
rect 8753 8132 8809 8188
rect 8809 8132 8813 8188
rect 8749 8128 8813 8132
rect 8829 8188 8893 8192
rect 8829 8132 8833 8188
rect 8833 8132 8889 8188
rect 8889 8132 8893 8188
rect 8829 8128 8893 8132
rect 8909 8188 8973 8192
rect 8909 8132 8913 8188
rect 8913 8132 8969 8188
rect 8969 8132 8973 8188
rect 8909 8128 8973 8132
rect 8989 8188 9053 8192
rect 8989 8132 8993 8188
rect 8993 8132 9049 8188
rect 9049 8132 9053 8188
rect 8989 8128 9053 8132
rect 13947 8188 14011 8192
rect 13947 8132 13951 8188
rect 13951 8132 14007 8188
rect 14007 8132 14011 8188
rect 13947 8128 14011 8132
rect 14027 8188 14091 8192
rect 14027 8132 14031 8188
rect 14031 8132 14087 8188
rect 14087 8132 14091 8188
rect 14027 8128 14091 8132
rect 14107 8188 14171 8192
rect 14107 8132 14111 8188
rect 14111 8132 14167 8188
rect 14167 8132 14171 8188
rect 14107 8128 14171 8132
rect 14187 8188 14251 8192
rect 14187 8132 14191 8188
rect 14191 8132 14247 8188
rect 14247 8132 14251 8188
rect 14187 8128 14251 8132
rect 19145 8188 19209 8192
rect 19145 8132 19149 8188
rect 19149 8132 19205 8188
rect 19205 8132 19209 8188
rect 19145 8128 19209 8132
rect 19225 8188 19289 8192
rect 19225 8132 19229 8188
rect 19229 8132 19285 8188
rect 19285 8132 19289 8188
rect 19225 8128 19289 8132
rect 19305 8188 19369 8192
rect 19305 8132 19309 8188
rect 19309 8132 19365 8188
rect 19365 8132 19369 8188
rect 19305 8128 19369 8132
rect 19385 8188 19449 8192
rect 19385 8132 19389 8188
rect 19389 8132 19445 8188
rect 19445 8132 19449 8188
rect 19385 8128 19449 8132
rect 6150 7644 6214 7648
rect 6150 7588 6154 7644
rect 6154 7588 6210 7644
rect 6210 7588 6214 7644
rect 6150 7584 6214 7588
rect 6230 7644 6294 7648
rect 6230 7588 6234 7644
rect 6234 7588 6290 7644
rect 6290 7588 6294 7644
rect 6230 7584 6294 7588
rect 6310 7644 6374 7648
rect 6310 7588 6314 7644
rect 6314 7588 6370 7644
rect 6370 7588 6374 7644
rect 6310 7584 6374 7588
rect 6390 7644 6454 7648
rect 6390 7588 6394 7644
rect 6394 7588 6450 7644
rect 6450 7588 6454 7644
rect 6390 7584 6454 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 16546 7644 16610 7648
rect 16546 7588 16550 7644
rect 16550 7588 16606 7644
rect 16606 7588 16610 7644
rect 16546 7584 16610 7588
rect 16626 7644 16690 7648
rect 16626 7588 16630 7644
rect 16630 7588 16686 7644
rect 16686 7588 16690 7644
rect 16626 7584 16690 7588
rect 16706 7644 16770 7648
rect 16706 7588 16710 7644
rect 16710 7588 16766 7644
rect 16766 7588 16770 7644
rect 16706 7584 16770 7588
rect 16786 7644 16850 7648
rect 16786 7588 16790 7644
rect 16790 7588 16846 7644
rect 16846 7588 16850 7644
rect 16786 7584 16850 7588
rect 21744 7644 21808 7648
rect 21744 7588 21748 7644
rect 21748 7588 21804 7644
rect 21804 7588 21808 7644
rect 21744 7584 21808 7588
rect 21824 7644 21888 7648
rect 21824 7588 21828 7644
rect 21828 7588 21884 7644
rect 21884 7588 21888 7644
rect 21824 7584 21888 7588
rect 21904 7644 21968 7648
rect 21904 7588 21908 7644
rect 21908 7588 21964 7644
rect 21964 7588 21968 7644
rect 21904 7584 21968 7588
rect 21984 7644 22048 7648
rect 21984 7588 21988 7644
rect 21988 7588 22044 7644
rect 22044 7588 22048 7644
rect 21984 7584 22048 7588
rect 3551 7100 3615 7104
rect 3551 7044 3555 7100
rect 3555 7044 3611 7100
rect 3611 7044 3615 7100
rect 3551 7040 3615 7044
rect 3631 7100 3695 7104
rect 3631 7044 3635 7100
rect 3635 7044 3691 7100
rect 3691 7044 3695 7100
rect 3631 7040 3695 7044
rect 3711 7100 3775 7104
rect 3711 7044 3715 7100
rect 3715 7044 3771 7100
rect 3771 7044 3775 7100
rect 3711 7040 3775 7044
rect 3791 7100 3855 7104
rect 3791 7044 3795 7100
rect 3795 7044 3851 7100
rect 3851 7044 3855 7100
rect 3791 7040 3855 7044
rect 8749 7100 8813 7104
rect 8749 7044 8753 7100
rect 8753 7044 8809 7100
rect 8809 7044 8813 7100
rect 8749 7040 8813 7044
rect 8829 7100 8893 7104
rect 8829 7044 8833 7100
rect 8833 7044 8889 7100
rect 8889 7044 8893 7100
rect 8829 7040 8893 7044
rect 8909 7100 8973 7104
rect 8909 7044 8913 7100
rect 8913 7044 8969 7100
rect 8969 7044 8973 7100
rect 8909 7040 8973 7044
rect 8989 7100 9053 7104
rect 8989 7044 8993 7100
rect 8993 7044 9049 7100
rect 9049 7044 9053 7100
rect 8989 7040 9053 7044
rect 13947 7100 14011 7104
rect 13947 7044 13951 7100
rect 13951 7044 14007 7100
rect 14007 7044 14011 7100
rect 13947 7040 14011 7044
rect 14027 7100 14091 7104
rect 14027 7044 14031 7100
rect 14031 7044 14087 7100
rect 14087 7044 14091 7100
rect 14027 7040 14091 7044
rect 14107 7100 14171 7104
rect 14107 7044 14111 7100
rect 14111 7044 14167 7100
rect 14167 7044 14171 7100
rect 14107 7040 14171 7044
rect 14187 7100 14251 7104
rect 14187 7044 14191 7100
rect 14191 7044 14247 7100
rect 14247 7044 14251 7100
rect 14187 7040 14251 7044
rect 19145 7100 19209 7104
rect 19145 7044 19149 7100
rect 19149 7044 19205 7100
rect 19205 7044 19209 7100
rect 19145 7040 19209 7044
rect 19225 7100 19289 7104
rect 19225 7044 19229 7100
rect 19229 7044 19285 7100
rect 19285 7044 19289 7100
rect 19225 7040 19289 7044
rect 19305 7100 19369 7104
rect 19305 7044 19309 7100
rect 19309 7044 19365 7100
rect 19365 7044 19369 7100
rect 19305 7040 19369 7044
rect 19385 7100 19449 7104
rect 19385 7044 19389 7100
rect 19389 7044 19445 7100
rect 19445 7044 19449 7100
rect 19385 7040 19449 7044
rect 6150 6556 6214 6560
rect 6150 6500 6154 6556
rect 6154 6500 6210 6556
rect 6210 6500 6214 6556
rect 6150 6496 6214 6500
rect 6230 6556 6294 6560
rect 6230 6500 6234 6556
rect 6234 6500 6290 6556
rect 6290 6500 6294 6556
rect 6230 6496 6294 6500
rect 6310 6556 6374 6560
rect 6310 6500 6314 6556
rect 6314 6500 6370 6556
rect 6370 6500 6374 6556
rect 6310 6496 6374 6500
rect 6390 6556 6454 6560
rect 6390 6500 6394 6556
rect 6394 6500 6450 6556
rect 6450 6500 6454 6556
rect 6390 6496 6454 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 16546 6556 16610 6560
rect 16546 6500 16550 6556
rect 16550 6500 16606 6556
rect 16606 6500 16610 6556
rect 16546 6496 16610 6500
rect 16626 6556 16690 6560
rect 16626 6500 16630 6556
rect 16630 6500 16686 6556
rect 16686 6500 16690 6556
rect 16626 6496 16690 6500
rect 16706 6556 16770 6560
rect 16706 6500 16710 6556
rect 16710 6500 16766 6556
rect 16766 6500 16770 6556
rect 16706 6496 16770 6500
rect 16786 6556 16850 6560
rect 16786 6500 16790 6556
rect 16790 6500 16846 6556
rect 16846 6500 16850 6556
rect 16786 6496 16850 6500
rect 21744 6556 21808 6560
rect 21744 6500 21748 6556
rect 21748 6500 21804 6556
rect 21804 6500 21808 6556
rect 21744 6496 21808 6500
rect 21824 6556 21888 6560
rect 21824 6500 21828 6556
rect 21828 6500 21884 6556
rect 21884 6500 21888 6556
rect 21824 6496 21888 6500
rect 21904 6556 21968 6560
rect 21904 6500 21908 6556
rect 21908 6500 21964 6556
rect 21964 6500 21968 6556
rect 21904 6496 21968 6500
rect 21984 6556 22048 6560
rect 21984 6500 21988 6556
rect 21988 6500 22044 6556
rect 22044 6500 22048 6556
rect 21984 6496 22048 6500
rect 3551 6012 3615 6016
rect 3551 5956 3555 6012
rect 3555 5956 3611 6012
rect 3611 5956 3615 6012
rect 3551 5952 3615 5956
rect 3631 6012 3695 6016
rect 3631 5956 3635 6012
rect 3635 5956 3691 6012
rect 3691 5956 3695 6012
rect 3631 5952 3695 5956
rect 3711 6012 3775 6016
rect 3711 5956 3715 6012
rect 3715 5956 3771 6012
rect 3771 5956 3775 6012
rect 3711 5952 3775 5956
rect 3791 6012 3855 6016
rect 3791 5956 3795 6012
rect 3795 5956 3851 6012
rect 3851 5956 3855 6012
rect 3791 5952 3855 5956
rect 8749 6012 8813 6016
rect 8749 5956 8753 6012
rect 8753 5956 8809 6012
rect 8809 5956 8813 6012
rect 8749 5952 8813 5956
rect 8829 6012 8893 6016
rect 8829 5956 8833 6012
rect 8833 5956 8889 6012
rect 8889 5956 8893 6012
rect 8829 5952 8893 5956
rect 8909 6012 8973 6016
rect 8909 5956 8913 6012
rect 8913 5956 8969 6012
rect 8969 5956 8973 6012
rect 8909 5952 8973 5956
rect 8989 6012 9053 6016
rect 8989 5956 8993 6012
rect 8993 5956 9049 6012
rect 9049 5956 9053 6012
rect 8989 5952 9053 5956
rect 13947 6012 14011 6016
rect 13947 5956 13951 6012
rect 13951 5956 14007 6012
rect 14007 5956 14011 6012
rect 13947 5952 14011 5956
rect 14027 6012 14091 6016
rect 14027 5956 14031 6012
rect 14031 5956 14087 6012
rect 14087 5956 14091 6012
rect 14027 5952 14091 5956
rect 14107 6012 14171 6016
rect 14107 5956 14111 6012
rect 14111 5956 14167 6012
rect 14167 5956 14171 6012
rect 14107 5952 14171 5956
rect 14187 6012 14251 6016
rect 14187 5956 14191 6012
rect 14191 5956 14247 6012
rect 14247 5956 14251 6012
rect 14187 5952 14251 5956
rect 19145 6012 19209 6016
rect 19145 5956 19149 6012
rect 19149 5956 19205 6012
rect 19205 5956 19209 6012
rect 19145 5952 19209 5956
rect 19225 6012 19289 6016
rect 19225 5956 19229 6012
rect 19229 5956 19285 6012
rect 19285 5956 19289 6012
rect 19225 5952 19289 5956
rect 19305 6012 19369 6016
rect 19305 5956 19309 6012
rect 19309 5956 19365 6012
rect 19365 5956 19369 6012
rect 19305 5952 19369 5956
rect 19385 6012 19449 6016
rect 19385 5956 19389 6012
rect 19389 5956 19445 6012
rect 19445 5956 19449 6012
rect 19385 5952 19449 5956
rect 6150 5468 6214 5472
rect 6150 5412 6154 5468
rect 6154 5412 6210 5468
rect 6210 5412 6214 5468
rect 6150 5408 6214 5412
rect 6230 5468 6294 5472
rect 6230 5412 6234 5468
rect 6234 5412 6290 5468
rect 6290 5412 6294 5468
rect 6230 5408 6294 5412
rect 6310 5468 6374 5472
rect 6310 5412 6314 5468
rect 6314 5412 6370 5468
rect 6370 5412 6374 5468
rect 6310 5408 6374 5412
rect 6390 5468 6454 5472
rect 6390 5412 6394 5468
rect 6394 5412 6450 5468
rect 6450 5412 6454 5468
rect 6390 5408 6454 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 16546 5468 16610 5472
rect 16546 5412 16550 5468
rect 16550 5412 16606 5468
rect 16606 5412 16610 5468
rect 16546 5408 16610 5412
rect 16626 5468 16690 5472
rect 16626 5412 16630 5468
rect 16630 5412 16686 5468
rect 16686 5412 16690 5468
rect 16626 5408 16690 5412
rect 16706 5468 16770 5472
rect 16706 5412 16710 5468
rect 16710 5412 16766 5468
rect 16766 5412 16770 5468
rect 16706 5408 16770 5412
rect 16786 5468 16850 5472
rect 16786 5412 16790 5468
rect 16790 5412 16846 5468
rect 16846 5412 16850 5468
rect 16786 5408 16850 5412
rect 21744 5468 21808 5472
rect 21744 5412 21748 5468
rect 21748 5412 21804 5468
rect 21804 5412 21808 5468
rect 21744 5408 21808 5412
rect 21824 5468 21888 5472
rect 21824 5412 21828 5468
rect 21828 5412 21884 5468
rect 21884 5412 21888 5468
rect 21824 5408 21888 5412
rect 21904 5468 21968 5472
rect 21904 5412 21908 5468
rect 21908 5412 21964 5468
rect 21964 5412 21968 5468
rect 21904 5408 21968 5412
rect 21984 5468 22048 5472
rect 21984 5412 21988 5468
rect 21988 5412 22044 5468
rect 22044 5412 22048 5468
rect 21984 5408 22048 5412
rect 7052 4992 7116 4996
rect 7052 4936 7066 4992
rect 7066 4936 7116 4992
rect 7052 4932 7116 4936
rect 3551 4924 3615 4928
rect 3551 4868 3555 4924
rect 3555 4868 3611 4924
rect 3611 4868 3615 4924
rect 3551 4864 3615 4868
rect 3631 4924 3695 4928
rect 3631 4868 3635 4924
rect 3635 4868 3691 4924
rect 3691 4868 3695 4924
rect 3631 4864 3695 4868
rect 3711 4924 3775 4928
rect 3711 4868 3715 4924
rect 3715 4868 3771 4924
rect 3771 4868 3775 4924
rect 3711 4864 3775 4868
rect 3791 4924 3855 4928
rect 3791 4868 3795 4924
rect 3795 4868 3851 4924
rect 3851 4868 3855 4924
rect 3791 4864 3855 4868
rect 8749 4924 8813 4928
rect 8749 4868 8753 4924
rect 8753 4868 8809 4924
rect 8809 4868 8813 4924
rect 8749 4864 8813 4868
rect 8829 4924 8893 4928
rect 8829 4868 8833 4924
rect 8833 4868 8889 4924
rect 8889 4868 8893 4924
rect 8829 4864 8893 4868
rect 8909 4924 8973 4928
rect 8909 4868 8913 4924
rect 8913 4868 8969 4924
rect 8969 4868 8973 4924
rect 8909 4864 8973 4868
rect 8989 4924 9053 4928
rect 8989 4868 8993 4924
rect 8993 4868 9049 4924
rect 9049 4868 9053 4924
rect 8989 4864 9053 4868
rect 13947 4924 14011 4928
rect 13947 4868 13951 4924
rect 13951 4868 14007 4924
rect 14007 4868 14011 4924
rect 13947 4864 14011 4868
rect 14027 4924 14091 4928
rect 14027 4868 14031 4924
rect 14031 4868 14087 4924
rect 14087 4868 14091 4924
rect 14027 4864 14091 4868
rect 14107 4924 14171 4928
rect 14107 4868 14111 4924
rect 14111 4868 14167 4924
rect 14167 4868 14171 4924
rect 14107 4864 14171 4868
rect 14187 4924 14251 4928
rect 14187 4868 14191 4924
rect 14191 4868 14247 4924
rect 14247 4868 14251 4924
rect 14187 4864 14251 4868
rect 19145 4924 19209 4928
rect 19145 4868 19149 4924
rect 19149 4868 19205 4924
rect 19205 4868 19209 4924
rect 19145 4864 19209 4868
rect 19225 4924 19289 4928
rect 19225 4868 19229 4924
rect 19229 4868 19285 4924
rect 19285 4868 19289 4924
rect 19225 4864 19289 4868
rect 19305 4924 19369 4928
rect 19305 4868 19309 4924
rect 19309 4868 19365 4924
rect 19365 4868 19369 4924
rect 19305 4864 19369 4868
rect 19385 4924 19449 4928
rect 19385 4868 19389 4924
rect 19389 4868 19445 4924
rect 19445 4868 19449 4924
rect 19385 4864 19449 4868
rect 6150 4380 6214 4384
rect 6150 4324 6154 4380
rect 6154 4324 6210 4380
rect 6210 4324 6214 4380
rect 6150 4320 6214 4324
rect 6230 4380 6294 4384
rect 6230 4324 6234 4380
rect 6234 4324 6290 4380
rect 6290 4324 6294 4380
rect 6230 4320 6294 4324
rect 6310 4380 6374 4384
rect 6310 4324 6314 4380
rect 6314 4324 6370 4380
rect 6370 4324 6374 4380
rect 6310 4320 6374 4324
rect 6390 4380 6454 4384
rect 6390 4324 6394 4380
rect 6394 4324 6450 4380
rect 6450 4324 6454 4380
rect 6390 4320 6454 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 16546 4380 16610 4384
rect 16546 4324 16550 4380
rect 16550 4324 16606 4380
rect 16606 4324 16610 4380
rect 16546 4320 16610 4324
rect 16626 4380 16690 4384
rect 16626 4324 16630 4380
rect 16630 4324 16686 4380
rect 16686 4324 16690 4380
rect 16626 4320 16690 4324
rect 16706 4380 16770 4384
rect 16706 4324 16710 4380
rect 16710 4324 16766 4380
rect 16766 4324 16770 4380
rect 16706 4320 16770 4324
rect 16786 4380 16850 4384
rect 16786 4324 16790 4380
rect 16790 4324 16846 4380
rect 16846 4324 16850 4380
rect 16786 4320 16850 4324
rect 21744 4380 21808 4384
rect 21744 4324 21748 4380
rect 21748 4324 21804 4380
rect 21804 4324 21808 4380
rect 21744 4320 21808 4324
rect 21824 4380 21888 4384
rect 21824 4324 21828 4380
rect 21828 4324 21884 4380
rect 21884 4324 21888 4380
rect 21824 4320 21888 4324
rect 21904 4380 21968 4384
rect 21904 4324 21908 4380
rect 21908 4324 21964 4380
rect 21964 4324 21968 4380
rect 21904 4320 21968 4324
rect 21984 4380 22048 4384
rect 21984 4324 21988 4380
rect 21988 4324 22044 4380
rect 22044 4324 22048 4380
rect 21984 4320 22048 4324
rect 5580 3844 5644 3908
rect 3551 3836 3615 3840
rect 3551 3780 3555 3836
rect 3555 3780 3611 3836
rect 3611 3780 3615 3836
rect 3551 3776 3615 3780
rect 3631 3836 3695 3840
rect 3631 3780 3635 3836
rect 3635 3780 3691 3836
rect 3691 3780 3695 3836
rect 3631 3776 3695 3780
rect 3711 3836 3775 3840
rect 3711 3780 3715 3836
rect 3715 3780 3771 3836
rect 3771 3780 3775 3836
rect 3711 3776 3775 3780
rect 3791 3836 3855 3840
rect 3791 3780 3795 3836
rect 3795 3780 3851 3836
rect 3851 3780 3855 3836
rect 3791 3776 3855 3780
rect 8749 3836 8813 3840
rect 8749 3780 8753 3836
rect 8753 3780 8809 3836
rect 8809 3780 8813 3836
rect 8749 3776 8813 3780
rect 8829 3836 8893 3840
rect 8829 3780 8833 3836
rect 8833 3780 8889 3836
rect 8889 3780 8893 3836
rect 8829 3776 8893 3780
rect 8909 3836 8973 3840
rect 8909 3780 8913 3836
rect 8913 3780 8969 3836
rect 8969 3780 8973 3836
rect 8909 3776 8973 3780
rect 8989 3836 9053 3840
rect 8989 3780 8993 3836
rect 8993 3780 9049 3836
rect 9049 3780 9053 3836
rect 8989 3776 9053 3780
rect 13947 3836 14011 3840
rect 13947 3780 13951 3836
rect 13951 3780 14007 3836
rect 14007 3780 14011 3836
rect 13947 3776 14011 3780
rect 14027 3836 14091 3840
rect 14027 3780 14031 3836
rect 14031 3780 14087 3836
rect 14087 3780 14091 3836
rect 14027 3776 14091 3780
rect 14107 3836 14171 3840
rect 14107 3780 14111 3836
rect 14111 3780 14167 3836
rect 14167 3780 14171 3836
rect 14107 3776 14171 3780
rect 14187 3836 14251 3840
rect 14187 3780 14191 3836
rect 14191 3780 14247 3836
rect 14247 3780 14251 3836
rect 14187 3776 14251 3780
rect 19145 3836 19209 3840
rect 19145 3780 19149 3836
rect 19149 3780 19205 3836
rect 19205 3780 19209 3836
rect 19145 3776 19209 3780
rect 19225 3836 19289 3840
rect 19225 3780 19229 3836
rect 19229 3780 19285 3836
rect 19285 3780 19289 3836
rect 19225 3776 19289 3780
rect 19305 3836 19369 3840
rect 19305 3780 19309 3836
rect 19309 3780 19365 3836
rect 19365 3780 19369 3836
rect 19305 3776 19369 3780
rect 19385 3836 19449 3840
rect 19385 3780 19389 3836
rect 19389 3780 19445 3836
rect 19445 3780 19449 3836
rect 19385 3776 19449 3780
rect 8340 3572 8404 3636
rect 9260 3436 9324 3500
rect 6150 3292 6214 3296
rect 6150 3236 6154 3292
rect 6154 3236 6210 3292
rect 6210 3236 6214 3292
rect 6150 3232 6214 3236
rect 6230 3292 6294 3296
rect 6230 3236 6234 3292
rect 6234 3236 6290 3292
rect 6290 3236 6294 3292
rect 6230 3232 6294 3236
rect 6310 3292 6374 3296
rect 6310 3236 6314 3292
rect 6314 3236 6370 3292
rect 6370 3236 6374 3292
rect 6310 3232 6374 3236
rect 6390 3292 6454 3296
rect 6390 3236 6394 3292
rect 6394 3236 6450 3292
rect 6450 3236 6454 3292
rect 6390 3232 6454 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 16546 3292 16610 3296
rect 16546 3236 16550 3292
rect 16550 3236 16606 3292
rect 16606 3236 16610 3292
rect 16546 3232 16610 3236
rect 16626 3292 16690 3296
rect 16626 3236 16630 3292
rect 16630 3236 16686 3292
rect 16686 3236 16690 3292
rect 16626 3232 16690 3236
rect 16706 3292 16770 3296
rect 16706 3236 16710 3292
rect 16710 3236 16766 3292
rect 16766 3236 16770 3292
rect 16706 3232 16770 3236
rect 16786 3292 16850 3296
rect 16786 3236 16790 3292
rect 16790 3236 16846 3292
rect 16846 3236 16850 3292
rect 16786 3232 16850 3236
rect 21744 3292 21808 3296
rect 21744 3236 21748 3292
rect 21748 3236 21804 3292
rect 21804 3236 21808 3292
rect 21744 3232 21808 3236
rect 21824 3292 21888 3296
rect 21824 3236 21828 3292
rect 21828 3236 21884 3292
rect 21884 3236 21888 3292
rect 21824 3232 21888 3236
rect 21904 3292 21968 3296
rect 21904 3236 21908 3292
rect 21908 3236 21964 3292
rect 21964 3236 21968 3292
rect 21904 3232 21968 3236
rect 21984 3292 22048 3296
rect 21984 3236 21988 3292
rect 21988 3236 22044 3292
rect 22044 3236 22048 3292
rect 21984 3232 22048 3236
rect 8156 3028 8220 3092
rect 3551 2748 3615 2752
rect 3551 2692 3555 2748
rect 3555 2692 3611 2748
rect 3611 2692 3615 2748
rect 3551 2688 3615 2692
rect 3631 2748 3695 2752
rect 3631 2692 3635 2748
rect 3635 2692 3691 2748
rect 3691 2692 3695 2748
rect 3631 2688 3695 2692
rect 3711 2748 3775 2752
rect 3711 2692 3715 2748
rect 3715 2692 3771 2748
rect 3771 2692 3775 2748
rect 3711 2688 3775 2692
rect 3791 2748 3855 2752
rect 3791 2692 3795 2748
rect 3795 2692 3851 2748
rect 3851 2692 3855 2748
rect 3791 2688 3855 2692
rect 8749 2748 8813 2752
rect 8749 2692 8753 2748
rect 8753 2692 8809 2748
rect 8809 2692 8813 2748
rect 8749 2688 8813 2692
rect 8829 2748 8893 2752
rect 8829 2692 8833 2748
rect 8833 2692 8889 2748
rect 8889 2692 8893 2748
rect 8829 2688 8893 2692
rect 8909 2748 8973 2752
rect 8909 2692 8913 2748
rect 8913 2692 8969 2748
rect 8969 2692 8973 2748
rect 8909 2688 8973 2692
rect 8989 2748 9053 2752
rect 8989 2692 8993 2748
rect 8993 2692 9049 2748
rect 9049 2692 9053 2748
rect 8989 2688 9053 2692
rect 13947 2748 14011 2752
rect 13947 2692 13951 2748
rect 13951 2692 14007 2748
rect 14007 2692 14011 2748
rect 13947 2688 14011 2692
rect 14027 2748 14091 2752
rect 14027 2692 14031 2748
rect 14031 2692 14087 2748
rect 14087 2692 14091 2748
rect 14027 2688 14091 2692
rect 14107 2748 14171 2752
rect 14107 2692 14111 2748
rect 14111 2692 14167 2748
rect 14167 2692 14171 2748
rect 14107 2688 14171 2692
rect 14187 2748 14251 2752
rect 14187 2692 14191 2748
rect 14191 2692 14247 2748
rect 14247 2692 14251 2748
rect 14187 2688 14251 2692
rect 19145 2748 19209 2752
rect 19145 2692 19149 2748
rect 19149 2692 19205 2748
rect 19205 2692 19209 2748
rect 19145 2688 19209 2692
rect 19225 2748 19289 2752
rect 19225 2692 19229 2748
rect 19229 2692 19285 2748
rect 19285 2692 19289 2748
rect 19225 2688 19289 2692
rect 19305 2748 19369 2752
rect 19305 2692 19309 2748
rect 19309 2692 19365 2748
rect 19365 2692 19369 2748
rect 19305 2688 19369 2692
rect 19385 2748 19449 2752
rect 19385 2692 19389 2748
rect 19389 2692 19445 2748
rect 19445 2692 19449 2748
rect 19385 2688 19449 2692
rect 7052 2212 7116 2276
rect 6150 2204 6214 2208
rect 6150 2148 6154 2204
rect 6154 2148 6210 2204
rect 6210 2148 6214 2204
rect 6150 2144 6214 2148
rect 6230 2204 6294 2208
rect 6230 2148 6234 2204
rect 6234 2148 6290 2204
rect 6290 2148 6294 2204
rect 6230 2144 6294 2148
rect 6310 2204 6374 2208
rect 6310 2148 6314 2204
rect 6314 2148 6370 2204
rect 6370 2148 6374 2204
rect 6310 2144 6374 2148
rect 6390 2204 6454 2208
rect 6390 2148 6394 2204
rect 6394 2148 6450 2204
rect 6450 2148 6454 2204
rect 6390 2144 6454 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 16546 2204 16610 2208
rect 16546 2148 16550 2204
rect 16550 2148 16606 2204
rect 16606 2148 16610 2204
rect 16546 2144 16610 2148
rect 16626 2204 16690 2208
rect 16626 2148 16630 2204
rect 16630 2148 16686 2204
rect 16686 2148 16690 2204
rect 16626 2144 16690 2148
rect 16706 2204 16770 2208
rect 16706 2148 16710 2204
rect 16710 2148 16766 2204
rect 16766 2148 16770 2204
rect 16706 2144 16770 2148
rect 16786 2204 16850 2208
rect 16786 2148 16790 2204
rect 16790 2148 16846 2204
rect 16846 2148 16850 2204
rect 16786 2144 16850 2148
rect 21744 2204 21808 2208
rect 21744 2148 21748 2204
rect 21748 2148 21804 2204
rect 21804 2148 21808 2204
rect 21744 2144 21808 2148
rect 21824 2204 21888 2208
rect 21824 2148 21828 2204
rect 21828 2148 21884 2204
rect 21884 2148 21888 2204
rect 21824 2144 21888 2148
rect 21904 2204 21968 2208
rect 21904 2148 21908 2204
rect 21908 2148 21964 2204
rect 21964 2148 21968 2204
rect 21904 2144 21968 2148
rect 21984 2204 22048 2208
rect 21984 2148 21988 2204
rect 21988 2148 22044 2204
rect 22044 2148 22048 2204
rect 21984 2144 22048 2148
rect 9444 2136 9508 2140
rect 9444 2080 9458 2136
rect 9458 2080 9508 2136
rect 9444 2076 9508 2080
<< metal4 >>
rect 3543 20160 3863 20720
rect 3543 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3863 20160
rect 3543 19072 3863 20096
rect 3543 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3863 19072
rect 3543 17984 3863 19008
rect 3543 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3863 17984
rect 3543 16896 3863 17920
rect 3543 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3863 16896
rect 3543 15808 3863 16832
rect 3543 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3863 15808
rect 3543 14720 3863 15744
rect 3543 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3863 14720
rect 3543 13632 3863 14656
rect 3543 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3863 13632
rect 3543 12544 3863 13568
rect 6142 20704 6462 20720
rect 6142 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6462 20704
rect 6142 19616 6462 20640
rect 6142 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6462 19616
rect 6142 18528 6462 19552
rect 6142 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6462 18528
rect 6142 17440 6462 18464
rect 6142 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6462 17440
rect 6142 16352 6462 17376
rect 6142 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6462 16352
rect 6142 15264 6462 16288
rect 6142 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6462 15264
rect 6142 14176 6462 15200
rect 6142 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6462 14176
rect 6142 13088 6462 14112
rect 8741 20160 9061 20720
rect 8741 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9061 20160
rect 8741 19072 9061 20096
rect 8741 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9061 19072
rect 8741 17984 9061 19008
rect 8741 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9061 17984
rect 8741 16896 9061 17920
rect 8741 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9061 16896
rect 8741 15808 9061 16832
rect 8741 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9061 15808
rect 8741 14720 9061 15744
rect 8741 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9061 14720
rect 8339 13972 8405 13973
rect 8339 13908 8340 13972
rect 8404 13908 8405 13972
rect 8339 13907 8405 13908
rect 6142 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6462 13088
rect 5579 12612 5645 12613
rect 5579 12548 5580 12612
rect 5644 12548 5645 12612
rect 5579 12547 5645 12548
rect 3543 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3863 12544
rect 3543 11456 3863 12480
rect 3543 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3863 11456
rect 3543 10368 3863 11392
rect 3543 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3863 10368
rect 3543 9280 3863 10304
rect 3543 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3863 9280
rect 3543 8192 3863 9216
rect 3543 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3863 8192
rect 3543 7104 3863 8128
rect 3543 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3863 7104
rect 3543 6016 3863 7040
rect 3543 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3863 6016
rect 3543 4928 3863 5952
rect 3543 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3863 4928
rect 3543 3840 3863 4864
rect 5582 3909 5642 12547
rect 6142 12000 6462 13024
rect 6142 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6462 12000
rect 6142 10912 6462 11936
rect 6142 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6462 10912
rect 6142 9824 6462 10848
rect 8155 10164 8221 10165
rect 8155 10100 8156 10164
rect 8220 10100 8221 10164
rect 8155 10099 8221 10100
rect 6142 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6462 9824
rect 6142 8736 6462 9760
rect 6142 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6462 8736
rect 6142 7648 6462 8672
rect 6142 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6462 7648
rect 6142 6560 6462 7584
rect 6142 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6462 6560
rect 6142 5472 6462 6496
rect 6142 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6462 5472
rect 6142 4384 6462 5408
rect 7051 4996 7117 4997
rect 7051 4932 7052 4996
rect 7116 4932 7117 4996
rect 7051 4931 7117 4932
rect 6142 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6462 4384
rect 5579 3908 5645 3909
rect 5579 3844 5580 3908
rect 5644 3844 5645 3908
rect 5579 3843 5645 3844
rect 3543 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3863 3840
rect 3543 2752 3863 3776
rect 3543 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3863 2752
rect 3543 2128 3863 2688
rect 6142 3296 6462 4320
rect 6142 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6462 3296
rect 6142 2208 6462 3232
rect 7054 2277 7114 4931
rect 8158 3093 8218 10099
rect 8342 3637 8402 13907
rect 8741 13632 9061 14656
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 9259 13836 9325 13837
rect 9259 13772 9260 13836
rect 9324 13772 9325 13836
rect 9259 13771 9325 13772
rect 8741 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9061 13632
rect 8741 12544 9061 13568
rect 8741 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9061 12544
rect 8741 11456 9061 12480
rect 8741 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9061 11456
rect 8741 10368 9061 11392
rect 8741 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9061 10368
rect 8741 9280 9061 10304
rect 8741 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9061 9280
rect 8741 8192 9061 9216
rect 8741 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9061 8192
rect 8741 7104 9061 8128
rect 8741 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9061 7104
rect 8741 6016 9061 7040
rect 8741 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9061 6016
rect 8741 4928 9061 5952
rect 8741 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9061 4928
rect 8741 3840 9061 4864
rect 8741 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9061 3840
rect 8339 3636 8405 3637
rect 8339 3572 8340 3636
rect 8404 3572 8405 3636
rect 8339 3571 8405 3572
rect 8155 3092 8221 3093
rect 8155 3028 8156 3092
rect 8220 3028 8221 3092
rect 8155 3027 8221 3028
rect 8741 2752 9061 3776
rect 9262 3501 9322 13771
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 9443 8668 9509 8669
rect 9443 8604 9444 8668
rect 9508 8604 9509 8668
rect 9443 8603 9509 8604
rect 9259 3500 9325 3501
rect 9259 3436 9260 3500
rect 9324 3436 9325 3500
rect 9259 3435 9325 3436
rect 8741 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9061 2752
rect 7051 2276 7117 2277
rect 7051 2212 7052 2276
rect 7116 2212 7117 2276
rect 7051 2211 7117 2212
rect 6142 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6462 2208
rect 6142 2128 6462 2144
rect 8741 2128 9061 2688
rect 9446 2141 9506 8603
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 9443 2140 9509 2141
rect 9443 2076 9444 2140
rect 9508 2076 9509 2140
rect 11340 2128 11660 2144
rect 13939 20160 14259 20720
rect 13939 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14259 20160
rect 13939 19072 14259 20096
rect 13939 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14259 19072
rect 13939 17984 14259 19008
rect 13939 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14259 17984
rect 13939 16896 14259 17920
rect 13939 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14259 16896
rect 13939 15808 14259 16832
rect 13939 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14259 15808
rect 13939 14720 14259 15744
rect 13939 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14259 14720
rect 13939 13632 14259 14656
rect 13939 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14259 13632
rect 13939 12544 14259 13568
rect 13939 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14259 12544
rect 13939 11456 14259 12480
rect 13939 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14259 11456
rect 13939 10368 14259 11392
rect 13939 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14259 10368
rect 13939 9280 14259 10304
rect 13939 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14259 9280
rect 13939 8192 14259 9216
rect 13939 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14259 8192
rect 13939 7104 14259 8128
rect 13939 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14259 7104
rect 13939 6016 14259 7040
rect 13939 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14259 6016
rect 13939 4928 14259 5952
rect 13939 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14259 4928
rect 13939 3840 14259 4864
rect 13939 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14259 3840
rect 13939 2752 14259 3776
rect 13939 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14259 2752
rect 13939 2128 14259 2688
rect 16538 20704 16858 20720
rect 16538 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16858 20704
rect 16538 19616 16858 20640
rect 16538 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16858 19616
rect 16538 18528 16858 19552
rect 16538 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16858 18528
rect 16538 17440 16858 18464
rect 16538 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16858 17440
rect 16538 16352 16858 17376
rect 16538 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16858 16352
rect 16538 15264 16858 16288
rect 16538 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16858 15264
rect 16538 14176 16858 15200
rect 16538 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16858 14176
rect 16538 13088 16858 14112
rect 16538 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16858 13088
rect 16538 12000 16858 13024
rect 16538 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16858 12000
rect 16538 10912 16858 11936
rect 16538 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16858 10912
rect 16538 9824 16858 10848
rect 16538 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16858 9824
rect 16538 8736 16858 9760
rect 16538 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16858 8736
rect 16538 7648 16858 8672
rect 16538 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16858 7648
rect 16538 6560 16858 7584
rect 16538 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16858 6560
rect 16538 5472 16858 6496
rect 16538 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16858 5472
rect 16538 4384 16858 5408
rect 16538 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16858 4384
rect 16538 3296 16858 4320
rect 16538 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16858 3296
rect 16538 2208 16858 3232
rect 16538 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16858 2208
rect 16538 2128 16858 2144
rect 19137 20160 19457 20720
rect 19137 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19457 20160
rect 19137 19072 19457 20096
rect 19137 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19457 19072
rect 19137 17984 19457 19008
rect 19137 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19457 17984
rect 19137 16896 19457 17920
rect 19137 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19457 16896
rect 19137 15808 19457 16832
rect 19137 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19457 15808
rect 19137 14720 19457 15744
rect 19137 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19457 14720
rect 19137 13632 19457 14656
rect 19137 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19457 13632
rect 19137 12544 19457 13568
rect 19137 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19457 12544
rect 19137 11456 19457 12480
rect 19137 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19457 11456
rect 19137 10368 19457 11392
rect 19137 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19457 10368
rect 19137 9280 19457 10304
rect 19137 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19457 9280
rect 19137 8192 19457 9216
rect 19137 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19457 8192
rect 19137 7104 19457 8128
rect 19137 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19457 7104
rect 19137 6016 19457 7040
rect 19137 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19457 6016
rect 19137 4928 19457 5952
rect 19137 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19457 4928
rect 19137 3840 19457 4864
rect 19137 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19457 3840
rect 19137 2752 19457 3776
rect 19137 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19457 2752
rect 19137 2128 19457 2688
rect 21736 20704 22056 20720
rect 21736 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22056 20704
rect 21736 19616 22056 20640
rect 21736 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22056 19616
rect 21736 18528 22056 19552
rect 21736 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22056 18528
rect 21736 17440 22056 18464
rect 21736 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22056 17440
rect 21736 16352 22056 17376
rect 21736 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22056 16352
rect 21736 15264 22056 16288
rect 21736 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22056 15264
rect 21736 14176 22056 15200
rect 21736 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22056 14176
rect 21736 13088 22056 14112
rect 21736 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22056 13088
rect 21736 12000 22056 13024
rect 21736 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22056 12000
rect 21736 10912 22056 11936
rect 21736 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22056 10912
rect 21736 9824 22056 10848
rect 21736 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22056 9824
rect 21736 8736 22056 9760
rect 21736 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22056 8736
rect 21736 7648 22056 8672
rect 21736 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22056 7648
rect 21736 6560 22056 7584
rect 21736 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22056 6560
rect 21736 5472 22056 6496
rect 21736 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22056 5472
rect 21736 4384 22056 5408
rect 21736 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22056 4384
rect 21736 3296 22056 4320
rect 21736 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22056 3296
rect 21736 2208 22056 3232
rect 21736 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22056 2208
rect 21736 2128 22056 2144
rect 9443 2075 9509 2076
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 18400 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1649977179
transform -1 0 3128 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1649977179
transform -1 0 2668 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A
timestamp 1649977179
transform -1 0 2576 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1649977179
transform 1 0 2576 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1649977179
transform -1 0 1656 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11040 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform -1 0 11040 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18308 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 21068 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 17112 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform -1 0 17940 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16376 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 16744 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 12880 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18308 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 17480 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 21252 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18400 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15916 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 11040 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18584 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 21068 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 20884 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16284 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18676 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 19320 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15732 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16192 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15732 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21252 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18124 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18952 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 17572 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 19044 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 20884 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21068 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 21068 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 17572 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18492 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 17756 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18124 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18492 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13708 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 15640 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13156 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13616 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 16100 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 14996 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13156 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13524 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 12420 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13156 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13064 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11040 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11040 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13156 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13524 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 12880 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13524 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16192 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13156 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13432 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15824 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16192 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 12144 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15732 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 19320 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 18124 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform -1 0 20884 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 20884 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 19780 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 21252 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 20884 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 21252 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21252 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 20976 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21252 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18768 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 17296 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14536 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18124 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 21252 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 4508 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 5060 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 3864 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 4416 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 5520 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__S
timestamp 1649977179
transform -1 0 4324 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 2852 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 2024 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 3220 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 4048 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 4140 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1649977179
transform -1 0 1564 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 4324 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 5888 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 4784 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 3864 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 4784 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 4232 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 2944 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 3312 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 3956 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 3128 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_1__A1
timestamp 1649977179
transform -1 0 1840 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 7912 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 5888 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8464 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 7912 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 4140 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 10304 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 7544 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 6900 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8464 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 9108 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6440 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 6992 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 4968 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 3680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 3128 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 7636 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_29.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 9752 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 3956 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 6808 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 6532 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 7360 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 5612 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 6808 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 3864 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 3128 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 2944 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 2116 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 3404 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 3772 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 3128 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 5888 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 6532 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 9752 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 3312 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 4876 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 2944 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6072 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 8556 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6716 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 7268 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 10028 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 10488 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 7452 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 8556 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 7360 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 9568 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 7544 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 9108 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 9108 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 5888 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 6072 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 6532 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 4968 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 5888 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1649977179
transform -1 0 5244 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 10120 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9384 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 9568 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 9108 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 10120 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 11776 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11316 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9016 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 10764 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 12880 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 12512 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11684 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 11868 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 10396 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform -1 0 18032 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2300 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2668 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37
timestamp 1649977179
transform 1 0 4508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42
timestamp 1649977179
transform 1 0 4968 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48
timestamp 1649977179
transform 1 0 5520 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1649977179
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64
timestamp 1649977179
transform 1 0 6992 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72
timestamp 1649977179
transform 1 0 7728 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76
timestamp 1649977179
transform 1 0 8096 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1649977179
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_87
timestamp 1649977179
transform 1 0 9108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_98
timestamp 1649977179
transform 1 0 10120 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_104 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10672 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1649977179
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_129
timestamp 1649977179
transform 1 0 12972 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_133
timestamp 1649977179
transform 1 0 13340 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1649977179
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_149
timestamp 1649977179
transform 1 0 14812 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_156 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15456 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_177 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_180
timestamp 1649977179
transform 1 0 17664 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_184
timestamp 1649977179
transform 1 0 18032 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_188
timestamp 1649977179
transform 1 0 18400 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1649977179
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_215
timestamp 1649977179
transform 1 0 20884 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_219
timestamp 1649977179
transform 1 0 21252 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_6
timestamp 1649977179
transform 1 0 1656 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_12
timestamp 1649977179
transform 1 0 2208 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_18
timestamp 1649977179
transform 1 0 2760 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_22
timestamp 1649977179
transform 1 0 3128 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_34
timestamp 1649977179
transform 1 0 4232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_42
timestamp 1649977179
transform 1 0 4968 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_48
timestamp 1649977179
transform 1 0 5520 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1649977179
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_76
timestamp 1649977179
transform 1 0 8096 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_84
timestamp 1649977179
transform 1 0 8832 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_92
timestamp 1649977179
transform 1 0 9568 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1649977179
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_129
timestamp 1649977179
transform 1 0 12972 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_135
timestamp 1649977179
transform 1 0 13524 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_141
timestamp 1649977179
transform 1 0 14076 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_149
timestamp 1649977179
transform 1 0 14812 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_155
timestamp 1649977179
transform 1 0 15364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_161
timestamp 1649977179
transform 1 0 15916 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1649977179
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_178
timestamp 1649977179
transform 1 0 17480 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_183
timestamp 1649977179
transform 1 0 17940 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_187
timestamp 1649977179
transform 1 0 18308 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_205
timestamp 1649977179
transform 1 0 19964 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_219
timestamp 1649977179
transform 1 0 21252 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1649977179
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_32
timestamp 1649977179
transform 1 0 4048 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_36
timestamp 1649977179
transform 1 0 4416 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_49
timestamp 1649977179
transform 1 0 5612 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_60
timestamp 1649977179
transform 1 0 6624 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_64
timestamp 1649977179
transform 1 0 6992 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_74
timestamp 1649977179
transform 1 0 7912 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1649977179
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_90
timestamp 1649977179
transform 1 0 9384 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_108
timestamp 1649977179
transform 1 0 11040 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_126
timestamp 1649977179
transform 1 0 12696 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_130
timestamp 1649977179
transform 1 0 13064 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1649977179
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_157
timestamp 1649977179
transform 1 0 15548 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_161
timestamp 1649977179
transform 1 0 15916 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_169
timestamp 1649977179
transform 1 0 16652 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_188
timestamp 1649977179
transform 1 0 18400 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1649977179
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_213
timestamp 1649977179
transform 1 0 20700 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_217
timestamp 1649977179
transform 1 0 21068 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_221
timestamp 1649977179
transform 1 0 21436 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_23
timestamp 1649977179
transform 1 0 3220 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_27
timestamp 1649977179
transform 1 0 3588 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_30
timestamp 1649977179
transform 1 0 3864 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_34
timestamp 1649977179
transform 1 0 4232 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_38
timestamp 1649977179
transform 1 0 4600 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_42
timestamp 1649977179
transform 1 0 4968 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_53
timestamp 1649977179
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_63
timestamp 1649977179
transform 1 0 6900 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_67
timestamp 1649977179
transform 1 0 7268 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_74
timestamp 1649977179
transform 1 0 7912 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_83
timestamp 1649977179
transform 1 0 8740 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_94
timestamp 1649977179
transform 1 0 9752 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_106
timestamp 1649977179
transform 1 0 10856 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1649977179
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_141
timestamp 1649977179
transform 1 0 14076 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_159
timestamp 1649977179
transform 1 0 15732 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_163
timestamp 1649977179
transform 1 0 16100 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_185
timestamp 1649977179
transform 1 0 18124 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_203
timestamp 1649977179
transform 1 0 19780 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_221
timestamp 1649977179
transform 1 0 21436 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_21
timestamp 1649977179
transform 1 0 3036 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_25
timestamp 1649977179
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_31
timestamp 1649977179
transform 1 0 3956 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_35
timestamp 1649977179
transform 1 0 4324 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_39
timestamp 1649977179
transform 1 0 4692 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_45
timestamp 1649977179
transform 1 0 5244 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_56
timestamp 1649977179
transform 1 0 6256 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_69
timestamp 1649977179
transform 1 0 7452 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_77
timestamp 1649977179
transform 1 0 8188 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1649977179
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_96
timestamp 1649977179
transform 1 0 9936 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_100
timestamp 1649977179
transform 1 0 10304 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_108
timestamp 1649977179
transform 1 0 11040 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_126
timestamp 1649977179
transform 1 0 12696 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_130
timestamp 1649977179
transform 1 0 13064 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1649977179
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_143
timestamp 1649977179
transform 1 0 14260 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_147
timestamp 1649977179
transform 1 0 14628 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_164
timestamp 1649977179
transform 1 0 16192 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_168
timestamp 1649977179
transform 1 0 16560 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_172
timestamp 1649977179
transform 1 0 16928 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_176
timestamp 1649977179
transform 1 0 17296 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1649977179
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_213
timestamp 1649977179
transform 1 0 20700 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_217
timestamp 1649977179
transform 1 0 21068 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_221
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_5
timestamp 1649977179
transform 1 0 1564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_10
timestamp 1649977179
transform 1 0 2024 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_21
timestamp 1649977179
transform 1 0 3036 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_32
timestamp 1649977179
transform 1 0 4048 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_37
timestamp 1649977179
transform 1 0 4508 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_48
timestamp 1649977179
transform 1 0 5520 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1649977179
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_66
timestamp 1649977179
transform 1 0 7176 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_70
timestamp 1649977179
transform 1 0 7544 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_78
timestamp 1649977179
transform 1 0 8280 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_82
timestamp 1649977179
transform 1 0 8648 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_92
timestamp 1649977179
transform 1 0 9568 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1649977179
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_129
timestamp 1649977179
transform 1 0 12972 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_133
timestamp 1649977179
transform 1 0 13340 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_137
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_145
timestamp 1649977179
transform 1 0 14444 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_162
timestamp 1649977179
transform 1 0 16008 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1649977179
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_185
timestamp 1649977179
transform 1 0 18124 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_189
timestamp 1649977179
transform 1 0 18492 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_193
timestamp 1649977179
transform 1 0 18860 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_196
timestamp 1649977179
transform 1 0 19136 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_200
timestamp 1649977179
transform 1 0 19504 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_218
timestamp 1649977179
transform 1 0 21160 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_222
timestamp 1649977179
transform 1 0 21528 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_12
timestamp 1649977179
transform 1 0 2208 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_23
timestamp 1649977179
transform 1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_31
timestamp 1649977179
transform 1 0 3956 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_35
timestamp 1649977179
transform 1 0 4324 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_46
timestamp 1649977179
transform 1 0 5336 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_50
timestamp 1649977179
transform 1 0 5704 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_61
timestamp 1649977179
transform 1 0 6716 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_65
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_76
timestamp 1649977179
transform 1 0 8096 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1649977179
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_94
timestamp 1649977179
transform 1 0 9752 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_99
timestamp 1649977179
transform 1 0 10212 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_107
timestamp 1649977179
transform 1 0 10948 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_110
timestamp 1649977179
transform 1 0 11224 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_128
timestamp 1649977179
transform 1 0 12880 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_132
timestamp 1649977179
transform 1 0 13248 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_135
timestamp 1649977179
transform 1 0 13524 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_157
timestamp 1649977179
transform 1 0 15548 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_161
timestamp 1649977179
transform 1 0 15916 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_189
timestamp 1649977179
transform 1 0 18492 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_193
timestamp 1649977179
transform 1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_214
timestamp 1649977179
transform 1 0 20792 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_219
timestamp 1649977179
transform 1 0 21252 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_18
timestamp 1649977179
transform 1 0 2760 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_23
timestamp 1649977179
transform 1 0 3220 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_31
timestamp 1649977179
transform 1 0 3956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_35
timestamp 1649977179
transform 1 0 4324 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_43
timestamp 1649977179
transform 1 0 5060 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1649977179
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1649977179
transform 1 0 6532 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_70
timestamp 1649977179
transform 1 0 7544 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_76
timestamp 1649977179
transform 1 0 8096 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_87
timestamp 1649977179
transform 1 0 9108 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_92
timestamp 1649977179
transform 1 0 9568 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_104
timestamp 1649977179
transform 1 0 10672 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_133
timestamp 1649977179
transform 1 0 13340 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_153
timestamp 1649977179
transform 1 0 15180 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_157
timestamp 1649977179
transform 1 0 15548 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_165
timestamp 1649977179
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_185
timestamp 1649977179
transform 1 0 18124 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_189
timestamp 1649977179
transform 1 0 18492 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_197
timestamp 1649977179
transform 1 0 19228 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_215
timestamp 1649977179
transform 1 0 20884 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_219
timestamp 1649977179
transform 1 0 21252 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_8
timestamp 1649977179
transform 1 0 1840 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_19
timestamp 1649977179
transform 1 0 2852 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_23
timestamp 1649977179
transform 1 0 3220 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1649977179
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_38
timestamp 1649977179
transform 1 0 4600 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_42
timestamp 1649977179
transform 1 0 4968 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_65
timestamp 1649977179
transform 1 0 7084 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_73
timestamp 1649977179
transform 1 0 7820 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_78
timestamp 1649977179
transform 1 0 8280 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1649977179
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_94
timestamp 1649977179
transform 1 0 9752 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_99
timestamp 1649977179
transform 1 0 10212 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_111
timestamp 1649977179
transform 1 0 11316 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_117
timestamp 1649977179
transform 1 0 11868 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_134
timestamp 1649977179
transform 1 0 13432 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1649977179
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_163
timestamp 1649977179
transform 1 0 16100 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_167
timestamp 1649977179
transform 1 0 16468 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_186
timestamp 1649977179
transform 1 0 18216 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_190
timestamp 1649977179
transform 1 0 18584 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_199
timestamp 1649977179
transform 1 0 19412 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_217
timestamp 1649977179
transform 1 0 21068 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_221
timestamp 1649977179
transform 1 0 21436 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_7
timestamp 1649977179
transform 1 0 1748 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_12
timestamp 1649977179
transform 1 0 2208 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_16
timestamp 1649977179
transform 1 0 2576 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_22
timestamp 1649977179
transform 1 0 3128 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_26
timestamp 1649977179
transform 1 0 3496 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_37
timestamp 1649977179
transform 1 0 4508 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_48
timestamp 1649977179
transform 1 0 5520 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1649977179
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_63
timestamp 1649977179
transform 1 0 6900 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_74
timestamp 1649977179
transform 1 0 7912 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_82
timestamp 1649977179
transform 1 0 8648 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_94
timestamp 1649977179
transform 1 0 9752 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_106
timestamp 1649977179
transform 1 0 10856 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_129
timestamp 1649977179
transform 1 0 12972 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_133
timestamp 1649977179
transform 1 0 13340 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_155
timestamp 1649977179
transform 1 0 15364 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_161
timestamp 1649977179
transform 1 0 15916 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_165
timestamp 1649977179
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_193
timestamp 1649977179
transform 1 0 18860 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_211
timestamp 1649977179
transform 1 0 20516 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_215
timestamp 1649977179
transform 1 0 20884 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_219
timestamp 1649977179
transform 1 0 21252 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_15
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_19
timestamp 1649977179
transform 1 0 2852 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_22
timestamp 1649977179
transform 1 0 3128 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1649977179
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_31
timestamp 1649977179
transform 1 0 3956 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_42
timestamp 1649977179
transform 1 0 4968 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_53
timestamp 1649977179
transform 1 0 5980 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_57
timestamp 1649977179
transform 1 0 6348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_60
timestamp 1649977179
transform 1 0 6624 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_64
timestamp 1649977179
transform 1 0 6992 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_75
timestamp 1649977179
transform 1 0 8004 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_79
timestamp 1649977179
transform 1 0 8372 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1649977179
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_87
timestamp 1649977179
transform 1 0 9108 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_98
timestamp 1649977179
transform 1 0 10120 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_110
timestamp 1649977179
transform 1 0 11224 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_127
timestamp 1649977179
transform 1 0 12788 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_133
timestamp 1649977179
transform 1 0 13340 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_137
timestamp 1649977179
transform 1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_159
timestamp 1649977179
transform 1 0 15732 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_177
timestamp 1649977179
transform 1 0 17388 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_181
timestamp 1649977179
transform 1 0 17756 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_187
timestamp 1649977179
transform 1 0 18308 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1649977179
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_213
timestamp 1649977179
transform 1 0 20700 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_217
timestamp 1649977179
transform 1 0 21068 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_221
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_15
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_21
timestamp 1649977179
transform 1 0 3036 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_25
timestamp 1649977179
transform 1 0 3404 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_28
timestamp 1649977179
transform 1 0 3680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_39
timestamp 1649977179
transform 1 0 4692 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_50
timestamp 1649977179
transform 1 0 5704 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1649977179
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_63
timestamp 1649977179
transform 1 0 6900 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_74
timestamp 1649977179
transform 1 0 7912 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_85
timestamp 1649977179
transform 1 0 8924 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_89
timestamp 1649977179
transform 1 0 9292 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_99
timestamp 1649977179
transform 1 0 10212 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_107
timestamp 1649977179
transform 1 0 10948 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1649977179
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_131
timestamp 1649977179
transform 1 0 13156 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_149
timestamp 1649977179
transform 1 0 14812 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_153
timestamp 1649977179
transform 1 0 15180 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_157
timestamp 1649977179
transform 1 0 15548 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_160
timestamp 1649977179
transform 1 0 15824 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_185
timestamp 1649977179
transform 1 0 18124 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_203
timestamp 1649977179
transform 1 0 19780 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_221
timestamp 1649977179
transform 1 0 21436 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_13
timestamp 1649977179
transform 1 0 2300 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1649977179
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_32
timestamp 1649977179
transform 1 0 4048 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_43
timestamp 1649977179
transform 1 0 5060 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_49
timestamp 1649977179
transform 1 0 5612 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_53
timestamp 1649977179
transform 1 0 5980 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_56
timestamp 1649977179
transform 1 0 6256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_61
timestamp 1649977179
transform 1 0 6716 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_66
timestamp 1649977179
transform 1 0 7176 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_77
timestamp 1649977179
transform 1 0 8188 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_81
timestamp 1649977179
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_87
timestamp 1649977179
transform 1 0 9108 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_92
timestamp 1649977179
transform 1 0 9568 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_110
timestamp 1649977179
transform 1 0 11224 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_128
timestamp 1649977179
transform 1 0 12880 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_132
timestamp 1649977179
transform 1 0 13248 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_158
timestamp 1649977179
transform 1 0 15640 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_177
timestamp 1649977179
transform 1 0 17388 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_181
timestamp 1649977179
transform 1 0 17756 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_187
timestamp 1649977179
transform 1 0 18308 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_191
timestamp 1649977179
transform 1 0 18676 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1649977179
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_200
timestamp 1649977179
transform 1 0 19504 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_218
timestamp 1649977179
transform 1 0 21160 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_222
timestamp 1649977179
transform 1 0 21528 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_15
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_21
timestamp 1649977179
transform 1 0 3036 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_24
timestamp 1649977179
transform 1 0 3312 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_35
timestamp 1649977179
transform 1 0 4324 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_47
timestamp 1649977179
transform 1 0 5428 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_51
timestamp 1649977179
transform 1 0 5796 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1649977179
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_66
timestamp 1649977179
transform 1 0 7176 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_77
timestamp 1649977179
transform 1 0 8188 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_82
timestamp 1649977179
transform 1 0 8648 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_88
timestamp 1649977179
transform 1 0 9200 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_99
timestamp 1649977179
transform 1 0 10212 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1649977179
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_129
timestamp 1649977179
transform 1 0 12972 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_133
timestamp 1649977179
transform 1 0 13340 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_145
timestamp 1649977179
transform 1 0 14444 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_157
timestamp 1649977179
transform 1 0 15548 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_165
timestamp 1649977179
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_189
timestamp 1649977179
transform 1 0 18492 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_194
timestamp 1649977179
transform 1 0 18952 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_214
timestamp 1649977179
transform 1 0 20792 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_218
timestamp 1649977179
transform 1 0 21160 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_221
timestamp 1649977179
transform 1 0 21436 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_15
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_18
timestamp 1649977179
transform 1 0 2760 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_22
timestamp 1649977179
transform 1 0 3128 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1649977179
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_33
timestamp 1649977179
transform 1 0 4140 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_45
timestamp 1649977179
transform 1 0 5244 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_56
timestamp 1649977179
transform 1 0 6256 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_60
timestamp 1649977179
transform 1 0 6624 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_63
timestamp 1649977179
transform 1 0 6900 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_67
timestamp 1649977179
transform 1 0 7268 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_71
timestamp 1649977179
transform 1 0 7636 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1649977179
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_94
timestamp 1649977179
transform 1 0 9752 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_98
timestamp 1649977179
transform 1 0 10120 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_102
timestamp 1649977179
transform 1 0 10488 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_121
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_125
timestamp 1649977179
transform 1 0 12604 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_137
timestamp 1649977179
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_145
timestamp 1649977179
transform 1 0 14444 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_148
timestamp 1649977179
transform 1 0 14720 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_160
timestamp 1649977179
transform 1 0 15824 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_166
timestamp 1649977179
transform 1 0 16376 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_174
timestamp 1649977179
transform 1 0 17112 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_192
timestamp 1649977179
transform 1 0 18768 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_213
timestamp 1649977179
transform 1 0 20700 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_217
timestamp 1649977179
transform 1 0 21068 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_221
timestamp 1649977179
transform 1 0 21436 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_18
timestamp 1649977179
transform 1 0 2760 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_24
timestamp 1649977179
transform 1 0 3312 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_35
timestamp 1649977179
transform 1 0 4324 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_48
timestamp 1649977179
transform 1 0 5520 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 1649977179
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_61
timestamp 1649977179
transform 1 0 6716 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_72
timestamp 1649977179
transform 1 0 7728 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_77
timestamp 1649977179
transform 1 0 8188 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_90
timestamp 1649977179
transform 1 0 9384 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_94
timestamp 1649977179
transform 1 0 9752 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_99
timestamp 1649977179
transform 1 0 10212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_119
timestamp 1649977179
transform 1 0 12052 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_122
timestamp 1649977179
transform 1 0 12328 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_146
timestamp 1649977179
transform 1 0 14536 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_164
timestamp 1649977179
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_185
timestamp 1649977179
transform 1 0 18124 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_203
timestamp 1649977179
transform 1 0 19780 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_221
timestamp 1649977179
transform 1 0 21436 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_5
timestamp 1649977179
transform 1 0 1564 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_16
timestamp 1649977179
transform 1 0 2576 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_21
timestamp 1649977179
transform 1 0 3036 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1649977179
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_33
timestamp 1649977179
transform 1 0 4140 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_46
timestamp 1649977179
transform 1 0 5336 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_57
timestamp 1649977179
transform 1 0 6348 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_64
timestamp 1649977179
transform 1 0 6992 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_68
timestamp 1649977179
transform 1 0 7360 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_71
timestamp 1649977179
transform 1 0 7636 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1649977179
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_88
timestamp 1649977179
transform 1 0 9200 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_92
timestamp 1649977179
transform 1 0 9568 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_96
timestamp 1649977179
transform 1 0 9936 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_100
timestamp 1649977179
transform 1 0 10304 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_120
timestamp 1649977179
transform 1 0 12144 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1649977179
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_143
timestamp 1649977179
transform 1 0 14260 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_161
timestamp 1649977179
transform 1 0 15916 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_179
timestamp 1649977179
transform 1 0 17572 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_183
timestamp 1649977179
transform 1 0 17940 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_187
timestamp 1649977179
transform 1 0 18308 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_191
timestamp 1649977179
transform 1 0 18676 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1649977179
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_214
timestamp 1649977179
transform 1 0 20792 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_218
timestamp 1649977179
transform 1 0 21160 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_222
timestamp 1649977179
transform 1 0 21528 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_9
timestamp 1649977179
transform 1 0 1932 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_20
timestamp 1649977179
transform 1 0 2944 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_25
timestamp 1649977179
transform 1 0 3404 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_29
timestamp 1649977179
transform 1 0 3772 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_40
timestamp 1649977179
transform 1 0 4784 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1649977179
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_66
timestamp 1649977179
transform 1 0 7176 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_70
timestamp 1649977179
transform 1 0 7544 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_81
timestamp 1649977179
transform 1 0 8556 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_92
timestamp 1649977179
transform 1 0 9568 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1649977179
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_115
timestamp 1649977179
transform 1 0 11684 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_135
timestamp 1649977179
transform 1 0 13524 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_139
timestamp 1649977179
transform 1 0 13892 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_158
timestamp 1649977179
transform 1 0 15640 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_162
timestamp 1649977179
transform 1 0 16008 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1649977179
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_185
timestamp 1649977179
transform 1 0 18124 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_203
timestamp 1649977179
transform 1 0 19780 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_221
timestamp 1649977179
transform 1 0 21436 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_9
timestamp 1649977179
transform 1 0 1932 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_20
timestamp 1649977179
transform 1 0 2944 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_24
timestamp 1649977179
transform 1 0 3312 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_33
timestamp 1649977179
transform 1 0 4140 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_44
timestamp 1649977179
transform 1 0 5152 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_49
timestamp 1649977179
transform 1 0 5612 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_60
timestamp 1649977179
transform 1 0 6624 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_71
timestamp 1649977179
transform 1 0 7636 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1649977179
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_87
timestamp 1649977179
transform 1 0 9108 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_98
timestamp 1649977179
transform 1 0 10120 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_109
timestamp 1649977179
transform 1 0 11132 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_114
timestamp 1649977179
transform 1 0 11592 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_132
timestamp 1649977179
transform 1 0 13248 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_136
timestamp 1649977179
transform 1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_153
timestamp 1649977179
transform 1 0 15180 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_157
timestamp 1649977179
transform 1 0 15548 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_174
timestamp 1649977179
transform 1 0 17112 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_178
timestamp 1649977179
transform 1 0 17480 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_190
timestamp 1649977179
transform 1 0 18584 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_18_197
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_205
timestamp 1649977179
transform 1 0 19964 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_217
timestamp 1649977179
transform 1 0 21068 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_221
timestamp 1649977179
transform 1 0 21436 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_5
timestamp 1649977179
transform 1 0 1564 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_13
timestamp 1649977179
transform 1 0 2300 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_19
timestamp 1649977179
transform 1 0 2852 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1649977179
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_39
timestamp 1649977179
transform 1 0 4692 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_43
timestamp 1649977179
transform 1 0 5060 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1649977179
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_61
timestamp 1649977179
transform 1 0 6716 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_66
timestamp 1649977179
transform 1 0 7176 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_77
timestamp 1649977179
transform 1 0 8188 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_81
timestamp 1649977179
transform 1 0 8556 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_85
timestamp 1649977179
transform 1 0 8924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_88
timestamp 1649977179
transform 1 0 9200 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_92
timestamp 1649977179
transform 1 0 9568 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_103
timestamp 1649977179
transform 1 0 10580 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_107
timestamp 1649977179
transform 1 0 10948 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_117
timestamp 1649977179
transform 1 0 11868 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_129
timestamp 1649977179
transform 1 0 12972 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_134
timestamp 1649977179
transform 1 0 13432 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_146
timestamp 1649977179
transform 1 0 14536 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_158
timestamp 1649977179
transform 1 0 15640 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1649977179
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1649977179
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1649977179
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1649977179
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1649977179
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_5
timestamp 1649977179
transform 1 0 1564 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_16
timestamp 1649977179
transform 1 0 2576 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1649977179
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_31
timestamp 1649977179
transform 1 0 3956 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_42
timestamp 1649977179
transform 1 0 4968 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_47
timestamp 1649977179
transform 1 0 5428 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_60
timestamp 1649977179
transform 1 0 6624 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_64
timestamp 1649977179
transform 1 0 6992 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_68
timestamp 1649977179
transform 1 0 7360 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_81
timestamp 1649977179
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_88
timestamp 1649977179
transform 1 0 9200 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_92
timestamp 1649977179
transform 1 0 9568 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_97
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_108
timestamp 1649977179
transform 1 0 11040 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_113
timestamp 1649977179
transform 1 0 11500 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_117
timestamp 1649977179
transform 1 0 11868 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_128
timestamp 1649977179
transform 1 0 12880 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1649977179
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1649977179
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1649977179
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1649977179
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1649977179
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_221
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_7
timestamp 1649977179
transform 1 0 1748 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_12
timestamp 1649977179
transform 1 0 2208 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_18
timestamp 1649977179
transform 1 0 2760 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_22
timestamp 1649977179
transform 1 0 3128 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_33
timestamp 1649977179
transform 1 0 4140 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_38
timestamp 1649977179
transform 1 0 4600 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_50
timestamp 1649977179
transform 1 0 5704 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1649977179
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_62
timestamp 1649977179
transform 1 0 6808 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_72
timestamp 1649977179
transform 1 0 7728 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_83
timestamp 1649977179
transform 1 0 8740 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_87
timestamp 1649977179
transform 1 0 9108 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_99
timestamp 1649977179
transform 1 0 10212 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1649977179
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_122
timestamp 1649977179
transform 1 0 12328 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_133
timestamp 1649977179
transform 1 0 13340 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_145
timestamp 1649977179
transform 1 0 14444 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_157
timestamp 1649977179
transform 1 0 15548 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_165
timestamp 1649977179
transform 1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1649977179
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1649977179
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1649977179
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1649977179
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_7
timestamp 1649977179
transform 1 0 1748 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_19
timestamp 1649977179
transform 1 0 2852 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1649977179
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_38
timestamp 1649977179
transform 1 0 4600 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_42
timestamp 1649977179
transform 1 0 4968 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_46
timestamp 1649977179
transform 1 0 5336 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_49
timestamp 1649977179
transform 1 0 5612 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_53
timestamp 1649977179
transform 1 0 5980 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_56
timestamp 1649977179
transform 1 0 6256 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_68
timestamp 1649977179
transform 1 0 7360 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1649977179
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_87
timestamp 1649977179
transform 1 0 9108 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_98
timestamp 1649977179
transform 1 0 10120 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_106
timestamp 1649977179
transform 1 0 10856 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_112
timestamp 1649977179
transform 1 0 11408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_116
timestamp 1649977179
transform 1 0 11776 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_124
timestamp 1649977179
transform 1 0 12512 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_128
timestamp 1649977179
transform 1 0 12880 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1649977179
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1649977179
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1649977179
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1649977179
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1649977179
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1649977179
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_221
timestamp 1649977179
transform 1 0 21436 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_7
timestamp 1649977179
transform 1 0 1748 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_12
timestamp 1649977179
transform 1 0 2208 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_24
timestamp 1649977179
transform 1 0 3312 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_32
timestamp 1649977179
transform 1 0 4048 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_43
timestamp 1649977179
transform 1 0 5060 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1649977179
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_59
timestamp 1649977179
transform 1 0 6532 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_72
timestamp 1649977179
transform 1 0 7728 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_77
timestamp 1649977179
transform 1 0 8188 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_89
timestamp 1649977179
transform 1 0 9292 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_101
timestamp 1649977179
transform 1 0 10396 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_109
timestamp 1649977179
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1649977179
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1649977179
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1649977179
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1649977179
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1649977179
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1649977179
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1649977179
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1649977179
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1649977179
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_9
timestamp 1649977179
transform 1 0 1932 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_15
timestamp 1649977179
transform 1 0 2484 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_21
timestamp 1649977179
transform 1 0 3036 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_24_41
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_50
timestamp 1649977179
transform 1 0 5704 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_54
timestamp 1649977179
transform 1 0 6072 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_66
timestamp 1649977179
transform 1 0 7176 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_76
timestamp 1649977179
transform 1 0 8096 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_81
timestamp 1649977179
transform 1 0 8556 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1649977179
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1649977179
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1649977179
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1649977179
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1649977179
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1649977179
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1649977179
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1649977179
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1649977179
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1649977179
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_221
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_7
timestamp 1649977179
transform 1 0 1748 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_12
timestamp 1649977179
transform 1 0 2208 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_24
timestamp 1649977179
transform 1 0 3312 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_36
timestamp 1649977179
transform 1 0 4416 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_42
timestamp 1649977179
transform 1 0 4968 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_45
timestamp 1649977179
transform 1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1649977179
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1649977179
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1649977179
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1649977179
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1649977179
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1649977179
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1649977179
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1649977179
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1649977179
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1649977179
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1649977179
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1649977179
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1649977179
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1649977179
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1649977179
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_33
timestamp 1649977179
transform 1 0 4140 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_40
timestamp 1649977179
transform 1 0 4784 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_52
timestamp 1649977179
transform 1 0 5888 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_59
timestamp 1649977179
transform 1 0 6532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_67
timestamp 1649977179
transform 1 0 7268 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_75
timestamp 1649977179
transform 1 0 8004 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1649977179
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_94
timestamp 1649977179
transform 1 0 9752 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_99
timestamp 1649977179
transform 1 0 10212 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_103
timestamp 1649977179
transform 1 0 10580 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_115
timestamp 1649977179
transform 1 0 11684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_127
timestamp 1649977179
transform 1 0 12788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1649977179
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1649977179
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1649977179
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1649977179
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1649977179
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1649977179
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_221
timestamp 1649977179
transform 1 0 21436 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_8
timestamp 1649977179
transform 1 0 1840 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_16
timestamp 1649977179
transform 1 0 2576 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_24
timestamp 1649977179
transform 1 0 3312 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_31
timestamp 1649977179
transform 1 0 3956 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_39
timestamp 1649977179
transform 1 0 4692 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_48
timestamp 1649977179
transform 1 0 5520 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_65
timestamp 1649977179
transform 1 0 7084 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_73
timestamp 1649977179
transform 1 0 7820 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_85
timestamp 1649977179
transform 1 0 8924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_97
timestamp 1649977179
transform 1 0 10028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_109
timestamp 1649977179
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1649977179
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1649977179
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1649977179
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1649977179
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1649977179
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1649977179
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1649977179
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1649977179
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1649977179
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_7
timestamp 1649977179
transform 1 0 1748 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_12
timestamp 1649977179
transform 1 0 2208 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 1649977179
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_34
timestamp 1649977179
transform 1 0 4232 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_42
timestamp 1649977179
transform 1 0 4968 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_54
timestamp 1649977179
transform 1 0 6072 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_62
timestamp 1649977179
transform 1 0 6808 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_69
timestamp 1649977179
transform 1 0 7452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_81
timestamp 1649977179
transform 1 0 8556 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1649977179
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1649977179
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1649977179
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1649977179
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1649977179
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1649977179
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1649977179
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1649977179
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1649977179
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1649977179
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1649977179
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_221
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1649977179
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1649977179
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_43
timestamp 1649977179
transform 1 0 5060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1649977179
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1649977179
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1649977179
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1649977179
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1649977179
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1649977179
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1649977179
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1649977179
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1649977179
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1649977179
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1649977179
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1649977179
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1649977179
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1649977179
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1649977179
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1649977179
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1649977179
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1649977179
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1649977179
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1649977179
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1649977179
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1649977179
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1649977179
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1649977179
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1649977179
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1649977179
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1649977179
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1649977179
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1649977179
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1649977179
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1649977179
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1649977179
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1649977179
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_221
timestamp 1649977179
transform 1 0 21436 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1649977179
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_27
timestamp 1649977179
transform 1 0 3588 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_35
timestamp 1649977179
transform 1 0 4324 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_40
timestamp 1649977179
transform 1 0 4784 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_52
timestamp 1649977179
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_69
timestamp 1649977179
transform 1 0 7452 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_77
timestamp 1649977179
transform 1 0 8188 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_85
timestamp 1649977179
transform 1 0 8924 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_97
timestamp 1649977179
transform 1 0 10028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_109
timestamp 1649977179
transform 1 0 11132 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1649977179
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1649977179
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1649977179
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1649977179
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1649977179
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1649977179
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1649977179
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1649977179
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1649977179
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1649977179
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1649977179
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_35
timestamp 1649977179
transform 1 0 4324 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_40
timestamp 1649977179
transform 1 0 4784 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_52
timestamp 1649977179
transform 1 0 5888 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_64
timestamp 1649977179
transform 1 0 6992 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_72
timestamp 1649977179
transform 1 0 7728 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1649977179
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1649977179
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1649977179
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1649977179
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1649977179
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1649977179
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1649977179
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1649977179
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1649977179
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1649977179
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1649977179
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1649977179
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_27
timestamp 1649977179
transform 1 0 3588 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_29
timestamp 1649977179
transform 1 0 3772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_41
timestamp 1649977179
transform 1 0 4876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_53
timestamp 1649977179
transform 1 0 5980 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1649977179
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_81
timestamp 1649977179
transform 1 0 8556 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_85
timestamp 1649977179
transform 1 0 8924 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_97
timestamp 1649977179
transform 1 0 10028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_109
timestamp 1649977179
transform 1 0 11132 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1649977179
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_137
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_141
timestamp 1649977179
transform 1 0 14076 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_153
timestamp 1649977179
transform 1 0 15180 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_165
timestamp 1649977179
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1649977179
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_193
timestamp 1649977179
transform 1 0 18860 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_197
timestamp 1649977179
transform 1 0 19228 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_209
timestamp 1649977179
transform 1 0 20332 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_221
timestamp 1649977179
transform 1 0 21436 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 21896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 21896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 21896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 21896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 21896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 21896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 21896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 21896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 21896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 21896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 21896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 21896 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 21896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 21896 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 21896 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 21896 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 21896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 21896 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 21896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 21896 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 21896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 21896 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 21896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 21896 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 21896 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 21896 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 21896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 21896 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 21896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 21896 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 21896 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 21896 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 3680 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 8832 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 13984 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _035_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2944 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1649977179
transform -1 0 4876 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1649977179
transform -1 0 16376 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1649977179
transform 1 0 5336 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1649977179
transform -1 0 6900 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1649977179
transform 1 0 6900 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1649977179
transform 1 0 8372 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1649977179
transform 1 0 6716 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1649977179
transform 1 0 7912 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1649977179
transform 1 0 8280 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1649977179
transform -1 0 5428 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1649977179
transform -1 0 7176 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1649977179
transform 1 0 2760 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1649977179
transform 1 0 11316 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1649977179
transform 1 0 9752 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1649977179
transform 1 0 13156 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1649977179
transform 1 0 9936 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1649977179
transform 1 0 2760 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1649977179
transform 1 0 3864 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1649977179
transform 1 0 4324 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1649977179
transform 1 0 8004 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1649977179
transform -1 0 6900 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1649977179
transform 1 0 9936 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1649977179
transform -1 0 8648 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1649977179
transform 1 0 9936 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1649977179
transform 1 0 9292 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1649977179
transform -1 0 9568 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _066_
timestamp 1649977179
transform -1 0 6716 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _067_
timestamp 1649977179
transform 1 0 5336 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _068_
timestamp 1649977179
transform 1 0 7912 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _069_
timestamp 1649977179
transform -1 0 9200 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _070_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18584 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1649977179
transform -1 0 1932 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1649977179
transform 1 0 2392 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1649977179
transform -1 0 2208 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1649977179
transform -1 0 2208 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1649977179
transform -1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1649977179
transform -1 0 2484 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1649977179
transform -1 0 3036 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1649977179
transform -1 0 1932 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1649977179
transform -1 0 2208 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1649977179
transform -1 0 1840 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1649977179
transform -1 0 3956 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1649977179
transform -1 0 2208 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1649977179
transform -1 0 4232 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1649977179
transform -1 0 4968 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1649977179
transform -1 0 5060 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1649977179
transform -1 0 4876 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1649977179
transform -1 0 4784 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1649977179
transform -1 0 4784 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1649977179
transform -1 0 5888 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1649977179
transform 1 0 9016 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1649977179
transform 1 0 5152 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1649977179
transform 1 0 8280 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1649977179
transform 1 0 4600 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1649977179
transform 1 0 14996 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1649977179
transform -1 0 5520 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1649977179
transform -1 0 6072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1649977179
transform -1 0 6992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1649977179
transform -1 0 8096 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1649977179
transform -1 0 6072 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1649977179
transform 1 0 10304 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1649977179
transform 1 0 13156 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1649977179
transform 1 0 13708 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1649977179
transform 1 0 15548 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1649977179
transform 1 0 15088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1649977179
transform 1 0 2392 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1649977179
transform 1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1649977179
transform 1 0 1840 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1649977179
transform 1 0 1840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 11224 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21436 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 16192 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 12696 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19412 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 21160 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18216 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15732 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 11040 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 18492 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 19780 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 16100 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15180 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 17020 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20700 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15548 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 16008 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15548 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20700 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18400 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18952 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 15916 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19412 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 20792 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21068 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 20516 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 17388 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18124 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16100 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18492 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12052 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 15640 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12880 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11960 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 13892 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 14812 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13800 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 12972 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12972 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13340 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 10764 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13156 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 12880 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 11224 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11224 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 14076 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12972 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11224 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12788 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 16192 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12972 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11224 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11776 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14168 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15916 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 10672 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14260 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 18308 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18860 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 19780 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 18308 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21436 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20792 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21436 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 20792 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21160 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18768 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 17112 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 14536 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19964 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4692 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1649977179
transform 1 0 5152 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1649977179
transform 1 0 6716 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1649977179
transform -1 0 5336 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1649977179
transform 1 0 6256 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 5244 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5060 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1649977179
transform -1 0 3036 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1649977179
transform 1 0 3220 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 2392 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1649977179
transform -1 0 2208 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1649977179
transform -1 0 2484 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2668 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1649977179
transform 1 0 5796 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1649977179
transform -1 0 6256 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1649977179
transform -1 0 7452 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6624 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 6900 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_0_
timestamp 1649977179
transform -1 0 4508 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_1_
timestamp 1649977179
transform 1 0 4140 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_0_
timestamp 1649977179
transform 1 0 3864 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_1_
timestamp 1649977179
transform -1 0 2852 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l3_in_0_
timestamp 1649977179
transform -1 0 4600 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 4508 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1649977179
transform -1 0 10120 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 14812 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l1_in_0_
timestamp 1649977179
transform -1 0 5980 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8096 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 7820 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_0_
timestamp 1649977179
transform -1 0 9108 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 8648 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_0_
timestamp 1649977179
transform -1 0 6716 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8740 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 8648 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9108 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8924 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 8740 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_0_
timestamp 1649977179
transform -1 0 8096 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 8280 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_0_
timestamp 1649977179
transform -1 0 10120 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9384 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7176 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7084 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 7176 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5152 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1649977179
transform 1 0 4876 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1649977179
transform -1 0 5520 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 7360 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l1_in_0_
timestamp 1649977179
transform -1 0 5520 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l2_in_0_
timestamp 1649977179
transform -1 0 7728 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 9016 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_29.mux_l1_in_0_
timestamp 1649977179
transform -1 0 9384 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_29.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9384 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 8832 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5796 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1649977179
transform 1 0 7360 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1649977179
transform 1 0 5796 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5244 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1649977179
transform 1 0 4968 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4324 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3588 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1649977179
transform 1 0 4600 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1649977179
transform 1 0 4416 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4232 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1649977179
transform -1 0 3312 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1649977179
transform 1 0 3496 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 1932 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 3956 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1649977179
transform -1 0 2944 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1649977179
transform -1 0 2576 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 2116 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1649977179
transform 1 0 1932 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1649977179
transform 1 0 1748 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1748 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1649977179
transform -1 0 6256 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1649977179
transform 1 0 7820 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5520 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1649977179
transform -1 0 4324 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4508 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3496 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1649977179
transform 1 0 4140 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1649977179
transform -1 0 4140 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2484 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7360 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7084 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3496 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7820 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3312 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10396 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7360 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 4048 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7820 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 4876 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8740 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7728 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 5704 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7912 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6900 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 4784 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9292 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7268 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 5520 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5244 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1649977179
transform 1 0 4876 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4232 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2576 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6808 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 6532 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10212 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7728 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 7268 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10304 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9292 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 8004 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9384 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 7452 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1649977179
transform -1 0 10580 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1649977179
transform 1 0 12144 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 7820 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l1_in_0_
timestamp 1649977179
transform 1 0 12512 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l2_in_0_
timestamp 1649977179
transform 1 0 10396 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 7728 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l1_in_0_
timestamp 1649977179
transform 1 0 12052 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_39.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 8924 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20148 0 -1 3264
box -38 -48 1142 592
<< labels >>
flabel metal2 s 20074 0 20130 800 0 FreeSans 224 90 0 0 SC_IN_BOT
port 0 nsew signal input
flabel metal2 s 20442 0 20498 800 0 FreeSans 224 90 0 0 SC_OUT_BOT
port 1 nsew signal tristate
flabel metal4 s 6142 2128 6462 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 11340 2128 11660 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 16538 2128 16858 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 21736 2128 22056 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 3543 2128 3863 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal4 s 8741 2128 9061 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal4 s 13939 2128 14259 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal4 s 19137 2128 19457 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal2 s 2042 0 2098 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_42_
port 4 nsew signal input
flabel metal2 s 2410 0 2466 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_43_
port 5 nsew signal input
flabel metal2 s 2778 0 2834 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_44_
port 6 nsew signal input
flabel metal2 s 3146 0 3202 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_45_
port 7 nsew signal input
flabel metal2 s 3514 0 3570 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_46_
port 8 nsew signal input
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_47_
port 9 nsew signal input
flabel metal2 s 4250 0 4306 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_48_
port 10 nsew signal input
flabel metal2 s 4618 0 4674 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_49_
port 11 nsew signal input
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 bottom_right_grid_pin_1_
port 12 nsew signal input
flabel metal3 s 22200 5720 23000 5840 0 FreeSans 480 0 0 0 ccff_head
port 13 nsew signal input
flabel metal3 s 22200 17144 23000 17264 0 FreeSans 480 0 0 0 ccff_tail
port 14 nsew signal tristate
flabel metal3 s 0 4904 800 5024 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 15 nsew signal input
flabel metal3 s 0 8984 800 9104 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 16 nsew signal input
flabel metal3 s 0 9392 800 9512 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 17 nsew signal input
flabel metal3 s 0 9800 800 9920 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 18 nsew signal input
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 19 nsew signal input
flabel metal3 s 0 10616 800 10736 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 20 nsew signal input
flabel metal3 s 0 11024 800 11144 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 21 nsew signal input
flabel metal3 s 0 11432 800 11552 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 22 nsew signal input
flabel metal3 s 0 11840 800 11960 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 23 nsew signal input
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 24 nsew signal input
flabel metal3 s 0 12656 800 12776 0 FreeSans 480 0 0 0 chanx_left_in[19]
port 25 nsew signal input
flabel metal3 s 0 5312 800 5432 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 26 nsew signal input
flabel metal3 s 0 5720 800 5840 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 27 nsew signal input
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 28 nsew signal input
flabel metal3 s 0 6536 800 6656 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 29 nsew signal input
flabel metal3 s 0 6944 800 7064 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 30 nsew signal input
flabel metal3 s 0 7352 800 7472 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 31 nsew signal input
flabel metal3 s 0 7760 800 7880 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 32 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 33 nsew signal input
flabel metal3 s 0 8576 800 8696 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 34 nsew signal input
flabel metal3 s 0 13064 800 13184 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 35 nsew signal tristate
flabel metal3 s 0 17144 800 17264 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 36 nsew signal tristate
flabel metal3 s 0 17552 800 17672 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 37 nsew signal tristate
flabel metal3 s 0 17960 800 18080 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 38 nsew signal tristate
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 39 nsew signal tristate
flabel metal3 s 0 18776 800 18896 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 40 nsew signal tristate
flabel metal3 s 0 19184 800 19304 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 41 nsew signal tristate
flabel metal3 s 0 19592 800 19712 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 42 nsew signal tristate
flabel metal3 s 0 20000 800 20120 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 43 nsew signal tristate
flabel metal3 s 0 20408 800 20528 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 44 nsew signal tristate
flabel metal3 s 0 20816 800 20936 0 FreeSans 480 0 0 0 chanx_left_out[19]
port 45 nsew signal tristate
flabel metal3 s 0 13472 800 13592 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 46 nsew signal tristate
flabel metal3 s 0 13880 800 14000 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 47 nsew signal tristate
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 48 nsew signal tristate
flabel metal3 s 0 14696 800 14816 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 49 nsew signal tristate
flabel metal3 s 0 15104 800 15224 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 50 nsew signal tristate
flabel metal3 s 0 15512 800 15632 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 51 nsew signal tristate
flabel metal3 s 0 15920 800 16040 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 52 nsew signal tristate
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 53 nsew signal tristate
flabel metal3 s 0 16736 800 16856 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 54 nsew signal tristate
flabel metal2 s 4986 0 5042 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 55 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 56 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 57 nsew signal input
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 58 nsew signal input
flabel metal2 s 9770 0 9826 800 0 FreeSans 224 90 0 0 chany_bottom_in[13]
port 59 nsew signal input
flabel metal2 s 10138 0 10194 800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 60 nsew signal input
flabel metal2 s 10506 0 10562 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 61 nsew signal input
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 chany_bottom_in[16]
port 62 nsew signal input
flabel metal2 s 11242 0 11298 800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 63 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 64 nsew signal input
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 chany_bottom_in[19]
port 65 nsew signal input
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 66 nsew signal input
flabel metal2 s 5722 0 5778 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 67 nsew signal input
flabel metal2 s 6090 0 6146 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 68 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 69 nsew signal input
flabel metal2 s 6826 0 6882 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 70 nsew signal input
flabel metal2 s 7194 0 7250 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 71 nsew signal input
flabel metal2 s 7562 0 7618 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 72 nsew signal input
flabel metal2 s 7930 0 7986 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 73 nsew signal input
flabel metal2 s 8298 0 8354 800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 74 nsew signal input
flabel metal2 s 12346 0 12402 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 75 nsew signal tristate
flabel metal2 s 16026 0 16082 800 0 FreeSans 224 90 0 0 chany_bottom_out[10]
port 76 nsew signal tristate
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 chany_bottom_out[11]
port 77 nsew signal tristate
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 chany_bottom_out[12]
port 78 nsew signal tristate
flabel metal2 s 17130 0 17186 800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 79 nsew signal tristate
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 chany_bottom_out[14]
port 80 nsew signal tristate
flabel metal2 s 17866 0 17922 800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 81 nsew signal tristate
flabel metal2 s 18234 0 18290 800 0 FreeSans 224 90 0 0 chany_bottom_out[16]
port 82 nsew signal tristate
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 83 nsew signal tristate
flabel metal2 s 18970 0 19026 800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 84 nsew signal tristate
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 chany_bottom_out[19]
port 85 nsew signal tristate
flabel metal2 s 12714 0 12770 800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 86 nsew signal tristate
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 87 nsew signal tristate
flabel metal2 s 13450 0 13506 800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 88 nsew signal tristate
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 89 nsew signal tristate
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 90 nsew signal tristate
flabel metal2 s 14554 0 14610 800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 91 nsew signal tristate
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 92 nsew signal tristate
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 chany_bottom_out[8]
port 93 nsew signal tristate
flabel metal2 s 15658 0 15714 800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 94 nsew signal tristate
flabel metal3 s 0 1640 800 1760 0 FreeSans 480 0 0 0 left_bottom_grid_pin_34_
port 95 nsew signal input
flabel metal3 s 0 2048 800 2168 0 FreeSans 480 0 0 0 left_bottom_grid_pin_35_
port 96 nsew signal input
flabel metal3 s 0 2456 800 2576 0 FreeSans 480 0 0 0 left_bottom_grid_pin_36_
port 97 nsew signal input
flabel metal3 s 0 2864 800 2984 0 FreeSans 480 0 0 0 left_bottom_grid_pin_37_
port 98 nsew signal input
flabel metal3 s 0 3272 800 3392 0 FreeSans 480 0 0 0 left_bottom_grid_pin_38_
port 99 nsew signal input
flabel metal3 s 0 3680 800 3800 0 FreeSans 480 0 0 0 left_bottom_grid_pin_39_
port 100 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 left_bottom_grid_pin_40_
port 101 nsew signal input
flabel metal3 s 0 4496 800 4616 0 FreeSans 480 0 0 0 left_bottom_grid_pin_41_
port 102 nsew signal input
flabel metal3 s 0 21224 800 21344 0 FreeSans 480 0 0 0 left_top_grid_pin_1_
port 103 nsew signal input
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 prog_clk_0_S_in
port 104 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
