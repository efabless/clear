magic
tech sky130A
magscale 1 2
timestamp 1625784957
<< locali >>
rect 3157 20383 3191 20553
rect 12173 19771 12207 20009
rect 12633 19907 12667 20009
rect 2513 19159 2547 19397
rect 4261 19227 4295 19465
rect 15669 18071 15703 18309
rect 3617 17527 3651 17765
rect 6285 17595 6319 17697
rect 7113 17527 7147 17697
rect 3801 15895 3835 15997
rect 12357 15487 12391 15657
rect 8125 14807 8159 15113
rect 14473 14331 14507 14433
rect 4169 11543 4203 11781
rect 7113 11067 7147 11305
rect 7021 7191 7055 7497
<< viali >>
rect 3157 20553 3191 20587
rect 10885 20553 10919 20587
rect 12725 20553 12759 20587
rect 16773 20553 16807 20587
rect 2421 20485 2455 20519
rect 2973 20485 3007 20519
rect 7297 20485 7331 20519
rect 7849 20485 7883 20519
rect 12081 20485 12115 20519
rect 13093 20485 13127 20519
rect 13645 20485 13679 20519
rect 14749 20485 14783 20519
rect 16313 20485 16347 20519
rect 17693 20485 17727 20519
rect 18245 20485 18279 20519
rect 18797 20485 18831 20519
rect 20085 20485 20119 20519
rect 3525 20417 3559 20451
rect 4629 20417 4663 20451
rect 6101 20417 6135 20451
rect 9873 20417 9907 20451
rect 9965 20417 9999 20451
rect 11529 20417 11563 20451
rect 17233 20417 17267 20451
rect 1685 20349 1719 20383
rect 1869 20349 1903 20383
rect 3157 20349 3191 20383
rect 3341 20349 3375 20383
rect 4537 20349 4571 20383
rect 7481 20349 7515 20383
rect 8585 20349 8619 20383
rect 10609 20349 10643 20383
rect 12265 20349 12299 20383
rect 15761 20349 15795 20383
rect 20269 20349 20303 20383
rect 20821 20349 20855 20383
rect 21281 20349 21315 20383
rect 2237 20281 2271 20315
rect 2789 20281 2823 20315
rect 6837 20281 6871 20315
rect 8033 20281 8067 20315
rect 11345 20281 11379 20315
rect 12633 20281 12667 20315
rect 13277 20281 13311 20315
rect 13829 20281 13863 20315
rect 14933 20281 14967 20315
rect 15577 20281 15611 20315
rect 16129 20281 16163 20315
rect 16681 20281 16715 20315
rect 17877 20281 17911 20315
rect 18429 20281 18463 20315
rect 18981 20281 19015 20315
rect 4077 20213 4111 20247
rect 4445 20213 4479 20247
rect 5089 20213 5123 20247
rect 5457 20213 5491 20247
rect 5825 20213 5859 20247
rect 5917 20213 5951 20247
rect 6929 20213 6963 20247
rect 8401 20213 8435 20247
rect 9413 20213 9447 20247
rect 9781 20213 9815 20247
rect 10425 20213 10459 20247
rect 19349 20213 19383 20247
rect 21189 20213 21223 20247
rect 3065 20009 3099 20043
rect 4813 20009 4847 20043
rect 7205 20009 7239 20043
rect 8401 20009 8435 20043
rect 8493 20009 8527 20043
rect 12173 20009 12207 20043
rect 12541 20009 12575 20043
rect 12633 20009 12667 20043
rect 12817 20009 12851 20043
rect 13369 20009 13403 20043
rect 17693 20009 17727 20043
rect 18337 20009 18371 20043
rect 6662 19941 6696 19975
rect 11170 19941 11204 19975
rect 1777 19873 1811 19907
rect 2329 19873 2363 19907
rect 3157 19873 3191 19907
rect 4077 19873 4111 19907
rect 4905 19873 4939 19907
rect 6929 19873 6963 19907
rect 7389 19873 7423 19907
rect 9505 19873 9539 19907
rect 11437 19873 11471 19907
rect 11897 19873 11931 19907
rect 2973 19805 3007 19839
rect 4721 19805 4755 19839
rect 8585 19805 8619 19839
rect 15393 19941 15427 19975
rect 15945 19941 15979 19975
rect 16497 19941 16531 19975
rect 17049 19941 17083 19975
rect 19993 19941 20027 19975
rect 20545 19941 20579 19975
rect 21097 19941 21131 19975
rect 12357 19873 12391 19907
rect 12633 19873 12667 19907
rect 13185 19873 13219 19907
rect 13829 19873 13863 19907
rect 14657 19873 14691 19907
rect 15577 19873 15611 19907
rect 16129 19873 16163 19907
rect 16681 19873 16715 19907
rect 17233 19873 17267 19907
rect 17785 19873 17819 19907
rect 18153 19873 18187 19907
rect 18613 19873 18647 19907
rect 20177 19873 20211 19907
rect 20729 19873 20763 19907
rect 21281 19873 21315 19907
rect 19625 19805 19659 19839
rect 1593 19737 1627 19771
rect 2513 19737 2547 19771
rect 5549 19737 5583 19771
rect 10057 19737 10091 19771
rect 12081 19737 12115 19771
rect 12173 19737 12207 19771
rect 13645 19737 13679 19771
rect 19073 19737 19107 19771
rect 3525 19669 3559 19703
rect 5273 19669 5307 19703
rect 7665 19669 7699 19703
rect 8033 19669 8067 19703
rect 9321 19669 9355 19703
rect 14841 19669 14875 19703
rect 18797 19669 18831 19703
rect 4261 19465 4295 19499
rect 4721 19465 4755 19499
rect 13185 19465 13219 19499
rect 13829 19465 13863 19499
rect 14289 19465 14323 19499
rect 15485 19465 15519 19499
rect 17141 19465 17175 19499
rect 17785 19465 17819 19499
rect 18061 19465 18095 19499
rect 18521 19465 18555 19499
rect 19441 19465 19475 19499
rect 2513 19397 2547 19431
rect 1593 19261 1627 19295
rect 2145 19261 2179 19295
rect 1777 19193 1811 19227
rect 2329 19193 2363 19227
rect 4077 19261 4111 19295
rect 12725 19397 12759 19431
rect 16037 19397 16071 19431
rect 5834 19261 5868 19295
rect 6101 19261 6135 19295
rect 6653 19261 6687 19295
rect 8605 19261 8639 19295
rect 8861 19261 8895 19295
rect 9689 19261 9723 19295
rect 9956 19261 9990 19295
rect 11713 19261 11747 19295
rect 12081 19261 12115 19295
rect 12541 19261 12575 19295
rect 13001 19261 13035 19295
rect 14013 19261 14047 19295
rect 14473 19261 14507 19295
rect 14749 19261 14783 19295
rect 15301 19261 15335 19295
rect 15853 19261 15887 19295
rect 16497 19261 16531 19295
rect 17325 19261 17359 19295
rect 17601 19261 17635 19295
rect 18245 19261 18279 19295
rect 18705 19261 18739 19295
rect 18981 19261 19015 19295
rect 21373 19261 21407 19295
rect 3832 19193 3866 19227
rect 4261 19193 4295 19227
rect 7113 19193 7147 19227
rect 13461 19193 13495 19227
rect 20545 19193 20579 19227
rect 2513 19125 2547 19159
rect 2697 19125 2731 19159
rect 4353 19125 4387 19159
rect 7481 19125 7515 19159
rect 9413 19125 9447 19159
rect 11069 19125 11103 19159
rect 12265 19125 12299 19159
rect 14933 19125 14967 19159
rect 16313 19125 16347 19159
rect 19165 19125 19199 19159
rect 19901 19125 19935 19159
rect 2237 18921 2271 18955
rect 4077 18921 4111 18955
rect 6377 18921 6411 18955
rect 6837 18921 6871 18955
rect 7757 18921 7791 18955
rect 9321 18921 9355 18955
rect 12541 18921 12575 18955
rect 13185 18921 13219 18955
rect 14013 18921 14047 18955
rect 15025 18921 15059 18955
rect 17877 18921 17911 18955
rect 18337 18921 18371 18955
rect 21373 18921 21407 18955
rect 2329 18853 2363 18887
rect 7113 18853 7147 18887
rect 11437 18853 11471 18887
rect 13461 18853 13495 18887
rect 17150 18853 17184 18887
rect 1593 18785 1627 18819
rect 1777 18785 1811 18819
rect 2881 18785 2915 18819
rect 3341 18785 3375 18819
rect 4261 18785 4295 18819
rect 4721 18785 4755 18819
rect 4997 18785 5031 18819
rect 5264 18785 5298 18819
rect 6653 18785 6687 18819
rect 7849 18785 7883 18819
rect 8493 18785 8527 18819
rect 10445 18785 10479 18819
rect 11161 18785 11195 18819
rect 12173 18785 12207 18819
rect 13001 18785 13035 18819
rect 13829 18785 13863 18819
rect 15117 18785 15151 18819
rect 17417 18785 17451 18819
rect 17693 18785 17727 18819
rect 18153 18785 18187 18819
rect 18797 18785 18831 18819
rect 7573 18717 7607 18751
rect 10701 18717 10735 18751
rect 11989 18717 12023 18751
rect 12081 18717 12115 18751
rect 14381 18717 14415 18751
rect 14933 18717 14967 18751
rect 4537 18649 4571 18683
rect 18613 18649 18647 18683
rect 2697 18581 2731 18615
rect 3157 18581 3191 18615
rect 8217 18581 8251 18615
rect 10977 18581 11011 18615
rect 15485 18581 15519 18615
rect 16037 18581 16071 18615
rect 19165 18581 19199 18615
rect 1685 18377 1719 18411
rect 2237 18377 2271 18411
rect 8309 18377 8343 18411
rect 8861 18377 8895 18411
rect 12909 18377 12943 18411
rect 15761 18377 15795 18411
rect 17325 18377 17359 18411
rect 17969 18377 18003 18411
rect 7849 18309 7883 18343
rect 14105 18309 14139 18343
rect 15669 18309 15703 18343
rect 18705 18309 18739 18343
rect 5365 18241 5399 18275
rect 6469 18241 6503 18275
rect 7389 18241 7423 18275
rect 9781 18241 9815 18275
rect 9965 18241 9999 18275
rect 12081 18241 12115 18275
rect 13461 18241 13495 18275
rect 2329 18173 2363 18207
rect 2881 18173 2915 18207
rect 3148 18173 3182 18207
rect 8033 18173 8067 18207
rect 8493 18173 8527 18207
rect 9045 18173 9079 18207
rect 9689 18173 9723 18207
rect 10517 18173 10551 18207
rect 10977 18173 11011 18207
rect 15229 18173 15263 18207
rect 15485 18173 15519 18207
rect 1777 18105 1811 18139
rect 5181 18105 5215 18139
rect 5825 18105 5859 18139
rect 11253 18105 11287 18139
rect 12173 18105 12207 18139
rect 16313 18241 16347 18275
rect 16129 18173 16163 18207
rect 17141 18173 17175 18207
rect 17785 18173 17819 18207
rect 18245 18173 18279 18207
rect 4261 18037 4295 18071
rect 4813 18037 4847 18071
rect 5273 18037 5307 18071
rect 6837 18037 6871 18071
rect 7205 18037 7239 18071
rect 7297 18037 7331 18071
rect 9321 18037 9355 18071
rect 10333 18037 10367 18071
rect 10793 18037 10827 18071
rect 12265 18037 12299 18071
rect 12633 18037 12667 18071
rect 13277 18037 13311 18071
rect 13369 18037 13403 18071
rect 15669 18037 15703 18071
rect 16221 18037 16255 18071
rect 18429 18037 18463 18071
rect 4077 17833 4111 17867
rect 4813 17833 4847 17867
rect 9597 17833 9631 17867
rect 13829 17833 13863 17867
rect 15117 17833 15151 17867
rect 15577 17833 15611 17867
rect 16313 17833 16347 17867
rect 16865 17833 16899 17867
rect 1777 17765 1811 17799
rect 2329 17765 2363 17799
rect 3617 17765 3651 17799
rect 5948 17765 5982 17799
rect 7472 17765 7506 17799
rect 17969 17765 18003 17799
rect 19073 17765 19107 17799
rect 1593 17697 1627 17731
rect 3157 17697 3191 17731
rect 2881 17629 2915 17663
rect 3065 17629 3099 17663
rect 4261 17697 4295 17731
rect 6285 17697 6319 17731
rect 6653 17697 6687 17731
rect 7113 17697 7147 17731
rect 9689 17697 9723 17731
rect 10517 17697 10551 17731
rect 10977 17697 11011 17731
rect 11437 17697 11471 17731
rect 12826 17697 12860 17731
rect 13553 17697 13587 17731
rect 14013 17697 14047 17731
rect 15209 17697 15243 17731
rect 16221 17697 16255 17731
rect 17877 17697 17911 17731
rect 6193 17629 6227 17663
rect 6285 17561 6319 17595
rect 6469 17561 6503 17595
rect 2237 17493 2271 17527
rect 3525 17493 3559 17527
rect 3617 17493 3651 17527
rect 7205 17629 7239 17663
rect 9505 17629 9539 17663
rect 13093 17629 13127 17663
rect 15025 17629 15059 17663
rect 16405 17629 16439 17663
rect 17785 17629 17819 17663
rect 18797 17629 18831 17663
rect 11253 17561 11287 17595
rect 15853 17561 15887 17595
rect 7113 17493 7147 17527
rect 8585 17493 8619 17527
rect 10057 17493 10091 17527
rect 10333 17493 10367 17527
rect 10793 17493 10827 17527
rect 11713 17493 11747 17527
rect 13369 17493 13403 17527
rect 14381 17493 14415 17527
rect 18337 17493 18371 17527
rect 2237 17289 2271 17323
rect 4353 17289 4387 17323
rect 5365 17289 5399 17323
rect 6469 17289 6503 17323
rect 7021 17289 7055 17323
rect 10609 17289 10643 17323
rect 11713 17289 11747 17323
rect 13553 17289 13587 17323
rect 14197 17289 14231 17323
rect 16221 17289 16255 17323
rect 19533 17289 19567 17323
rect 10885 17221 10919 17255
rect 13829 17221 13863 17255
rect 19257 17221 19291 17255
rect 4905 17153 4939 17187
rect 5917 17153 5951 17187
rect 12909 17153 12943 17187
rect 13093 17153 13127 17187
rect 19993 17153 20027 17187
rect 20085 17153 20119 17187
rect 2329 17085 2363 17119
rect 4077 17085 4111 17119
rect 5825 17085 5859 17119
rect 8134 17085 8168 17119
rect 8401 17085 8435 17119
rect 9229 17085 9263 17119
rect 11069 17085 11103 17119
rect 14841 17085 14875 17119
rect 16497 17085 16531 17119
rect 17877 17085 17911 17119
rect 19901 17085 19935 17119
rect 1593 17017 1627 17051
rect 1777 17017 1811 17051
rect 3832 17017 3866 17051
rect 4813 17017 4847 17051
rect 9496 17017 9530 17051
rect 15108 17017 15142 17051
rect 18144 17017 18178 17051
rect 2697 16949 2731 16983
rect 4721 16949 4755 16983
rect 5733 16949 5767 16983
rect 8953 16949 8987 16983
rect 12357 16949 12391 16983
rect 13185 16949 13219 16983
rect 17325 16949 17359 16983
rect 2145 16745 2179 16779
rect 2605 16745 2639 16779
rect 3157 16745 3191 16779
rect 4261 16745 4295 16779
rect 5733 16745 5767 16779
rect 6653 16745 6687 16779
rect 7205 16745 7239 16779
rect 7481 16745 7515 16779
rect 8493 16745 8527 16779
rect 9321 16745 9355 16779
rect 9689 16745 9723 16779
rect 9781 16745 9815 16779
rect 13645 16745 13679 16779
rect 13921 16745 13955 16779
rect 15761 16745 15795 16779
rect 17509 16745 17543 16779
rect 19165 16745 19199 16779
rect 5089 16677 5123 16711
rect 11060 16677 11094 16711
rect 14381 16677 14415 16711
rect 18030 16677 18064 16711
rect 1593 16609 1627 16643
rect 1777 16609 1811 16643
rect 2329 16609 2363 16643
rect 2789 16609 2823 16643
rect 4077 16609 4111 16643
rect 5181 16609 5215 16643
rect 5925 16609 5959 16643
rect 6377 16609 6411 16643
rect 7849 16609 7883 16643
rect 7941 16609 7975 16643
rect 8677 16609 8711 16643
rect 10517 16609 10551 16643
rect 10793 16609 10827 16643
rect 12633 16609 12667 16643
rect 13185 16609 13219 16643
rect 13277 16609 13311 16643
rect 15393 16609 15427 16643
rect 16385 16609 16419 16643
rect 19993 16609 20027 16643
rect 5273 16541 5307 16575
rect 8125 16541 8159 16575
rect 9965 16541 9999 16575
rect 13001 16541 13035 16575
rect 15209 16541 15243 16575
rect 15301 16541 15335 16575
rect 16129 16541 16163 16575
rect 17785 16541 17819 16575
rect 12173 16473 12207 16507
rect 4721 16405 4755 16439
rect 6193 16405 6227 16439
rect 10333 16405 10367 16439
rect 12449 16405 12483 16439
rect 19625 16405 19659 16439
rect 2145 16201 2179 16235
rect 2605 16201 2639 16235
rect 3065 16201 3099 16235
rect 3525 16201 3559 16235
rect 6009 16201 6043 16235
rect 7113 16201 7147 16235
rect 10057 16201 10091 16235
rect 11897 16201 11931 16235
rect 15209 16201 15243 16235
rect 17877 16201 17911 16235
rect 19901 16201 19935 16235
rect 3985 16133 4019 16167
rect 6653 16133 6687 16167
rect 13369 16133 13403 16167
rect 1593 16065 1627 16099
rect 8309 16065 8343 16099
rect 11161 16065 11195 16099
rect 12541 16065 12575 16099
rect 15945 16065 15979 16099
rect 17233 16065 17267 16099
rect 2329 15997 2363 16031
rect 2789 15997 2823 16031
rect 3249 15997 3283 16031
rect 3709 15997 3743 16031
rect 3801 15997 3835 16031
rect 4169 15997 4203 16031
rect 4629 15997 4663 16031
rect 4896 15997 4930 16031
rect 6837 15997 6871 16031
rect 7297 15997 7331 16031
rect 8677 15997 8711 16031
rect 8933 15997 8967 16031
rect 12265 15997 12299 16031
rect 13093 15997 13127 16031
rect 13829 15997 13863 16031
rect 17509 15997 17543 16031
rect 19358 15997 19392 16031
rect 19625 15997 19659 16031
rect 1777 15929 1811 15963
rect 8033 15929 8067 15963
rect 10977 15929 11011 15963
rect 14096 15929 14130 15963
rect 16129 15929 16163 15963
rect 3801 15861 3835 15895
rect 7665 15861 7699 15895
rect 8125 15861 8159 15895
rect 10609 15861 10643 15895
rect 11069 15861 11103 15895
rect 12357 15861 12391 15895
rect 12909 15861 12943 15895
rect 16037 15861 16071 15895
rect 16497 15861 16531 15895
rect 17417 15861 17451 15895
rect 18245 15861 18279 15895
rect 2145 15657 2179 15691
rect 4077 15657 4111 15691
rect 4537 15657 4571 15691
rect 6193 15657 6227 15691
rect 9321 15657 9355 15691
rect 9781 15657 9815 15691
rect 12357 15657 12391 15691
rect 17141 15657 17175 15691
rect 6920 15589 6954 15623
rect 11998 15589 12032 15623
rect 1593 15521 1627 15555
rect 1777 15521 1811 15555
rect 2329 15521 2363 15555
rect 2605 15521 2639 15555
rect 3249 15521 3283 15555
rect 4261 15521 4295 15555
rect 5661 15521 5695 15555
rect 8493 15521 8527 15555
rect 9689 15521 9723 15555
rect 10333 15521 10367 15555
rect 12265 15521 12299 15555
rect 13645 15589 13679 15623
rect 18061 15589 18095 15623
rect 19165 15589 19199 15623
rect 12909 15521 12943 15555
rect 13737 15521 13771 15555
rect 15301 15521 15335 15555
rect 15761 15521 15795 15555
rect 16028 15521 16062 15555
rect 5917 15453 5951 15487
rect 6653 15453 6687 15487
rect 9873 15453 9907 15487
rect 12357 15453 12391 15487
rect 13829 15453 13863 15487
rect 17877 15453 17911 15487
rect 17969 15453 18003 15487
rect 18705 15453 18739 15487
rect 3065 15385 3099 15419
rect 12541 15385 12575 15419
rect 14933 15385 14967 15419
rect 2789 15317 2823 15351
rect 8033 15317 8067 15351
rect 8309 15317 8343 15351
rect 10517 15317 10551 15351
rect 10885 15317 10919 15351
rect 13277 15317 13311 15351
rect 14381 15317 14415 15351
rect 15485 15317 15519 15351
rect 18429 15317 18463 15351
rect 1685 15113 1719 15147
rect 2145 15113 2179 15147
rect 5365 15113 5399 15147
rect 8125 15113 8159 15147
rect 8309 15113 8343 15147
rect 12817 15113 12851 15147
rect 13093 15113 13127 15147
rect 14749 15113 14783 15147
rect 16589 15113 16623 15147
rect 3985 15045 4019 15079
rect 4813 14977 4847 15011
rect 5917 14977 5951 15011
rect 6837 14977 6871 15011
rect 8033 14977 8067 15011
rect 2329 14909 2363 14943
rect 2605 14909 2639 14943
rect 2872 14909 2906 14943
rect 4721 14909 4755 14943
rect 5825 14909 5859 14943
rect 1777 14841 1811 14875
rect 4629 14841 4663 14875
rect 6929 14841 6963 14875
rect 11713 15045 11747 15079
rect 12265 14977 12299 15011
rect 12357 14977 12391 15011
rect 15301 14977 15335 15011
rect 15945 14977 15979 15011
rect 17969 14977 18003 15011
rect 9689 14909 9723 14943
rect 11345 14909 11379 14943
rect 12449 14909 12483 14943
rect 14206 14909 14240 14943
rect 14473 14909 14507 14943
rect 18225 14909 18259 14943
rect 9444 14841 9478 14875
rect 11078 14841 11112 14875
rect 4261 14773 4295 14807
rect 5733 14773 5767 14807
rect 7021 14773 7055 14807
rect 7389 14773 7423 14807
rect 8125 14773 8159 14807
rect 9965 14773 9999 14807
rect 15117 14773 15151 14807
rect 15209 14773 15243 14807
rect 16129 14773 16163 14807
rect 16221 14773 16255 14807
rect 16957 14773 16991 14807
rect 17509 14773 17543 14807
rect 19349 14773 19383 14807
rect 2237 14569 2271 14603
rect 3249 14569 3283 14603
rect 5457 14569 5491 14603
rect 8217 14569 8251 14603
rect 9137 14569 9171 14603
rect 9873 14569 9907 14603
rect 12265 14569 12299 14603
rect 12725 14569 12759 14603
rect 13645 14569 13679 14603
rect 14013 14569 14047 14603
rect 14749 14569 14783 14603
rect 15117 14569 15151 14603
rect 15393 14569 15427 14603
rect 17969 14569 18003 14603
rect 18061 14569 18095 14603
rect 18429 14569 18463 14603
rect 4344 14501 4378 14535
rect 6101 14501 6135 14535
rect 13553 14501 13587 14535
rect 17049 14501 17083 14535
rect 1777 14433 1811 14467
rect 2329 14433 2363 14467
rect 3157 14433 3191 14467
rect 6377 14433 6411 14467
rect 6644 14433 6678 14467
rect 8033 14433 8067 14467
rect 8493 14433 8527 14467
rect 9965 14433 9999 14467
rect 10609 14433 10643 14467
rect 10876 14433 10910 14467
rect 12633 14433 12667 14467
rect 14473 14433 14507 14467
rect 14565 14433 14599 14467
rect 16506 14433 16540 14467
rect 16773 14433 16807 14467
rect 3433 14365 3467 14399
rect 4077 14365 4111 14399
rect 9781 14365 9815 14399
rect 12817 14365 12851 14399
rect 13461 14365 13495 14399
rect 17877 14365 17911 14399
rect 8677 14297 8711 14331
rect 10333 14297 10367 14331
rect 14473 14297 14507 14331
rect 1685 14229 1719 14263
rect 2789 14229 2823 14263
rect 7757 14229 7791 14263
rect 11989 14229 12023 14263
rect 2145 14025 2179 14059
rect 2605 14025 2639 14059
rect 3801 14025 3835 14059
rect 4721 14025 4755 14059
rect 6653 14025 6687 14059
rect 7665 14025 7699 14059
rect 9781 14025 9815 14059
rect 13921 14025 13955 14059
rect 16313 14025 16347 14059
rect 4261 13957 4295 13991
rect 8125 13957 8159 13991
rect 17417 13957 17451 13991
rect 3157 13889 3191 13923
rect 7297 13889 7331 13923
rect 15301 13889 15335 13923
rect 15669 13889 15703 13923
rect 15853 13889 15887 13923
rect 1593 13821 1627 13855
rect 1777 13821 1811 13855
rect 2329 13821 2363 13855
rect 2789 13821 2823 13855
rect 3617 13821 3651 13855
rect 4077 13821 4111 13855
rect 6101 13821 6135 13855
rect 9505 13821 9539 13855
rect 10894 13821 10928 13855
rect 11161 13821 11195 13855
rect 13645 13821 13679 13855
rect 15034 13821 15068 13855
rect 18909 13821 18943 13855
rect 19165 13821 19199 13855
rect 5834 13753 5868 13787
rect 7021 13753 7055 13787
rect 7113 13753 7147 13787
rect 9249 13753 9283 13787
rect 15945 13753 15979 13787
rect 12357 13685 12391 13719
rect 17785 13685 17819 13719
rect 2237 13481 2271 13515
rect 2513 13481 2547 13515
rect 4353 13481 4387 13515
rect 4813 13481 4847 13515
rect 5365 13481 5399 13515
rect 5825 13481 5859 13515
rect 8493 13481 8527 13515
rect 9321 13481 9355 13515
rect 10885 13481 10919 13515
rect 11897 13481 11931 13515
rect 12357 13481 12391 13515
rect 13185 13481 13219 13515
rect 15485 13481 15519 13515
rect 16129 13481 16163 13515
rect 16589 13481 16623 13515
rect 3433 13413 3467 13447
rect 4721 13413 4755 13447
rect 6377 13413 6411 13447
rect 9689 13413 9723 13447
rect 9781 13413 9815 13447
rect 11253 13413 11287 13447
rect 15025 13413 15059 13447
rect 17325 13413 17359 13447
rect 17877 13413 17911 13447
rect 1593 13345 1627 13379
rect 2053 13345 2087 13379
rect 2697 13345 2731 13379
rect 2973 13345 3007 13379
rect 3893 13345 3927 13379
rect 5733 13345 5767 13379
rect 7021 13345 7055 13379
rect 7757 13345 7791 13379
rect 8401 13345 8435 13379
rect 12265 13345 12299 13379
rect 13553 13345 13587 13379
rect 14565 13345 14599 13379
rect 17969 13345 18003 13379
rect 4997 13277 5031 13311
rect 5917 13277 5951 13311
rect 8677 13277 8711 13311
rect 9873 13277 9907 13311
rect 11345 13277 11379 13311
rect 11437 13277 11471 13311
rect 12449 13277 12483 13311
rect 13645 13277 13679 13311
rect 13737 13277 13771 13311
rect 17785 13277 17819 13311
rect 1777 13209 1811 13243
rect 3157 13209 3191 13243
rect 6837 13209 6871 13243
rect 10333 13209 10367 13243
rect 8033 13141 8067 13175
rect 18337 13141 18371 13175
rect 1501 12937 1535 12971
rect 1777 12937 1811 12971
rect 2237 12937 2271 12971
rect 6745 12937 6779 12971
rect 9137 12937 9171 12971
rect 13553 12937 13587 12971
rect 15025 12937 15059 12971
rect 18613 12937 18647 12971
rect 9873 12869 9907 12903
rect 10609 12869 10643 12903
rect 10977 12869 11011 12903
rect 6009 12801 6043 12835
rect 7297 12801 7331 12835
rect 13277 12801 13311 12835
rect 14013 12801 14047 12835
rect 14197 12801 14231 12835
rect 16405 12801 16439 12835
rect 17785 12801 17819 12835
rect 17877 12801 17911 12835
rect 19165 12801 19199 12835
rect 1961 12733 1995 12767
rect 2421 12733 2455 12767
rect 4353 12733 4387 12767
rect 5753 12733 5787 12767
rect 7757 12733 7791 12767
rect 8013 12733 8047 12767
rect 9597 12733 9631 12767
rect 13010 12733 13044 12767
rect 14749 12733 14783 12767
rect 17141 12733 17175 12767
rect 17969 12733 18003 12767
rect 18981 12733 19015 12767
rect 4108 12665 4142 12699
rect 7113 12665 7147 12699
rect 13921 12665 13955 12699
rect 16138 12665 16172 12699
rect 19073 12665 19107 12699
rect 2973 12597 3007 12631
rect 4629 12597 4663 12631
rect 7205 12597 7239 12631
rect 9413 12597 9447 12631
rect 11253 12597 11287 12631
rect 11897 12597 11931 12631
rect 14565 12597 14599 12631
rect 17325 12597 17359 12631
rect 18337 12597 18371 12631
rect 1777 12393 1811 12427
rect 2421 12393 2455 12427
rect 2697 12393 2731 12427
rect 3341 12393 3375 12427
rect 5457 12393 5491 12427
rect 7573 12393 7607 12427
rect 9229 12393 9263 12427
rect 10517 12393 10551 12427
rect 12633 12393 12667 12427
rect 16221 12393 16255 12427
rect 18981 12393 19015 12427
rect 7030 12325 7064 12359
rect 10057 12325 10091 12359
rect 13001 12325 13035 12359
rect 17592 12325 17626 12359
rect 1961 12257 1995 12291
rect 2237 12257 2271 12291
rect 2881 12257 2915 12291
rect 3157 12257 3191 12291
rect 4333 12257 4367 12291
rect 7297 12257 7331 12291
rect 7941 12257 7975 12291
rect 8769 12257 8803 12291
rect 10149 12257 10183 12291
rect 10793 12257 10827 12291
rect 11345 12257 11379 12291
rect 11897 12257 11931 12291
rect 11989 12257 12023 12291
rect 13829 12257 13863 12291
rect 14832 12257 14866 12291
rect 16589 12257 16623 12291
rect 17325 12257 17359 12291
rect 21106 12257 21140 12291
rect 21373 12257 21407 12291
rect 1501 12189 1535 12223
rect 4077 12189 4111 12223
rect 8033 12189 8067 12223
rect 8217 12189 8251 12223
rect 9965 12189 9999 12223
rect 11805 12189 11839 12223
rect 13093 12189 13127 12223
rect 13185 12189 13219 12223
rect 14565 12189 14599 12223
rect 16681 12189 16715 12223
rect 16773 12189 16807 12223
rect 12357 12121 12391 12155
rect 15945 12121 15979 12155
rect 18705 12121 18739 12155
rect 5917 12053 5951 12087
rect 8585 12053 8619 12087
rect 13645 12053 13679 12087
rect 19993 12053 20027 12087
rect 1777 11849 1811 11883
rect 2237 11849 2271 11883
rect 3341 11849 3375 11883
rect 5365 11849 5399 11883
rect 5917 11849 5951 11883
rect 7941 11849 7975 11883
rect 11069 11849 11103 11883
rect 12817 11849 12851 11883
rect 14841 11849 14875 11883
rect 15853 11849 15887 11883
rect 21189 11849 21223 11883
rect 4169 11781 4203 11815
rect 6653 11781 6687 11815
rect 17693 11781 17727 11815
rect 3893 11713 3927 11747
rect 1961 11645 1995 11679
rect 2421 11645 2455 11679
rect 2697 11645 2731 11679
rect 3709 11577 3743 11611
rect 4905 11713 4939 11747
rect 7113 11713 7147 11747
rect 7297 11713 7331 11747
rect 8493 11713 8527 11747
rect 12173 11713 12207 11747
rect 13277 11713 13311 11747
rect 14289 11713 14323 11747
rect 15301 11713 15335 11747
rect 16313 11713 16347 11747
rect 19073 11713 19107 11747
rect 6101 11645 6135 11679
rect 8401 11645 8435 11679
rect 9689 11645 9723 11679
rect 9956 11645 9990 11679
rect 13461 11645 13495 11679
rect 15393 11645 15427 11679
rect 16957 11645 16991 11679
rect 18806 11645 18840 11679
rect 20913 11645 20947 11679
rect 21373 11645 21407 11679
rect 7021 11577 7055 11611
rect 8309 11577 8343 11611
rect 12357 11577 12391 11611
rect 12449 11577 12483 11611
rect 15485 11577 15519 11611
rect 1409 11509 1443 11543
rect 2881 11509 2915 11543
rect 3801 11509 3835 11543
rect 4169 11509 4203 11543
rect 4353 11509 4387 11543
rect 4721 11509 4755 11543
rect 4813 11509 4847 11543
rect 11805 11509 11839 11543
rect 13369 11509 13403 11543
rect 13829 11509 13863 11543
rect 14381 11509 14415 11543
rect 14473 11509 14507 11543
rect 1593 11305 1627 11339
rect 1869 11305 1903 11339
rect 3433 11305 3467 11339
rect 4445 11305 4479 11339
rect 5089 11305 5123 11339
rect 7113 11305 7147 11339
rect 7205 11305 7239 11339
rect 9321 11305 9355 11339
rect 13553 11305 13587 11339
rect 14013 11305 14047 11339
rect 15945 11305 15979 11339
rect 6285 11237 6319 11271
rect 1409 11169 1443 11203
rect 2053 11169 2087 11203
rect 2789 11169 2823 11203
rect 6193 11169 6227 11203
rect 2881 11101 2915 11135
rect 3065 11101 3099 11135
rect 4169 11101 4203 11135
rect 4353 11101 4387 11135
rect 6469 11101 6503 11135
rect 6929 11101 6963 11135
rect 10508 11237 10542 11271
rect 14810 11237 14844 11271
rect 16488 11237 16522 11271
rect 8318 11169 8352 11203
rect 12173 11169 12207 11203
rect 12440 11169 12474 11203
rect 14565 11169 14599 11203
rect 16221 11169 16255 11203
rect 8585 11101 8619 11135
rect 10241 11101 10275 11135
rect 5825 11033 5859 11067
rect 7113 11033 7147 11067
rect 2421 10965 2455 10999
rect 4813 10965 4847 10999
rect 11621 10965 11655 10999
rect 17601 10965 17635 10999
rect 2513 10761 2547 10795
rect 2789 10761 2823 10795
rect 8033 10761 8067 10795
rect 9781 10761 9815 10795
rect 11345 10761 11379 10795
rect 13277 10761 13311 10795
rect 14933 10761 14967 10795
rect 17141 10693 17175 10727
rect 1961 10625 1995 10659
rect 4169 10625 4203 10659
rect 4905 10625 4939 10659
rect 4997 10625 5031 10659
rect 6653 10625 6687 10659
rect 9045 10625 9079 10659
rect 9229 10625 9263 10659
rect 15577 10625 15611 10659
rect 18521 10625 18555 10659
rect 2145 10557 2179 10591
rect 6909 10557 6943 10591
rect 9597 10557 9631 10591
rect 11897 10557 11931 10591
rect 13553 10557 13587 10591
rect 13820 10557 13854 10591
rect 2053 10489 2087 10523
rect 3924 10489 3958 10523
rect 12142 10489 12176 10523
rect 15669 10489 15703 10523
rect 18254 10489 18288 10523
rect 1409 10421 1443 10455
rect 4445 10421 4479 10455
rect 4813 10421 4847 10455
rect 5457 10421 5491 10455
rect 5825 10421 5859 10455
rect 8585 10421 8619 10455
rect 8953 10421 8987 10455
rect 15761 10421 15795 10455
rect 16129 10421 16163 10455
rect 16589 10421 16623 10455
rect 1593 10217 1627 10251
rect 4813 10217 4847 10251
rect 6653 10217 6687 10251
rect 7757 10217 7791 10251
rect 8217 10217 8251 10251
rect 11529 10217 11563 10251
rect 11897 10217 11931 10251
rect 12449 10217 12483 10251
rect 15209 10217 15243 10251
rect 16957 10217 16991 10251
rect 17325 10217 17359 10251
rect 16865 10149 16899 10183
rect 1409 10081 1443 10115
rect 2982 10081 3016 10115
rect 4445 10081 4479 10115
rect 5540 10081 5574 10115
rect 8125 10081 8159 10115
rect 10434 10081 10468 10115
rect 10701 10081 10735 10115
rect 11437 10081 11471 10115
rect 3249 10013 3283 10047
rect 4169 10013 4203 10047
rect 4353 10013 4387 10047
rect 5273 10013 5307 10047
rect 7113 10013 7147 10047
rect 8309 10013 8343 10047
rect 11253 10013 11287 10047
rect 16773 10013 16807 10047
rect 9321 9945 9355 9979
rect 1869 9877 1903 9911
rect 9321 9673 9355 9707
rect 11069 9673 11103 9707
rect 1593 9605 1627 9639
rect 2973 9605 3007 9639
rect 4721 9605 4755 9639
rect 6653 9605 6687 9639
rect 9597 9605 9631 9639
rect 2697 9537 2731 9571
rect 3617 9537 3651 9571
rect 7205 9537 7239 9571
rect 7941 9537 7975 9571
rect 10149 9537 10183 9571
rect 1409 9469 1443 9503
rect 1869 9469 1903 9503
rect 3341 9469 3375 9503
rect 4445 9469 4479 9503
rect 7021 9469 7055 9503
rect 10057 9469 10091 9503
rect 8186 9401 8220 9435
rect 2053 9333 2087 9367
rect 3433 9333 3467 9367
rect 3985 9333 4019 9367
rect 7113 9333 7147 9367
rect 9965 9333 9999 9367
rect 3157 9129 3191 9163
rect 5365 9129 5399 9163
rect 7113 9129 7147 9163
rect 9781 9129 9815 9163
rect 1409 9061 1443 9095
rect 1777 8993 1811 9027
rect 2421 8993 2455 9027
rect 2697 8993 2731 9027
rect 3893 8993 3927 9027
rect 5273 8993 5307 9027
rect 7481 8993 7515 9027
rect 7573 8993 7607 9027
rect 5457 8925 5491 8959
rect 7665 8925 7699 8959
rect 1961 8857 1995 8891
rect 2237 8857 2271 8891
rect 2881 8857 2915 8891
rect 4905 8789 4939 8823
rect 9413 8789 9447 8823
rect 1777 8585 1811 8619
rect 3709 8585 3743 8619
rect 9045 8517 9079 8551
rect 8401 8449 8435 8483
rect 8585 8449 8619 8483
rect 1961 8381 1995 8415
rect 2329 8381 2363 8415
rect 4077 8381 4111 8415
rect 6653 8381 6687 8415
rect 6920 8381 6954 8415
rect 2574 8313 2608 8347
rect 4322 8313 4356 8347
rect 8677 8313 8711 8347
rect 1409 8245 1443 8279
rect 5457 8245 5491 8279
rect 8033 8245 8067 8279
rect 1593 8041 1627 8075
rect 2053 8041 2087 8075
rect 2789 8041 2823 8075
rect 7389 8041 7423 8075
rect 9321 8041 9355 8075
rect 9781 8041 9815 8075
rect 3249 7973 3283 8007
rect 5190 7973 5224 8007
rect 5978 7973 6012 8007
rect 1409 7905 1443 7939
rect 2237 7905 2271 7939
rect 3157 7905 3191 7939
rect 5733 7905 5767 7939
rect 8502 7905 8536 7939
rect 8769 7905 8803 7939
rect 9689 7905 9723 7939
rect 3433 7837 3467 7871
rect 5457 7837 5491 7871
rect 9873 7837 9907 7871
rect 4077 7701 4111 7735
rect 7113 7701 7147 7735
rect 3617 7497 3651 7531
rect 6745 7497 6779 7531
rect 7021 7497 7055 7531
rect 8861 7497 8895 7531
rect 18613 7497 18647 7531
rect 19257 7497 19291 7531
rect 2053 7429 2087 7463
rect 4261 7361 4295 7395
rect 5181 7361 5215 7395
rect 1409 7293 1443 7327
rect 1869 7293 1903 7327
rect 2697 7293 2731 7327
rect 2329 7225 2363 7259
rect 3985 7225 4019 7259
rect 5641 7225 5675 7259
rect 7297 7361 7331 7395
rect 8309 7361 8343 7395
rect 7481 7293 7515 7327
rect 18797 7293 18831 7327
rect 19073 7293 19107 7327
rect 8401 7225 8435 7259
rect 9137 7225 9171 7259
rect 1593 7157 1627 7191
rect 3249 7157 3283 7191
rect 4077 7157 4111 7191
rect 4629 7157 4663 7191
rect 4997 7157 5031 7191
rect 5089 7157 5123 7191
rect 7021 7157 7055 7191
rect 7389 7157 7423 7191
rect 7849 7157 7883 7191
rect 8493 7157 8527 7191
rect 9505 7157 9539 7191
rect 4353 6953 4387 6987
rect 4721 6953 4755 6987
rect 7757 6953 7791 6987
rect 7665 6885 7699 6919
rect 1409 6817 1443 6851
rect 1869 6817 1903 6851
rect 4813 6817 4847 6851
rect 8309 6817 8343 6851
rect 19809 6817 19843 6851
rect 20269 6817 20303 6851
rect 4905 6749 4939 6783
rect 7941 6749 7975 6783
rect 1593 6681 1627 6715
rect 7297 6681 7331 6715
rect 19993 6681 20027 6715
rect 3985 6613 4019 6647
rect 20269 6409 20303 6443
rect 1409 6205 1443 6239
rect 1869 6205 1903 6239
rect 20085 6205 20119 6239
rect 20545 6205 20579 6239
rect 1593 6069 1627 6103
rect 20545 5865 20579 5899
rect 1409 5729 1443 5763
rect 1869 5729 1903 5763
rect 20729 5729 20763 5763
rect 21005 5661 21039 5695
rect 1593 5593 1627 5627
rect 1593 5321 1627 5355
rect 20821 5321 20855 5355
rect 1409 5117 1443 5151
rect 2237 5117 2271 5151
rect 21005 5117 21039 5151
rect 21281 5117 21315 5151
rect 1869 4981 1903 5015
rect 2329 4709 2363 4743
rect 1409 4641 1443 4675
rect 1869 4641 1903 4675
rect 1593 4505 1627 4539
rect 2053 4505 2087 4539
rect 1869 4097 1903 4131
rect 1685 3961 1719 3995
rect 2513 3961 2547 3995
rect 2145 3893 2179 3927
rect 1777 3689 1811 3723
rect 2421 3621 2455 3655
rect 1685 3553 1719 3587
rect 2237 3553 2271 3587
rect 2697 3485 2731 3519
rect 3157 3349 3191 3383
rect 1685 3145 1719 3179
rect 2421 3077 2455 3111
rect 2973 3077 3007 3111
rect 3249 3009 3283 3043
rect 1777 2941 1811 2975
rect 2789 2941 2823 2975
rect 2237 2873 2271 2907
rect 3985 2873 4019 2907
rect 3617 2805 3651 2839
rect 2329 2601 2363 2635
rect 2973 2533 3007 2567
rect 12265 2533 12299 2567
rect 12633 2533 12667 2567
rect 1685 2465 1719 2499
rect 2237 2465 2271 2499
rect 2789 2465 2823 2499
rect 3893 2465 3927 2499
rect 3249 2397 3283 2431
rect 1869 2329 1903 2363
rect 12081 2329 12115 2363
<< metal1 >>
rect 3970 20816 3976 20868
rect 4028 20856 4034 20868
rect 7834 20856 7840 20868
rect 4028 20828 7840 20856
rect 4028 20816 4034 20828
rect 7834 20816 7840 20828
rect 7892 20816 7898 20868
rect 9398 20816 9404 20868
rect 9456 20856 9462 20868
rect 10134 20856 10140 20868
rect 9456 20828 10140 20856
rect 9456 20816 9462 20828
rect 10134 20816 10140 20828
rect 10192 20816 10198 20868
rect 4062 20748 4068 20800
rect 4120 20788 4126 20800
rect 7282 20788 7288 20800
rect 4120 20760 7288 20788
rect 4120 20748 4126 20760
rect 7282 20748 7288 20760
rect 7340 20748 7346 20800
rect 8938 20748 8944 20800
rect 8996 20788 9002 20800
rect 10042 20788 10048 20800
rect 8996 20760 10048 20788
rect 8996 20748 9002 20760
rect 10042 20748 10048 20760
rect 10100 20748 10106 20800
rect 1104 20698 21896 20720
rect 1104 20646 4447 20698
rect 4499 20646 4511 20698
rect 4563 20646 4575 20698
rect 4627 20646 4639 20698
rect 4691 20646 11378 20698
rect 11430 20646 11442 20698
rect 11494 20646 11506 20698
rect 11558 20646 11570 20698
rect 11622 20646 18308 20698
rect 18360 20646 18372 20698
rect 18424 20646 18436 20698
rect 18488 20646 18500 20698
rect 18552 20646 21896 20698
rect 1104 20624 21896 20646
rect 3145 20587 3203 20593
rect 3145 20553 3157 20587
rect 3191 20584 3203 20587
rect 7558 20584 7564 20596
rect 3191 20556 7564 20584
rect 3191 20553 3203 20556
rect 3145 20547 3203 20553
rect 7558 20544 7564 20556
rect 7616 20544 7622 20596
rect 7650 20544 7656 20596
rect 7708 20584 7714 20596
rect 7708 20556 8432 20584
rect 7708 20544 7714 20556
rect 2409 20519 2467 20525
rect 2409 20485 2421 20519
rect 2455 20516 2467 20519
rect 2774 20516 2780 20528
rect 2455 20488 2780 20516
rect 2455 20485 2467 20488
rect 2409 20479 2467 20485
rect 2774 20476 2780 20488
rect 2832 20476 2838 20528
rect 2961 20519 3019 20525
rect 2961 20485 2973 20519
rect 3007 20516 3019 20519
rect 7098 20516 7104 20528
rect 3007 20488 7104 20516
rect 3007 20485 3019 20488
rect 2961 20479 3019 20485
rect 7098 20476 7104 20488
rect 7156 20476 7162 20528
rect 7282 20516 7288 20528
rect 7243 20488 7288 20516
rect 7282 20476 7288 20488
rect 7340 20476 7346 20528
rect 7834 20516 7840 20528
rect 7795 20488 7840 20516
rect 7834 20476 7840 20488
rect 7892 20476 7898 20528
rect 8404 20516 8432 20556
rect 8478 20544 8484 20596
rect 8536 20584 8542 20596
rect 10873 20587 10931 20593
rect 10873 20584 10885 20587
rect 8536 20556 10885 20584
rect 8536 20544 8542 20556
rect 10873 20553 10885 20556
rect 10919 20553 10931 20587
rect 10873 20547 10931 20553
rect 12713 20587 12771 20593
rect 12713 20553 12725 20587
rect 12759 20584 12771 20587
rect 14458 20584 14464 20596
rect 12759 20556 14464 20584
rect 12759 20553 12771 20556
rect 12713 20547 12771 20553
rect 14458 20544 14464 20556
rect 14516 20544 14522 20596
rect 16761 20587 16819 20593
rect 16761 20553 16773 20587
rect 16807 20584 16819 20587
rect 19518 20584 19524 20596
rect 16807 20556 19524 20584
rect 16807 20553 16819 20556
rect 16761 20547 16819 20553
rect 19518 20544 19524 20556
rect 19576 20544 19582 20596
rect 11330 20516 11336 20528
rect 8404 20488 9812 20516
rect 1578 20408 1584 20460
rect 1636 20448 1642 20460
rect 3513 20451 3571 20457
rect 1636 20420 3372 20448
rect 1636 20408 1642 20420
rect 198 20340 204 20392
rect 256 20380 262 20392
rect 1302 20380 1308 20392
rect 256 20352 1308 20380
rect 256 20340 262 20352
rect 1302 20340 1308 20352
rect 1360 20380 1366 20392
rect 3344 20389 3372 20420
rect 3513 20417 3525 20451
rect 3559 20448 3571 20451
rect 4154 20448 4160 20460
rect 3559 20420 4160 20448
rect 3559 20417 3571 20420
rect 3513 20411 3571 20417
rect 4154 20408 4160 20420
rect 4212 20408 4218 20460
rect 4617 20451 4675 20457
rect 4617 20448 4629 20451
rect 4448 20420 4629 20448
rect 1673 20383 1731 20389
rect 1673 20380 1685 20383
rect 1360 20352 1685 20380
rect 1360 20340 1366 20352
rect 1673 20349 1685 20352
rect 1719 20349 1731 20383
rect 1673 20343 1731 20349
rect 1857 20383 1915 20389
rect 1857 20349 1869 20383
rect 1903 20380 1915 20383
rect 3145 20383 3203 20389
rect 3145 20380 3157 20383
rect 1903 20352 3157 20380
rect 1903 20349 1915 20352
rect 1857 20343 1915 20349
rect 3145 20349 3157 20352
rect 3191 20349 3203 20383
rect 3145 20343 3203 20349
rect 3329 20383 3387 20389
rect 3329 20349 3341 20383
rect 3375 20380 3387 20383
rect 3602 20380 3608 20392
rect 3375 20352 3608 20380
rect 3375 20349 3387 20352
rect 3329 20343 3387 20349
rect 3602 20340 3608 20352
rect 3660 20340 3666 20392
rect 4246 20340 4252 20392
rect 4304 20380 4310 20392
rect 4448 20380 4476 20420
rect 4617 20417 4629 20420
rect 4663 20417 4675 20451
rect 6086 20448 6092 20460
rect 6047 20420 6092 20448
rect 4617 20411 4675 20417
rect 6086 20408 6092 20420
rect 6144 20408 6150 20460
rect 6546 20408 6552 20460
rect 6604 20448 6610 20460
rect 9674 20448 9680 20460
rect 6604 20420 9680 20448
rect 6604 20408 6610 20420
rect 9674 20408 9680 20420
rect 9732 20408 9738 20460
rect 4304 20352 4476 20380
rect 4525 20383 4583 20389
rect 4304 20340 4310 20352
rect 4525 20349 4537 20383
rect 4571 20380 4583 20383
rect 4982 20380 4988 20392
rect 4571 20352 4988 20380
rect 4571 20349 4583 20352
rect 4525 20343 4583 20349
rect 4982 20340 4988 20352
rect 5040 20340 5046 20392
rect 6730 20340 6736 20392
rect 6788 20380 6794 20392
rect 7469 20383 7527 20389
rect 7469 20380 7481 20383
rect 6788 20352 7481 20380
rect 6788 20340 6794 20352
rect 7469 20349 7481 20352
rect 7515 20349 7527 20383
rect 7469 20343 7527 20349
rect 7650 20340 7656 20392
rect 7708 20380 7714 20392
rect 8573 20383 8631 20389
rect 8573 20380 8585 20383
rect 7708 20352 8585 20380
rect 7708 20340 7714 20352
rect 8573 20349 8585 20352
rect 8619 20349 8631 20383
rect 8573 20343 8631 20349
rect 658 20272 664 20324
rect 716 20312 722 20324
rect 2222 20312 2228 20324
rect 716 20284 2228 20312
rect 716 20272 722 20284
rect 2222 20272 2228 20284
rect 2280 20272 2286 20324
rect 2777 20315 2835 20321
rect 2777 20281 2789 20315
rect 2823 20312 2835 20315
rect 2823 20284 2857 20312
rect 2823 20281 2835 20284
rect 2777 20275 2835 20281
rect 1118 20204 1124 20256
rect 1176 20244 1182 20256
rect 2792 20244 2820 20275
rect 3694 20272 3700 20324
rect 3752 20312 3758 20324
rect 6822 20312 6828 20324
rect 3752 20284 6828 20312
rect 3752 20272 3758 20284
rect 6822 20272 6828 20284
rect 6880 20272 6886 20324
rect 7006 20272 7012 20324
rect 7064 20312 7070 20324
rect 8021 20315 8079 20321
rect 8021 20312 8033 20315
rect 7064 20284 8033 20312
rect 7064 20272 7070 20284
rect 8021 20281 8033 20284
rect 8067 20281 8079 20315
rect 9306 20312 9312 20324
rect 8021 20275 8079 20281
rect 8312 20284 9312 20312
rect 3418 20244 3424 20256
rect 1176 20216 3424 20244
rect 1176 20204 1182 20216
rect 3418 20204 3424 20216
rect 3476 20204 3482 20256
rect 4062 20244 4068 20256
rect 4023 20216 4068 20244
rect 4062 20204 4068 20216
rect 4120 20204 4126 20256
rect 4433 20247 4491 20253
rect 4433 20213 4445 20247
rect 4479 20244 4491 20247
rect 4614 20244 4620 20256
rect 4479 20216 4620 20244
rect 4479 20213 4491 20216
rect 4433 20207 4491 20213
rect 4614 20204 4620 20216
rect 4672 20204 4678 20256
rect 5074 20244 5080 20256
rect 5035 20216 5080 20244
rect 5074 20204 5080 20216
rect 5132 20204 5138 20256
rect 5442 20244 5448 20256
rect 5403 20216 5448 20244
rect 5442 20204 5448 20216
rect 5500 20204 5506 20256
rect 5810 20244 5816 20256
rect 5771 20216 5816 20244
rect 5810 20204 5816 20216
rect 5868 20204 5874 20256
rect 5905 20247 5963 20253
rect 5905 20213 5917 20247
rect 5951 20244 5963 20247
rect 6546 20244 6552 20256
rect 5951 20216 6552 20244
rect 5951 20213 5963 20216
rect 5905 20207 5963 20213
rect 6546 20204 6552 20216
rect 6604 20204 6610 20256
rect 6917 20247 6975 20253
rect 6917 20213 6929 20247
rect 6963 20244 6975 20247
rect 8312 20244 8340 20284
rect 9306 20272 9312 20284
rect 9364 20272 9370 20324
rect 6963 20216 8340 20244
rect 8389 20247 8447 20253
rect 6963 20213 6975 20216
rect 6917 20207 6975 20213
rect 8389 20213 8401 20247
rect 8435 20244 8447 20247
rect 8478 20244 8484 20256
rect 8435 20216 8484 20244
rect 8435 20213 8447 20216
rect 8389 20207 8447 20213
rect 8478 20204 8484 20216
rect 8536 20204 8542 20256
rect 9401 20247 9459 20253
rect 9401 20213 9413 20247
rect 9447 20244 9459 20247
rect 9674 20244 9680 20256
rect 9447 20216 9680 20244
rect 9447 20213 9459 20216
rect 9401 20207 9459 20213
rect 9674 20204 9680 20216
rect 9732 20204 9738 20256
rect 9784 20253 9812 20488
rect 9876 20488 11336 20516
rect 9876 20457 9904 20488
rect 11330 20476 11336 20488
rect 11388 20476 11394 20528
rect 11606 20476 11612 20528
rect 11664 20516 11670 20528
rect 12069 20519 12127 20525
rect 12069 20516 12081 20519
rect 11664 20488 12081 20516
rect 11664 20476 11670 20488
rect 12069 20485 12081 20488
rect 12115 20485 12127 20519
rect 13078 20516 13084 20528
rect 13039 20488 13084 20516
rect 12069 20479 12127 20485
rect 13078 20476 13084 20488
rect 13136 20476 13142 20528
rect 13538 20476 13544 20528
rect 13596 20516 13602 20528
rect 13633 20519 13691 20525
rect 13633 20516 13645 20519
rect 13596 20488 13645 20516
rect 13596 20476 13602 20488
rect 13633 20485 13645 20488
rect 13679 20485 13691 20519
rect 13633 20479 13691 20485
rect 13998 20476 14004 20528
rect 14056 20516 14062 20528
rect 14737 20519 14795 20525
rect 14737 20516 14749 20519
rect 14056 20488 14749 20516
rect 14056 20476 14062 20488
rect 14737 20485 14749 20488
rect 14783 20485 14795 20519
rect 14737 20479 14795 20485
rect 16301 20519 16359 20525
rect 16301 20485 16313 20519
rect 16347 20516 16359 20519
rect 17678 20516 17684 20528
rect 16347 20488 17540 20516
rect 17639 20488 17684 20516
rect 16347 20485 16359 20488
rect 16301 20479 16359 20485
rect 9861 20451 9919 20457
rect 9861 20417 9873 20451
rect 9907 20417 9919 20451
rect 9861 20411 9919 20417
rect 9950 20408 9956 20460
rect 10008 20448 10014 20460
rect 11517 20451 11575 20457
rect 10008 20420 10053 20448
rect 10008 20408 10014 20420
rect 11517 20417 11529 20451
rect 11563 20448 11575 20451
rect 14918 20448 14924 20460
rect 11563 20420 14924 20448
rect 11563 20417 11575 20420
rect 11517 20411 11575 20417
rect 14918 20408 14924 20420
rect 14976 20408 14982 20460
rect 16574 20408 16580 20460
rect 16632 20448 16638 20460
rect 17221 20451 17279 20457
rect 17221 20448 17233 20451
rect 16632 20420 17233 20448
rect 16632 20408 16638 20420
rect 17221 20417 17233 20420
rect 17267 20417 17279 20451
rect 17512 20448 17540 20488
rect 17678 20476 17684 20488
rect 17736 20476 17742 20528
rect 18138 20476 18144 20528
rect 18196 20516 18202 20528
rect 18233 20519 18291 20525
rect 18233 20516 18245 20519
rect 18196 20488 18245 20516
rect 18196 20476 18202 20488
rect 18233 20485 18245 20488
rect 18279 20485 18291 20519
rect 18233 20479 18291 20485
rect 18598 20476 18604 20528
rect 18656 20516 18662 20528
rect 18785 20519 18843 20525
rect 18785 20516 18797 20519
rect 18656 20488 18797 20516
rect 18656 20476 18662 20488
rect 18785 20485 18797 20488
rect 18831 20485 18843 20519
rect 18785 20479 18843 20485
rect 19058 20476 19064 20528
rect 19116 20516 19122 20528
rect 20073 20519 20131 20525
rect 20073 20516 20085 20519
rect 19116 20488 20085 20516
rect 19116 20476 19122 20488
rect 20073 20485 20085 20488
rect 20119 20485 20131 20519
rect 20073 20479 20131 20485
rect 21358 20448 21364 20460
rect 17512 20420 21364 20448
rect 17221 20411 17279 20417
rect 21358 20408 21364 20420
rect 21416 20408 21422 20460
rect 10042 20340 10048 20392
rect 10100 20380 10106 20392
rect 10597 20383 10655 20389
rect 10597 20380 10609 20383
rect 10100 20352 10609 20380
rect 10100 20340 10106 20352
rect 10597 20349 10609 20352
rect 10643 20380 10655 20383
rect 10962 20380 10968 20392
rect 10643 20352 10968 20380
rect 10643 20349 10655 20352
rect 10597 20343 10655 20349
rect 10962 20340 10968 20352
rect 11020 20340 11026 20392
rect 12253 20383 12311 20389
rect 12253 20380 12265 20383
rect 11256 20352 12265 20380
rect 10134 20272 10140 20324
rect 10192 20312 10198 20324
rect 11256 20312 11284 20352
rect 12253 20349 12265 20352
rect 12299 20380 12311 20383
rect 12802 20380 12808 20392
rect 12299 20352 12808 20380
rect 12299 20349 12311 20352
rect 12253 20343 12311 20349
rect 12802 20340 12808 20352
rect 12860 20340 12866 20392
rect 14274 20380 14280 20392
rect 13096 20352 14280 20380
rect 10192 20284 11284 20312
rect 11333 20315 11391 20321
rect 10192 20272 10198 20284
rect 11333 20281 11345 20315
rect 11379 20312 11391 20315
rect 12621 20315 12679 20321
rect 11379 20284 12572 20312
rect 11379 20281 11391 20284
rect 11333 20275 11391 20281
rect 9769 20247 9827 20253
rect 9769 20213 9781 20247
rect 9815 20244 9827 20247
rect 10042 20244 10048 20256
rect 9815 20216 10048 20244
rect 9815 20213 9827 20216
rect 9769 20207 9827 20213
rect 10042 20204 10048 20216
rect 10100 20204 10106 20256
rect 10410 20244 10416 20256
rect 10371 20216 10416 20244
rect 10410 20204 10416 20216
rect 10468 20204 10474 20256
rect 10502 20204 10508 20256
rect 10560 20244 10566 20256
rect 12250 20244 12256 20256
rect 10560 20216 12256 20244
rect 10560 20204 10566 20216
rect 12250 20204 12256 20216
rect 12308 20204 12314 20256
rect 12544 20244 12572 20284
rect 12621 20281 12633 20315
rect 12667 20312 12679 20315
rect 13096 20312 13124 20352
rect 14274 20340 14280 20352
rect 14332 20340 14338 20392
rect 15749 20383 15807 20389
rect 15749 20349 15761 20383
rect 15795 20380 15807 20383
rect 15795 20352 19104 20380
rect 15795 20349 15807 20352
rect 15749 20343 15807 20349
rect 13262 20312 13268 20324
rect 12667 20284 13124 20312
rect 13223 20284 13268 20312
rect 12667 20281 12679 20284
rect 12621 20275 12679 20281
rect 13262 20272 13268 20284
rect 13320 20272 13326 20324
rect 13814 20312 13820 20324
rect 13775 20284 13820 20312
rect 13814 20272 13820 20284
rect 13872 20272 13878 20324
rect 13906 20272 13912 20324
rect 13964 20312 13970 20324
rect 14921 20315 14979 20321
rect 14921 20312 14933 20315
rect 13964 20284 14933 20312
rect 13964 20272 13970 20284
rect 14921 20281 14933 20284
rect 14967 20281 14979 20315
rect 15562 20312 15568 20324
rect 15523 20284 15568 20312
rect 14921 20275 14979 20281
rect 15562 20272 15568 20284
rect 15620 20272 15626 20324
rect 16114 20312 16120 20324
rect 16075 20284 16120 20312
rect 16114 20272 16120 20284
rect 16172 20272 16178 20324
rect 16669 20315 16727 20321
rect 16669 20281 16681 20315
rect 16715 20281 16727 20315
rect 16669 20275 16727 20281
rect 17865 20315 17923 20321
rect 17865 20281 17877 20315
rect 17911 20312 17923 20315
rect 18046 20312 18052 20324
rect 17911 20284 18052 20312
rect 17911 20281 17923 20284
rect 17865 20275 17923 20281
rect 13630 20244 13636 20256
rect 12544 20216 13636 20244
rect 13630 20204 13636 20216
rect 13688 20204 13694 20256
rect 16684 20244 16712 20275
rect 18046 20272 18052 20284
rect 18104 20272 18110 20324
rect 18417 20315 18475 20321
rect 18417 20281 18429 20315
rect 18463 20312 18475 20315
rect 18598 20312 18604 20324
rect 18463 20284 18604 20312
rect 18463 20281 18475 20284
rect 18417 20275 18475 20281
rect 18598 20272 18604 20284
rect 18656 20272 18662 20324
rect 18966 20312 18972 20324
rect 18927 20284 18972 20312
rect 18966 20272 18972 20284
rect 19024 20272 19030 20324
rect 19076 20312 19104 20352
rect 19334 20340 19340 20392
rect 19392 20380 19398 20392
rect 20257 20383 20315 20389
rect 20257 20380 20269 20383
rect 19392 20352 20269 20380
rect 19392 20340 19398 20352
rect 20257 20349 20269 20352
rect 20303 20349 20315 20383
rect 20257 20343 20315 20349
rect 20809 20383 20867 20389
rect 20809 20349 20821 20383
rect 20855 20380 20867 20383
rect 21269 20383 21327 20389
rect 21269 20380 21281 20383
rect 20855 20352 21281 20380
rect 20855 20349 20867 20352
rect 20809 20343 20867 20349
rect 21269 20349 21281 20352
rect 21315 20380 21327 20383
rect 22738 20380 22744 20392
rect 21315 20352 22744 20380
rect 21315 20349 21327 20352
rect 21269 20343 21327 20349
rect 22738 20340 22744 20352
rect 22796 20340 22802 20392
rect 21818 20312 21824 20324
rect 19076 20284 21824 20312
rect 21818 20272 21824 20284
rect 21876 20272 21882 20324
rect 18874 20244 18880 20256
rect 16684 20216 18880 20244
rect 18874 20204 18880 20216
rect 18932 20204 18938 20256
rect 19242 20204 19248 20256
rect 19300 20244 19306 20256
rect 19337 20247 19395 20253
rect 19337 20244 19349 20247
rect 19300 20216 19349 20244
rect 19300 20204 19306 20216
rect 19337 20213 19349 20216
rect 19383 20213 19395 20247
rect 21174 20244 21180 20256
rect 21135 20216 21180 20244
rect 19337 20207 19395 20213
rect 21174 20204 21180 20216
rect 21232 20204 21238 20256
rect 1104 20154 21896 20176
rect 1104 20102 7912 20154
rect 7964 20102 7976 20154
rect 8028 20102 8040 20154
rect 8092 20102 8104 20154
rect 8156 20102 14843 20154
rect 14895 20102 14907 20154
rect 14959 20102 14971 20154
rect 15023 20102 15035 20154
rect 15087 20102 21896 20154
rect 1104 20080 21896 20102
rect 3053 20043 3111 20049
rect 3053 20009 3065 20043
rect 3099 20040 3111 20043
rect 4062 20040 4068 20052
rect 3099 20012 4068 20040
rect 3099 20009 3111 20012
rect 3053 20003 3111 20009
rect 4062 20000 4068 20012
rect 4120 20000 4126 20052
rect 4801 20043 4859 20049
rect 4801 20009 4813 20043
rect 4847 20040 4859 20043
rect 5442 20040 5448 20052
rect 4847 20012 5448 20040
rect 4847 20009 4859 20012
rect 4801 20003 4859 20009
rect 5442 20000 5448 20012
rect 5500 20000 5506 20052
rect 5994 20000 6000 20052
rect 6052 20040 6058 20052
rect 7193 20043 7251 20049
rect 7193 20040 7205 20043
rect 6052 20012 7205 20040
rect 6052 20000 6058 20012
rect 7193 20009 7205 20012
rect 7239 20009 7251 20043
rect 7193 20003 7251 20009
rect 7282 20000 7288 20052
rect 7340 20040 7346 20052
rect 8386 20040 8392 20052
rect 7340 20012 8392 20040
rect 7340 20000 7346 20012
rect 8386 20000 8392 20012
rect 8444 20000 8450 20052
rect 8481 20043 8539 20049
rect 8481 20009 8493 20043
rect 8527 20040 8539 20043
rect 10410 20040 10416 20052
rect 8527 20012 10416 20040
rect 8527 20009 8539 20012
rect 8481 20003 8539 20009
rect 10410 20000 10416 20012
rect 10468 20000 10474 20052
rect 10502 20000 10508 20052
rect 10560 20040 10566 20052
rect 12161 20043 12219 20049
rect 12161 20040 12173 20043
rect 10560 20012 12173 20040
rect 10560 20000 10566 20012
rect 12161 20009 12173 20012
rect 12207 20009 12219 20043
rect 12161 20003 12219 20009
rect 12529 20043 12587 20049
rect 12529 20009 12541 20043
rect 12575 20040 12587 20043
rect 12621 20043 12679 20049
rect 12621 20040 12633 20043
rect 12575 20012 12633 20040
rect 12575 20009 12587 20012
rect 12529 20003 12587 20009
rect 12621 20009 12633 20012
rect 12667 20009 12679 20043
rect 12802 20040 12808 20052
rect 12763 20012 12808 20040
rect 12621 20003 12679 20009
rect 12802 20000 12808 20012
rect 12860 20000 12866 20052
rect 13357 20043 13415 20049
rect 13357 20009 13369 20043
rect 13403 20040 13415 20043
rect 13906 20040 13912 20052
rect 13403 20012 13912 20040
rect 13403 20009 13415 20012
rect 13357 20003 13415 20009
rect 13906 20000 13912 20012
rect 13964 20000 13970 20052
rect 16114 20000 16120 20052
rect 16172 20040 16178 20052
rect 16172 20012 17172 20040
rect 16172 20000 16178 20012
rect 1302 19932 1308 19984
rect 1360 19972 1366 19984
rect 5074 19972 5080 19984
rect 1360 19944 5080 19972
rect 1360 19932 1366 19944
rect 5074 19932 5080 19944
rect 5132 19932 5138 19984
rect 6086 19932 6092 19984
rect 6144 19972 6150 19984
rect 6650 19975 6708 19981
rect 6650 19972 6662 19975
rect 6144 19944 6662 19972
rect 6144 19932 6150 19944
rect 6650 19941 6662 19944
rect 6696 19941 6708 19975
rect 6650 19935 6708 19941
rect 7558 19932 7564 19984
rect 7616 19972 7622 19984
rect 10870 19972 10876 19984
rect 7616 19944 10876 19972
rect 7616 19932 7622 19944
rect 10870 19932 10876 19944
rect 10928 19932 10934 19984
rect 11054 19932 11060 19984
rect 11112 19972 11118 19984
rect 11158 19975 11216 19981
rect 11158 19972 11170 19975
rect 11112 19944 11170 19972
rect 11112 19932 11118 19944
rect 11158 19941 11170 19944
rect 11204 19941 11216 19975
rect 15378 19972 15384 19984
rect 15339 19944 15384 19972
rect 11158 19935 11216 19941
rect 15378 19932 15384 19944
rect 15436 19932 15442 19984
rect 15838 19932 15844 19984
rect 15896 19972 15902 19984
rect 15933 19975 15991 19981
rect 15933 19972 15945 19975
rect 15896 19944 15945 19972
rect 15896 19932 15902 19944
rect 15933 19941 15945 19944
rect 15979 19941 15991 19975
rect 15933 19935 15991 19941
rect 16298 19932 16304 19984
rect 16356 19972 16362 19984
rect 16485 19975 16543 19981
rect 16485 19972 16497 19975
rect 16356 19944 16497 19972
rect 16356 19932 16362 19944
rect 16485 19941 16497 19944
rect 16531 19941 16543 19975
rect 16485 19935 16543 19941
rect 16758 19932 16764 19984
rect 16816 19972 16822 19984
rect 17037 19975 17095 19981
rect 17037 19972 17049 19975
rect 16816 19944 17049 19972
rect 16816 19932 16822 19944
rect 17037 19941 17049 19944
rect 17083 19941 17095 19975
rect 17144 19972 17172 20012
rect 17218 20000 17224 20052
rect 17276 20040 17282 20052
rect 17681 20043 17739 20049
rect 17681 20040 17693 20043
rect 17276 20012 17693 20040
rect 17276 20000 17282 20012
rect 17681 20009 17693 20012
rect 17727 20009 17739 20043
rect 17681 20003 17739 20009
rect 18325 20043 18383 20049
rect 18325 20009 18337 20043
rect 18371 20040 18383 20043
rect 18966 20040 18972 20052
rect 18371 20012 18972 20040
rect 18371 20009 18383 20012
rect 18325 20003 18383 20009
rect 18966 20000 18972 20012
rect 19024 20000 19030 20052
rect 19150 19972 19156 19984
rect 17144 19944 19156 19972
rect 17037 19935 17095 19941
rect 19150 19932 19156 19944
rect 19208 19932 19214 19984
rect 19978 19972 19984 19984
rect 19939 19944 19984 19972
rect 19978 19932 19984 19944
rect 20036 19932 20042 19984
rect 20438 19932 20444 19984
rect 20496 19972 20502 19984
rect 20533 19975 20591 19981
rect 20533 19972 20545 19975
rect 20496 19944 20545 19972
rect 20496 19932 20502 19944
rect 20533 19941 20545 19944
rect 20579 19941 20591 19975
rect 20533 19935 20591 19941
rect 20898 19932 20904 19984
rect 20956 19972 20962 19984
rect 21085 19975 21143 19981
rect 21085 19972 21097 19975
rect 20956 19944 21097 19972
rect 20956 19932 20962 19944
rect 21085 19941 21097 19944
rect 21131 19941 21143 19975
rect 21085 19935 21143 19941
rect 1765 19907 1823 19913
rect 1765 19873 1777 19907
rect 1811 19904 1823 19907
rect 2038 19904 2044 19916
rect 1811 19876 2044 19904
rect 1811 19873 1823 19876
rect 1765 19867 1823 19873
rect 2038 19864 2044 19876
rect 2096 19864 2102 19916
rect 2317 19907 2375 19913
rect 2317 19873 2329 19907
rect 2363 19904 2375 19907
rect 2498 19904 2504 19916
rect 2363 19876 2504 19904
rect 2363 19873 2375 19876
rect 2317 19867 2375 19873
rect 2498 19864 2504 19876
rect 2556 19864 2562 19916
rect 3145 19907 3203 19913
rect 3145 19873 3157 19907
rect 3191 19904 3203 19907
rect 4065 19907 4123 19913
rect 4065 19904 4077 19907
rect 3191 19876 4077 19904
rect 3191 19873 3203 19876
rect 3145 19867 3203 19873
rect 4065 19873 4077 19876
rect 4111 19873 4123 19907
rect 4065 19867 4123 19873
rect 4893 19907 4951 19913
rect 4893 19873 4905 19907
rect 4939 19904 4951 19907
rect 6362 19904 6368 19916
rect 4939 19876 6368 19904
rect 4939 19873 4951 19876
rect 4893 19867 4951 19873
rect 6362 19864 6368 19876
rect 6420 19864 6426 19916
rect 6822 19864 6828 19916
rect 6880 19904 6886 19916
rect 6917 19907 6975 19913
rect 6917 19904 6929 19907
rect 6880 19876 6929 19904
rect 6880 19864 6886 19876
rect 6917 19873 6929 19876
rect 6963 19873 6975 19907
rect 7377 19907 7435 19913
rect 7377 19904 7389 19907
rect 6917 19867 6975 19873
rect 7024 19876 7389 19904
rect 2961 19839 3019 19845
rect 2961 19805 2973 19839
rect 3007 19805 3019 19839
rect 2961 19799 3019 19805
rect 4709 19839 4767 19845
rect 4709 19805 4721 19839
rect 4755 19836 4767 19839
rect 4755 19808 5580 19836
rect 4755 19805 4767 19808
rect 4709 19799 4767 19805
rect 1578 19768 1584 19780
rect 1539 19740 1584 19768
rect 1578 19728 1584 19740
rect 1636 19728 1642 19780
rect 2501 19771 2559 19777
rect 2501 19737 2513 19771
rect 2547 19768 2559 19771
rect 2976 19768 3004 19799
rect 5552 19780 5580 19808
rect 3142 19768 3148 19780
rect 2547 19740 2774 19768
rect 2976 19740 3148 19768
rect 2547 19737 2559 19740
rect 2501 19731 2559 19737
rect 2746 19700 2774 19740
rect 3142 19728 3148 19740
rect 3200 19728 3206 19780
rect 5350 19768 5356 19780
rect 3252 19740 5356 19768
rect 3252 19700 3280 19740
rect 5350 19728 5356 19740
rect 5408 19728 5414 19780
rect 5534 19768 5540 19780
rect 5447 19740 5540 19768
rect 5534 19728 5540 19740
rect 5592 19728 5598 19780
rect 2746 19672 3280 19700
rect 3513 19703 3571 19709
rect 3513 19669 3525 19703
rect 3559 19700 3571 19703
rect 5166 19700 5172 19712
rect 3559 19672 5172 19700
rect 3559 19669 3571 19672
rect 3513 19663 3571 19669
rect 5166 19660 5172 19672
rect 5224 19660 5230 19712
rect 5261 19703 5319 19709
rect 5261 19669 5273 19703
rect 5307 19700 5319 19703
rect 7024 19700 7052 19876
rect 7377 19873 7389 19876
rect 7423 19873 7435 19907
rect 7377 19867 7435 19873
rect 8662 19864 8668 19916
rect 8720 19904 8726 19916
rect 9493 19907 9551 19913
rect 9493 19904 9505 19907
rect 8720 19876 9505 19904
rect 8720 19864 8726 19876
rect 9493 19873 9505 19876
rect 9539 19873 9551 19907
rect 9493 19867 9551 19873
rect 9582 19864 9588 19916
rect 9640 19904 9646 19916
rect 10686 19904 10692 19916
rect 9640 19876 10692 19904
rect 9640 19864 9646 19876
rect 10686 19864 10692 19876
rect 10744 19864 10750 19916
rect 11330 19864 11336 19916
rect 11388 19904 11394 19916
rect 11425 19907 11483 19913
rect 11425 19904 11437 19907
rect 11388 19876 11437 19904
rect 11388 19864 11394 19876
rect 11425 19873 11437 19876
rect 11471 19873 11483 19907
rect 11425 19867 11483 19873
rect 11885 19907 11943 19913
rect 11885 19873 11897 19907
rect 11931 19873 11943 19907
rect 12342 19904 12348 19916
rect 12303 19876 12348 19904
rect 11885 19867 11943 19873
rect 8573 19839 8631 19845
rect 8573 19805 8585 19839
rect 8619 19805 8631 19839
rect 8573 19799 8631 19805
rect 8588 19768 8616 19799
rect 8846 19796 8852 19848
rect 8904 19836 8910 19848
rect 8904 19808 10180 19836
rect 8904 19796 8910 19808
rect 8754 19768 8760 19780
rect 8588 19740 8760 19768
rect 8754 19728 8760 19740
rect 8812 19768 8818 19780
rect 10045 19771 10103 19777
rect 10045 19768 10057 19771
rect 8812 19740 10057 19768
rect 8812 19728 8818 19740
rect 10045 19737 10057 19740
rect 10091 19737 10103 19771
rect 10045 19731 10103 19737
rect 5307 19672 7052 19700
rect 5307 19669 5319 19672
rect 5261 19663 5319 19669
rect 7282 19660 7288 19712
rect 7340 19700 7346 19712
rect 7650 19700 7656 19712
rect 7340 19672 7656 19700
rect 7340 19660 7346 19672
rect 7650 19660 7656 19672
rect 7708 19660 7714 19712
rect 7742 19660 7748 19712
rect 7800 19700 7806 19712
rect 8021 19703 8079 19709
rect 8021 19700 8033 19703
rect 7800 19672 8033 19700
rect 7800 19660 7806 19672
rect 8021 19669 8033 19672
rect 8067 19669 8079 19703
rect 8021 19663 8079 19669
rect 8202 19660 8208 19712
rect 8260 19700 8266 19712
rect 9309 19703 9367 19709
rect 9309 19700 9321 19703
rect 8260 19672 9321 19700
rect 8260 19660 8266 19672
rect 9309 19669 9321 19672
rect 9355 19669 9367 19703
rect 10152 19700 10180 19808
rect 11790 19700 11796 19712
rect 10152 19672 11796 19700
rect 9309 19663 9367 19669
rect 11790 19660 11796 19672
rect 11848 19660 11854 19712
rect 11900 19700 11928 19867
rect 12342 19864 12348 19876
rect 12400 19864 12406 19916
rect 12621 19907 12679 19913
rect 12621 19873 12633 19907
rect 12667 19904 12679 19907
rect 13173 19907 13231 19913
rect 13173 19904 13185 19907
rect 12667 19876 13185 19904
rect 12667 19873 12679 19876
rect 12621 19867 12679 19873
rect 13173 19873 13185 19876
rect 13219 19873 13231 19907
rect 13173 19867 13231 19873
rect 13817 19907 13875 19913
rect 13817 19873 13829 19907
rect 13863 19873 13875 19907
rect 13817 19867 13875 19873
rect 13832 19836 13860 19867
rect 14182 19864 14188 19916
rect 14240 19904 14246 19916
rect 14645 19907 14703 19913
rect 14645 19904 14657 19907
rect 14240 19876 14657 19904
rect 14240 19864 14246 19876
rect 14645 19873 14657 19876
rect 14691 19873 14703 19907
rect 14645 19867 14703 19873
rect 15194 19864 15200 19916
rect 15252 19904 15258 19916
rect 15565 19907 15623 19913
rect 15565 19904 15577 19907
rect 15252 19876 15577 19904
rect 15252 19864 15258 19876
rect 15565 19873 15577 19876
rect 15611 19873 15623 19907
rect 16114 19904 16120 19916
rect 16075 19876 16120 19904
rect 15565 19867 15623 19873
rect 16114 19864 16120 19876
rect 16172 19864 16178 19916
rect 16666 19904 16672 19916
rect 16627 19876 16672 19904
rect 16666 19864 16672 19876
rect 16724 19864 16730 19916
rect 17218 19904 17224 19916
rect 17179 19876 17224 19904
rect 17218 19864 17224 19876
rect 17276 19864 17282 19916
rect 17770 19904 17776 19916
rect 17731 19876 17776 19904
rect 17770 19864 17776 19876
rect 17828 19864 17834 19916
rect 18138 19904 18144 19916
rect 18099 19876 18144 19904
rect 18138 19864 18144 19876
rect 18196 19864 18202 19916
rect 18601 19907 18659 19913
rect 18601 19873 18613 19907
rect 18647 19904 18659 19907
rect 18690 19904 18696 19916
rect 18647 19876 18696 19904
rect 18647 19873 18659 19876
rect 18601 19867 18659 19873
rect 18690 19864 18696 19876
rect 18748 19864 18754 19916
rect 19702 19864 19708 19916
rect 19760 19904 19766 19916
rect 20165 19907 20223 19913
rect 20165 19904 20177 19907
rect 19760 19876 20177 19904
rect 19760 19864 19766 19876
rect 20165 19873 20177 19876
rect 20211 19873 20223 19907
rect 20165 19867 20223 19873
rect 20717 19907 20775 19913
rect 20717 19873 20729 19907
rect 20763 19873 20775 19907
rect 20717 19867 20775 19873
rect 21269 19907 21327 19913
rect 21269 19873 21281 19907
rect 21315 19873 21327 19907
rect 21269 19867 21327 19873
rect 12084 19808 13860 19836
rect 12084 19777 12112 19808
rect 13998 19796 14004 19848
rect 14056 19836 14062 19848
rect 19426 19836 19432 19848
rect 14056 19808 19432 19836
rect 14056 19796 14062 19808
rect 19426 19796 19432 19808
rect 19484 19836 19490 19848
rect 19613 19839 19671 19845
rect 19613 19836 19625 19839
rect 19484 19808 19625 19836
rect 19484 19796 19490 19808
rect 19613 19805 19625 19808
rect 19659 19805 19671 19839
rect 19613 19799 19671 19805
rect 19978 19796 19984 19848
rect 20036 19836 20042 19848
rect 20732 19836 20760 19867
rect 20036 19808 20760 19836
rect 20036 19796 20042 19808
rect 12069 19771 12127 19777
rect 12069 19737 12081 19771
rect 12115 19737 12127 19771
rect 12069 19731 12127 19737
rect 12161 19771 12219 19777
rect 12161 19737 12173 19771
rect 12207 19768 12219 19771
rect 13630 19768 13636 19780
rect 12207 19740 13492 19768
rect 13591 19740 13636 19768
rect 12207 19737 12219 19740
rect 12161 19731 12219 19737
rect 13170 19700 13176 19712
rect 11900 19672 13176 19700
rect 13170 19660 13176 19672
rect 13228 19660 13234 19712
rect 13464 19700 13492 19740
rect 13630 19728 13636 19740
rect 13688 19728 13694 19780
rect 19061 19771 19119 19777
rect 19061 19768 19073 19771
rect 14752 19740 19073 19768
rect 14752 19700 14780 19740
rect 19061 19737 19073 19740
rect 19107 19768 19119 19771
rect 19242 19768 19248 19780
rect 19107 19740 19248 19768
rect 19107 19737 19119 19740
rect 19061 19731 19119 19737
rect 19242 19728 19248 19740
rect 19300 19728 19306 19780
rect 19794 19728 19800 19780
rect 19852 19768 19858 19780
rect 21284 19768 21312 19867
rect 19852 19740 21312 19768
rect 19852 19728 19858 19740
rect 13464 19672 14780 19700
rect 14829 19703 14887 19709
rect 14829 19669 14841 19703
rect 14875 19700 14887 19703
rect 15286 19700 15292 19712
rect 14875 19672 15292 19700
rect 14875 19669 14887 19672
rect 14829 19663 14887 19669
rect 15286 19660 15292 19672
rect 15344 19660 15350 19712
rect 18785 19703 18843 19709
rect 18785 19669 18797 19703
rect 18831 19700 18843 19703
rect 18966 19700 18972 19712
rect 18831 19672 18972 19700
rect 18831 19669 18843 19672
rect 18785 19663 18843 19669
rect 18966 19660 18972 19672
rect 19024 19660 19030 19712
rect 1104 19610 21896 19632
rect 1104 19558 4447 19610
rect 4499 19558 4511 19610
rect 4563 19558 4575 19610
rect 4627 19558 4639 19610
rect 4691 19558 11378 19610
rect 11430 19558 11442 19610
rect 11494 19558 11506 19610
rect 11558 19558 11570 19610
rect 11622 19558 18308 19610
rect 18360 19558 18372 19610
rect 18424 19558 18436 19610
rect 18488 19558 18500 19610
rect 18552 19558 21896 19610
rect 1104 19536 21896 19558
rect 3418 19456 3424 19508
rect 3476 19496 3482 19508
rect 4246 19496 4252 19508
rect 3476 19468 4108 19496
rect 4159 19468 4252 19496
rect 3476 19456 3482 19468
rect 2222 19388 2228 19440
rect 2280 19428 2286 19440
rect 2501 19431 2559 19437
rect 2501 19428 2513 19431
rect 2280 19400 2513 19428
rect 2280 19388 2286 19400
rect 2501 19397 2513 19400
rect 2547 19397 2559 19431
rect 2501 19391 2559 19397
rect 4080 19360 4108 19468
rect 4246 19456 4252 19468
rect 4304 19496 4310 19508
rect 4709 19499 4767 19505
rect 4709 19496 4721 19499
rect 4304 19468 4721 19496
rect 4304 19456 4310 19468
rect 4709 19465 4721 19468
rect 4755 19465 4767 19499
rect 4709 19459 4767 19465
rect 5166 19456 5172 19508
rect 5224 19496 5230 19508
rect 6454 19496 6460 19508
rect 5224 19468 6460 19496
rect 5224 19456 5230 19468
rect 6454 19456 6460 19468
rect 6512 19456 6518 19508
rect 6822 19496 6828 19508
rect 6564 19468 6828 19496
rect 6564 19428 6592 19468
rect 6822 19456 6828 19468
rect 6880 19456 6886 19508
rect 7098 19456 7104 19508
rect 7156 19496 7162 19508
rect 7156 19468 10732 19496
rect 7156 19456 7162 19468
rect 6288 19400 6592 19428
rect 4080 19332 4200 19360
rect 1578 19292 1584 19304
rect 1539 19264 1584 19292
rect 1578 19252 1584 19264
rect 1636 19252 1642 19304
rect 2133 19295 2191 19301
rect 2133 19261 2145 19295
rect 2179 19292 2191 19295
rect 2774 19292 2780 19304
rect 2179 19264 2780 19292
rect 2179 19261 2191 19264
rect 2133 19255 2191 19261
rect 2774 19252 2780 19264
rect 2832 19252 2838 19304
rect 4062 19292 4068 19304
rect 4023 19264 4068 19292
rect 4062 19252 4068 19264
rect 4120 19252 4126 19304
rect 4172 19292 4200 19332
rect 6288 19304 6316 19400
rect 6638 19388 6644 19440
rect 6696 19388 6702 19440
rect 6656 19360 6684 19388
rect 10704 19360 10732 19468
rect 10870 19456 10876 19508
rect 10928 19496 10934 19508
rect 13078 19496 13084 19508
rect 10928 19468 13084 19496
rect 10928 19456 10934 19468
rect 13078 19456 13084 19468
rect 13136 19456 13142 19508
rect 13173 19499 13231 19505
rect 13173 19465 13185 19499
rect 13219 19496 13231 19499
rect 13262 19496 13268 19508
rect 13219 19468 13268 19496
rect 13219 19465 13231 19468
rect 13173 19459 13231 19465
rect 13262 19456 13268 19468
rect 13320 19456 13326 19508
rect 13814 19496 13820 19508
rect 13775 19468 13820 19496
rect 13814 19456 13820 19468
rect 13872 19456 13878 19508
rect 14274 19496 14280 19508
rect 14235 19468 14280 19496
rect 14274 19456 14280 19468
rect 14332 19456 14338 19508
rect 15473 19499 15531 19505
rect 15473 19465 15485 19499
rect 15519 19496 15531 19499
rect 16114 19496 16120 19508
rect 15519 19468 16120 19496
rect 15519 19465 15531 19468
rect 15473 19459 15531 19465
rect 16114 19456 16120 19468
rect 16172 19456 16178 19508
rect 17129 19499 17187 19505
rect 17129 19465 17141 19499
rect 17175 19496 17187 19499
rect 17218 19496 17224 19508
rect 17175 19468 17224 19496
rect 17175 19465 17187 19468
rect 17129 19459 17187 19465
rect 17218 19456 17224 19468
rect 17276 19456 17282 19508
rect 17770 19496 17776 19508
rect 17731 19468 17776 19496
rect 17770 19456 17776 19468
rect 17828 19456 17834 19508
rect 18046 19496 18052 19508
rect 18007 19468 18052 19496
rect 18046 19456 18052 19468
rect 18104 19456 18110 19508
rect 18509 19499 18567 19505
rect 18509 19465 18521 19499
rect 18555 19496 18567 19499
rect 18598 19496 18604 19508
rect 18555 19468 18604 19496
rect 18555 19465 18567 19468
rect 18509 19459 18567 19465
rect 18598 19456 18604 19468
rect 18656 19456 18662 19508
rect 19426 19496 19432 19508
rect 19387 19468 19432 19496
rect 19426 19456 19432 19468
rect 19484 19456 19490 19508
rect 11146 19388 11152 19440
rect 11204 19428 11210 19440
rect 11330 19428 11336 19440
rect 11204 19400 11336 19428
rect 11204 19388 11210 19400
rect 11330 19388 11336 19400
rect 11388 19388 11394 19440
rect 12526 19388 12532 19440
rect 12584 19388 12590 19440
rect 12713 19431 12771 19437
rect 12713 19397 12725 19431
rect 12759 19397 12771 19431
rect 12713 19391 12771 19397
rect 12544 19360 12572 19388
rect 6656 19332 6776 19360
rect 10704 19332 12572 19360
rect 4172 19264 4936 19292
rect 1765 19227 1823 19233
rect 1765 19193 1777 19227
rect 1811 19193 1823 19227
rect 1765 19187 1823 19193
rect 1780 19156 1808 19187
rect 2222 19184 2228 19236
rect 2280 19224 2286 19236
rect 2317 19227 2375 19233
rect 2317 19224 2329 19227
rect 2280 19196 2329 19224
rect 2280 19184 2286 19196
rect 2317 19193 2329 19196
rect 2363 19193 2375 19227
rect 3820 19227 3878 19233
rect 2317 19187 2375 19193
rect 2608 19196 3280 19224
rect 2406 19156 2412 19168
rect 1780 19128 2412 19156
rect 2406 19116 2412 19128
rect 2464 19116 2470 19168
rect 2501 19159 2559 19165
rect 2501 19125 2513 19159
rect 2547 19156 2559 19159
rect 2608 19156 2636 19196
rect 2547 19128 2636 19156
rect 2685 19159 2743 19165
rect 2547 19125 2559 19128
rect 2501 19119 2559 19125
rect 2685 19125 2697 19159
rect 2731 19156 2743 19159
rect 3142 19156 3148 19168
rect 2731 19128 3148 19156
rect 2731 19125 2743 19128
rect 2685 19119 2743 19125
rect 3142 19116 3148 19128
rect 3200 19116 3206 19168
rect 3252 19156 3280 19196
rect 3820 19193 3832 19227
rect 3866 19224 3878 19227
rect 4249 19227 4307 19233
rect 4249 19224 4261 19227
rect 3866 19196 4261 19224
rect 3866 19193 3878 19196
rect 3820 19187 3878 19193
rect 4249 19193 4261 19196
rect 4295 19193 4307 19227
rect 4908 19224 4936 19264
rect 5534 19252 5540 19304
rect 5592 19292 5598 19304
rect 5822 19295 5880 19301
rect 5822 19292 5834 19295
rect 5592 19264 5834 19292
rect 5592 19252 5598 19264
rect 5822 19261 5834 19264
rect 5868 19261 5880 19295
rect 5822 19255 5880 19261
rect 6089 19295 6147 19301
rect 6089 19261 6101 19295
rect 6135 19292 6147 19295
rect 6270 19292 6276 19304
rect 6135 19264 6276 19292
rect 6135 19261 6147 19264
rect 6089 19255 6147 19261
rect 6270 19252 6276 19264
rect 6328 19252 6334 19304
rect 6362 19252 6368 19304
rect 6420 19292 6426 19304
rect 6641 19295 6699 19301
rect 6641 19292 6653 19295
rect 6420 19264 6653 19292
rect 6420 19252 6426 19264
rect 6641 19261 6653 19264
rect 6687 19261 6699 19295
rect 6748 19292 6776 19332
rect 8593 19295 8651 19301
rect 6748 19264 8064 19292
rect 6641 19255 6699 19261
rect 7101 19227 7159 19233
rect 7101 19224 7113 19227
rect 4908 19196 7113 19224
rect 4249 19187 4307 19193
rect 7101 19193 7113 19196
rect 7147 19193 7159 19227
rect 7101 19187 7159 19193
rect 4341 19159 4399 19165
rect 4341 19156 4353 19159
rect 3252 19128 4353 19156
rect 4341 19125 4353 19128
rect 4387 19125 4399 19159
rect 4341 19119 4399 19125
rect 4430 19116 4436 19168
rect 4488 19156 4494 19168
rect 7282 19156 7288 19168
rect 4488 19128 7288 19156
rect 4488 19116 4494 19128
rect 7282 19116 7288 19128
rect 7340 19116 7346 19168
rect 7466 19156 7472 19168
rect 7427 19128 7472 19156
rect 7466 19116 7472 19128
rect 7524 19116 7530 19168
rect 8036 19156 8064 19264
rect 8593 19261 8605 19295
rect 8639 19292 8651 19295
rect 8754 19292 8760 19304
rect 8639 19264 8760 19292
rect 8639 19261 8651 19264
rect 8593 19255 8651 19261
rect 8754 19252 8760 19264
rect 8812 19252 8818 19304
rect 8849 19295 8907 19301
rect 8849 19261 8861 19295
rect 8895 19292 8907 19295
rect 9214 19292 9220 19304
rect 8895 19264 9220 19292
rect 8895 19261 8907 19264
rect 8849 19255 8907 19261
rect 9214 19252 9220 19264
rect 9272 19292 9278 19304
rect 9950 19301 9956 19304
rect 9677 19295 9735 19301
rect 9677 19292 9689 19295
rect 9272 19264 9689 19292
rect 9272 19252 9278 19264
rect 9677 19261 9689 19264
rect 9723 19261 9735 19295
rect 9944 19292 9956 19301
rect 9911 19264 9956 19292
rect 9677 19255 9735 19261
rect 9944 19255 9956 19264
rect 9950 19252 9956 19255
rect 10008 19252 10014 19304
rect 10962 19252 10968 19304
rect 11020 19292 11026 19304
rect 11701 19295 11759 19301
rect 11701 19292 11713 19295
rect 11020 19264 11713 19292
rect 11020 19252 11026 19264
rect 11701 19261 11713 19264
rect 11747 19261 11759 19295
rect 12066 19292 12072 19304
rect 12027 19264 12072 19292
rect 11701 19255 11759 19261
rect 12066 19252 12072 19264
rect 12124 19252 12130 19304
rect 12526 19292 12532 19304
rect 12487 19264 12532 19292
rect 12526 19252 12532 19264
rect 12584 19252 12590 19304
rect 12728 19292 12756 19391
rect 12802 19388 12808 19440
rect 12860 19428 12866 19440
rect 13446 19428 13452 19440
rect 12860 19400 13452 19428
rect 12860 19388 12866 19400
rect 13446 19388 13452 19400
rect 13504 19388 13510 19440
rect 16025 19431 16083 19437
rect 16025 19397 16037 19431
rect 16071 19428 16083 19431
rect 16666 19428 16672 19440
rect 16071 19400 16672 19428
rect 16071 19397 16083 19400
rect 16025 19391 16083 19397
rect 16666 19388 16672 19400
rect 16724 19388 16730 19440
rect 15562 19320 15568 19372
rect 15620 19360 15626 19372
rect 15620 19332 19932 19360
rect 15620 19320 15626 19332
rect 12989 19295 13047 19301
rect 12989 19292 13001 19295
rect 12728 19264 13001 19292
rect 12989 19261 13001 19264
rect 13035 19261 13047 19295
rect 13998 19292 14004 19304
rect 12989 19255 13047 19261
rect 13188 19264 13584 19292
rect 13959 19264 14004 19292
rect 8110 19184 8116 19236
rect 8168 19224 8174 19236
rect 10410 19224 10416 19236
rect 8168 19196 10416 19224
rect 8168 19184 8174 19196
rect 10410 19184 10416 19196
rect 10468 19184 10474 19236
rect 9306 19156 9312 19168
rect 8036 19128 9312 19156
rect 9306 19116 9312 19128
rect 9364 19116 9370 19168
rect 9401 19159 9459 19165
rect 9401 19125 9413 19159
rect 9447 19156 9459 19159
rect 9674 19156 9680 19168
rect 9447 19128 9680 19156
rect 9447 19125 9459 19128
rect 9401 19119 9459 19125
rect 9674 19116 9680 19128
rect 9732 19116 9738 19168
rect 11054 19156 11060 19168
rect 11015 19128 11060 19156
rect 11054 19116 11060 19128
rect 11112 19116 11118 19168
rect 12253 19159 12311 19165
rect 12253 19125 12265 19159
rect 12299 19156 12311 19159
rect 13188 19156 13216 19264
rect 13354 19184 13360 19236
rect 13412 19224 13418 19236
rect 13449 19227 13507 19233
rect 13449 19224 13461 19227
rect 13412 19196 13461 19224
rect 13412 19184 13418 19196
rect 13449 19193 13461 19196
rect 13495 19193 13507 19227
rect 13556 19224 13584 19264
rect 13998 19252 14004 19264
rect 14056 19252 14062 19304
rect 14461 19295 14519 19301
rect 14461 19261 14473 19295
rect 14507 19261 14519 19295
rect 14461 19255 14519 19261
rect 14737 19295 14795 19301
rect 14737 19261 14749 19295
rect 14783 19261 14795 19295
rect 15286 19292 15292 19304
rect 15247 19264 15292 19292
rect 14737 19255 14795 19261
rect 14476 19224 14504 19255
rect 13556 19196 14504 19224
rect 13449 19187 13507 19193
rect 12299 19128 13216 19156
rect 12299 19125 12311 19128
rect 12253 19119 12311 19125
rect 13262 19116 13268 19168
rect 13320 19156 13326 19168
rect 14752 19156 14780 19255
rect 15286 19252 15292 19264
rect 15344 19252 15350 19304
rect 15841 19295 15899 19301
rect 15841 19261 15853 19295
rect 15887 19292 15899 19295
rect 16482 19292 16488 19304
rect 15887 19264 16344 19292
rect 16443 19264 16488 19292
rect 15887 19261 15899 19264
rect 15841 19255 15899 19261
rect 13320 19128 14780 19156
rect 14921 19159 14979 19165
rect 13320 19116 13326 19128
rect 14921 19125 14933 19159
rect 14967 19156 14979 19159
rect 15194 19156 15200 19168
rect 14967 19128 15200 19156
rect 14967 19125 14979 19128
rect 14921 19119 14979 19125
rect 15194 19116 15200 19128
rect 15252 19116 15258 19168
rect 16316 19165 16344 19264
rect 16482 19252 16488 19264
rect 16540 19252 16546 19304
rect 17310 19292 17316 19304
rect 17271 19264 17316 19292
rect 17310 19252 17316 19264
rect 17368 19252 17374 19304
rect 17589 19295 17647 19301
rect 17589 19261 17601 19295
rect 17635 19292 17647 19295
rect 17862 19292 17868 19304
rect 17635 19264 17868 19292
rect 17635 19261 17647 19264
rect 17589 19255 17647 19261
rect 17862 19252 17868 19264
rect 17920 19252 17926 19304
rect 17954 19252 17960 19304
rect 18012 19292 18018 19304
rect 18233 19295 18291 19301
rect 18233 19292 18245 19295
rect 18012 19264 18245 19292
rect 18012 19252 18018 19264
rect 18233 19261 18245 19264
rect 18279 19261 18291 19295
rect 18233 19255 18291 19261
rect 18322 19252 18328 19304
rect 18380 19292 18386 19304
rect 18693 19295 18751 19301
rect 18693 19292 18705 19295
rect 18380 19264 18705 19292
rect 18380 19252 18386 19264
rect 18693 19261 18705 19264
rect 18739 19261 18751 19295
rect 18966 19292 18972 19304
rect 18927 19264 18972 19292
rect 18693 19255 18751 19261
rect 18966 19252 18972 19264
rect 19024 19252 19030 19304
rect 16301 19159 16359 19165
rect 16301 19125 16313 19159
rect 16347 19125 16359 19159
rect 16301 19119 16359 19125
rect 19153 19159 19211 19165
rect 19153 19125 19165 19159
rect 19199 19156 19211 19159
rect 19334 19156 19340 19168
rect 19199 19128 19340 19156
rect 19199 19125 19211 19128
rect 19153 19119 19211 19125
rect 19334 19116 19340 19128
rect 19392 19116 19398 19168
rect 19904 19165 19932 19332
rect 21358 19292 21364 19304
rect 21271 19264 21364 19292
rect 21358 19252 21364 19264
rect 21416 19292 21422 19304
rect 22278 19292 22284 19304
rect 21416 19264 22284 19292
rect 21416 19252 21422 19264
rect 22278 19252 22284 19264
rect 22336 19252 22342 19304
rect 20533 19227 20591 19233
rect 20533 19193 20545 19227
rect 20579 19224 20591 19227
rect 20714 19224 20720 19236
rect 20579 19196 20720 19224
rect 20579 19193 20591 19196
rect 20533 19187 20591 19193
rect 20714 19184 20720 19196
rect 20772 19184 20778 19236
rect 19889 19159 19947 19165
rect 19889 19125 19901 19159
rect 19935 19156 19947 19159
rect 20806 19156 20812 19168
rect 19935 19128 20812 19156
rect 19935 19125 19947 19128
rect 19889 19119 19947 19125
rect 20806 19116 20812 19128
rect 20864 19116 20870 19168
rect 1104 19066 21896 19088
rect 1104 19014 7912 19066
rect 7964 19014 7976 19066
rect 8028 19014 8040 19066
rect 8092 19014 8104 19066
rect 8156 19014 14843 19066
rect 14895 19014 14907 19066
rect 14959 19014 14971 19066
rect 15023 19014 15035 19066
rect 15087 19014 21896 19066
rect 1104 18992 21896 19014
rect 2225 18955 2283 18961
rect 2225 18921 2237 18955
rect 2271 18952 2283 18955
rect 2866 18952 2872 18964
rect 2271 18924 2872 18952
rect 2271 18921 2283 18924
rect 2225 18915 2283 18921
rect 2866 18912 2872 18924
rect 2924 18912 2930 18964
rect 4065 18955 4123 18961
rect 4065 18921 4077 18955
rect 4111 18921 4123 18955
rect 4065 18915 4123 18921
rect 2317 18887 2375 18893
rect 2317 18853 2329 18887
rect 2363 18884 2375 18887
rect 4080 18884 4108 18915
rect 4522 18912 4528 18964
rect 4580 18952 4586 18964
rect 5902 18952 5908 18964
rect 4580 18924 5908 18952
rect 4580 18912 4586 18924
rect 5902 18912 5908 18924
rect 5960 18912 5966 18964
rect 6086 18912 6092 18964
rect 6144 18952 6150 18964
rect 6365 18955 6423 18961
rect 6365 18952 6377 18955
rect 6144 18924 6377 18952
rect 6144 18912 6150 18924
rect 6365 18921 6377 18924
rect 6411 18921 6423 18955
rect 6365 18915 6423 18921
rect 6730 18912 6736 18964
rect 6788 18952 6794 18964
rect 6825 18955 6883 18961
rect 6825 18952 6837 18955
rect 6788 18924 6837 18952
rect 6788 18912 6794 18924
rect 6825 18921 6837 18924
rect 6871 18921 6883 18955
rect 7742 18952 7748 18964
rect 7703 18924 7748 18952
rect 6825 18915 6883 18921
rect 7742 18912 7748 18924
rect 7800 18912 7806 18964
rect 9309 18955 9367 18961
rect 9309 18921 9321 18955
rect 9355 18952 9367 18955
rect 9950 18952 9956 18964
rect 9355 18924 9956 18952
rect 9355 18921 9367 18924
rect 9309 18915 9367 18921
rect 9950 18912 9956 18924
rect 10008 18912 10014 18964
rect 11146 18952 11152 18964
rect 10244 18924 11152 18952
rect 5994 18884 6000 18896
rect 2363 18856 4108 18884
rect 4724 18856 6000 18884
rect 2363 18853 2375 18856
rect 2317 18847 2375 18853
rect 1578 18816 1584 18828
rect 1539 18788 1584 18816
rect 1578 18776 1584 18788
rect 1636 18776 1642 18828
rect 1765 18819 1823 18825
rect 1765 18785 1777 18819
rect 1811 18816 1823 18819
rect 2130 18816 2136 18828
rect 1811 18788 2136 18816
rect 1811 18785 1823 18788
rect 1765 18779 1823 18785
rect 2130 18776 2136 18788
rect 2188 18776 2194 18828
rect 2869 18819 2927 18825
rect 2869 18785 2881 18819
rect 2915 18785 2927 18819
rect 2869 18779 2927 18785
rect 3329 18819 3387 18825
rect 3329 18785 3341 18819
rect 3375 18816 3387 18819
rect 4062 18816 4068 18828
rect 3375 18788 4068 18816
rect 3375 18785 3387 18788
rect 3329 18779 3387 18785
rect 2884 18748 2912 18779
rect 4062 18776 4068 18788
rect 4120 18776 4126 18828
rect 4246 18816 4252 18828
rect 4207 18788 4252 18816
rect 4246 18776 4252 18788
rect 4304 18776 4310 18828
rect 4724 18825 4752 18856
rect 5994 18844 6000 18856
rect 6052 18844 6058 18896
rect 7098 18884 7104 18896
rect 6472 18856 7104 18884
rect 4709 18819 4767 18825
rect 4709 18785 4721 18819
rect 4755 18785 4767 18819
rect 4709 18779 4767 18785
rect 4985 18819 5043 18825
rect 4985 18785 4997 18819
rect 5031 18816 5043 18819
rect 5074 18816 5080 18828
rect 5031 18788 5080 18816
rect 5031 18785 5043 18788
rect 4985 18779 5043 18785
rect 5074 18776 5080 18788
rect 5132 18776 5138 18828
rect 5258 18825 5264 18828
rect 5252 18816 5264 18825
rect 5219 18788 5264 18816
rect 5252 18779 5264 18788
rect 5258 18776 5264 18779
rect 5316 18776 5322 18828
rect 5718 18776 5724 18828
rect 5776 18816 5782 18828
rect 6472 18816 6500 18856
rect 7098 18844 7104 18856
rect 7156 18844 7162 18896
rect 7558 18844 7564 18896
rect 7616 18884 7622 18896
rect 10244 18884 10272 18924
rect 11146 18912 11152 18924
rect 11204 18912 11210 18964
rect 12158 18912 12164 18964
rect 12216 18912 12222 18964
rect 12434 18912 12440 18964
rect 12492 18952 12498 18964
rect 12529 18955 12587 18961
rect 12529 18952 12541 18955
rect 12492 18924 12541 18952
rect 12492 18912 12498 18924
rect 12529 18921 12541 18924
rect 12575 18921 12587 18955
rect 12529 18915 12587 18921
rect 13173 18955 13231 18961
rect 13173 18921 13185 18955
rect 13219 18952 13231 18955
rect 13262 18952 13268 18964
rect 13219 18924 13268 18952
rect 13219 18921 13231 18924
rect 13173 18915 13231 18921
rect 13262 18912 13268 18924
rect 13320 18912 13326 18964
rect 13998 18952 14004 18964
rect 13959 18924 14004 18952
rect 13998 18912 14004 18924
rect 14056 18912 14062 18964
rect 14274 18912 14280 18964
rect 14332 18952 14338 18964
rect 15013 18955 15071 18961
rect 15013 18952 15025 18955
rect 14332 18924 15025 18952
rect 14332 18912 14338 18924
rect 15013 18921 15025 18924
rect 15059 18921 15071 18955
rect 17862 18952 17868 18964
rect 17823 18924 17868 18952
rect 15013 18915 15071 18921
rect 17862 18912 17868 18924
rect 17920 18912 17926 18964
rect 18322 18952 18328 18964
rect 18283 18924 18328 18952
rect 18322 18912 18328 18924
rect 18380 18912 18386 18964
rect 21358 18952 21364 18964
rect 21319 18924 21364 18952
rect 21358 18912 21364 18924
rect 21416 18912 21422 18964
rect 7616 18856 10272 18884
rect 7616 18844 7622 18856
rect 10318 18844 10324 18896
rect 10376 18884 10382 18896
rect 11425 18887 11483 18893
rect 11425 18884 11437 18887
rect 10376 18856 11437 18884
rect 10376 18844 10382 18856
rect 6638 18816 6644 18828
rect 5776 18788 6500 18816
rect 6599 18788 6644 18816
rect 5776 18776 5782 18788
rect 6638 18776 6644 18788
rect 6696 18776 6702 18828
rect 7837 18819 7895 18825
rect 7392 18788 7788 18816
rect 2884 18720 4936 18748
rect 2314 18640 2320 18692
rect 2372 18680 2378 18692
rect 4525 18683 4583 18689
rect 4525 18680 4537 18683
rect 2372 18652 4537 18680
rect 2372 18640 2378 18652
rect 4525 18649 4537 18652
rect 4571 18649 4583 18683
rect 4525 18643 4583 18649
rect 2682 18612 2688 18624
rect 2643 18584 2688 18612
rect 2682 18572 2688 18584
rect 2740 18572 2746 18624
rect 2958 18572 2964 18624
rect 3016 18612 3022 18624
rect 3145 18615 3203 18621
rect 3145 18612 3157 18615
rect 3016 18584 3157 18612
rect 3016 18572 3022 18584
rect 3145 18581 3157 18584
rect 3191 18581 3203 18615
rect 4908 18612 4936 18720
rect 6178 18708 6184 18760
rect 6236 18748 6242 18760
rect 7392 18748 7420 18788
rect 6236 18720 7420 18748
rect 6236 18708 6242 18720
rect 7466 18708 7472 18760
rect 7524 18748 7530 18760
rect 7561 18751 7619 18757
rect 7561 18748 7573 18751
rect 7524 18720 7573 18748
rect 7524 18708 7530 18720
rect 7561 18717 7573 18720
rect 7607 18717 7619 18751
rect 7760 18748 7788 18788
rect 7837 18785 7849 18819
rect 7883 18816 7895 18819
rect 8481 18819 8539 18825
rect 8481 18816 8493 18819
rect 7883 18788 8493 18816
rect 7883 18785 7895 18788
rect 7837 18779 7895 18785
rect 8481 18785 8493 18788
rect 8527 18785 8539 18819
rect 8481 18779 8539 18785
rect 9306 18776 9312 18828
rect 9364 18816 9370 18828
rect 10134 18816 10140 18828
rect 9364 18788 10140 18816
rect 9364 18776 9370 18788
rect 10134 18776 10140 18788
rect 10192 18776 10198 18828
rect 10433 18819 10491 18825
rect 10433 18785 10445 18819
rect 10479 18816 10491 18819
rect 10594 18816 10600 18828
rect 10479 18788 10600 18816
rect 10479 18785 10491 18788
rect 10433 18779 10491 18785
rect 10594 18776 10600 18788
rect 10652 18776 10658 18828
rect 11164 18825 11192 18856
rect 11425 18853 11437 18856
rect 11471 18853 11483 18887
rect 12176 18884 12204 18912
rect 13449 18887 13507 18893
rect 13449 18884 13461 18887
rect 12176 18856 13461 18884
rect 11425 18847 11483 18853
rect 13449 18853 13461 18856
rect 13495 18884 13507 18887
rect 13538 18884 13544 18896
rect 13495 18856 13544 18884
rect 13495 18853 13507 18856
rect 13449 18847 13507 18853
rect 13538 18844 13544 18856
rect 13596 18844 13602 18896
rect 16298 18884 16304 18896
rect 14936 18856 16304 18884
rect 11149 18819 11207 18825
rect 11149 18785 11161 18819
rect 11195 18785 11207 18819
rect 12158 18816 12164 18828
rect 12119 18788 12164 18816
rect 11149 18779 11207 18785
rect 12158 18776 12164 18788
rect 12216 18776 12222 18828
rect 12986 18816 12992 18828
rect 12947 18788 12992 18816
rect 12986 18776 12992 18788
rect 13044 18776 13050 18828
rect 13814 18816 13820 18828
rect 13775 18788 13820 18816
rect 13814 18776 13820 18788
rect 13872 18776 13878 18828
rect 8662 18748 8668 18760
rect 7760 18720 8668 18748
rect 7561 18711 7619 18717
rect 8662 18708 8668 18720
rect 8720 18708 8726 18760
rect 10689 18751 10747 18757
rect 10689 18717 10701 18751
rect 10735 18748 10747 18751
rect 11330 18748 11336 18760
rect 10735 18720 11336 18748
rect 10735 18717 10747 18720
rect 10689 18711 10747 18717
rect 8846 18680 8852 18692
rect 7033 18652 8852 18680
rect 7033 18612 7061 18652
rect 8846 18640 8852 18652
rect 8904 18640 8910 18692
rect 4908 18584 7061 18612
rect 3145 18575 3203 18581
rect 8018 18572 8024 18624
rect 8076 18612 8082 18624
rect 8205 18615 8263 18621
rect 8205 18612 8217 18615
rect 8076 18584 8217 18612
rect 8076 18572 8082 18584
rect 8205 18581 8217 18584
rect 8251 18581 8263 18615
rect 8205 18575 8263 18581
rect 9214 18572 9220 18624
rect 9272 18612 9278 18624
rect 10704 18612 10732 18711
rect 11330 18708 11336 18720
rect 11388 18708 11394 18760
rect 11974 18748 11980 18760
rect 11935 18720 11980 18748
rect 11974 18708 11980 18720
rect 12032 18708 12038 18760
rect 12069 18751 12127 18757
rect 12069 18717 12081 18751
rect 12115 18748 12127 18751
rect 12710 18748 12716 18760
rect 12115 18720 12716 18748
rect 12115 18717 12127 18720
rect 12069 18711 12127 18717
rect 12710 18708 12716 18720
rect 12768 18708 12774 18760
rect 14366 18748 14372 18760
rect 14327 18720 14372 18748
rect 14366 18708 14372 18720
rect 14424 18708 14430 18760
rect 14936 18757 14964 18856
rect 16298 18844 16304 18856
rect 16356 18884 16362 18896
rect 17138 18887 17196 18893
rect 17138 18884 17150 18887
rect 16356 18856 17150 18884
rect 16356 18844 16362 18856
rect 17138 18853 17150 18856
rect 17184 18853 17196 18887
rect 17138 18847 17196 18853
rect 15105 18819 15163 18825
rect 15105 18785 15117 18819
rect 15151 18816 15163 18819
rect 16390 18816 16396 18828
rect 15151 18788 16396 18816
rect 15151 18785 15163 18788
rect 15105 18779 15163 18785
rect 16390 18776 16396 18788
rect 16448 18776 16454 18828
rect 16758 18776 16764 18828
rect 16816 18816 16822 18828
rect 17405 18819 17463 18825
rect 17405 18816 17417 18819
rect 16816 18788 17417 18816
rect 16816 18776 16822 18788
rect 17405 18785 17417 18788
rect 17451 18785 17463 18819
rect 17678 18816 17684 18828
rect 17639 18788 17684 18816
rect 17405 18779 17463 18785
rect 17678 18776 17684 18788
rect 17736 18776 17742 18828
rect 18141 18819 18199 18825
rect 18141 18785 18153 18819
rect 18187 18816 18199 18819
rect 18598 18816 18604 18828
rect 18187 18788 18604 18816
rect 18187 18785 18199 18788
rect 18141 18779 18199 18785
rect 18598 18776 18604 18788
rect 18656 18776 18662 18828
rect 18782 18816 18788 18828
rect 18743 18788 18788 18816
rect 18782 18776 18788 18788
rect 18840 18776 18846 18828
rect 14921 18751 14979 18757
rect 14921 18717 14933 18751
rect 14967 18717 14979 18751
rect 14921 18711 14979 18717
rect 17494 18708 17500 18760
rect 17552 18748 17558 18760
rect 21174 18748 21180 18760
rect 17552 18720 21180 18748
rect 17552 18708 17558 18720
rect 21174 18708 21180 18720
rect 21232 18708 21238 18760
rect 12250 18640 12256 18692
rect 12308 18680 12314 18692
rect 14734 18680 14740 18692
rect 12308 18652 14740 18680
rect 12308 18640 12314 18652
rect 14734 18640 14740 18652
rect 14792 18640 14798 18692
rect 18138 18640 18144 18692
rect 18196 18680 18202 18692
rect 18601 18683 18659 18689
rect 18601 18680 18613 18683
rect 18196 18652 18613 18680
rect 18196 18640 18202 18652
rect 18601 18649 18613 18652
rect 18647 18649 18659 18683
rect 18601 18643 18659 18649
rect 10962 18612 10968 18624
rect 9272 18584 10732 18612
rect 10923 18584 10968 18612
rect 9272 18572 9278 18584
rect 10962 18572 10968 18584
rect 11020 18572 11026 18624
rect 11698 18572 11704 18624
rect 11756 18612 11762 18624
rect 13354 18612 13360 18624
rect 11756 18584 13360 18612
rect 11756 18572 11762 18584
rect 13354 18572 13360 18584
rect 13412 18572 13418 18624
rect 15473 18615 15531 18621
rect 15473 18581 15485 18615
rect 15519 18612 15531 18615
rect 15838 18612 15844 18624
rect 15519 18584 15844 18612
rect 15519 18581 15531 18584
rect 15473 18575 15531 18581
rect 15838 18572 15844 18584
rect 15896 18572 15902 18624
rect 16022 18612 16028 18624
rect 15983 18584 16028 18612
rect 16022 18572 16028 18584
rect 16080 18572 16086 18624
rect 19150 18612 19156 18624
rect 19063 18584 19156 18612
rect 19150 18572 19156 18584
rect 19208 18612 19214 18624
rect 20530 18612 20536 18624
rect 19208 18584 20536 18612
rect 19208 18572 19214 18584
rect 20530 18572 20536 18584
rect 20588 18572 20594 18624
rect 1104 18522 21896 18544
rect 1104 18470 4447 18522
rect 4499 18470 4511 18522
rect 4563 18470 4575 18522
rect 4627 18470 4639 18522
rect 4691 18470 11378 18522
rect 11430 18470 11442 18522
rect 11494 18470 11506 18522
rect 11558 18470 11570 18522
rect 11622 18470 18308 18522
rect 18360 18470 18372 18522
rect 18424 18470 18436 18522
rect 18488 18470 18500 18522
rect 18552 18470 21896 18522
rect 1104 18448 21896 18470
rect 1670 18408 1676 18420
rect 1631 18380 1676 18408
rect 1670 18368 1676 18380
rect 1728 18368 1734 18420
rect 2225 18411 2283 18417
rect 2225 18377 2237 18411
rect 2271 18408 2283 18411
rect 3050 18408 3056 18420
rect 2271 18380 3056 18408
rect 2271 18377 2283 18380
rect 2225 18371 2283 18377
rect 3050 18368 3056 18380
rect 3108 18368 3114 18420
rect 4890 18368 4896 18420
rect 4948 18408 4954 18420
rect 6362 18408 6368 18420
rect 4948 18380 6368 18408
rect 4948 18368 4954 18380
rect 6362 18368 6368 18380
rect 6420 18368 6426 18420
rect 6638 18368 6644 18420
rect 6696 18408 6702 18420
rect 8297 18411 8355 18417
rect 8297 18408 8309 18411
rect 6696 18380 8309 18408
rect 6696 18368 6702 18380
rect 8297 18377 8309 18380
rect 8343 18377 8355 18411
rect 8846 18408 8852 18420
rect 8807 18380 8852 18408
rect 8297 18371 8355 18377
rect 8846 18368 8852 18380
rect 8904 18368 8910 18420
rect 11698 18408 11704 18420
rect 8956 18380 11704 18408
rect 4062 18300 4068 18352
rect 4120 18340 4126 18352
rect 7837 18343 7895 18349
rect 7837 18340 7849 18343
rect 4120 18312 7849 18340
rect 4120 18300 4126 18312
rect 7837 18309 7849 18312
rect 7883 18309 7895 18343
rect 7837 18303 7895 18309
rect 4798 18232 4804 18284
rect 4856 18272 4862 18284
rect 5258 18272 5264 18284
rect 4856 18244 5264 18272
rect 4856 18232 4862 18244
rect 5258 18232 5264 18244
rect 5316 18272 5322 18284
rect 5353 18275 5411 18281
rect 5353 18272 5365 18275
rect 5316 18244 5365 18272
rect 5316 18232 5322 18244
rect 5353 18241 5365 18244
rect 5399 18241 5411 18275
rect 5353 18235 5411 18241
rect 5442 18232 5448 18284
rect 5500 18272 5506 18284
rect 6457 18275 6515 18281
rect 6457 18272 6469 18275
rect 5500 18244 6469 18272
rect 5500 18232 5506 18244
rect 6457 18241 6469 18244
rect 6503 18272 6515 18275
rect 6822 18272 6828 18284
rect 6503 18244 6828 18272
rect 6503 18241 6515 18244
rect 6457 18235 6515 18241
rect 6822 18232 6828 18244
rect 6880 18232 6886 18284
rect 7374 18272 7380 18284
rect 7335 18244 7380 18272
rect 7374 18232 7380 18244
rect 7432 18232 7438 18284
rect 8956 18272 8984 18380
rect 11698 18368 11704 18380
rect 11756 18368 11762 18420
rect 12710 18368 12716 18420
rect 12768 18408 12774 18420
rect 12897 18411 12955 18417
rect 12897 18408 12909 18411
rect 12768 18380 12909 18408
rect 12768 18368 12774 18380
rect 12897 18377 12909 18380
rect 12943 18377 12955 18411
rect 12897 18371 12955 18377
rect 13814 18368 13820 18420
rect 13872 18408 13878 18420
rect 15749 18411 15807 18417
rect 15749 18408 15761 18411
rect 13872 18380 15761 18408
rect 13872 18368 13878 18380
rect 15749 18377 15761 18380
rect 15795 18377 15807 18411
rect 17310 18408 17316 18420
rect 17271 18380 17316 18408
rect 15749 18371 15807 18377
rect 17310 18368 17316 18380
rect 17368 18368 17374 18420
rect 17954 18408 17960 18420
rect 17915 18380 17960 18408
rect 17954 18368 17960 18380
rect 18012 18368 18018 18420
rect 12802 18340 12808 18352
rect 12084 18312 12808 18340
rect 9766 18272 9772 18284
rect 7484 18244 8984 18272
rect 9727 18244 9772 18272
rect 2314 18204 2320 18216
rect 2275 18176 2320 18204
rect 2314 18164 2320 18176
rect 2372 18164 2378 18216
rect 3142 18213 3148 18216
rect 2869 18207 2927 18213
rect 2869 18173 2881 18207
rect 2915 18173 2927 18207
rect 2869 18167 2927 18173
rect 3136 18167 3148 18213
rect 3200 18204 3206 18216
rect 3200 18176 3236 18204
rect 1765 18139 1823 18145
rect 1765 18105 1777 18139
rect 1811 18136 1823 18139
rect 2498 18136 2504 18148
rect 1811 18108 2504 18136
rect 1811 18105 1823 18108
rect 1765 18099 1823 18105
rect 2498 18096 2504 18108
rect 2556 18096 2562 18148
rect 2884 18136 2912 18167
rect 3142 18164 3148 18167
rect 3200 18164 3206 18176
rect 3602 18164 3608 18216
rect 3660 18204 3666 18216
rect 7484 18204 7512 18244
rect 9766 18232 9772 18244
rect 9824 18232 9830 18284
rect 9953 18275 10011 18281
rect 9953 18241 9965 18275
rect 9999 18272 10011 18275
rect 11054 18272 11060 18284
rect 9999 18244 11060 18272
rect 9999 18241 10011 18244
rect 9953 18235 10011 18241
rect 11054 18232 11060 18244
rect 11112 18232 11118 18284
rect 12084 18281 12112 18312
rect 12802 18300 12808 18312
rect 12860 18340 12866 18352
rect 14093 18343 14151 18349
rect 14093 18340 14105 18343
rect 12860 18312 14105 18340
rect 12860 18300 12866 18312
rect 14093 18309 14105 18312
rect 14139 18309 14151 18343
rect 14093 18303 14151 18309
rect 15657 18343 15715 18349
rect 15657 18309 15669 18343
rect 15703 18340 15715 18343
rect 17494 18340 17500 18352
rect 15703 18312 17500 18340
rect 15703 18309 15715 18312
rect 15657 18303 15715 18309
rect 17494 18300 17500 18312
rect 17552 18300 17558 18352
rect 18046 18300 18052 18352
rect 18104 18340 18110 18352
rect 18693 18343 18751 18349
rect 18693 18340 18705 18343
rect 18104 18312 18705 18340
rect 18104 18300 18110 18312
rect 18693 18309 18705 18312
rect 18739 18309 18751 18343
rect 18693 18303 18751 18309
rect 12069 18275 12127 18281
rect 12069 18241 12081 18275
rect 12115 18241 12127 18275
rect 12069 18235 12127 18241
rect 12710 18232 12716 18284
rect 12768 18272 12774 18284
rect 13449 18275 13507 18281
rect 13449 18272 13461 18275
rect 12768 18244 13461 18272
rect 12768 18232 12774 18244
rect 13449 18241 13461 18244
rect 13495 18241 13507 18275
rect 16022 18272 16028 18284
rect 13449 18235 13507 18241
rect 15396 18244 16028 18272
rect 8018 18204 8024 18216
rect 3660 18176 7512 18204
rect 7979 18176 8024 18204
rect 3660 18164 3666 18176
rect 8018 18164 8024 18176
rect 8076 18164 8082 18216
rect 8481 18207 8539 18213
rect 8481 18173 8493 18207
rect 8527 18173 8539 18207
rect 8481 18167 8539 18173
rect 9033 18207 9091 18213
rect 9033 18173 9045 18207
rect 9079 18204 9091 18207
rect 9674 18204 9680 18216
rect 9079 18176 9352 18204
rect 9635 18176 9680 18204
rect 9079 18173 9091 18176
rect 9033 18167 9091 18173
rect 3878 18136 3884 18148
rect 2884 18108 3884 18136
rect 3878 18096 3884 18108
rect 3936 18096 3942 18148
rect 4890 18136 4896 18148
rect 4080 18108 4896 18136
rect 1946 18028 1952 18080
rect 2004 18068 2010 18080
rect 4080 18068 4108 18108
rect 4890 18096 4896 18108
rect 4948 18096 4954 18148
rect 5169 18139 5227 18145
rect 5169 18105 5181 18139
rect 5215 18136 5227 18139
rect 5813 18139 5871 18145
rect 5813 18136 5825 18139
rect 5215 18108 5825 18136
rect 5215 18105 5227 18108
rect 5169 18099 5227 18105
rect 5813 18105 5825 18108
rect 5859 18105 5871 18139
rect 8496 18136 8524 18167
rect 5813 18099 5871 18105
rect 5920 18108 8524 18136
rect 2004 18040 4108 18068
rect 2004 18028 2010 18040
rect 4154 18028 4160 18080
rect 4212 18068 4218 18080
rect 4249 18071 4307 18077
rect 4249 18068 4261 18071
rect 4212 18040 4261 18068
rect 4212 18028 4218 18040
rect 4249 18037 4261 18040
rect 4295 18037 4307 18071
rect 4249 18031 4307 18037
rect 4801 18071 4859 18077
rect 4801 18037 4813 18071
rect 4847 18068 4859 18071
rect 4982 18068 4988 18080
rect 4847 18040 4988 18068
rect 4847 18037 4859 18040
rect 4801 18031 4859 18037
rect 4982 18028 4988 18040
rect 5040 18028 5046 18080
rect 5258 18028 5264 18080
rect 5316 18068 5322 18080
rect 5316 18040 5361 18068
rect 5316 18028 5322 18040
rect 5534 18028 5540 18080
rect 5592 18068 5598 18080
rect 5920 18068 5948 18108
rect 5592 18040 5948 18068
rect 5592 18028 5598 18040
rect 6270 18028 6276 18080
rect 6328 18068 6334 18080
rect 6825 18071 6883 18077
rect 6825 18068 6837 18071
rect 6328 18040 6837 18068
rect 6328 18028 6334 18040
rect 6825 18037 6837 18040
rect 6871 18037 6883 18071
rect 7190 18068 7196 18080
rect 7151 18040 7196 18068
rect 6825 18031 6883 18037
rect 7190 18028 7196 18040
rect 7248 18028 7254 18080
rect 7282 18028 7288 18080
rect 7340 18068 7346 18080
rect 9324 18077 9352 18176
rect 9674 18164 9680 18176
rect 9732 18164 9738 18216
rect 9858 18164 9864 18216
rect 9916 18204 9922 18216
rect 10505 18207 10563 18213
rect 10505 18204 10517 18207
rect 9916 18176 10517 18204
rect 9916 18164 9922 18176
rect 10505 18173 10517 18176
rect 10551 18173 10563 18207
rect 10505 18167 10563 18173
rect 10520 18136 10548 18167
rect 10778 18164 10784 18216
rect 10836 18204 10842 18216
rect 10965 18207 11023 18213
rect 10965 18204 10977 18207
rect 10836 18176 10977 18204
rect 10836 18164 10842 18176
rect 10965 18173 10977 18176
rect 11011 18204 11023 18207
rect 11698 18204 11704 18216
rect 11011 18176 11704 18204
rect 11011 18173 11023 18176
rect 10965 18167 11023 18173
rect 11698 18164 11704 18176
rect 11756 18164 11762 18216
rect 12894 18164 12900 18216
rect 12952 18204 12958 18216
rect 13998 18204 14004 18216
rect 12952 18176 14004 18204
rect 12952 18164 12958 18176
rect 13998 18164 14004 18176
rect 14056 18164 14062 18216
rect 15217 18207 15275 18213
rect 15217 18173 15229 18207
rect 15263 18204 15275 18207
rect 15396 18204 15424 18244
rect 16022 18232 16028 18244
rect 16080 18272 16086 18284
rect 16301 18275 16359 18281
rect 16301 18272 16313 18275
rect 16080 18244 16313 18272
rect 16080 18232 16086 18244
rect 16301 18241 16313 18244
rect 16347 18241 16359 18275
rect 16301 18235 16359 18241
rect 16666 18232 16672 18284
rect 16724 18272 16730 18284
rect 16724 18244 18276 18272
rect 16724 18232 16730 18244
rect 15263 18176 15424 18204
rect 15473 18207 15531 18213
rect 15263 18173 15275 18176
rect 15217 18167 15275 18173
rect 15473 18173 15485 18207
rect 15519 18173 15531 18207
rect 15473 18167 15531 18173
rect 11241 18139 11299 18145
rect 11241 18136 11253 18139
rect 10520 18108 11253 18136
rect 11241 18105 11253 18108
rect 11287 18105 11299 18139
rect 11241 18099 11299 18105
rect 12161 18139 12219 18145
rect 12161 18105 12173 18139
rect 12207 18136 12219 18139
rect 15488 18136 15516 18167
rect 15838 18164 15844 18216
rect 15896 18204 15902 18216
rect 16117 18207 16175 18213
rect 16117 18204 16129 18207
rect 15896 18176 16129 18204
rect 15896 18164 15902 18176
rect 16117 18173 16129 18176
rect 16163 18173 16175 18207
rect 17126 18204 17132 18216
rect 17087 18176 17132 18204
rect 16117 18167 16175 18173
rect 17126 18164 17132 18176
rect 17184 18164 17190 18216
rect 17773 18207 17831 18213
rect 17773 18173 17785 18207
rect 17819 18204 17831 18207
rect 18138 18204 18144 18216
rect 17819 18176 18144 18204
rect 17819 18173 17831 18176
rect 17773 18167 17831 18173
rect 18138 18164 18144 18176
rect 18196 18164 18202 18216
rect 18248 18213 18276 18244
rect 18233 18207 18291 18213
rect 18233 18173 18245 18207
rect 18279 18173 18291 18207
rect 18233 18167 18291 18173
rect 16758 18136 16764 18148
rect 12207 18108 13584 18136
rect 15488 18108 16764 18136
rect 12207 18105 12219 18108
rect 12161 18099 12219 18105
rect 9309 18071 9367 18077
rect 7340 18040 7385 18068
rect 7340 18028 7346 18040
rect 9309 18037 9321 18071
rect 9355 18037 9367 18071
rect 10318 18068 10324 18080
rect 10279 18040 10324 18068
rect 9309 18031 9367 18037
rect 10318 18028 10324 18040
rect 10376 18028 10382 18080
rect 10778 18068 10784 18080
rect 10739 18040 10784 18068
rect 10778 18028 10784 18040
rect 10836 18028 10842 18080
rect 11054 18028 11060 18080
rect 11112 18068 11118 18080
rect 12253 18071 12311 18077
rect 12253 18068 12265 18071
rect 11112 18040 12265 18068
rect 11112 18028 11118 18040
rect 12253 18037 12265 18040
rect 12299 18037 12311 18071
rect 12253 18031 12311 18037
rect 12434 18028 12440 18080
rect 12492 18068 12498 18080
rect 12621 18071 12679 18077
rect 12621 18068 12633 18071
rect 12492 18040 12633 18068
rect 12492 18028 12498 18040
rect 12621 18037 12633 18040
rect 12667 18037 12679 18071
rect 13262 18068 13268 18080
rect 13223 18040 13268 18068
rect 12621 18031 12679 18037
rect 13262 18028 13268 18040
rect 13320 18028 13326 18080
rect 13354 18028 13360 18080
rect 13412 18068 13418 18080
rect 13556 18068 13584 18108
rect 16758 18096 16764 18108
rect 16816 18136 16822 18148
rect 16816 18108 18460 18136
rect 16816 18096 16822 18108
rect 15657 18071 15715 18077
rect 15657 18068 15669 18071
rect 13412 18040 13457 18068
rect 13556 18040 15669 18068
rect 13412 18028 13418 18040
rect 15657 18037 15669 18040
rect 15703 18037 15715 18071
rect 15657 18031 15715 18037
rect 16206 18028 16212 18080
rect 16264 18068 16270 18080
rect 18432 18077 18460 18108
rect 18417 18071 18475 18077
rect 16264 18040 16309 18068
rect 16264 18028 16270 18040
rect 18417 18037 18429 18071
rect 18463 18037 18475 18071
rect 18417 18031 18475 18037
rect 1104 17978 21896 18000
rect 1104 17926 7912 17978
rect 7964 17926 7976 17978
rect 8028 17926 8040 17978
rect 8092 17926 8104 17978
rect 8156 17926 14843 17978
rect 14895 17926 14907 17978
rect 14959 17926 14971 17978
rect 15023 17926 15035 17978
rect 15087 17926 21896 17978
rect 1104 17904 21896 17926
rect 4065 17867 4123 17873
rect 4065 17864 4077 17867
rect 1780 17836 4077 17864
rect 1780 17805 1808 17836
rect 4065 17833 4077 17836
rect 4111 17833 4123 17867
rect 4798 17864 4804 17876
rect 4759 17836 4804 17864
rect 4065 17827 4123 17833
rect 4798 17824 4804 17836
rect 4856 17824 4862 17876
rect 4890 17824 4896 17876
rect 4948 17864 4954 17876
rect 7558 17864 7564 17876
rect 4948 17836 7564 17864
rect 4948 17824 4954 17836
rect 7558 17824 7564 17836
rect 7616 17824 7622 17876
rect 9585 17867 9643 17873
rect 9585 17833 9597 17867
rect 9631 17864 9643 17867
rect 10318 17864 10324 17876
rect 9631 17836 10324 17864
rect 9631 17833 9643 17836
rect 9585 17827 9643 17833
rect 10318 17824 10324 17836
rect 10376 17824 10382 17876
rect 10502 17824 10508 17876
rect 10560 17864 10566 17876
rect 13817 17867 13875 17873
rect 13817 17864 13829 17867
rect 10560 17836 13829 17864
rect 10560 17824 10566 17836
rect 13817 17833 13829 17836
rect 13863 17833 13875 17867
rect 13817 17827 13875 17833
rect 14734 17824 14740 17876
rect 14792 17864 14798 17876
rect 15105 17867 15163 17873
rect 15105 17864 15117 17867
rect 14792 17836 15117 17864
rect 14792 17824 14798 17836
rect 15105 17833 15117 17836
rect 15151 17864 15163 17867
rect 15378 17864 15384 17876
rect 15151 17836 15384 17864
rect 15151 17833 15163 17836
rect 15105 17827 15163 17833
rect 15378 17824 15384 17836
rect 15436 17824 15442 17876
rect 15565 17867 15623 17873
rect 15565 17833 15577 17867
rect 15611 17864 15623 17867
rect 16301 17867 16359 17873
rect 16301 17864 16313 17867
rect 15611 17836 16313 17864
rect 15611 17833 15623 17836
rect 15565 17827 15623 17833
rect 16301 17833 16313 17836
rect 16347 17833 16359 17867
rect 16301 17827 16359 17833
rect 16390 17824 16396 17876
rect 16448 17864 16454 17876
rect 16853 17867 16911 17873
rect 16853 17864 16865 17867
rect 16448 17836 16865 17864
rect 16448 17824 16454 17836
rect 16853 17833 16865 17836
rect 16899 17833 16911 17867
rect 16853 17827 16911 17833
rect 1765 17799 1823 17805
rect 1765 17765 1777 17799
rect 1811 17765 1823 17799
rect 1765 17759 1823 17765
rect 2317 17799 2375 17805
rect 2317 17765 2329 17799
rect 2363 17796 2375 17799
rect 2682 17796 2688 17808
rect 2363 17768 2688 17796
rect 2363 17765 2375 17768
rect 2317 17759 2375 17765
rect 2682 17756 2688 17768
rect 2740 17756 2746 17808
rect 2866 17756 2872 17808
rect 2924 17756 2930 17808
rect 3605 17799 3663 17805
rect 3605 17765 3617 17799
rect 3651 17796 3663 17799
rect 5534 17796 5540 17808
rect 3651 17768 5540 17796
rect 3651 17765 3663 17768
rect 3605 17759 3663 17765
rect 5534 17756 5540 17768
rect 5592 17756 5598 17808
rect 5626 17756 5632 17808
rect 5684 17796 5690 17808
rect 5994 17805 6000 17808
rect 5936 17799 6000 17805
rect 5936 17796 5948 17799
rect 5684 17768 5948 17796
rect 5684 17756 5690 17768
rect 5936 17765 5948 17768
rect 5982 17765 6000 17799
rect 5936 17759 6000 17765
rect 5994 17756 6000 17759
rect 6052 17756 6058 17808
rect 6454 17756 6460 17808
rect 6512 17796 6518 17808
rect 7466 17805 7472 17808
rect 7460 17796 7472 17805
rect 6512 17768 6684 17796
rect 7427 17768 7472 17796
rect 6512 17756 6518 17768
rect 1581 17731 1639 17737
rect 1581 17697 1593 17731
rect 1627 17728 1639 17731
rect 2884 17728 2912 17756
rect 3142 17728 3148 17740
rect 1627 17700 2912 17728
rect 3103 17700 3148 17728
rect 1627 17697 1639 17700
rect 1581 17691 1639 17697
rect 3142 17688 3148 17700
rect 3200 17688 3206 17740
rect 6656 17737 6684 17768
rect 7460 17759 7472 17768
rect 7466 17756 7472 17759
rect 7524 17756 7530 17808
rect 17957 17799 18015 17805
rect 17957 17796 17969 17799
rect 7576 17768 17969 17796
rect 4249 17731 4307 17737
rect 4249 17697 4261 17731
rect 4295 17728 4307 17731
rect 6273 17731 6331 17737
rect 6273 17728 6285 17731
rect 4295 17700 6285 17728
rect 4295 17697 4307 17700
rect 4249 17691 4307 17697
rect 6273 17697 6285 17700
rect 6319 17697 6331 17731
rect 6273 17691 6331 17697
rect 6641 17731 6699 17737
rect 6641 17697 6653 17731
rect 6687 17697 6699 17731
rect 6641 17691 6699 17697
rect 7101 17731 7159 17737
rect 7101 17697 7113 17731
rect 7147 17728 7159 17731
rect 7576 17728 7604 17768
rect 17957 17765 17969 17768
rect 18003 17796 18015 17799
rect 19061 17799 19119 17805
rect 19061 17796 19073 17799
rect 18003 17768 19073 17796
rect 18003 17765 18015 17768
rect 17957 17759 18015 17765
rect 19061 17765 19073 17768
rect 19107 17765 19119 17799
rect 19061 17759 19119 17765
rect 7147 17700 7604 17728
rect 9677 17731 9735 17737
rect 7147 17697 7159 17700
rect 7101 17691 7159 17697
rect 9677 17697 9689 17731
rect 9723 17728 9735 17731
rect 9858 17728 9864 17740
rect 9723 17700 9864 17728
rect 9723 17697 9735 17700
rect 9677 17691 9735 17697
rect 9858 17688 9864 17700
rect 9916 17688 9922 17740
rect 10134 17688 10140 17740
rect 10192 17728 10198 17740
rect 10318 17728 10324 17740
rect 10192 17700 10324 17728
rect 10192 17688 10198 17700
rect 10318 17688 10324 17700
rect 10376 17728 10382 17740
rect 10505 17731 10563 17737
rect 10505 17728 10517 17731
rect 10376 17700 10517 17728
rect 10376 17688 10382 17700
rect 10505 17697 10517 17700
rect 10551 17697 10563 17731
rect 10505 17691 10563 17697
rect 10965 17731 11023 17737
rect 10965 17697 10977 17731
rect 11011 17697 11023 17731
rect 10965 17691 11023 17697
rect 2866 17660 2872 17672
rect 2827 17632 2872 17660
rect 2866 17620 2872 17632
rect 2924 17620 2930 17672
rect 3053 17663 3111 17669
rect 3053 17629 3065 17663
rect 3099 17660 3111 17663
rect 4338 17660 4344 17672
rect 3099 17632 4344 17660
rect 3099 17629 3111 17632
rect 3053 17623 3111 17629
rect 4338 17620 4344 17632
rect 4396 17620 4402 17672
rect 6178 17660 6184 17672
rect 6139 17632 6184 17660
rect 6178 17620 6184 17632
rect 6236 17660 6242 17672
rect 7193 17663 7251 17669
rect 7193 17660 7205 17663
rect 6236 17632 7205 17660
rect 6236 17620 6242 17632
rect 7193 17629 7205 17632
rect 7239 17629 7251 17663
rect 7193 17623 7251 17629
rect 9493 17663 9551 17669
rect 9493 17629 9505 17663
rect 9539 17660 9551 17663
rect 10042 17660 10048 17672
rect 9539 17632 10048 17660
rect 9539 17629 9551 17632
rect 9493 17623 9551 17629
rect 10042 17620 10048 17632
rect 10100 17620 10106 17672
rect 10980 17660 11008 17691
rect 11238 17688 11244 17740
rect 11296 17728 11302 17740
rect 11425 17731 11483 17737
rect 11425 17728 11437 17731
rect 11296 17700 11437 17728
rect 11296 17688 11302 17700
rect 11425 17697 11437 17700
rect 11471 17697 11483 17731
rect 11425 17691 11483 17697
rect 12802 17688 12808 17740
rect 12860 17737 12866 17740
rect 12860 17728 12872 17737
rect 13538 17728 13544 17740
rect 12860 17700 12905 17728
rect 13499 17700 13544 17728
rect 12860 17691 12872 17700
rect 12860 17688 12866 17691
rect 13538 17688 13544 17700
rect 13596 17688 13602 17740
rect 13998 17728 14004 17740
rect 13959 17700 14004 17728
rect 13998 17688 14004 17700
rect 14056 17688 14062 17740
rect 15197 17731 15255 17737
rect 15197 17697 15209 17731
rect 15243 17728 15255 17731
rect 15286 17728 15292 17740
rect 15243 17700 15292 17728
rect 15243 17697 15255 17700
rect 15197 17691 15255 17697
rect 15286 17688 15292 17700
rect 15344 17688 15350 17740
rect 15746 17688 15752 17740
rect 15804 17728 15810 17740
rect 16209 17731 16267 17737
rect 16209 17728 16221 17731
rect 15804 17700 16221 17728
rect 15804 17688 15810 17700
rect 16209 17697 16221 17700
rect 16255 17697 16267 17731
rect 17865 17731 17923 17737
rect 17865 17728 17877 17731
rect 16209 17691 16267 17697
rect 16500 17700 17877 17728
rect 11330 17660 11336 17672
rect 10980 17632 11336 17660
rect 11330 17620 11336 17632
rect 11388 17620 11394 17672
rect 13081 17663 13139 17669
rect 13081 17629 13093 17663
rect 13127 17660 13139 17663
rect 14366 17660 14372 17672
rect 13127 17632 14372 17660
rect 13127 17629 13139 17632
rect 13081 17623 13139 17629
rect 14366 17620 14372 17632
rect 14424 17620 14430 17672
rect 15013 17663 15071 17669
rect 15013 17629 15025 17663
rect 15059 17629 15071 17663
rect 15013 17623 15071 17629
rect 2682 17552 2688 17604
rect 2740 17592 2746 17604
rect 6273 17595 6331 17601
rect 2740 17564 5304 17592
rect 2740 17552 2746 17564
rect 2222 17524 2228 17536
rect 2183 17496 2228 17524
rect 2222 17484 2228 17496
rect 2280 17484 2286 17536
rect 3513 17527 3571 17533
rect 3513 17493 3525 17527
rect 3559 17524 3571 17527
rect 3605 17527 3663 17533
rect 3605 17524 3617 17527
rect 3559 17496 3617 17524
rect 3559 17493 3571 17496
rect 3513 17487 3571 17493
rect 3605 17493 3617 17496
rect 3651 17493 3663 17527
rect 5276 17524 5304 17564
rect 6273 17561 6285 17595
rect 6319 17592 6331 17595
rect 6457 17595 6515 17601
rect 6457 17592 6469 17595
rect 6319 17564 6469 17592
rect 6319 17561 6331 17564
rect 6273 17555 6331 17561
rect 6457 17561 6469 17564
rect 6503 17561 6515 17595
rect 6457 17555 6515 17561
rect 9030 17552 9036 17604
rect 9088 17592 9094 17604
rect 9088 17564 10456 17592
rect 9088 17552 9094 17564
rect 7101 17527 7159 17533
rect 7101 17524 7113 17527
rect 5276 17496 7113 17524
rect 3605 17487 3663 17493
rect 7101 17493 7113 17496
rect 7147 17493 7159 17527
rect 7101 17487 7159 17493
rect 8110 17484 8116 17536
rect 8168 17524 8174 17536
rect 8573 17527 8631 17533
rect 8573 17524 8585 17527
rect 8168 17496 8585 17524
rect 8168 17484 8174 17496
rect 8573 17493 8585 17496
rect 8619 17493 8631 17527
rect 8573 17487 8631 17493
rect 9766 17484 9772 17536
rect 9824 17524 9830 17536
rect 10045 17527 10103 17533
rect 10045 17524 10057 17527
rect 9824 17496 10057 17524
rect 9824 17484 9830 17496
rect 10045 17493 10057 17496
rect 10091 17493 10103 17527
rect 10045 17487 10103 17493
rect 10134 17484 10140 17536
rect 10192 17524 10198 17536
rect 10321 17527 10379 17533
rect 10321 17524 10333 17527
rect 10192 17496 10333 17524
rect 10192 17484 10198 17496
rect 10321 17493 10333 17496
rect 10367 17493 10379 17527
rect 10428 17524 10456 17564
rect 10502 17552 10508 17604
rect 10560 17592 10566 17604
rect 11241 17595 11299 17601
rect 11241 17592 11253 17595
rect 10560 17564 11253 17592
rect 10560 17552 10566 17564
rect 11241 17561 11253 17564
rect 11287 17561 11299 17595
rect 15028 17592 15056 17623
rect 16298 17620 16304 17672
rect 16356 17660 16362 17672
rect 16393 17663 16451 17669
rect 16393 17660 16405 17663
rect 16356 17632 16405 17660
rect 16356 17620 16362 17632
rect 16393 17629 16405 17632
rect 16439 17629 16451 17663
rect 16393 17623 16451 17629
rect 15194 17592 15200 17604
rect 15028 17564 15200 17592
rect 11241 17555 11299 17561
rect 15194 17552 15200 17564
rect 15252 17552 15258 17604
rect 15841 17595 15899 17601
rect 15841 17561 15853 17595
rect 15887 17592 15899 17595
rect 16206 17592 16212 17604
rect 15887 17564 16212 17592
rect 15887 17561 15899 17564
rect 15841 17555 15899 17561
rect 16206 17552 16212 17564
rect 16264 17552 16270 17604
rect 10781 17527 10839 17533
rect 10781 17524 10793 17527
rect 10428 17496 10793 17524
rect 10321 17487 10379 17493
rect 10781 17493 10793 17496
rect 10827 17493 10839 17527
rect 10781 17487 10839 17493
rect 11701 17527 11759 17533
rect 11701 17493 11713 17527
rect 11747 17524 11759 17527
rect 12710 17524 12716 17536
rect 11747 17496 12716 17524
rect 11747 17493 11759 17496
rect 11701 17487 11759 17493
rect 12710 17484 12716 17496
rect 12768 17484 12774 17536
rect 13357 17527 13415 17533
rect 13357 17493 13369 17527
rect 13403 17524 13415 17527
rect 13538 17524 13544 17536
rect 13403 17496 13544 17524
rect 13403 17493 13415 17496
rect 13357 17487 13415 17493
rect 13538 17484 13544 17496
rect 13596 17484 13602 17536
rect 13630 17484 13636 17536
rect 13688 17524 13694 17536
rect 14369 17527 14427 17533
rect 14369 17524 14381 17527
rect 13688 17496 14381 17524
rect 13688 17484 13694 17496
rect 14369 17493 14381 17496
rect 14415 17493 14427 17527
rect 14369 17487 14427 17493
rect 14458 17484 14464 17536
rect 14516 17524 14522 17536
rect 16500 17524 16528 17700
rect 17865 17697 17877 17700
rect 17911 17697 17923 17731
rect 17865 17691 17923 17697
rect 17773 17663 17831 17669
rect 17773 17629 17785 17663
rect 17819 17629 17831 17663
rect 17773 17623 17831 17629
rect 18785 17663 18843 17669
rect 18785 17629 18797 17663
rect 18831 17660 18843 17663
rect 19886 17660 19892 17672
rect 18831 17632 19892 17660
rect 18831 17629 18843 17632
rect 18785 17623 18843 17629
rect 17788 17592 17816 17623
rect 19886 17620 19892 17632
rect 19944 17620 19950 17672
rect 17954 17592 17960 17604
rect 17788 17564 17960 17592
rect 17954 17552 17960 17564
rect 18012 17552 18018 17604
rect 14516 17496 16528 17524
rect 18325 17527 18383 17533
rect 14516 17484 14522 17496
rect 18325 17493 18337 17527
rect 18371 17524 18383 17527
rect 18966 17524 18972 17536
rect 18371 17496 18972 17524
rect 18371 17493 18383 17496
rect 18325 17487 18383 17493
rect 18966 17484 18972 17496
rect 19024 17484 19030 17536
rect 1104 17434 21896 17456
rect 1104 17382 4447 17434
rect 4499 17382 4511 17434
rect 4563 17382 4575 17434
rect 4627 17382 4639 17434
rect 4691 17382 11378 17434
rect 11430 17382 11442 17434
rect 11494 17382 11506 17434
rect 11558 17382 11570 17434
rect 11622 17382 18308 17434
rect 18360 17382 18372 17434
rect 18424 17382 18436 17434
rect 18488 17382 18500 17434
rect 18552 17382 21896 17434
rect 1104 17360 21896 17382
rect 2225 17323 2283 17329
rect 2225 17289 2237 17323
rect 2271 17320 2283 17323
rect 2774 17320 2780 17332
rect 2271 17292 2780 17320
rect 2271 17289 2283 17292
rect 2225 17283 2283 17289
rect 2774 17280 2780 17292
rect 2832 17280 2838 17332
rect 4338 17320 4344 17332
rect 4299 17292 4344 17320
rect 4338 17280 4344 17292
rect 4396 17280 4402 17332
rect 5258 17280 5264 17332
rect 5316 17320 5322 17332
rect 5353 17323 5411 17329
rect 5353 17320 5365 17323
rect 5316 17292 5365 17320
rect 5316 17280 5322 17292
rect 5353 17289 5365 17292
rect 5399 17289 5411 17323
rect 5353 17283 5411 17289
rect 6362 17280 6368 17332
rect 6420 17320 6426 17332
rect 6457 17323 6515 17329
rect 6457 17320 6469 17323
rect 6420 17292 6469 17320
rect 6420 17280 6426 17292
rect 6457 17289 6469 17292
rect 6503 17289 6515 17323
rect 6457 17283 6515 17289
rect 7009 17323 7067 17329
rect 7009 17289 7021 17323
rect 7055 17320 7067 17323
rect 7374 17320 7380 17332
rect 7055 17292 7380 17320
rect 7055 17289 7067 17292
rect 7009 17283 7067 17289
rect 7374 17280 7380 17292
rect 7432 17280 7438 17332
rect 7484 17292 8432 17320
rect 5442 17212 5448 17264
rect 5500 17252 5506 17264
rect 7484 17252 7512 17292
rect 5500 17224 7512 17252
rect 8404 17252 8432 17292
rect 8570 17280 8576 17332
rect 8628 17320 8634 17332
rect 10594 17320 10600 17332
rect 8628 17292 10180 17320
rect 10555 17292 10600 17320
rect 8628 17280 8634 17292
rect 9122 17252 9128 17264
rect 8404 17224 9128 17252
rect 5500 17212 5506 17224
rect 9122 17212 9128 17224
rect 9180 17212 9186 17264
rect 10152 17252 10180 17292
rect 10594 17280 10600 17292
rect 10652 17280 10658 17332
rect 11698 17320 11704 17332
rect 11659 17292 11704 17320
rect 11698 17280 11704 17292
rect 11756 17280 11762 17332
rect 12250 17280 12256 17332
rect 12308 17320 12314 17332
rect 12434 17320 12440 17332
rect 12308 17292 12440 17320
rect 12308 17280 12314 17292
rect 12434 17280 12440 17292
rect 12492 17280 12498 17332
rect 12618 17280 12624 17332
rect 12676 17320 12682 17332
rect 13170 17320 13176 17332
rect 12676 17292 13176 17320
rect 12676 17280 12682 17292
rect 13170 17280 13176 17292
rect 13228 17280 13234 17332
rect 13354 17280 13360 17332
rect 13412 17320 13418 17332
rect 13541 17323 13599 17329
rect 13541 17320 13553 17323
rect 13412 17292 13553 17320
rect 13412 17280 13418 17292
rect 13541 17289 13553 17292
rect 13587 17289 13599 17323
rect 13541 17283 13599 17289
rect 13998 17280 14004 17332
rect 14056 17320 14062 17332
rect 14185 17323 14243 17329
rect 14185 17320 14197 17323
rect 14056 17292 14197 17320
rect 14056 17280 14062 17292
rect 14185 17289 14197 17292
rect 14231 17289 14243 17323
rect 14185 17283 14243 17289
rect 16209 17323 16267 17329
rect 16209 17289 16221 17323
rect 16255 17320 16267 17323
rect 16298 17320 16304 17332
rect 16255 17292 16304 17320
rect 16255 17289 16267 17292
rect 16209 17283 16267 17289
rect 16298 17280 16304 17292
rect 16356 17280 16362 17332
rect 18138 17280 18144 17332
rect 18196 17320 18202 17332
rect 19521 17323 19579 17329
rect 19521 17320 19533 17323
rect 18196 17292 19533 17320
rect 18196 17280 18202 17292
rect 19521 17289 19533 17292
rect 19567 17289 19579 17323
rect 19521 17283 19579 17289
rect 10873 17255 10931 17261
rect 10873 17252 10885 17255
rect 10152 17224 10885 17252
rect 10873 17221 10885 17224
rect 10919 17221 10931 17255
rect 10873 17215 10931 17221
rect 11238 17212 11244 17264
rect 11296 17252 11302 17264
rect 13817 17255 13875 17261
rect 13817 17252 13829 17255
rect 11296 17224 13829 17252
rect 11296 17212 11302 17224
rect 13817 17221 13829 17224
rect 13863 17221 13875 17255
rect 13817 17215 13875 17221
rect 19245 17255 19303 17261
rect 19245 17221 19257 17255
rect 19291 17252 19303 17255
rect 19334 17252 19340 17264
rect 19291 17224 19340 17252
rect 19291 17221 19303 17224
rect 19245 17215 19303 17221
rect 19334 17212 19340 17224
rect 19392 17252 19398 17264
rect 19392 17224 20116 17252
rect 19392 17212 19398 17224
rect 4154 17144 4160 17196
rect 4212 17184 4218 17196
rect 4893 17187 4951 17193
rect 4893 17184 4905 17187
rect 4212 17156 4905 17184
rect 4212 17144 4218 17156
rect 4893 17153 4905 17156
rect 4939 17153 4951 17187
rect 4893 17147 4951 17153
rect 5626 17144 5632 17196
rect 5684 17184 5690 17196
rect 5905 17187 5963 17193
rect 5905 17184 5917 17187
rect 5684 17156 5917 17184
rect 5684 17144 5690 17156
rect 5905 17153 5917 17156
rect 5951 17153 5963 17187
rect 5905 17147 5963 17153
rect 11882 17144 11888 17196
rect 11940 17184 11946 17196
rect 12434 17184 12440 17196
rect 11940 17156 12440 17184
rect 11940 17144 11946 17156
rect 12434 17144 12440 17156
rect 12492 17144 12498 17196
rect 12802 17144 12808 17196
rect 12860 17184 12866 17196
rect 12897 17187 12955 17193
rect 12897 17184 12909 17187
rect 12860 17156 12909 17184
rect 12860 17144 12866 17156
rect 12897 17153 12909 17156
rect 12943 17153 12955 17187
rect 12897 17147 12955 17153
rect 13078 17144 13084 17196
rect 13136 17184 13142 17196
rect 13136 17156 13181 17184
rect 13136 17144 13142 17156
rect 18966 17144 18972 17196
rect 19024 17184 19030 17196
rect 20088 17193 20116 17224
rect 19981 17187 20039 17193
rect 19981 17184 19993 17187
rect 19024 17156 19993 17184
rect 19024 17144 19030 17156
rect 19981 17153 19993 17156
rect 20027 17153 20039 17187
rect 19981 17147 20039 17153
rect 20073 17187 20131 17193
rect 20073 17153 20085 17187
rect 20119 17153 20131 17187
rect 20073 17147 20131 17153
rect 2317 17119 2375 17125
rect 2317 17085 2329 17119
rect 2363 17116 2375 17119
rect 2958 17116 2964 17128
rect 2363 17088 2964 17116
rect 2363 17085 2375 17088
rect 2317 17079 2375 17085
rect 2958 17076 2964 17088
rect 3016 17076 3022 17128
rect 4062 17116 4068 17128
rect 4023 17088 4068 17116
rect 4062 17076 4068 17088
rect 4120 17076 4126 17128
rect 5813 17119 5871 17125
rect 5813 17085 5825 17119
rect 5859 17116 5871 17119
rect 7742 17116 7748 17128
rect 5859 17088 7748 17116
rect 5859 17085 5871 17088
rect 5813 17079 5871 17085
rect 7742 17076 7748 17088
rect 7800 17076 7806 17128
rect 8110 17076 8116 17128
rect 8168 17125 8174 17128
rect 8168 17116 8180 17125
rect 8389 17119 8447 17125
rect 8168 17088 8213 17116
rect 8168 17079 8180 17088
rect 8389 17085 8401 17119
rect 8435 17116 8447 17119
rect 9214 17116 9220 17128
rect 8435 17088 9220 17116
rect 8435 17085 8447 17088
rect 8389 17079 8447 17085
rect 8168 17076 8174 17079
rect 9214 17076 9220 17088
rect 9272 17116 9278 17128
rect 11057 17119 11115 17125
rect 9272 17088 10364 17116
rect 9272 17076 9278 17088
rect 1578 17048 1584 17060
rect 1539 17020 1584 17048
rect 1578 17008 1584 17020
rect 1636 17008 1642 17060
rect 1762 17048 1768 17060
rect 1723 17020 1768 17048
rect 1762 17008 1768 17020
rect 1820 17008 1826 17060
rect 3820 17051 3878 17057
rect 3820 17017 3832 17051
rect 3866 17048 3878 17051
rect 4154 17048 4160 17060
rect 3866 17020 4160 17048
rect 3866 17017 3878 17020
rect 3820 17011 3878 17017
rect 4154 17008 4160 17020
rect 4212 17008 4218 17060
rect 4801 17051 4859 17057
rect 4801 17017 4813 17051
rect 4847 17048 4859 17051
rect 6178 17048 6184 17060
rect 4847 17020 6184 17048
rect 4847 17017 4859 17020
rect 4801 17011 4859 17017
rect 6178 17008 6184 17020
rect 6236 17008 6242 17060
rect 9484 17051 9542 17057
rect 9484 17017 9496 17051
rect 9530 17048 9542 17051
rect 10042 17048 10048 17060
rect 9530 17020 10048 17048
rect 9530 17017 9542 17020
rect 9484 17011 9542 17017
rect 10042 17008 10048 17020
rect 10100 17008 10106 17060
rect 2685 16983 2743 16989
rect 2685 16949 2697 16983
rect 2731 16980 2743 16983
rect 2866 16980 2872 16992
rect 2731 16952 2872 16980
rect 2731 16949 2743 16952
rect 2685 16943 2743 16949
rect 2866 16940 2872 16952
rect 2924 16940 2930 16992
rect 3326 16940 3332 16992
rect 3384 16980 3390 16992
rect 4709 16983 4767 16989
rect 4709 16980 4721 16983
rect 3384 16952 4721 16980
rect 3384 16940 3390 16952
rect 4709 16949 4721 16952
rect 4755 16980 4767 16983
rect 5626 16980 5632 16992
rect 4755 16952 5632 16980
rect 4755 16949 4767 16952
rect 4709 16943 4767 16949
rect 5626 16940 5632 16952
rect 5684 16940 5690 16992
rect 5721 16983 5779 16989
rect 5721 16949 5733 16983
rect 5767 16980 5779 16983
rect 6362 16980 6368 16992
rect 5767 16952 6368 16980
rect 5767 16949 5779 16952
rect 5721 16943 5779 16949
rect 6362 16940 6368 16952
rect 6420 16940 6426 16992
rect 8941 16983 8999 16989
rect 8941 16949 8953 16983
rect 8987 16980 8999 16983
rect 9674 16980 9680 16992
rect 8987 16952 9680 16980
rect 8987 16949 8999 16952
rect 8941 16943 8999 16949
rect 9674 16940 9680 16952
rect 9732 16940 9738 16992
rect 10336 16980 10364 17088
rect 11057 17085 11069 17119
rect 11103 17116 11115 17119
rect 11146 17116 11152 17128
rect 11103 17088 11152 17116
rect 11103 17085 11115 17088
rect 11057 17079 11115 17085
rect 11146 17076 11152 17088
rect 11204 17076 11210 17128
rect 14366 17076 14372 17128
rect 14424 17116 14430 17128
rect 14829 17119 14887 17125
rect 14829 17116 14841 17119
rect 14424 17088 14841 17116
rect 14424 17076 14430 17088
rect 14829 17085 14841 17088
rect 14875 17085 14887 17119
rect 14829 17079 14887 17085
rect 15378 17076 15384 17128
rect 15436 17116 15442 17128
rect 16485 17119 16543 17125
rect 16485 17116 16497 17119
rect 15436 17088 16497 17116
rect 15436 17076 15442 17088
rect 16485 17085 16497 17088
rect 16531 17085 16543 17119
rect 16485 17079 16543 17085
rect 17770 17076 17776 17128
rect 17828 17116 17834 17128
rect 17865 17119 17923 17125
rect 17865 17116 17877 17119
rect 17828 17088 17877 17116
rect 17828 17076 17834 17088
rect 17865 17085 17877 17088
rect 17911 17085 17923 17119
rect 19886 17116 19892 17128
rect 19847 17088 19892 17116
rect 17865 17079 17923 17085
rect 19886 17076 19892 17088
rect 19944 17076 19950 17128
rect 10410 17008 10416 17060
rect 10468 17048 10474 17060
rect 13906 17048 13912 17060
rect 10468 17020 12940 17048
rect 10468 17008 10474 17020
rect 11882 16980 11888 16992
rect 10336 16952 11888 16980
rect 11882 16940 11888 16952
rect 11940 16940 11946 16992
rect 12342 16980 12348 16992
rect 12303 16952 12348 16980
rect 12342 16940 12348 16952
rect 12400 16940 12406 16992
rect 12912 16980 12940 17020
rect 13096 17020 13912 17048
rect 13096 16980 13124 17020
rect 13906 17008 13912 17020
rect 13964 17008 13970 17060
rect 15096 17051 15154 17057
rect 15096 17017 15108 17051
rect 15142 17048 15154 17051
rect 15194 17048 15200 17060
rect 15142 17020 15200 17048
rect 15142 17017 15154 17020
rect 15096 17011 15154 17017
rect 15194 17008 15200 17020
rect 15252 17008 15258 17060
rect 15286 17008 15292 17060
rect 15344 17048 15350 17060
rect 15470 17048 15476 17060
rect 15344 17020 15476 17048
rect 15344 17008 15350 17020
rect 15470 17008 15476 17020
rect 15528 17048 15534 17060
rect 15528 17020 17448 17048
rect 15528 17008 15534 17020
rect 12912 16952 13124 16980
rect 13173 16983 13231 16989
rect 13173 16949 13185 16983
rect 13219 16980 13231 16983
rect 13446 16980 13452 16992
rect 13219 16952 13452 16980
rect 13219 16949 13231 16952
rect 13173 16943 13231 16949
rect 13446 16940 13452 16952
rect 13504 16940 13510 16992
rect 17310 16980 17316 16992
rect 17271 16952 17316 16980
rect 17310 16940 17316 16952
rect 17368 16940 17374 16992
rect 17420 16980 17448 17020
rect 17954 17008 17960 17060
rect 18012 17048 18018 17060
rect 18132 17051 18190 17057
rect 18132 17048 18144 17051
rect 18012 17020 18144 17048
rect 18012 17008 18018 17020
rect 18132 17017 18144 17020
rect 18178 17048 18190 17051
rect 19150 17048 19156 17060
rect 18178 17020 19156 17048
rect 18178 17017 18190 17020
rect 18132 17011 18190 17017
rect 19150 17008 19156 17020
rect 19208 17008 19214 17060
rect 18046 16980 18052 16992
rect 17420 16952 18052 16980
rect 18046 16940 18052 16952
rect 18104 16940 18110 16992
rect 1104 16890 21896 16912
rect 1104 16838 7912 16890
rect 7964 16838 7976 16890
rect 8028 16838 8040 16890
rect 8092 16838 8104 16890
rect 8156 16838 14843 16890
rect 14895 16838 14907 16890
rect 14959 16838 14971 16890
rect 15023 16838 15035 16890
rect 15087 16838 21896 16890
rect 1104 16816 21896 16838
rect 1762 16736 1768 16788
rect 1820 16776 1826 16788
rect 2133 16779 2191 16785
rect 2133 16776 2145 16779
rect 1820 16748 2145 16776
rect 1820 16736 1826 16748
rect 2133 16745 2145 16748
rect 2179 16745 2191 16779
rect 2133 16739 2191 16745
rect 2498 16736 2504 16788
rect 2556 16776 2562 16788
rect 2593 16779 2651 16785
rect 2593 16776 2605 16779
rect 2556 16748 2605 16776
rect 2556 16736 2562 16748
rect 2593 16745 2605 16748
rect 2639 16745 2651 16779
rect 3142 16776 3148 16788
rect 3103 16748 3148 16776
rect 2593 16739 2651 16745
rect 3142 16736 3148 16748
rect 3200 16736 3206 16788
rect 4246 16776 4252 16788
rect 4207 16748 4252 16776
rect 4246 16736 4252 16748
rect 4304 16736 4310 16788
rect 4890 16736 4896 16788
rect 4948 16776 4954 16788
rect 5721 16779 5779 16785
rect 5721 16776 5733 16779
rect 4948 16748 5733 16776
rect 4948 16736 4954 16748
rect 5721 16745 5733 16748
rect 5767 16745 5779 16779
rect 5902 16776 5908 16788
rect 5721 16739 5779 16745
rect 5828 16748 5908 16776
rect 3050 16708 3056 16720
rect 2332 16680 3056 16708
rect 1578 16640 1584 16652
rect 1539 16612 1584 16640
rect 1578 16600 1584 16612
rect 1636 16600 1642 16652
rect 1762 16640 1768 16652
rect 1723 16612 1768 16640
rect 1762 16600 1768 16612
rect 1820 16600 1826 16652
rect 2332 16649 2360 16680
rect 3050 16668 3056 16680
rect 3108 16668 3114 16720
rect 5077 16711 5135 16717
rect 5077 16677 5089 16711
rect 5123 16708 5135 16711
rect 5534 16708 5540 16720
rect 5123 16680 5540 16708
rect 5123 16677 5135 16680
rect 5077 16671 5135 16677
rect 5534 16668 5540 16680
rect 5592 16668 5598 16720
rect 2317 16643 2375 16649
rect 2317 16609 2329 16643
rect 2363 16609 2375 16643
rect 2317 16603 2375 16609
rect 2777 16643 2835 16649
rect 2777 16609 2789 16643
rect 2823 16640 2835 16643
rect 3510 16640 3516 16652
rect 2823 16612 3516 16640
rect 2823 16609 2835 16612
rect 2777 16603 2835 16609
rect 3510 16600 3516 16612
rect 3568 16600 3574 16652
rect 4065 16643 4123 16649
rect 4065 16609 4077 16643
rect 4111 16640 4123 16643
rect 4982 16640 4988 16652
rect 4111 16612 4988 16640
rect 4111 16609 4123 16612
rect 4065 16603 4123 16609
rect 4982 16600 4988 16612
rect 5040 16600 5046 16652
rect 5166 16640 5172 16652
rect 5127 16612 5172 16640
rect 5166 16600 5172 16612
rect 5224 16600 5230 16652
rect 5828 16640 5856 16748
rect 5902 16736 5908 16748
rect 5960 16776 5966 16788
rect 6641 16779 6699 16785
rect 6641 16776 6653 16779
rect 5960 16748 6653 16776
rect 5960 16736 5966 16748
rect 6641 16745 6653 16748
rect 6687 16745 6699 16779
rect 7190 16776 7196 16788
rect 7151 16748 7196 16776
rect 6641 16739 6699 16745
rect 7190 16736 7196 16748
rect 7248 16736 7254 16788
rect 7282 16736 7288 16788
rect 7340 16776 7346 16788
rect 7469 16779 7527 16785
rect 7469 16776 7481 16779
rect 7340 16748 7481 16776
rect 7340 16736 7346 16748
rect 7469 16745 7481 16748
rect 7515 16745 7527 16779
rect 7469 16739 7527 16745
rect 7742 16736 7748 16788
rect 7800 16776 7806 16788
rect 8481 16779 8539 16785
rect 8481 16776 8493 16779
rect 7800 16748 8493 16776
rect 7800 16736 7806 16748
rect 8481 16745 8493 16748
rect 8527 16745 8539 16779
rect 8481 16739 8539 16745
rect 9309 16779 9367 16785
rect 9309 16745 9321 16779
rect 9355 16745 9367 16779
rect 9674 16776 9680 16788
rect 9635 16748 9680 16776
rect 9309 16739 9367 16745
rect 9324 16708 9352 16739
rect 9674 16736 9680 16748
rect 9732 16736 9738 16788
rect 9766 16736 9772 16788
rect 9824 16776 9830 16788
rect 9824 16748 9869 16776
rect 10152 16748 11652 16776
rect 9824 16736 9830 16748
rect 6196 16680 9352 16708
rect 5913 16643 5971 16649
rect 5913 16640 5925 16643
rect 5828 16612 5925 16640
rect 5913 16609 5925 16612
rect 5959 16609 5971 16643
rect 6196 16640 6224 16680
rect 5913 16603 5971 16609
rect 6012 16612 6224 16640
rect 6365 16643 6423 16649
rect 5258 16572 5264 16584
rect 5219 16544 5264 16572
rect 5258 16532 5264 16544
rect 5316 16532 5322 16584
rect 5350 16532 5356 16584
rect 5408 16572 5414 16584
rect 6012 16572 6040 16612
rect 6365 16609 6377 16643
rect 6411 16640 6423 16643
rect 6454 16640 6460 16652
rect 6411 16612 6460 16640
rect 6411 16609 6423 16612
rect 6365 16603 6423 16609
rect 6454 16600 6460 16612
rect 6512 16600 6518 16652
rect 6638 16600 6644 16652
rect 6696 16640 6702 16652
rect 7837 16643 7895 16649
rect 7837 16640 7849 16643
rect 6696 16612 7849 16640
rect 6696 16600 6702 16612
rect 7837 16609 7849 16612
rect 7883 16609 7895 16643
rect 7837 16603 7895 16609
rect 7929 16643 7987 16649
rect 7929 16609 7941 16643
rect 7975 16640 7987 16643
rect 8294 16640 8300 16652
rect 7975 16612 8300 16640
rect 7975 16609 7987 16612
rect 7929 16603 7987 16609
rect 5408 16544 6040 16572
rect 5408 16532 5414 16544
rect 2774 16464 2780 16516
rect 2832 16504 2838 16516
rect 7006 16504 7012 16516
rect 2832 16476 7012 16504
rect 2832 16464 2838 16476
rect 7006 16464 7012 16476
rect 7064 16464 7070 16516
rect 7852 16504 7880 16603
rect 8294 16600 8300 16612
rect 8352 16600 8358 16652
rect 8662 16640 8668 16652
rect 8623 16612 8668 16640
rect 8662 16600 8668 16612
rect 8720 16600 8726 16652
rect 10152 16640 10180 16748
rect 10226 16668 10232 16720
rect 10284 16708 10290 16720
rect 11048 16711 11106 16717
rect 10284 16680 10916 16708
rect 10284 16668 10290 16680
rect 8772 16612 10180 16640
rect 8113 16575 8171 16581
rect 8113 16541 8125 16575
rect 8159 16572 8171 16575
rect 8202 16572 8208 16584
rect 8159 16544 8208 16572
rect 8159 16541 8171 16544
rect 8113 16535 8171 16541
rect 8202 16532 8208 16544
rect 8260 16532 8266 16584
rect 8772 16572 8800 16612
rect 10410 16600 10416 16652
rect 10468 16640 10474 16652
rect 10505 16643 10563 16649
rect 10505 16640 10517 16643
rect 10468 16612 10517 16640
rect 10468 16600 10474 16612
rect 10505 16609 10517 16612
rect 10551 16609 10563 16643
rect 10505 16603 10563 16609
rect 10686 16600 10692 16652
rect 10744 16640 10750 16652
rect 10781 16643 10839 16649
rect 10781 16640 10793 16643
rect 10744 16612 10793 16640
rect 10744 16600 10750 16612
rect 10781 16609 10793 16612
rect 10827 16609 10839 16643
rect 10888 16640 10916 16680
rect 11048 16677 11060 16711
rect 11094 16708 11106 16711
rect 11238 16708 11244 16720
rect 11094 16680 11244 16708
rect 11094 16677 11106 16680
rect 11048 16671 11106 16677
rect 11238 16668 11244 16680
rect 11296 16668 11302 16720
rect 11624 16708 11652 16748
rect 13262 16736 13268 16788
rect 13320 16776 13326 16788
rect 13633 16779 13691 16785
rect 13633 16776 13645 16779
rect 13320 16748 13645 16776
rect 13320 16736 13326 16748
rect 13633 16745 13645 16748
rect 13679 16745 13691 16779
rect 13906 16776 13912 16788
rect 13867 16748 13912 16776
rect 13633 16739 13691 16745
rect 13906 16736 13912 16748
rect 13964 16736 13970 16788
rect 15746 16776 15752 16788
rect 15707 16748 15752 16776
rect 15746 16736 15752 16748
rect 15804 16736 15810 16788
rect 17497 16779 17555 16785
rect 17497 16745 17509 16779
rect 17543 16745 17555 16779
rect 19150 16776 19156 16788
rect 19111 16748 19156 16776
rect 17497 16739 17555 16745
rect 14369 16711 14427 16717
rect 14369 16708 14381 16711
rect 11624 16680 14381 16708
rect 14369 16677 14381 16680
rect 14415 16677 14427 16711
rect 14369 16671 14427 16677
rect 15396 16680 17172 16708
rect 12621 16643 12679 16649
rect 12621 16640 12633 16643
rect 10888 16612 12633 16640
rect 10781 16603 10839 16609
rect 12621 16609 12633 16612
rect 12667 16609 12679 16643
rect 13170 16640 13176 16652
rect 13131 16612 13176 16640
rect 12621 16603 12679 16609
rect 13170 16600 13176 16612
rect 13228 16600 13234 16652
rect 13265 16643 13323 16649
rect 13265 16609 13277 16643
rect 13311 16609 13323 16643
rect 13265 16603 13323 16609
rect 8680 16544 8800 16572
rect 9953 16575 10011 16581
rect 8680 16504 8708 16544
rect 9953 16541 9965 16575
rect 9999 16572 10011 16575
rect 10594 16572 10600 16584
rect 9999 16544 10600 16572
rect 9999 16541 10011 16544
rect 9953 16535 10011 16541
rect 10594 16532 10600 16544
rect 10652 16532 10658 16584
rect 12802 16532 12808 16584
rect 12860 16572 12866 16584
rect 12989 16575 13047 16581
rect 12989 16572 13001 16575
rect 12860 16544 13001 16572
rect 12860 16532 12866 16544
rect 12989 16541 13001 16544
rect 13035 16541 13047 16575
rect 13280 16572 13308 16603
rect 13354 16600 13360 16652
rect 13412 16640 13418 16652
rect 15396 16649 15424 16680
rect 15381 16643 15439 16649
rect 15381 16640 15393 16643
rect 13412 16612 15393 16640
rect 13412 16600 13418 16612
rect 15381 16609 15393 16612
rect 15427 16609 15439 16643
rect 15381 16603 15439 16609
rect 15930 16600 15936 16652
rect 15988 16640 15994 16652
rect 16373 16643 16431 16649
rect 16373 16640 16385 16643
rect 15988 16612 16385 16640
rect 15988 16600 15994 16612
rect 16373 16609 16385 16612
rect 16419 16609 16431 16643
rect 17144 16640 17172 16680
rect 17218 16668 17224 16720
rect 17276 16708 17282 16720
rect 17512 16708 17540 16739
rect 19150 16736 19156 16748
rect 19208 16736 19214 16788
rect 18018 16711 18076 16717
rect 18018 16708 18030 16711
rect 17276 16680 18030 16708
rect 17276 16668 17282 16680
rect 18018 16677 18030 16680
rect 18064 16677 18076 16711
rect 18018 16671 18076 16677
rect 18138 16668 18144 16720
rect 18196 16668 18202 16720
rect 18156 16640 18184 16668
rect 19981 16643 20039 16649
rect 19981 16640 19993 16643
rect 17144 16612 19993 16640
rect 16373 16603 16431 16609
rect 19981 16609 19993 16612
rect 20027 16609 20039 16643
rect 19981 16603 20039 16609
rect 14458 16572 14464 16584
rect 13280 16544 14464 16572
rect 12989 16535 13047 16541
rect 14458 16532 14464 16544
rect 14516 16532 14522 16584
rect 15194 16572 15200 16584
rect 15155 16544 15200 16572
rect 15194 16532 15200 16544
rect 15252 16532 15258 16584
rect 15286 16532 15292 16584
rect 15344 16572 15350 16584
rect 16117 16575 16175 16581
rect 15344 16544 15389 16572
rect 15344 16532 15350 16544
rect 16117 16541 16129 16575
rect 16163 16541 16175 16575
rect 17770 16572 17776 16584
rect 16117 16535 16175 16541
rect 17328 16544 17776 16572
rect 7852 16476 8708 16504
rect 11974 16464 11980 16516
rect 12032 16504 12038 16516
rect 12161 16507 12219 16513
rect 12161 16504 12173 16507
rect 12032 16476 12173 16504
rect 12032 16464 12038 16476
rect 12161 16473 12173 16476
rect 12207 16473 12219 16507
rect 12161 16467 12219 16473
rect 4154 16396 4160 16448
rect 4212 16436 4218 16448
rect 4709 16439 4767 16445
rect 4709 16436 4721 16439
rect 4212 16408 4721 16436
rect 4212 16396 4218 16408
rect 4709 16405 4721 16408
rect 4755 16405 4767 16439
rect 6178 16436 6184 16448
rect 6139 16408 6184 16436
rect 4709 16399 4767 16405
rect 6178 16396 6184 16408
rect 6236 16396 6242 16448
rect 10318 16436 10324 16448
rect 10279 16408 10324 16436
rect 10318 16396 10324 16408
rect 10376 16396 10382 16448
rect 11882 16396 11888 16448
rect 11940 16436 11946 16448
rect 12437 16439 12495 16445
rect 12437 16436 12449 16439
rect 11940 16408 12449 16436
rect 11940 16396 11946 16408
rect 12437 16405 12449 16408
rect 12483 16405 12495 16439
rect 12437 16399 12495 16405
rect 12802 16396 12808 16448
rect 12860 16436 12866 16448
rect 15378 16436 15384 16448
rect 12860 16408 15384 16436
rect 12860 16396 12866 16408
rect 15378 16396 15384 16408
rect 15436 16396 15442 16448
rect 16132 16436 16160 16535
rect 16758 16436 16764 16448
rect 16132 16408 16764 16436
rect 16758 16396 16764 16408
rect 16816 16436 16822 16448
rect 17328 16436 17356 16544
rect 17770 16532 17776 16544
rect 17828 16532 17834 16584
rect 16816 16408 17356 16436
rect 16816 16396 16822 16408
rect 17586 16396 17592 16448
rect 17644 16436 17650 16448
rect 19613 16439 19671 16445
rect 19613 16436 19625 16439
rect 17644 16408 19625 16436
rect 17644 16396 17650 16408
rect 19613 16405 19625 16408
rect 19659 16436 19671 16439
rect 19886 16436 19892 16448
rect 19659 16408 19892 16436
rect 19659 16405 19671 16408
rect 19613 16399 19671 16405
rect 19886 16396 19892 16408
rect 19944 16396 19950 16448
rect 1104 16346 21896 16368
rect 1104 16294 4447 16346
rect 4499 16294 4511 16346
rect 4563 16294 4575 16346
rect 4627 16294 4639 16346
rect 4691 16294 11378 16346
rect 11430 16294 11442 16346
rect 11494 16294 11506 16346
rect 11558 16294 11570 16346
rect 11622 16294 18308 16346
rect 18360 16294 18372 16346
rect 18424 16294 18436 16346
rect 18488 16294 18500 16346
rect 18552 16294 21896 16346
rect 1104 16272 21896 16294
rect 1762 16192 1768 16244
rect 1820 16232 1826 16244
rect 2133 16235 2191 16241
rect 2133 16232 2145 16235
rect 1820 16204 2145 16232
rect 1820 16192 1826 16204
rect 2133 16201 2145 16204
rect 2179 16201 2191 16235
rect 2133 16195 2191 16201
rect 2314 16192 2320 16244
rect 2372 16232 2378 16244
rect 2593 16235 2651 16241
rect 2593 16232 2605 16235
rect 2372 16204 2605 16232
rect 2372 16192 2378 16204
rect 2593 16201 2605 16204
rect 2639 16201 2651 16235
rect 3050 16232 3056 16244
rect 3011 16204 3056 16232
rect 2593 16195 2651 16201
rect 3050 16192 3056 16204
rect 3108 16192 3114 16244
rect 3510 16232 3516 16244
rect 3471 16204 3516 16232
rect 3510 16192 3516 16204
rect 3568 16192 3574 16244
rect 4982 16192 4988 16244
rect 5040 16232 5046 16244
rect 5994 16232 6000 16244
rect 5040 16204 5672 16232
rect 5955 16204 6000 16232
rect 5040 16192 5046 16204
rect 3973 16167 4031 16173
rect 3973 16133 3985 16167
rect 4019 16133 4031 16167
rect 5644 16164 5672 16204
rect 5994 16192 6000 16204
rect 6052 16192 6058 16244
rect 6546 16192 6552 16244
rect 6604 16232 6610 16244
rect 7101 16235 7159 16241
rect 7101 16232 7113 16235
rect 6604 16204 7113 16232
rect 6604 16192 6610 16204
rect 7101 16201 7113 16204
rect 7147 16201 7159 16235
rect 10042 16232 10048 16244
rect 10003 16204 10048 16232
rect 7101 16195 7159 16201
rect 10042 16192 10048 16204
rect 10100 16192 10106 16244
rect 11146 16192 11152 16244
rect 11204 16192 11210 16244
rect 11885 16235 11943 16241
rect 11885 16201 11897 16235
rect 11931 16232 11943 16235
rect 12158 16232 12164 16244
rect 11931 16204 12164 16232
rect 11931 16201 11943 16204
rect 11885 16195 11943 16201
rect 12158 16192 12164 16204
rect 12216 16192 12222 16244
rect 15194 16232 15200 16244
rect 13740 16204 14780 16232
rect 15155 16204 15200 16232
rect 6641 16167 6699 16173
rect 6641 16164 6653 16167
rect 5644 16136 6653 16164
rect 3973 16127 4031 16133
rect 6641 16133 6653 16136
rect 6687 16133 6699 16167
rect 11164 16164 11192 16192
rect 13357 16167 13415 16173
rect 13357 16164 13369 16167
rect 11164 16136 13369 16164
rect 6641 16127 6699 16133
rect 13357 16133 13369 16136
rect 13403 16133 13415 16167
rect 13357 16127 13415 16133
rect 1578 16096 1584 16108
rect 1539 16068 1584 16096
rect 1578 16056 1584 16068
rect 1636 16056 1642 16108
rect 3988 16096 4016 16127
rect 8294 16096 8300 16108
rect 2792 16068 4016 16096
rect 8255 16068 8300 16096
rect 2314 16028 2320 16040
rect 2275 16000 2320 16028
rect 2314 15988 2320 16000
rect 2372 15988 2378 16040
rect 2792 16037 2820 16068
rect 8294 16056 8300 16068
rect 8352 16096 8358 16108
rect 8352 16068 8800 16096
rect 8352 16056 8358 16068
rect 2777 16031 2835 16037
rect 2777 15997 2789 16031
rect 2823 15997 2835 16031
rect 2777 15991 2835 15997
rect 3237 16031 3295 16037
rect 3237 15997 3249 16031
rect 3283 15997 3295 16031
rect 3237 15991 3295 15997
rect 3697 16031 3755 16037
rect 3697 15997 3709 16031
rect 3743 16028 3755 16031
rect 3789 16031 3847 16037
rect 3789 16028 3801 16031
rect 3743 16000 3801 16028
rect 3743 15997 3755 16000
rect 3697 15991 3755 15997
rect 3789 15997 3801 16000
rect 3835 15997 3847 16031
rect 4154 16028 4160 16040
rect 4115 16000 4160 16028
rect 3789 15991 3847 15997
rect 1762 15960 1768 15972
rect 1723 15932 1768 15960
rect 1762 15920 1768 15932
rect 1820 15920 1826 15972
rect 3252 15960 3280 15991
rect 4154 15988 4160 16000
rect 4212 15988 4218 16040
rect 4614 16028 4620 16040
rect 4575 16000 4620 16028
rect 4614 15988 4620 16000
rect 4672 15988 4678 16040
rect 4884 16031 4942 16037
rect 4884 15997 4896 16031
rect 4930 16028 4942 16031
rect 5258 16028 5264 16040
rect 4930 16000 5264 16028
rect 4930 15997 4942 16000
rect 4884 15991 4942 15997
rect 5258 15988 5264 16000
rect 5316 15988 5322 16040
rect 6822 16028 6828 16040
rect 6783 16000 6828 16028
rect 6822 15988 6828 16000
rect 6880 15988 6886 16040
rect 7098 15988 7104 16040
rect 7156 16028 7162 16040
rect 7285 16031 7343 16037
rect 7285 16028 7297 16031
rect 7156 16000 7297 16028
rect 7156 15988 7162 16000
rect 7285 15997 7297 16000
rect 7331 15997 7343 16031
rect 7285 15991 7343 15997
rect 8665 16031 8723 16037
rect 8665 15997 8677 16031
rect 8711 15997 8723 16031
rect 8772 16028 8800 16068
rect 10870 16056 10876 16108
rect 10928 16096 10934 16108
rect 11149 16099 11207 16105
rect 11149 16096 11161 16099
rect 10928 16068 11161 16096
rect 10928 16056 10934 16068
rect 11149 16065 11161 16068
rect 11195 16065 11207 16099
rect 11149 16059 11207 16065
rect 11238 16056 11244 16108
rect 11296 16096 11302 16108
rect 12529 16099 12587 16105
rect 12529 16096 12541 16099
rect 11296 16068 12541 16096
rect 11296 16056 11302 16068
rect 12529 16065 12541 16068
rect 12575 16096 12587 16099
rect 12710 16096 12716 16108
rect 12575 16068 12716 16096
rect 12575 16065 12587 16068
rect 12529 16059 12587 16065
rect 12710 16056 12716 16068
rect 12768 16056 12774 16108
rect 8921 16031 8979 16037
rect 8921 16028 8933 16031
rect 8772 16000 8933 16028
rect 8665 15991 8723 15997
rect 8921 15997 8933 16000
rect 8967 15997 8979 16031
rect 8921 15991 8979 15997
rect 5350 15960 5356 15972
rect 3252 15932 5356 15960
rect 5350 15920 5356 15932
rect 5408 15920 5414 15972
rect 8021 15963 8079 15969
rect 8021 15929 8033 15963
rect 8067 15960 8079 15963
rect 8202 15960 8208 15972
rect 8067 15932 8208 15960
rect 8067 15929 8079 15932
rect 8021 15923 8079 15929
rect 8202 15920 8208 15932
rect 8260 15920 8266 15972
rect 8680 15960 8708 15991
rect 10410 15988 10416 16040
rect 10468 16028 10474 16040
rect 11698 16028 11704 16040
rect 10468 16000 11704 16028
rect 10468 15988 10474 16000
rect 11698 15988 11704 16000
rect 11756 15988 11762 16040
rect 12253 16031 12311 16037
rect 12253 15997 12265 16031
rect 12299 16028 12311 16031
rect 12342 16028 12348 16040
rect 12299 16000 12348 16028
rect 12299 15997 12311 16000
rect 12253 15991 12311 15997
rect 12342 15988 12348 16000
rect 12400 15988 12406 16040
rect 13081 16031 13139 16037
rect 13081 15997 13093 16031
rect 13127 16028 13139 16031
rect 13740 16028 13768 16204
rect 14752 16164 14780 16204
rect 15194 16192 15200 16204
rect 15252 16192 15258 16244
rect 17678 16192 17684 16244
rect 17736 16232 17742 16244
rect 17865 16235 17923 16241
rect 17865 16232 17877 16235
rect 17736 16204 17877 16232
rect 17736 16192 17742 16204
rect 17865 16201 17877 16204
rect 17911 16201 17923 16235
rect 19886 16232 19892 16244
rect 19847 16204 19892 16232
rect 17865 16195 17923 16201
rect 19886 16192 19892 16204
rect 19944 16192 19950 16244
rect 16666 16164 16672 16176
rect 14752 16136 16672 16164
rect 16666 16124 16672 16136
rect 16724 16124 16730 16176
rect 15930 16096 15936 16108
rect 15891 16068 15936 16096
rect 15930 16056 15936 16068
rect 15988 16056 15994 16108
rect 17218 16096 17224 16108
rect 17179 16068 17224 16096
rect 17218 16056 17224 16068
rect 17276 16056 17282 16108
rect 13127 16000 13768 16028
rect 13817 16031 13875 16037
rect 13127 15997 13139 16000
rect 13081 15991 13139 15997
rect 13817 15997 13829 16031
rect 13863 16028 13875 16031
rect 14366 16028 14372 16040
rect 13863 16000 14372 16028
rect 13863 15997 13875 16000
rect 13817 15991 13875 15997
rect 9214 15960 9220 15972
rect 8680 15932 9220 15960
rect 9214 15920 9220 15932
rect 9272 15920 9278 15972
rect 10965 15963 11023 15969
rect 10965 15929 10977 15963
rect 11011 15960 11023 15963
rect 11882 15960 11888 15972
rect 11011 15932 11888 15960
rect 11011 15929 11023 15932
rect 10965 15923 11023 15929
rect 11882 15920 11888 15932
rect 11940 15920 11946 15972
rect 3789 15895 3847 15901
rect 3789 15861 3801 15895
rect 3835 15892 3847 15895
rect 6270 15892 6276 15904
rect 3835 15864 6276 15892
rect 3835 15861 3847 15864
rect 3789 15855 3847 15861
rect 6270 15852 6276 15864
rect 6328 15852 6334 15904
rect 7650 15892 7656 15904
rect 7611 15864 7656 15892
rect 7650 15852 7656 15864
rect 7708 15852 7714 15904
rect 8113 15895 8171 15901
rect 8113 15861 8125 15895
rect 8159 15892 8171 15895
rect 9306 15892 9312 15904
rect 8159 15864 9312 15892
rect 8159 15861 8171 15864
rect 8113 15855 8171 15861
rect 9306 15852 9312 15864
rect 9364 15852 9370 15904
rect 10594 15892 10600 15904
rect 10555 15864 10600 15892
rect 10594 15852 10600 15864
rect 10652 15852 10658 15904
rect 11054 15852 11060 15904
rect 11112 15892 11118 15904
rect 11112 15864 11157 15892
rect 11112 15852 11118 15864
rect 12250 15852 12256 15904
rect 12308 15892 12314 15904
rect 12345 15895 12403 15901
rect 12345 15892 12357 15895
rect 12308 15864 12357 15892
rect 12308 15852 12314 15864
rect 12345 15861 12357 15864
rect 12391 15861 12403 15895
rect 12894 15892 12900 15904
rect 12807 15864 12900 15892
rect 12345 15855 12403 15861
rect 12894 15852 12900 15864
rect 12952 15892 12958 15904
rect 13832 15892 13860 15991
rect 14366 15988 14372 16000
rect 14424 15988 14430 16040
rect 17310 15988 17316 16040
rect 17368 16028 17374 16040
rect 17497 16031 17555 16037
rect 17497 16028 17509 16031
rect 17368 16000 17509 16028
rect 17368 15988 17374 16000
rect 17497 15997 17509 16000
rect 17543 15997 17555 16031
rect 17497 15991 17555 15997
rect 19334 15988 19340 16040
rect 19392 16037 19398 16040
rect 19392 16028 19404 16037
rect 19613 16031 19671 16037
rect 19392 16000 19437 16028
rect 19392 15991 19404 16000
rect 19613 15997 19625 16031
rect 19659 15997 19671 16031
rect 19613 15991 19671 15997
rect 19392 15988 19398 15991
rect 14090 15969 14096 15972
rect 14084 15923 14096 15969
rect 14148 15960 14154 15972
rect 14148 15932 14184 15960
rect 14090 15920 14096 15923
rect 14148 15920 14154 15932
rect 14550 15920 14556 15972
rect 14608 15960 14614 15972
rect 16117 15963 16175 15969
rect 16117 15960 16129 15963
rect 14608 15932 16129 15960
rect 14608 15920 14614 15932
rect 16117 15929 16129 15932
rect 16163 15929 16175 15963
rect 16574 15960 16580 15972
rect 16117 15923 16175 15929
rect 16408 15932 16580 15960
rect 12952 15864 13860 15892
rect 12952 15852 12958 15864
rect 15286 15852 15292 15904
rect 15344 15892 15350 15904
rect 16025 15895 16083 15901
rect 16025 15892 16037 15895
rect 15344 15864 16037 15892
rect 15344 15852 15350 15864
rect 16025 15861 16037 15864
rect 16071 15892 16083 15895
rect 16408 15892 16436 15932
rect 16574 15920 16580 15932
rect 16632 15960 16638 15972
rect 17586 15960 17592 15972
rect 16632 15932 17592 15960
rect 16632 15920 16638 15932
rect 17586 15920 17592 15932
rect 17644 15920 17650 15972
rect 17770 15920 17776 15972
rect 17828 15960 17834 15972
rect 19628 15960 19656 15991
rect 17828 15932 19656 15960
rect 17828 15920 17834 15932
rect 16071 15864 16436 15892
rect 16485 15895 16543 15901
rect 16071 15861 16083 15864
rect 16025 15855 16083 15861
rect 16485 15861 16497 15895
rect 16531 15892 16543 15895
rect 17405 15895 17463 15901
rect 17405 15892 17417 15895
rect 16531 15864 17417 15892
rect 16531 15861 16543 15864
rect 16485 15855 16543 15861
rect 17405 15861 17417 15864
rect 17451 15861 17463 15895
rect 18230 15892 18236 15904
rect 18191 15864 18236 15892
rect 17405 15855 17463 15861
rect 18230 15852 18236 15864
rect 18288 15852 18294 15904
rect 1104 15802 21896 15824
rect 1104 15750 7912 15802
rect 7964 15750 7976 15802
rect 8028 15750 8040 15802
rect 8092 15750 8104 15802
rect 8156 15750 14843 15802
rect 14895 15750 14907 15802
rect 14959 15750 14971 15802
rect 15023 15750 15035 15802
rect 15087 15750 21896 15802
rect 1104 15728 21896 15750
rect 2130 15688 2136 15700
rect 2091 15660 2136 15688
rect 2130 15648 2136 15660
rect 2188 15648 2194 15700
rect 4065 15691 4123 15697
rect 4065 15688 4077 15691
rect 2332 15660 4077 15688
rect 1578 15552 1584 15564
rect 1539 15524 1584 15552
rect 1578 15512 1584 15524
rect 1636 15512 1642 15564
rect 1765 15555 1823 15561
rect 1765 15521 1777 15555
rect 1811 15552 1823 15555
rect 1854 15552 1860 15564
rect 1811 15524 1860 15552
rect 1811 15521 1823 15524
rect 1765 15515 1823 15521
rect 1854 15512 1860 15524
rect 1912 15512 1918 15564
rect 2332 15561 2360 15660
rect 4065 15657 4077 15660
rect 4111 15657 4123 15691
rect 4065 15651 4123 15657
rect 4525 15691 4583 15697
rect 4525 15657 4537 15691
rect 4571 15688 4583 15691
rect 5258 15688 5264 15700
rect 4571 15660 5264 15688
rect 4571 15657 4583 15660
rect 4525 15651 4583 15657
rect 5258 15648 5264 15660
rect 5316 15648 5322 15700
rect 5534 15648 5540 15700
rect 5592 15688 5598 15700
rect 6181 15691 6239 15697
rect 6181 15688 6193 15691
rect 5592 15660 6193 15688
rect 5592 15648 5598 15660
rect 6181 15657 6193 15660
rect 6227 15657 6239 15691
rect 7650 15688 7656 15700
rect 6181 15651 6239 15657
rect 6288 15660 7656 15688
rect 6288 15620 6316 15660
rect 7650 15648 7656 15660
rect 7708 15648 7714 15700
rect 9306 15688 9312 15700
rect 9267 15660 9312 15688
rect 9306 15648 9312 15660
rect 9364 15648 9370 15700
rect 9769 15691 9827 15697
rect 9769 15657 9781 15691
rect 9815 15688 9827 15691
rect 10962 15688 10968 15700
rect 9815 15660 10968 15688
rect 9815 15657 9827 15660
rect 9769 15651 9827 15657
rect 10962 15648 10968 15660
rect 11020 15648 11026 15700
rect 12345 15691 12403 15697
rect 11900 15660 12296 15688
rect 3252 15592 6316 15620
rect 6908 15623 6966 15629
rect 2317 15555 2375 15561
rect 2317 15521 2329 15555
rect 2363 15521 2375 15555
rect 2590 15552 2596 15564
rect 2551 15524 2596 15552
rect 2317 15515 2375 15521
rect 2590 15512 2596 15524
rect 2648 15512 2654 15564
rect 3252 15561 3280 15592
rect 6908 15589 6920 15623
rect 6954 15620 6966 15623
rect 7374 15620 7380 15632
rect 6954 15592 7380 15620
rect 6954 15589 6966 15592
rect 6908 15583 6966 15589
rect 7374 15580 7380 15592
rect 7432 15580 7438 15632
rect 11900 15620 11928 15660
rect 9692 15592 11928 15620
rect 9692 15564 9720 15592
rect 11974 15580 11980 15632
rect 12032 15629 12038 15632
rect 12032 15620 12044 15629
rect 12268 15620 12296 15660
rect 12345 15657 12357 15691
rect 12391 15688 12403 15691
rect 12894 15688 12900 15700
rect 12391 15660 12900 15688
rect 12391 15657 12403 15660
rect 12345 15651 12403 15657
rect 12894 15648 12900 15660
rect 12952 15648 12958 15700
rect 15286 15688 15292 15700
rect 13556 15660 15292 15688
rect 12032 15592 12077 15620
rect 12268 15592 12388 15620
rect 12032 15583 12044 15592
rect 12032 15580 12038 15583
rect 3237 15555 3295 15561
rect 3237 15521 3249 15555
rect 3283 15521 3295 15555
rect 3237 15515 3295 15521
rect 4249 15555 4307 15561
rect 4249 15521 4261 15555
rect 4295 15521 4307 15555
rect 4249 15515 4307 15521
rect 5649 15555 5707 15561
rect 5649 15521 5661 15555
rect 5695 15552 5707 15555
rect 5810 15552 5816 15564
rect 5695 15524 5816 15552
rect 5695 15521 5707 15524
rect 5649 15515 5707 15521
rect 2314 15376 2320 15428
rect 2372 15416 2378 15428
rect 3053 15419 3111 15425
rect 3053 15416 3065 15419
rect 2372 15388 3065 15416
rect 2372 15376 2378 15388
rect 3053 15385 3065 15388
rect 3099 15385 3111 15419
rect 3053 15379 3111 15385
rect 2774 15348 2780 15360
rect 2735 15320 2780 15348
rect 2774 15308 2780 15320
rect 2832 15308 2838 15360
rect 4264 15348 4292 15515
rect 5810 15512 5816 15524
rect 5868 15512 5874 15564
rect 7190 15512 7196 15564
rect 7248 15552 7254 15564
rect 8481 15555 8539 15561
rect 8481 15552 8493 15555
rect 7248 15524 8493 15552
rect 7248 15512 7254 15524
rect 8481 15521 8493 15524
rect 8527 15521 8539 15555
rect 9674 15552 9680 15564
rect 9635 15524 9680 15552
rect 8481 15515 8539 15521
rect 5905 15487 5963 15493
rect 5905 15453 5917 15487
rect 5951 15484 5963 15487
rect 5994 15484 6000 15496
rect 5951 15456 6000 15484
rect 5951 15453 5963 15456
rect 5905 15447 5963 15453
rect 5994 15444 6000 15456
rect 6052 15484 6058 15496
rect 6454 15484 6460 15496
rect 6052 15456 6460 15484
rect 6052 15444 6058 15456
rect 6454 15444 6460 15456
rect 6512 15484 6518 15496
rect 6641 15487 6699 15493
rect 6641 15484 6653 15487
rect 6512 15456 6653 15484
rect 6512 15444 6518 15456
rect 6641 15453 6653 15456
rect 6687 15453 6699 15487
rect 8496 15484 8524 15515
rect 9674 15512 9680 15524
rect 9732 15512 9738 15564
rect 10042 15552 10048 15564
rect 9784 15524 10048 15552
rect 9784 15484 9812 15524
rect 10042 15512 10048 15524
rect 10100 15512 10106 15564
rect 10321 15555 10379 15561
rect 10321 15521 10333 15555
rect 10367 15521 10379 15555
rect 10321 15515 10379 15521
rect 8496 15456 9812 15484
rect 6641 15447 6699 15453
rect 9858 15444 9864 15496
rect 9916 15484 9922 15496
rect 9916 15456 9961 15484
rect 9916 15444 9922 15456
rect 8754 15376 8760 15428
rect 8812 15416 8818 15428
rect 10336 15416 10364 15515
rect 10686 15512 10692 15564
rect 10744 15552 10750 15564
rect 12253 15555 12311 15561
rect 12253 15552 12265 15555
rect 10744 15524 12265 15552
rect 10744 15512 10750 15524
rect 12253 15521 12265 15524
rect 12299 15521 12311 15555
rect 12360 15552 12388 15592
rect 12434 15580 12440 15632
rect 12492 15620 12498 15632
rect 13556 15620 13584 15660
rect 15286 15648 15292 15660
rect 15344 15648 15350 15700
rect 15930 15648 15936 15700
rect 15988 15688 15994 15700
rect 17129 15691 17187 15697
rect 17129 15688 17141 15691
rect 15988 15660 17141 15688
rect 15988 15648 15994 15660
rect 17129 15657 17141 15660
rect 17175 15657 17187 15691
rect 17129 15651 17187 15657
rect 12492 15592 13584 15620
rect 13633 15623 13691 15629
rect 12492 15580 12498 15592
rect 13633 15589 13645 15623
rect 13679 15620 13691 15623
rect 14734 15620 14740 15632
rect 13679 15592 14740 15620
rect 13679 15589 13691 15592
rect 13633 15583 13691 15589
rect 14734 15580 14740 15592
rect 14792 15580 14798 15632
rect 16758 15620 16764 15632
rect 15764 15592 16764 15620
rect 12897 15555 12955 15561
rect 12897 15552 12909 15555
rect 12360 15524 12909 15552
rect 12253 15515 12311 15521
rect 12897 15521 12909 15524
rect 12943 15521 12955 15555
rect 12897 15515 12955 15521
rect 12268 15484 12296 15515
rect 13078 15512 13084 15564
rect 13136 15552 13142 15564
rect 13725 15555 13783 15561
rect 13136 15524 13676 15552
rect 13136 15512 13142 15524
rect 12345 15487 12403 15493
rect 12345 15484 12357 15487
rect 12268 15456 12357 15484
rect 12345 15453 12357 15456
rect 12391 15453 12403 15487
rect 12345 15447 12403 15453
rect 8812 15388 10364 15416
rect 8812 15376 8818 15388
rect 12250 15376 12256 15428
rect 12308 15416 12314 15428
rect 12529 15419 12587 15425
rect 12529 15416 12541 15419
rect 12308 15388 12541 15416
rect 12308 15376 12314 15388
rect 12529 15385 12541 15388
rect 12575 15385 12587 15419
rect 12529 15379 12587 15385
rect 13078 15376 13084 15428
rect 13136 15416 13142 15428
rect 13538 15416 13544 15428
rect 13136 15388 13544 15416
rect 13136 15376 13142 15388
rect 13538 15376 13544 15388
rect 13596 15376 13602 15428
rect 13648 15360 13676 15524
rect 13725 15521 13737 15555
rect 13771 15552 13783 15555
rect 13998 15552 14004 15564
rect 13771 15524 14004 15552
rect 13771 15521 13783 15524
rect 13725 15515 13783 15521
rect 13998 15512 14004 15524
rect 14056 15512 14062 15564
rect 14642 15512 14648 15564
rect 14700 15552 14706 15564
rect 15764 15561 15792 15592
rect 16758 15580 16764 15592
rect 16816 15580 16822 15632
rect 17954 15580 17960 15632
rect 18012 15620 18018 15632
rect 18049 15623 18107 15629
rect 18049 15620 18061 15623
rect 18012 15592 18061 15620
rect 18012 15580 18018 15592
rect 18049 15589 18061 15592
rect 18095 15589 18107 15623
rect 18049 15583 18107 15589
rect 18138 15580 18144 15632
rect 18196 15620 18202 15632
rect 19153 15623 19211 15629
rect 19153 15620 19165 15623
rect 18196 15592 19165 15620
rect 18196 15580 18202 15592
rect 19153 15589 19165 15592
rect 19199 15589 19211 15623
rect 19153 15583 19211 15589
rect 16022 15561 16028 15564
rect 15289 15555 15347 15561
rect 15289 15552 15301 15555
rect 14700 15524 15301 15552
rect 14700 15512 14706 15524
rect 15289 15521 15301 15524
rect 15335 15521 15347 15555
rect 15289 15515 15347 15521
rect 15749 15555 15807 15561
rect 15749 15521 15761 15555
rect 15795 15521 15807 15555
rect 16016 15552 16028 15561
rect 15983 15524 16028 15552
rect 15749 15515 15807 15521
rect 16016 15515 16028 15524
rect 16022 15512 16028 15515
rect 16080 15512 16086 15564
rect 18156 15552 18184 15580
rect 17972 15524 18184 15552
rect 17972 15493 18000 15524
rect 13817 15487 13875 15493
rect 13817 15484 13829 15487
rect 13740 15456 13829 15484
rect 13740 15428 13768 15456
rect 13817 15453 13829 15456
rect 13863 15453 13875 15487
rect 13817 15447 13875 15453
rect 17865 15487 17923 15493
rect 17865 15453 17877 15487
rect 17911 15453 17923 15487
rect 17865 15447 17923 15453
rect 17957 15487 18015 15493
rect 17957 15453 17969 15487
rect 18003 15453 18015 15487
rect 17957 15447 18015 15453
rect 13722 15376 13728 15428
rect 13780 15376 13786 15428
rect 13906 15376 13912 15428
rect 13964 15416 13970 15428
rect 14550 15416 14556 15428
rect 13964 15388 14556 15416
rect 13964 15376 13970 15388
rect 14550 15376 14556 15388
rect 14608 15416 14614 15428
rect 14921 15419 14979 15425
rect 14921 15416 14933 15419
rect 14608 15388 14933 15416
rect 14608 15376 14614 15388
rect 14921 15385 14933 15388
rect 14967 15385 14979 15419
rect 17880 15416 17908 15447
rect 18138 15444 18144 15496
rect 18196 15484 18202 15496
rect 18693 15487 18751 15493
rect 18693 15484 18705 15487
rect 18196 15456 18705 15484
rect 18196 15444 18202 15456
rect 18693 15453 18705 15456
rect 18739 15453 18751 15487
rect 18693 15447 18751 15453
rect 18046 15416 18052 15428
rect 17880 15388 18052 15416
rect 14921 15379 14979 15385
rect 18046 15376 18052 15388
rect 18104 15416 18110 15428
rect 18230 15416 18236 15428
rect 18104 15388 18236 15416
rect 18104 15376 18110 15388
rect 18230 15376 18236 15388
rect 18288 15376 18294 15428
rect 6638 15348 6644 15360
rect 4264 15320 6644 15348
rect 6638 15308 6644 15320
rect 6696 15308 6702 15360
rect 6914 15308 6920 15360
rect 6972 15348 6978 15360
rect 8021 15351 8079 15357
rect 8021 15348 8033 15351
rect 6972 15320 8033 15348
rect 6972 15308 6978 15320
rect 8021 15317 8033 15320
rect 8067 15317 8079 15351
rect 8021 15311 8079 15317
rect 8297 15351 8355 15357
rect 8297 15317 8309 15351
rect 8343 15348 8355 15351
rect 8386 15348 8392 15360
rect 8343 15320 8392 15348
rect 8343 15317 8355 15320
rect 8297 15311 8355 15317
rect 8386 15308 8392 15320
rect 8444 15308 8450 15360
rect 9306 15308 9312 15360
rect 9364 15348 9370 15360
rect 9950 15348 9956 15360
rect 9364 15320 9956 15348
rect 9364 15308 9370 15320
rect 9950 15308 9956 15320
rect 10008 15308 10014 15360
rect 10226 15308 10232 15360
rect 10284 15348 10290 15360
rect 10505 15351 10563 15357
rect 10505 15348 10517 15351
rect 10284 15320 10517 15348
rect 10284 15308 10290 15320
rect 10505 15317 10517 15320
rect 10551 15317 10563 15351
rect 10505 15311 10563 15317
rect 10873 15351 10931 15357
rect 10873 15317 10885 15351
rect 10919 15348 10931 15351
rect 10962 15348 10968 15360
rect 10919 15320 10968 15348
rect 10919 15317 10931 15320
rect 10873 15311 10931 15317
rect 10962 15308 10968 15320
rect 11020 15308 11026 15360
rect 13262 15348 13268 15360
rect 13223 15320 13268 15348
rect 13262 15308 13268 15320
rect 13320 15308 13326 15360
rect 13630 15348 13636 15360
rect 13543 15320 13636 15348
rect 13630 15308 13636 15320
rect 13688 15348 13694 15360
rect 13814 15348 13820 15360
rect 13688 15320 13820 15348
rect 13688 15308 13694 15320
rect 13814 15308 13820 15320
rect 13872 15348 13878 15360
rect 14369 15351 14427 15357
rect 14369 15348 14381 15351
rect 13872 15320 14381 15348
rect 13872 15308 13878 15320
rect 14369 15317 14381 15320
rect 14415 15348 14427 15351
rect 15102 15348 15108 15360
rect 14415 15320 15108 15348
rect 14415 15317 14427 15320
rect 14369 15311 14427 15317
rect 15102 15308 15108 15320
rect 15160 15308 15166 15360
rect 15473 15351 15531 15357
rect 15473 15317 15485 15351
rect 15519 15348 15531 15351
rect 16666 15348 16672 15360
rect 15519 15320 16672 15348
rect 15519 15317 15531 15320
rect 15473 15311 15531 15317
rect 16666 15308 16672 15320
rect 16724 15308 16730 15360
rect 17954 15308 17960 15360
rect 18012 15348 18018 15360
rect 18417 15351 18475 15357
rect 18417 15348 18429 15351
rect 18012 15320 18429 15348
rect 18012 15308 18018 15320
rect 18417 15317 18429 15320
rect 18463 15317 18475 15351
rect 18417 15311 18475 15317
rect 1104 15258 21896 15280
rect 1104 15206 4447 15258
rect 4499 15206 4511 15258
rect 4563 15206 4575 15258
rect 4627 15206 4639 15258
rect 4691 15206 11378 15258
rect 11430 15206 11442 15258
rect 11494 15206 11506 15258
rect 11558 15206 11570 15258
rect 11622 15206 18308 15258
rect 18360 15206 18372 15258
rect 18424 15206 18436 15258
rect 18488 15206 18500 15258
rect 18552 15206 21896 15258
rect 1104 15184 21896 15206
rect 1670 15144 1676 15156
rect 1631 15116 1676 15144
rect 1670 15104 1676 15116
rect 1728 15104 1734 15156
rect 1762 15104 1768 15156
rect 1820 15144 1826 15156
rect 2133 15147 2191 15153
rect 2133 15144 2145 15147
rect 1820 15116 2145 15144
rect 1820 15104 1826 15116
rect 2133 15113 2145 15116
rect 2179 15113 2191 15147
rect 2133 15107 2191 15113
rect 5166 15104 5172 15156
rect 5224 15144 5230 15156
rect 5353 15147 5411 15153
rect 5353 15144 5365 15147
rect 5224 15116 5365 15144
rect 5224 15104 5230 15116
rect 5353 15113 5365 15116
rect 5399 15113 5411 15147
rect 8113 15147 8171 15153
rect 8113 15144 8125 15147
rect 5353 15107 5411 15113
rect 6656 15116 8125 15144
rect 3973 15079 4031 15085
rect 3973 15045 3985 15079
rect 4019 15045 4031 15079
rect 3973 15039 4031 15045
rect 3988 15008 4016 15039
rect 5258 15036 5264 15088
rect 5316 15076 5322 15088
rect 6656 15076 6684 15116
rect 8113 15113 8125 15116
rect 8159 15113 8171 15147
rect 8294 15144 8300 15156
rect 8255 15116 8300 15144
rect 8113 15107 8171 15113
rect 8294 15104 8300 15116
rect 8352 15104 8358 15156
rect 10134 15144 10140 15156
rect 8404 15116 10140 15144
rect 8404 15076 8432 15116
rect 10134 15104 10140 15116
rect 10192 15104 10198 15156
rect 10410 15104 10416 15156
rect 10468 15144 10474 15156
rect 12066 15144 12072 15156
rect 10468 15116 12072 15144
rect 10468 15104 10474 15116
rect 12066 15104 12072 15116
rect 12124 15104 12130 15156
rect 12526 15104 12532 15156
rect 12584 15144 12590 15156
rect 12805 15147 12863 15153
rect 12805 15144 12817 15147
rect 12584 15116 12817 15144
rect 12584 15104 12590 15116
rect 12805 15113 12817 15116
rect 12851 15113 12863 15147
rect 12805 15107 12863 15113
rect 13081 15147 13139 15153
rect 13081 15113 13093 15147
rect 13127 15144 13139 15147
rect 14090 15144 14096 15156
rect 13127 15116 14096 15144
rect 13127 15113 13139 15116
rect 13081 15107 13139 15113
rect 11698 15076 11704 15088
rect 5316 15048 6684 15076
rect 6748 15048 8432 15076
rect 11659 15048 11704 15076
rect 5316 15036 5322 15048
rect 4338 15008 4344 15020
rect 3988 14980 4344 15008
rect 4338 14968 4344 14980
rect 4396 15008 4402 15020
rect 4801 15011 4859 15017
rect 4801 15008 4813 15011
rect 4396 14980 4813 15008
rect 4396 14968 4402 14980
rect 4801 14977 4813 14980
rect 4847 14977 4859 15011
rect 5902 15008 5908 15020
rect 5863 14980 5908 15008
rect 4801 14971 4859 14977
rect 5902 14968 5908 14980
rect 5960 14968 5966 15020
rect 2314 14940 2320 14952
rect 2275 14912 2320 14940
rect 2314 14900 2320 14912
rect 2372 14900 2378 14952
rect 2866 14949 2872 14952
rect 2593 14943 2651 14949
rect 2593 14909 2605 14943
rect 2639 14909 2651 14943
rect 2593 14903 2651 14909
rect 2860 14903 2872 14949
rect 2924 14940 2930 14952
rect 4709 14943 4767 14949
rect 2924 14912 2960 14940
rect 1762 14872 1768 14884
rect 1723 14844 1768 14872
rect 1762 14832 1768 14844
rect 1820 14832 1826 14884
rect 2608 14872 2636 14903
rect 2866 14900 2872 14903
rect 2924 14900 2930 14912
rect 4709 14909 4721 14943
rect 4755 14940 4767 14943
rect 4890 14940 4896 14952
rect 4755 14912 4896 14940
rect 4755 14909 4767 14912
rect 4709 14903 4767 14909
rect 4890 14900 4896 14912
rect 4948 14900 4954 14952
rect 5813 14943 5871 14949
rect 5813 14909 5825 14943
rect 5859 14940 5871 14943
rect 6748 14940 6776 15048
rect 11698 15036 11704 15048
rect 11756 15036 11762 15088
rect 13096 15076 13124 15107
rect 14090 15104 14096 15116
rect 14148 15104 14154 15156
rect 14734 15144 14740 15156
rect 14695 15116 14740 15144
rect 14734 15104 14740 15116
rect 14792 15104 14798 15156
rect 16577 15147 16635 15153
rect 16577 15113 16589 15147
rect 16623 15144 16635 15147
rect 17126 15144 17132 15156
rect 16623 15116 17132 15144
rect 16623 15113 16635 15116
rect 16577 15107 16635 15113
rect 17126 15104 17132 15116
rect 17184 15104 17190 15156
rect 12268 15048 13124 15076
rect 6825 15011 6883 15017
rect 6825 14977 6837 15011
rect 6871 15008 6883 15011
rect 6914 15008 6920 15020
rect 6871 14980 6920 15008
rect 6871 14977 6883 14980
rect 6825 14971 6883 14977
rect 6914 14968 6920 14980
rect 6972 14968 6978 15020
rect 8021 15011 8079 15017
rect 8021 14977 8033 15011
rect 8067 15008 8079 15011
rect 8202 15008 8208 15020
rect 8067 14980 8208 15008
rect 8067 14977 8079 14980
rect 8021 14971 8079 14977
rect 8202 14968 8208 14980
rect 8260 14968 8266 15020
rect 10318 15008 10324 15020
rect 9600 14980 10324 15008
rect 9600 14940 9628 14980
rect 10318 14968 10324 14980
rect 10376 14968 10382 15020
rect 12268 15017 12296 15048
rect 12253 15011 12311 15017
rect 12253 14977 12265 15011
rect 12299 14977 12311 15011
rect 12253 14971 12311 14977
rect 12345 15011 12403 15017
rect 12345 14977 12357 15011
rect 12391 15008 12403 15011
rect 13262 15008 13268 15020
rect 12391 14980 13268 15008
rect 12391 14977 12403 14980
rect 12345 14971 12403 14977
rect 13262 14968 13268 14980
rect 13320 14968 13326 15020
rect 14734 14968 14740 15020
rect 14792 15008 14798 15020
rect 15289 15011 15347 15017
rect 15289 15008 15301 15011
rect 14792 14980 15301 15008
rect 14792 14968 14798 14980
rect 15289 14977 15301 14980
rect 15335 14977 15347 15011
rect 15289 14971 15347 14977
rect 15378 14968 15384 15020
rect 15436 15008 15442 15020
rect 15933 15011 15991 15017
rect 15933 15008 15945 15011
rect 15436 14980 15945 15008
rect 15436 14968 15442 14980
rect 15933 14977 15945 14980
rect 15979 15008 15991 15011
rect 16022 15008 16028 15020
rect 15979 14980 16028 15008
rect 15979 14977 15991 14980
rect 15933 14971 15991 14977
rect 16022 14968 16028 14980
rect 16080 14968 16086 15020
rect 17770 14968 17776 15020
rect 17828 15008 17834 15020
rect 17957 15011 18015 15017
rect 17957 15008 17969 15011
rect 17828 14980 17969 15008
rect 17828 14968 17834 14980
rect 17957 14977 17969 14980
rect 18003 14977 18015 15011
rect 17957 14971 18015 14977
rect 5859 14912 6776 14940
rect 6932 14912 9628 14940
rect 9677 14943 9735 14949
rect 5859 14909 5871 14912
rect 5813 14903 5871 14909
rect 4062 14872 4068 14884
rect 2608 14844 4068 14872
rect 4062 14832 4068 14844
rect 4120 14832 4126 14884
rect 6932 14881 6960 14912
rect 9677 14909 9689 14943
rect 9723 14940 9735 14943
rect 9950 14940 9956 14952
rect 9723 14912 9956 14940
rect 9723 14909 9735 14912
rect 9677 14903 9735 14909
rect 9950 14900 9956 14912
rect 10008 14900 10014 14952
rect 11330 14940 11336 14952
rect 11291 14912 11336 14940
rect 11330 14900 11336 14912
rect 11388 14900 11394 14952
rect 12434 14900 12440 14952
rect 12492 14940 12498 14952
rect 12492 14912 12537 14940
rect 12492 14900 12498 14912
rect 13722 14900 13728 14952
rect 13780 14940 13786 14952
rect 14194 14943 14252 14949
rect 14194 14940 14206 14943
rect 13780 14912 14206 14940
rect 13780 14900 13786 14912
rect 14194 14909 14206 14912
rect 14240 14909 14252 14943
rect 14194 14903 14252 14909
rect 14366 14900 14372 14952
rect 14424 14940 14430 14952
rect 14461 14943 14519 14949
rect 14461 14940 14473 14943
rect 14424 14912 14473 14940
rect 14424 14900 14430 14912
rect 14461 14909 14473 14912
rect 14507 14909 14519 14943
rect 14461 14903 14519 14909
rect 18046 14900 18052 14952
rect 18104 14940 18110 14952
rect 18213 14943 18271 14949
rect 18213 14940 18225 14943
rect 18104 14912 18225 14940
rect 18104 14900 18110 14912
rect 18213 14909 18225 14912
rect 18259 14909 18271 14943
rect 18213 14903 18271 14909
rect 4617 14875 4675 14881
rect 4617 14841 4629 14875
rect 4663 14872 4675 14875
rect 6917 14875 6975 14881
rect 4663 14844 6132 14872
rect 4663 14841 4675 14844
rect 4617 14835 4675 14841
rect 4246 14804 4252 14816
rect 4207 14776 4252 14804
rect 4246 14764 4252 14776
rect 4304 14764 4310 14816
rect 5258 14764 5264 14816
rect 5316 14804 5322 14816
rect 5721 14807 5779 14813
rect 5721 14804 5733 14807
rect 5316 14776 5733 14804
rect 5316 14764 5322 14776
rect 5721 14773 5733 14776
rect 5767 14773 5779 14807
rect 6104 14804 6132 14844
rect 6917 14841 6929 14875
rect 6963 14841 6975 14875
rect 6917 14835 6975 14841
rect 7190 14832 7196 14884
rect 7248 14872 7254 14884
rect 8570 14872 8576 14884
rect 7248 14844 8576 14872
rect 7248 14832 7254 14844
rect 8570 14832 8576 14844
rect 8628 14832 8634 14884
rect 9432 14875 9490 14881
rect 9432 14841 9444 14875
rect 9478 14872 9490 14875
rect 9858 14872 9864 14884
rect 9478 14844 9864 14872
rect 9478 14841 9490 14844
rect 9432 14835 9490 14841
rect 9858 14832 9864 14844
rect 9916 14832 9922 14884
rect 10870 14872 10876 14884
rect 9968 14844 10876 14872
rect 6546 14804 6552 14816
rect 6104 14776 6552 14804
rect 5721 14767 5779 14773
rect 6546 14764 6552 14776
rect 6604 14804 6610 14816
rect 7009 14807 7067 14813
rect 7009 14804 7021 14807
rect 6604 14776 7021 14804
rect 6604 14764 6610 14776
rect 7009 14773 7021 14776
rect 7055 14773 7067 14807
rect 7009 14767 7067 14773
rect 7098 14764 7104 14816
rect 7156 14804 7162 14816
rect 7377 14807 7435 14813
rect 7377 14804 7389 14807
rect 7156 14776 7389 14804
rect 7156 14764 7162 14776
rect 7377 14773 7389 14776
rect 7423 14773 7435 14807
rect 7377 14767 7435 14773
rect 8113 14807 8171 14813
rect 8113 14773 8125 14807
rect 8159 14804 8171 14807
rect 9674 14804 9680 14816
rect 8159 14776 9680 14804
rect 8159 14773 8171 14776
rect 8113 14767 8171 14773
rect 9674 14764 9680 14776
rect 9732 14764 9738 14816
rect 9968 14813 9996 14844
rect 10870 14832 10876 14844
rect 10928 14832 10934 14884
rect 10962 14832 10968 14884
rect 11020 14872 11026 14884
rect 11066 14875 11124 14881
rect 11066 14872 11078 14875
rect 11020 14844 11078 14872
rect 11020 14832 11026 14844
rect 11066 14841 11078 14844
rect 11112 14872 11124 14875
rect 11238 14872 11244 14884
rect 11112 14844 11244 14872
rect 11112 14841 11124 14844
rect 11066 14835 11124 14841
rect 11238 14832 11244 14844
rect 11296 14832 11302 14884
rect 11348 14844 12480 14872
rect 9953 14807 10011 14813
rect 9953 14773 9965 14807
rect 9999 14773 10011 14807
rect 9953 14767 10011 14773
rect 10042 14764 10048 14816
rect 10100 14804 10106 14816
rect 11348 14804 11376 14844
rect 10100 14776 11376 14804
rect 12452 14804 12480 14844
rect 12526 14832 12532 14884
rect 12584 14872 12590 14884
rect 13170 14872 13176 14884
rect 12584 14844 13176 14872
rect 12584 14832 12590 14844
rect 13170 14832 13176 14844
rect 13228 14872 13234 14884
rect 13228 14844 15240 14872
rect 13228 14832 13234 14844
rect 14458 14804 14464 14816
rect 12452 14776 14464 14804
rect 10100 14764 10106 14776
rect 14458 14764 14464 14776
rect 14516 14804 14522 14816
rect 15212 14813 15240 14844
rect 15105 14807 15163 14813
rect 15105 14804 15117 14807
rect 14516 14776 15117 14804
rect 14516 14764 14522 14776
rect 15105 14773 15117 14776
rect 15151 14773 15163 14807
rect 15105 14767 15163 14773
rect 15197 14807 15255 14813
rect 15197 14773 15209 14807
rect 15243 14804 15255 14807
rect 15838 14804 15844 14816
rect 15243 14776 15844 14804
rect 15243 14773 15255 14776
rect 15197 14767 15255 14773
rect 15838 14764 15844 14776
rect 15896 14764 15902 14816
rect 16114 14804 16120 14816
rect 16075 14776 16120 14804
rect 16114 14764 16120 14776
rect 16172 14764 16178 14816
rect 16206 14764 16212 14816
rect 16264 14804 16270 14816
rect 16942 14804 16948 14816
rect 16264 14776 16309 14804
rect 16903 14776 16948 14804
rect 16264 14764 16270 14776
rect 16942 14764 16948 14776
rect 17000 14764 17006 14816
rect 17494 14804 17500 14816
rect 17455 14776 17500 14804
rect 17494 14764 17500 14776
rect 17552 14804 17558 14816
rect 17862 14804 17868 14816
rect 17552 14776 17868 14804
rect 17552 14764 17558 14776
rect 17862 14764 17868 14776
rect 17920 14764 17926 14816
rect 19058 14764 19064 14816
rect 19116 14804 19122 14816
rect 19337 14807 19395 14813
rect 19337 14804 19349 14807
rect 19116 14776 19349 14804
rect 19116 14764 19122 14776
rect 19337 14773 19349 14776
rect 19383 14773 19395 14807
rect 19337 14767 19395 14773
rect 1104 14714 21896 14736
rect 1104 14662 7912 14714
rect 7964 14662 7976 14714
rect 8028 14662 8040 14714
rect 8092 14662 8104 14714
rect 8156 14662 14843 14714
rect 14895 14662 14907 14714
rect 14959 14662 14971 14714
rect 15023 14662 15035 14714
rect 15087 14662 21896 14714
rect 1104 14640 21896 14662
rect 2222 14600 2228 14612
rect 2183 14572 2228 14600
rect 2222 14560 2228 14572
rect 2280 14560 2286 14612
rect 3237 14603 3295 14609
rect 3237 14569 3249 14603
rect 3283 14600 3295 14603
rect 4246 14600 4252 14612
rect 3283 14572 4252 14600
rect 3283 14569 3295 14572
rect 3237 14563 3295 14569
rect 4246 14560 4252 14572
rect 4304 14560 4310 14612
rect 5445 14603 5503 14609
rect 5445 14569 5457 14603
rect 5491 14600 5503 14603
rect 7374 14600 7380 14612
rect 5491 14572 7380 14600
rect 5491 14569 5503 14572
rect 5445 14563 5503 14569
rect 4338 14541 4344 14544
rect 4332 14532 4344 14541
rect 4299 14504 4344 14532
rect 4332 14495 4344 14504
rect 4338 14492 4344 14495
rect 4396 14492 4402 14544
rect 1765 14467 1823 14473
rect 1765 14433 1777 14467
rect 1811 14464 1823 14467
rect 1946 14464 1952 14476
rect 1811 14436 1952 14464
rect 1811 14433 1823 14436
rect 1765 14427 1823 14433
rect 1946 14424 1952 14436
rect 2004 14424 2010 14476
rect 2222 14424 2228 14476
rect 2280 14464 2286 14476
rect 2317 14467 2375 14473
rect 2317 14464 2329 14467
rect 2280 14436 2329 14464
rect 2280 14424 2286 14436
rect 2317 14433 2329 14436
rect 2363 14433 2375 14467
rect 3142 14464 3148 14476
rect 3103 14436 3148 14464
rect 2317 14427 2375 14433
rect 3142 14424 3148 14436
rect 3200 14424 3206 14476
rect 5460 14464 5488 14563
rect 7374 14560 7380 14572
rect 7432 14560 7438 14612
rect 8205 14603 8263 14609
rect 8205 14569 8217 14603
rect 8251 14569 8263 14603
rect 8205 14563 8263 14569
rect 6089 14535 6147 14541
rect 6089 14501 6101 14535
rect 6135 14532 6147 14535
rect 7006 14532 7012 14544
rect 6135 14504 7012 14532
rect 6135 14501 6147 14504
rect 6089 14495 6147 14501
rect 7006 14492 7012 14504
rect 7064 14492 7070 14544
rect 8220 14532 8248 14563
rect 8662 14560 8668 14612
rect 8720 14600 8726 14612
rect 9125 14603 9183 14609
rect 9125 14600 9137 14603
rect 8720 14572 9137 14600
rect 8720 14560 8726 14572
rect 9125 14569 9137 14572
rect 9171 14569 9183 14603
rect 9125 14563 9183 14569
rect 9861 14603 9919 14609
rect 9861 14569 9873 14603
rect 9907 14600 9919 14603
rect 10594 14600 10600 14612
rect 9907 14572 10600 14600
rect 9907 14569 9919 14572
rect 9861 14563 9919 14569
rect 10594 14560 10600 14572
rect 10652 14560 10658 14612
rect 11054 14560 11060 14612
rect 11112 14600 11118 14612
rect 12253 14603 12311 14609
rect 12253 14600 12265 14603
rect 11112 14572 12265 14600
rect 11112 14560 11118 14572
rect 12253 14569 12265 14572
rect 12299 14569 12311 14603
rect 12253 14563 12311 14569
rect 12713 14603 12771 14609
rect 12713 14569 12725 14603
rect 12759 14600 12771 14603
rect 12802 14600 12808 14612
rect 12759 14572 12808 14600
rect 12759 14569 12771 14572
rect 12713 14563 12771 14569
rect 12158 14532 12164 14544
rect 8220 14504 12164 14532
rect 12158 14492 12164 14504
rect 12216 14492 12222 14544
rect 12728 14532 12756 14563
rect 12802 14560 12808 14572
rect 12860 14560 12866 14612
rect 13446 14560 13452 14612
rect 13504 14600 13510 14612
rect 13633 14603 13691 14609
rect 13633 14600 13645 14603
rect 13504 14572 13645 14600
rect 13504 14560 13510 14572
rect 13633 14569 13645 14572
rect 13679 14569 13691 14603
rect 13998 14600 14004 14612
rect 13959 14572 14004 14600
rect 13633 14563 13691 14569
rect 13998 14560 14004 14572
rect 14056 14560 14062 14612
rect 14642 14560 14648 14612
rect 14700 14600 14706 14612
rect 14737 14603 14795 14609
rect 14737 14600 14749 14603
rect 14700 14572 14749 14600
rect 14700 14560 14706 14572
rect 14737 14569 14749 14572
rect 14783 14569 14795 14603
rect 14737 14563 14795 14569
rect 15105 14603 15163 14609
rect 15105 14569 15117 14603
rect 15151 14600 15163 14603
rect 15194 14600 15200 14612
rect 15151 14572 15200 14600
rect 15151 14569 15163 14572
rect 15105 14563 15163 14569
rect 15194 14560 15200 14572
rect 15252 14560 15258 14612
rect 15378 14600 15384 14612
rect 15339 14572 15384 14600
rect 15378 14560 15384 14572
rect 15436 14560 15442 14612
rect 17402 14600 17408 14612
rect 15488 14572 17408 14600
rect 13538 14532 13544 14544
rect 12268 14504 12756 14532
rect 13499 14504 13544 14532
rect 12268 14476 12296 14504
rect 13538 14492 13544 14504
rect 13596 14492 13602 14544
rect 15212 14532 15240 14560
rect 15488 14532 15516 14572
rect 17402 14560 17408 14572
rect 17460 14560 17466 14612
rect 17954 14600 17960 14612
rect 17915 14572 17960 14600
rect 17954 14560 17960 14572
rect 18012 14560 18018 14612
rect 18049 14603 18107 14609
rect 18049 14569 18061 14603
rect 18095 14600 18107 14603
rect 18138 14600 18144 14612
rect 18095 14572 18144 14600
rect 18095 14569 18107 14572
rect 18049 14563 18107 14569
rect 18138 14560 18144 14572
rect 18196 14560 18202 14612
rect 18417 14603 18475 14609
rect 18417 14569 18429 14603
rect 18463 14600 18475 14603
rect 18598 14600 18604 14612
rect 18463 14572 18604 14600
rect 18463 14569 18475 14572
rect 18417 14563 18475 14569
rect 18598 14560 18604 14572
rect 18656 14560 18662 14612
rect 16942 14532 16948 14544
rect 13832 14504 14780 14532
rect 15212 14504 15516 14532
rect 15580 14504 16948 14532
rect 3436 14436 5488 14464
rect 6365 14467 6423 14473
rect 3436 14405 3464 14436
rect 6365 14433 6377 14467
rect 6411 14464 6423 14467
rect 6454 14464 6460 14476
rect 6411 14436 6460 14464
rect 6411 14433 6423 14436
rect 6365 14427 6423 14433
rect 6454 14424 6460 14436
rect 6512 14424 6518 14476
rect 6632 14467 6690 14473
rect 6632 14433 6644 14467
rect 6678 14464 6690 14467
rect 6914 14464 6920 14476
rect 6678 14436 6920 14464
rect 6678 14433 6690 14436
rect 6632 14427 6690 14433
rect 6914 14424 6920 14436
rect 6972 14424 6978 14476
rect 7558 14424 7564 14476
rect 7616 14464 7622 14476
rect 8021 14467 8079 14473
rect 8021 14464 8033 14467
rect 7616 14436 8033 14464
rect 7616 14424 7622 14436
rect 8021 14433 8033 14436
rect 8067 14433 8079 14467
rect 8021 14427 8079 14433
rect 8481 14467 8539 14473
rect 8481 14433 8493 14467
rect 8527 14464 8539 14467
rect 8846 14464 8852 14476
rect 8527 14436 8852 14464
rect 8527 14433 8539 14436
rect 8481 14427 8539 14433
rect 3421 14399 3479 14405
rect 3421 14365 3433 14399
rect 3467 14365 3479 14399
rect 4062 14396 4068 14408
rect 4023 14368 4068 14396
rect 3421 14359 3479 14365
rect 4062 14356 4068 14368
rect 4120 14356 4126 14408
rect 5000 14300 5580 14328
rect 1670 14260 1676 14272
rect 1631 14232 1676 14260
rect 1670 14220 1676 14232
rect 1728 14220 1734 14272
rect 2774 14220 2780 14272
rect 2832 14260 2838 14272
rect 2832 14232 2877 14260
rect 2832 14220 2838 14232
rect 3602 14220 3608 14272
rect 3660 14260 3666 14272
rect 5000 14260 5028 14300
rect 3660 14232 5028 14260
rect 5552 14260 5580 14300
rect 6730 14260 6736 14272
rect 5552 14232 6736 14260
rect 3660 14220 3666 14232
rect 6730 14220 6736 14232
rect 6788 14220 6794 14272
rect 7742 14260 7748 14272
rect 7703 14232 7748 14260
rect 7742 14220 7748 14232
rect 7800 14220 7806 14272
rect 8036 14260 8064 14427
rect 8846 14424 8852 14436
rect 8904 14464 8910 14476
rect 9214 14464 9220 14476
rect 8904 14436 9220 14464
rect 8904 14424 8910 14436
rect 9214 14424 9220 14436
rect 9272 14424 9278 14476
rect 9950 14464 9956 14476
rect 9911 14436 9956 14464
rect 9950 14424 9956 14436
rect 10008 14424 10014 14476
rect 10597 14467 10655 14473
rect 10597 14433 10609 14467
rect 10643 14464 10655 14467
rect 10686 14464 10692 14476
rect 10643 14436 10692 14464
rect 10643 14433 10655 14436
rect 10597 14427 10655 14433
rect 10686 14424 10692 14436
rect 10744 14424 10750 14476
rect 10870 14473 10876 14476
rect 10864 14464 10876 14473
rect 10831 14436 10876 14464
rect 10864 14427 10876 14436
rect 10870 14424 10876 14427
rect 10928 14424 10934 14476
rect 11238 14424 11244 14476
rect 11296 14464 11302 14476
rect 11296 14436 12204 14464
rect 11296 14424 11302 14436
rect 12176 14408 12204 14436
rect 12250 14424 12256 14476
rect 12308 14424 12314 14476
rect 12621 14467 12679 14473
rect 12621 14433 12633 14467
rect 12667 14464 12679 14467
rect 12710 14464 12716 14476
rect 12667 14436 12716 14464
rect 12667 14433 12679 14436
rect 12621 14427 12679 14433
rect 12710 14424 12716 14436
rect 12768 14424 12774 14476
rect 13832 14464 13860 14504
rect 14752 14476 14780 14504
rect 13464 14436 13860 14464
rect 14461 14467 14519 14473
rect 9769 14399 9827 14405
rect 9769 14365 9781 14399
rect 9815 14396 9827 14399
rect 12158 14396 12164 14408
rect 9815 14368 10640 14396
rect 12071 14368 12164 14396
rect 9815 14365 9827 14368
rect 9769 14359 9827 14365
rect 8665 14331 8723 14337
rect 8665 14297 8677 14331
rect 8711 14328 8723 14331
rect 10042 14328 10048 14340
rect 8711 14300 10048 14328
rect 8711 14297 8723 14300
rect 8665 14291 8723 14297
rect 10042 14288 10048 14300
rect 10100 14288 10106 14340
rect 10321 14331 10379 14337
rect 10321 14297 10333 14331
rect 10367 14328 10379 14331
rect 10410 14328 10416 14340
rect 10367 14300 10416 14328
rect 10367 14297 10379 14300
rect 10321 14291 10379 14297
rect 10410 14288 10416 14300
rect 10468 14288 10474 14340
rect 10134 14260 10140 14272
rect 8036 14232 10140 14260
rect 10134 14220 10140 14232
rect 10192 14220 10198 14272
rect 10612 14260 10640 14368
rect 12158 14356 12164 14368
rect 12216 14396 12222 14408
rect 13464 14405 13492 14436
rect 14461 14433 14473 14467
rect 14507 14464 14519 14467
rect 14553 14467 14611 14473
rect 14553 14464 14565 14467
rect 14507 14436 14565 14464
rect 14507 14433 14519 14436
rect 14461 14427 14519 14433
rect 14553 14433 14565 14436
rect 14599 14433 14611 14467
rect 14553 14427 14611 14433
rect 14734 14424 14740 14476
rect 14792 14424 14798 14476
rect 12805 14399 12863 14405
rect 12805 14396 12817 14399
rect 12216 14368 12817 14396
rect 12216 14356 12222 14368
rect 12805 14365 12817 14368
rect 12851 14365 12863 14399
rect 12805 14359 12863 14365
rect 13449 14399 13507 14405
rect 13449 14365 13461 14399
rect 13495 14365 13507 14399
rect 13449 14359 13507 14365
rect 13538 14356 13544 14408
rect 13596 14396 13602 14408
rect 15580 14396 15608 14504
rect 16942 14492 16948 14504
rect 17000 14532 17006 14544
rect 17037 14535 17095 14541
rect 17037 14532 17049 14535
rect 17000 14504 17049 14532
rect 17000 14492 17006 14504
rect 17037 14501 17049 14504
rect 17083 14501 17095 14535
rect 17037 14495 17095 14501
rect 15654 14424 15660 14476
rect 15712 14464 15718 14476
rect 16494 14467 16552 14473
rect 16494 14464 16506 14467
rect 15712 14436 16506 14464
rect 15712 14424 15718 14436
rect 16494 14433 16506 14436
rect 16540 14433 16552 14467
rect 16758 14464 16764 14476
rect 16719 14436 16764 14464
rect 16494 14427 16552 14433
rect 16758 14424 16764 14436
rect 16816 14424 16822 14476
rect 13596 14368 15608 14396
rect 17865 14399 17923 14405
rect 13596 14356 13602 14368
rect 17865 14365 17877 14399
rect 17911 14396 17923 14399
rect 19058 14396 19064 14408
rect 17911 14368 19064 14396
rect 17911 14365 17923 14368
rect 17865 14359 17923 14365
rect 19058 14356 19064 14368
rect 19116 14356 19122 14408
rect 13170 14288 13176 14340
rect 13228 14328 13234 14340
rect 14461 14331 14519 14337
rect 14461 14328 14473 14331
rect 13228 14300 14473 14328
rect 13228 14288 13234 14300
rect 14461 14297 14473 14300
rect 14507 14297 14519 14331
rect 14461 14291 14519 14297
rect 11974 14260 11980 14272
rect 10612 14232 11980 14260
rect 11974 14220 11980 14232
rect 12032 14220 12038 14272
rect 12066 14220 12072 14272
rect 12124 14260 12130 14272
rect 14274 14260 14280 14272
rect 12124 14232 14280 14260
rect 12124 14220 12130 14232
rect 14274 14220 14280 14232
rect 14332 14220 14338 14272
rect 14366 14220 14372 14272
rect 14424 14260 14430 14272
rect 15194 14260 15200 14272
rect 14424 14232 15200 14260
rect 14424 14220 14430 14232
rect 15194 14220 15200 14232
rect 15252 14260 15258 14272
rect 15470 14260 15476 14272
rect 15252 14232 15476 14260
rect 15252 14220 15258 14232
rect 15470 14220 15476 14232
rect 15528 14220 15534 14272
rect 1104 14170 21896 14192
rect 1104 14118 4447 14170
rect 4499 14118 4511 14170
rect 4563 14118 4575 14170
rect 4627 14118 4639 14170
rect 4691 14118 11378 14170
rect 11430 14118 11442 14170
rect 11494 14118 11506 14170
rect 11558 14118 11570 14170
rect 11622 14118 18308 14170
rect 18360 14118 18372 14170
rect 18424 14118 18436 14170
rect 18488 14118 18500 14170
rect 18552 14118 21896 14170
rect 1104 14096 21896 14118
rect 2038 14016 2044 14068
rect 2096 14056 2102 14068
rect 2133 14059 2191 14065
rect 2133 14056 2145 14059
rect 2096 14028 2145 14056
rect 2096 14016 2102 14028
rect 2133 14025 2145 14028
rect 2179 14025 2191 14059
rect 2133 14019 2191 14025
rect 2314 14016 2320 14068
rect 2372 14056 2378 14068
rect 2593 14059 2651 14065
rect 2593 14056 2605 14059
rect 2372 14028 2605 14056
rect 2372 14016 2378 14028
rect 2593 14025 2605 14028
rect 2639 14025 2651 14059
rect 2593 14019 2651 14025
rect 3789 14059 3847 14065
rect 3789 14025 3801 14059
rect 3835 14056 3847 14059
rect 4338 14056 4344 14068
rect 3835 14028 4344 14056
rect 3835 14025 3847 14028
rect 3789 14019 3847 14025
rect 4338 14016 4344 14028
rect 4396 14016 4402 14068
rect 4709 14059 4767 14065
rect 4709 14025 4721 14059
rect 4755 14056 4767 14059
rect 5902 14056 5908 14068
rect 4755 14028 5908 14056
rect 4755 14025 4767 14028
rect 4709 14019 4767 14025
rect 5902 14016 5908 14028
rect 5960 14016 5966 14068
rect 6638 14056 6644 14068
rect 6599 14028 6644 14056
rect 6638 14016 6644 14028
rect 6696 14016 6702 14068
rect 6730 14016 6736 14068
rect 6788 14056 6794 14068
rect 7653 14059 7711 14065
rect 7653 14056 7665 14059
rect 6788 14028 7665 14056
rect 6788 14016 6794 14028
rect 7653 14025 7665 14028
rect 7699 14025 7711 14059
rect 9674 14056 9680 14068
rect 7653 14019 7711 14025
rect 8036 14028 9680 14056
rect 4249 13991 4307 13997
rect 4249 13957 4261 13991
rect 4295 13988 4307 13991
rect 5074 13988 5080 14000
rect 4295 13960 5080 13988
rect 4295 13957 4307 13960
rect 4249 13951 4307 13957
rect 5074 13948 5080 13960
rect 5132 13948 5138 14000
rect 6086 13948 6092 14000
rect 6144 13988 6150 14000
rect 8036 13988 8064 14028
rect 9674 14016 9680 14028
rect 9732 14016 9738 14068
rect 9769 14059 9827 14065
rect 9769 14025 9781 14059
rect 9815 14056 9827 14059
rect 9858 14056 9864 14068
rect 9815 14028 9864 14056
rect 9815 14025 9827 14028
rect 9769 14019 9827 14025
rect 9858 14016 9864 14028
rect 9916 14016 9922 14068
rect 12066 14056 12072 14068
rect 9968 14028 12072 14056
rect 6144 13960 8064 13988
rect 8113 13991 8171 13997
rect 6144 13948 6150 13960
rect 8113 13957 8125 13991
rect 8159 13988 8171 13991
rect 8202 13988 8208 14000
rect 8159 13960 8208 13988
rect 8159 13957 8171 13960
rect 8113 13951 8171 13957
rect 8202 13948 8208 13960
rect 8260 13948 8266 14000
rect 9490 13948 9496 14000
rect 9548 13948 9554 14000
rect 3142 13920 3148 13932
rect 3103 13892 3148 13920
rect 3142 13880 3148 13892
rect 3200 13880 3206 13932
rect 3528 13892 5028 13920
rect 1578 13852 1584 13864
rect 1539 13824 1584 13852
rect 1578 13812 1584 13824
rect 1636 13812 1642 13864
rect 1762 13852 1768 13864
rect 1723 13824 1768 13852
rect 1762 13812 1768 13824
rect 1820 13812 1826 13864
rect 2314 13852 2320 13864
rect 2275 13824 2320 13852
rect 2314 13812 2320 13824
rect 2372 13812 2378 13864
rect 2777 13855 2835 13861
rect 2777 13821 2789 13855
rect 2823 13852 2835 13855
rect 3528 13852 3556 13892
rect 2823 13824 3556 13852
rect 2823 13821 2835 13824
rect 2777 13815 2835 13821
rect 3602 13812 3608 13864
rect 3660 13852 3666 13864
rect 4062 13852 4068 13864
rect 3660 13824 3705 13852
rect 4023 13824 4068 13852
rect 3660 13812 3666 13824
rect 4062 13812 4068 13824
rect 4120 13812 4126 13864
rect 5000 13716 5028 13892
rect 6914 13880 6920 13932
rect 6972 13920 6978 13932
rect 7285 13923 7343 13929
rect 7285 13920 7297 13923
rect 6972 13892 7297 13920
rect 6972 13880 6978 13892
rect 7285 13889 7297 13892
rect 7331 13920 7343 13923
rect 7742 13920 7748 13932
rect 7331 13892 7748 13920
rect 7331 13889 7343 13892
rect 7285 13883 7343 13889
rect 7742 13880 7748 13892
rect 7800 13880 7806 13932
rect 9501 13920 9529 13948
rect 9968 13920 9996 14028
rect 12066 14016 12072 14028
rect 12124 14016 12130 14068
rect 13722 14016 13728 14068
rect 13780 14056 13786 14068
rect 13909 14059 13967 14065
rect 13909 14056 13921 14059
rect 13780 14028 13921 14056
rect 13780 14016 13786 14028
rect 13909 14025 13921 14028
rect 13955 14025 13967 14059
rect 13909 14019 13967 14025
rect 14016 14028 15332 14056
rect 13262 13948 13268 14000
rect 13320 13988 13326 14000
rect 14016 13988 14044 14028
rect 13320 13960 14044 13988
rect 13320 13948 13326 13960
rect 12710 13920 12716 13932
rect 9501 13892 9996 13920
rect 11072 13892 12716 13920
rect 5994 13812 6000 13864
rect 6052 13852 6058 13864
rect 6089 13855 6147 13861
rect 6089 13852 6101 13855
rect 6052 13824 6101 13852
rect 6052 13812 6058 13824
rect 6089 13821 6101 13824
rect 6135 13821 6147 13855
rect 6089 13815 6147 13821
rect 9398 13812 9404 13864
rect 9456 13852 9462 13864
rect 9493 13855 9551 13861
rect 9493 13852 9505 13855
rect 9456 13824 9505 13852
rect 9456 13812 9462 13824
rect 9493 13821 9505 13824
rect 9539 13821 9551 13855
rect 10882 13855 10940 13861
rect 10882 13852 10894 13855
rect 9493 13815 9551 13821
rect 9646 13824 10894 13852
rect 9646 13796 9674 13824
rect 10882 13821 10894 13824
rect 10928 13821 10940 13855
rect 11072 13852 11100 13892
rect 12710 13880 12716 13892
rect 12768 13920 12774 13932
rect 14274 13920 14280 13932
rect 12768 13892 14280 13920
rect 12768 13880 12774 13892
rect 14274 13880 14280 13892
rect 14332 13880 14338 13932
rect 15304 13929 15332 14028
rect 16114 14016 16120 14068
rect 16172 14056 16178 14068
rect 16301 14059 16359 14065
rect 16301 14056 16313 14059
rect 16172 14028 16313 14056
rect 16172 14016 16178 14028
rect 16301 14025 16313 14028
rect 16347 14025 16359 14059
rect 20714 14056 20720 14068
rect 16301 14019 16359 14025
rect 17144 14028 20720 14056
rect 15289 13923 15347 13929
rect 15289 13889 15301 13923
rect 15335 13889 15347 13923
rect 15654 13920 15660 13932
rect 15615 13892 15660 13920
rect 15289 13883 15347 13889
rect 15654 13880 15660 13892
rect 15712 13880 15718 13932
rect 15838 13920 15844 13932
rect 15799 13892 15844 13920
rect 15838 13880 15844 13892
rect 15896 13880 15902 13932
rect 10882 13815 10940 13821
rect 10980 13824 11100 13852
rect 11149 13855 11207 13861
rect 5534 13744 5540 13796
rect 5592 13784 5598 13796
rect 5822 13787 5880 13793
rect 5822 13784 5834 13787
rect 5592 13756 5834 13784
rect 5592 13744 5598 13756
rect 5822 13753 5834 13756
rect 5868 13753 5880 13787
rect 7006 13784 7012 13796
rect 6967 13756 7012 13784
rect 5822 13747 5880 13753
rect 7006 13744 7012 13756
rect 7064 13744 7070 13796
rect 7098 13744 7104 13796
rect 7156 13784 7162 13796
rect 7156 13756 7201 13784
rect 7156 13744 7162 13756
rect 9122 13744 9128 13796
rect 9180 13784 9186 13796
rect 9237 13787 9295 13793
rect 9237 13784 9249 13787
rect 9180 13756 9249 13784
rect 9180 13744 9186 13756
rect 9237 13753 9249 13756
rect 9283 13753 9295 13787
rect 9237 13747 9295 13753
rect 9628 13744 9634 13796
rect 9686 13744 9692 13796
rect 10594 13744 10600 13796
rect 10652 13784 10658 13796
rect 10980 13784 11008 13824
rect 11149 13821 11161 13855
rect 11195 13852 11207 13855
rect 13262 13852 13268 13864
rect 11195 13824 13268 13852
rect 11195 13821 11207 13824
rect 11149 13815 11207 13821
rect 13262 13812 13268 13824
rect 13320 13812 13326 13864
rect 13633 13855 13691 13861
rect 13633 13821 13645 13855
rect 13679 13852 13691 13855
rect 13679 13824 14688 13852
rect 13679 13821 13691 13824
rect 13633 13815 13691 13821
rect 14660 13784 14688 13824
rect 14734 13812 14740 13864
rect 14792 13852 14798 13864
rect 15022 13855 15080 13861
rect 15022 13852 15034 13855
rect 14792 13824 15034 13852
rect 14792 13812 14798 13824
rect 15022 13821 15034 13824
rect 15068 13821 15080 13855
rect 17144 13852 17172 14028
rect 20714 14016 20720 14028
rect 20772 14016 20778 14068
rect 17402 13988 17408 14000
rect 17363 13960 17408 13988
rect 17402 13948 17408 13960
rect 17460 13988 17466 14000
rect 18046 13988 18052 14000
rect 17460 13960 18052 13988
rect 17460 13948 17466 13960
rect 18046 13948 18052 13960
rect 18104 13948 18110 14000
rect 15022 13815 15080 13821
rect 15120 13824 17172 13852
rect 18897 13855 18955 13861
rect 15120 13784 15148 13824
rect 18897 13821 18909 13855
rect 18943 13852 18955 13855
rect 19058 13852 19064 13864
rect 18943 13824 19064 13852
rect 18943 13821 18955 13824
rect 18897 13815 18955 13821
rect 19058 13812 19064 13824
rect 19116 13812 19122 13864
rect 19153 13855 19211 13861
rect 19153 13821 19165 13855
rect 19199 13852 19211 13855
rect 19242 13852 19248 13864
rect 19199 13824 19248 13852
rect 19199 13821 19211 13824
rect 19153 13815 19211 13821
rect 19242 13812 19248 13824
rect 19300 13812 19306 13864
rect 15933 13787 15991 13793
rect 15933 13784 15945 13787
rect 10652 13756 11008 13784
rect 11072 13756 13584 13784
rect 14660 13756 15148 13784
rect 15764 13756 15945 13784
rect 10652 13744 10658 13756
rect 6822 13716 6828 13728
rect 5000 13688 6828 13716
rect 6822 13676 6828 13688
rect 6880 13676 6886 13728
rect 7466 13676 7472 13728
rect 7524 13716 7530 13728
rect 11072 13716 11100 13756
rect 7524 13688 11100 13716
rect 12345 13719 12403 13725
rect 7524 13676 7530 13688
rect 12345 13685 12357 13719
rect 12391 13716 12403 13719
rect 12526 13716 12532 13728
rect 12391 13688 12532 13716
rect 12391 13685 12403 13688
rect 12345 13679 12403 13685
rect 12526 13676 12532 13688
rect 12584 13716 12590 13728
rect 13170 13716 13176 13728
rect 12584 13688 13176 13716
rect 12584 13676 12590 13688
rect 13170 13676 13176 13688
rect 13228 13676 13234 13728
rect 13556 13716 13584 13756
rect 15470 13716 15476 13728
rect 13556 13688 15476 13716
rect 15470 13676 15476 13688
rect 15528 13716 15534 13728
rect 15764 13716 15792 13756
rect 15933 13753 15945 13756
rect 15979 13753 15991 13787
rect 15933 13747 15991 13753
rect 17770 13716 17776 13728
rect 15528 13688 15792 13716
rect 17731 13688 17776 13716
rect 15528 13676 15534 13688
rect 17770 13676 17776 13688
rect 17828 13676 17834 13728
rect 1104 13626 21896 13648
rect 1104 13574 7912 13626
rect 7964 13574 7976 13626
rect 8028 13574 8040 13626
rect 8092 13574 8104 13626
rect 8156 13574 14843 13626
rect 14895 13574 14907 13626
rect 14959 13574 14971 13626
rect 15023 13574 15035 13626
rect 15087 13574 21896 13626
rect 1104 13552 21896 13574
rect 2225 13515 2283 13521
rect 2225 13481 2237 13515
rect 2271 13512 2283 13515
rect 2314 13512 2320 13524
rect 2271 13484 2320 13512
rect 2271 13481 2283 13484
rect 2225 13475 2283 13481
rect 2314 13472 2320 13484
rect 2372 13472 2378 13524
rect 2501 13515 2559 13521
rect 2501 13481 2513 13515
rect 2547 13512 2559 13515
rect 2590 13512 2596 13524
rect 2547 13484 2596 13512
rect 2547 13481 2559 13484
rect 2501 13475 2559 13481
rect 2590 13472 2596 13484
rect 2648 13472 2654 13524
rect 4341 13515 4399 13521
rect 4341 13512 4353 13515
rect 2746 13484 4353 13512
rect 2746 13444 2774 13484
rect 4341 13481 4353 13484
rect 4387 13481 4399 13515
rect 4341 13475 4399 13481
rect 4801 13515 4859 13521
rect 4801 13481 4813 13515
rect 4847 13512 4859 13515
rect 5353 13515 5411 13521
rect 5353 13512 5365 13515
rect 4847 13484 5365 13512
rect 4847 13481 4859 13484
rect 4801 13475 4859 13481
rect 5353 13481 5365 13484
rect 5399 13481 5411 13515
rect 5353 13475 5411 13481
rect 5813 13515 5871 13521
rect 5813 13481 5825 13515
rect 5859 13512 5871 13515
rect 8386 13512 8392 13524
rect 5859 13484 8392 13512
rect 5859 13481 5871 13484
rect 5813 13475 5871 13481
rect 8386 13472 8392 13484
rect 8444 13472 8450 13524
rect 8481 13515 8539 13521
rect 8481 13481 8493 13515
rect 8527 13512 8539 13515
rect 9309 13515 9367 13521
rect 9309 13512 9321 13515
rect 8527 13484 9321 13512
rect 8527 13481 8539 13484
rect 8481 13475 8539 13481
rect 9309 13481 9321 13484
rect 9355 13481 9367 13515
rect 9309 13475 9367 13481
rect 9950 13472 9956 13524
rect 10008 13512 10014 13524
rect 10873 13515 10931 13521
rect 10873 13512 10885 13515
rect 10008 13484 10885 13512
rect 10008 13472 10014 13484
rect 10873 13481 10885 13484
rect 10919 13481 10931 13515
rect 11882 13512 11888 13524
rect 11843 13484 11888 13512
rect 10873 13475 10931 13481
rect 11882 13472 11888 13484
rect 11940 13472 11946 13524
rect 12342 13512 12348 13524
rect 12303 13484 12348 13512
rect 12342 13472 12348 13484
rect 12400 13472 12406 13524
rect 12434 13472 12440 13524
rect 12492 13512 12498 13524
rect 13173 13515 13231 13521
rect 13173 13512 13185 13515
rect 12492 13484 13185 13512
rect 12492 13472 12498 13484
rect 13173 13481 13185 13484
rect 13219 13481 13231 13515
rect 15470 13512 15476 13524
rect 15431 13484 15476 13512
rect 13173 13475 13231 13481
rect 15470 13472 15476 13484
rect 15528 13472 15534 13524
rect 16117 13515 16175 13521
rect 16117 13481 16129 13515
rect 16163 13512 16175 13515
rect 16206 13512 16212 13524
rect 16163 13484 16212 13512
rect 16163 13481 16175 13484
rect 16117 13475 16175 13481
rect 16206 13472 16212 13484
rect 16264 13472 16270 13524
rect 16574 13512 16580 13524
rect 16535 13484 16580 13512
rect 16574 13472 16580 13484
rect 16632 13472 16638 13524
rect 2056 13416 2774 13444
rect 1486 13336 1492 13388
rect 1544 13376 1550 13388
rect 2056 13385 2084 13416
rect 3142 13404 3148 13456
rect 3200 13444 3206 13456
rect 3421 13447 3479 13453
rect 3421 13444 3433 13447
rect 3200 13416 3433 13444
rect 3200 13404 3206 13416
rect 3421 13413 3433 13416
rect 3467 13413 3479 13447
rect 3421 13407 3479 13413
rect 4709 13447 4767 13453
rect 4709 13413 4721 13447
rect 4755 13444 4767 13447
rect 6365 13447 6423 13453
rect 6365 13444 6377 13447
rect 4755 13416 6377 13444
rect 4755 13413 4767 13416
rect 4709 13407 4767 13413
rect 6365 13413 6377 13416
rect 6411 13413 6423 13447
rect 8938 13444 8944 13456
rect 6365 13407 6423 13413
rect 6932 13416 8944 13444
rect 1581 13379 1639 13385
rect 1581 13376 1593 13379
rect 1544 13348 1593 13376
rect 1544 13336 1550 13348
rect 1581 13345 1593 13348
rect 1627 13345 1639 13379
rect 1581 13339 1639 13345
rect 2041 13379 2099 13385
rect 2041 13345 2053 13379
rect 2087 13345 2099 13379
rect 2041 13339 2099 13345
rect 2685 13379 2743 13385
rect 2685 13345 2697 13379
rect 2731 13376 2743 13379
rect 2774 13376 2780 13388
rect 2731 13348 2780 13376
rect 2731 13345 2743 13348
rect 2685 13339 2743 13345
rect 2774 13336 2780 13348
rect 2832 13336 2838 13388
rect 2866 13336 2872 13388
rect 2924 13376 2930 13388
rect 2961 13379 3019 13385
rect 2961 13376 2973 13379
rect 2924 13348 2973 13376
rect 2924 13336 2930 13348
rect 2961 13345 2973 13348
rect 3007 13376 3019 13379
rect 3881 13379 3939 13385
rect 3881 13376 3893 13379
rect 3007 13348 3893 13376
rect 3007 13345 3019 13348
rect 2961 13339 3019 13345
rect 3881 13345 3893 13348
rect 3927 13345 3939 13379
rect 3881 13339 3939 13345
rect 5721 13379 5779 13385
rect 5721 13345 5733 13379
rect 5767 13376 5779 13379
rect 6932 13376 6960 13416
rect 8938 13404 8944 13416
rect 8996 13444 9002 13456
rect 9677 13447 9735 13453
rect 9677 13444 9689 13447
rect 8996 13416 9689 13444
rect 8996 13404 9002 13416
rect 9677 13413 9689 13416
rect 9723 13413 9735 13447
rect 9677 13407 9735 13413
rect 9769 13447 9827 13453
rect 9769 13413 9781 13447
rect 9815 13444 9827 13447
rect 10778 13444 10784 13456
rect 9815 13416 10784 13444
rect 9815 13413 9827 13416
rect 9769 13407 9827 13413
rect 10778 13404 10784 13416
rect 10836 13404 10842 13456
rect 11241 13447 11299 13453
rect 11241 13413 11253 13447
rect 11287 13444 11299 13447
rect 15013 13447 15071 13453
rect 15013 13444 15025 13447
rect 11287 13416 15025 13444
rect 11287 13413 11299 13416
rect 11241 13407 11299 13413
rect 15013 13413 15025 13416
rect 15059 13413 15071 13447
rect 15013 13407 15071 13413
rect 17218 13404 17224 13456
rect 17276 13444 17282 13456
rect 17313 13447 17371 13453
rect 17313 13444 17325 13447
rect 17276 13416 17325 13444
rect 17276 13404 17282 13416
rect 17313 13413 17325 13416
rect 17359 13444 17371 13447
rect 17865 13447 17923 13453
rect 17865 13444 17877 13447
rect 17359 13416 17877 13444
rect 17359 13413 17371 13416
rect 17313 13407 17371 13413
rect 17865 13413 17877 13416
rect 17911 13413 17923 13447
rect 17865 13407 17923 13413
rect 5767 13348 6960 13376
rect 7009 13379 7067 13385
rect 5767 13345 5779 13348
rect 5721 13339 5779 13345
rect 7009 13345 7021 13379
rect 7055 13345 7067 13379
rect 7009 13339 7067 13345
rect 7745 13379 7803 13385
rect 7745 13345 7757 13379
rect 7791 13376 7803 13379
rect 8389 13379 8447 13385
rect 8389 13376 8401 13379
rect 7791 13348 8401 13376
rect 7791 13345 7803 13348
rect 7745 13339 7803 13345
rect 8389 13345 8401 13348
rect 8435 13345 8447 13379
rect 10226 13376 10232 13388
rect 8389 13339 8447 13345
rect 8496 13348 10232 13376
rect 4985 13311 5043 13317
rect 4985 13277 4997 13311
rect 5031 13308 5043 13311
rect 5534 13308 5540 13320
rect 5031 13280 5540 13308
rect 5031 13277 5043 13280
rect 4985 13271 5043 13277
rect 5534 13268 5540 13280
rect 5592 13268 5598 13320
rect 5902 13268 5908 13320
rect 5960 13308 5966 13320
rect 5960 13280 6005 13308
rect 5960 13268 5966 13280
rect 6454 13268 6460 13320
rect 6512 13308 6518 13320
rect 7024 13308 7052 13339
rect 8496 13308 8524 13348
rect 10226 13336 10232 13348
rect 10284 13336 10290 13388
rect 10870 13336 10876 13388
rect 10928 13376 10934 13388
rect 10928 13348 11468 13376
rect 10928 13336 10934 13348
rect 6512 13280 6940 13308
rect 7024 13280 8524 13308
rect 8665 13311 8723 13317
rect 6512 13268 6518 13280
rect 1765 13243 1823 13249
rect 1765 13209 1777 13243
rect 1811 13240 1823 13243
rect 3145 13243 3203 13249
rect 1811 13212 2774 13240
rect 1811 13209 1823 13212
rect 1765 13203 1823 13209
rect 2746 13172 2774 13212
rect 3145 13209 3157 13243
rect 3191 13240 3203 13243
rect 6638 13240 6644 13252
rect 3191 13212 6644 13240
rect 3191 13209 3203 13212
rect 3145 13203 3203 13209
rect 6638 13200 6644 13212
rect 6696 13200 6702 13252
rect 6825 13243 6883 13249
rect 6825 13209 6837 13243
rect 6871 13240 6883 13243
rect 6912 13240 6940 13280
rect 8665 13277 8677 13311
rect 8711 13308 8723 13311
rect 9490 13308 9496 13320
rect 8711 13280 9496 13308
rect 8711 13277 8723 13280
rect 8665 13271 8723 13277
rect 6871 13212 6940 13240
rect 6871 13209 6883 13212
rect 6825 13203 6883 13209
rect 8202 13200 8208 13252
rect 8260 13240 8266 13252
rect 8680 13240 8708 13271
rect 9490 13268 9496 13280
rect 9548 13268 9554 13320
rect 11440 13317 11468 13348
rect 11790 13336 11796 13388
rect 11848 13376 11854 13388
rect 12253 13379 12311 13385
rect 12253 13376 12265 13379
rect 11848 13348 12265 13376
rect 11848 13336 11854 13348
rect 12253 13345 12265 13348
rect 12299 13345 12311 13379
rect 12253 13339 12311 13345
rect 13541 13379 13599 13385
rect 13541 13345 13553 13379
rect 13587 13376 13599 13379
rect 14553 13379 14611 13385
rect 14553 13376 14565 13379
rect 13587 13348 14565 13376
rect 13587 13345 13599 13348
rect 13541 13339 13599 13345
rect 14553 13345 14565 13348
rect 14599 13345 14611 13379
rect 17954 13376 17960 13388
rect 17915 13348 17960 13376
rect 14553 13339 14611 13345
rect 17954 13336 17960 13348
rect 18012 13336 18018 13388
rect 9861 13311 9919 13317
rect 9861 13277 9873 13311
rect 9907 13277 9919 13311
rect 9861 13271 9919 13277
rect 11333 13311 11391 13317
rect 11333 13277 11345 13311
rect 11379 13277 11391 13311
rect 11333 13271 11391 13277
rect 11425 13311 11483 13317
rect 11425 13277 11437 13311
rect 11471 13277 11483 13311
rect 11425 13271 11483 13277
rect 8260 13212 8708 13240
rect 8260 13200 8266 13212
rect 9122 13200 9128 13252
rect 9180 13240 9186 13252
rect 9876 13240 9904 13271
rect 9180 13212 9904 13240
rect 9180 13200 9186 13212
rect 10134 13200 10140 13252
rect 10192 13240 10198 13252
rect 10321 13243 10379 13249
rect 10321 13240 10333 13243
rect 10192 13212 10333 13240
rect 10192 13200 10198 13212
rect 10321 13209 10333 13212
rect 10367 13209 10379 13243
rect 10321 13203 10379 13209
rect 6730 13172 6736 13184
rect 2746 13144 6736 13172
rect 6730 13132 6736 13144
rect 6788 13132 6794 13184
rect 6914 13132 6920 13184
rect 6972 13172 6978 13184
rect 8021 13175 8079 13181
rect 8021 13172 8033 13175
rect 6972 13144 8033 13172
rect 6972 13132 6978 13144
rect 8021 13141 8033 13144
rect 8067 13141 8079 13175
rect 8021 13135 8079 13141
rect 8110 13132 8116 13184
rect 8168 13172 8174 13184
rect 11348 13172 11376 13271
rect 12158 13268 12164 13320
rect 12216 13308 12222 13320
rect 12437 13311 12495 13317
rect 12437 13308 12449 13311
rect 12216 13280 12449 13308
rect 12216 13268 12222 13280
rect 12437 13277 12449 13280
rect 12483 13277 12495 13311
rect 13630 13308 13636 13320
rect 13591 13280 13636 13308
rect 12437 13271 12495 13277
rect 13630 13268 13636 13280
rect 13688 13268 13694 13320
rect 13722 13268 13728 13320
rect 13780 13308 13786 13320
rect 17770 13308 17776 13320
rect 13780 13280 13825 13308
rect 17731 13280 17776 13308
rect 13780 13268 13786 13280
rect 17770 13268 17776 13280
rect 17828 13268 17834 13320
rect 8168 13144 11376 13172
rect 8168 13132 8174 13144
rect 13998 13132 14004 13184
rect 14056 13172 14062 13184
rect 17586 13172 17592 13184
rect 14056 13144 17592 13172
rect 14056 13132 14062 13144
rect 17586 13132 17592 13144
rect 17644 13132 17650 13184
rect 18325 13175 18383 13181
rect 18325 13141 18337 13175
rect 18371 13172 18383 13175
rect 18966 13172 18972 13184
rect 18371 13144 18972 13172
rect 18371 13141 18383 13144
rect 18325 13135 18383 13141
rect 18966 13132 18972 13144
rect 19024 13132 19030 13184
rect 1104 13082 21896 13104
rect 1104 13030 4447 13082
rect 4499 13030 4511 13082
rect 4563 13030 4575 13082
rect 4627 13030 4639 13082
rect 4691 13030 11378 13082
rect 11430 13030 11442 13082
rect 11494 13030 11506 13082
rect 11558 13030 11570 13082
rect 11622 13030 18308 13082
rect 18360 13030 18372 13082
rect 18424 13030 18436 13082
rect 18488 13030 18500 13082
rect 18552 13030 21896 13082
rect 1104 13008 21896 13030
rect 1486 12968 1492 12980
rect 1447 12940 1492 12968
rect 1486 12928 1492 12940
rect 1544 12928 1550 12980
rect 1765 12971 1823 12977
rect 1765 12937 1777 12971
rect 1811 12968 1823 12971
rect 1854 12968 1860 12980
rect 1811 12940 1860 12968
rect 1811 12937 1823 12940
rect 1765 12931 1823 12937
rect 1854 12928 1860 12940
rect 1912 12928 1918 12980
rect 2225 12971 2283 12977
rect 2225 12937 2237 12971
rect 2271 12968 2283 12971
rect 2406 12968 2412 12980
rect 2271 12940 2412 12968
rect 2271 12937 2283 12940
rect 2225 12931 2283 12937
rect 2406 12928 2412 12940
rect 2464 12928 2470 12980
rect 6733 12971 6791 12977
rect 6733 12968 6745 12971
rect 4724 12940 6745 12968
rect 4724 12912 4752 12940
rect 6733 12937 6745 12940
rect 6779 12937 6791 12971
rect 6733 12931 6791 12937
rect 6822 12928 6828 12980
rect 6880 12968 6886 12980
rect 9122 12968 9128 12980
rect 6880 12940 8800 12968
rect 9083 12940 9128 12968
rect 6880 12928 6886 12940
rect 4706 12860 4712 12912
rect 4764 12860 4770 12912
rect 5994 12832 6000 12844
rect 4264 12804 4936 12832
rect 5955 12804 6000 12832
rect 1949 12767 2007 12773
rect 1949 12733 1961 12767
rect 1995 12733 2007 12767
rect 2406 12764 2412 12776
rect 2367 12736 2412 12764
rect 1949 12727 2007 12733
rect 1964 12696 1992 12727
rect 2406 12724 2412 12736
rect 2464 12724 2470 12776
rect 2590 12724 2596 12776
rect 2648 12764 2654 12776
rect 4264 12764 4292 12804
rect 2648 12736 4292 12764
rect 4341 12767 4399 12773
rect 2648 12724 2654 12736
rect 4341 12733 4353 12767
rect 4387 12764 4399 12767
rect 4798 12764 4804 12776
rect 4387 12736 4804 12764
rect 4387 12733 4399 12736
rect 4341 12727 4399 12733
rect 4798 12724 4804 12736
rect 4856 12724 4862 12776
rect 4908 12764 4936 12804
rect 5994 12792 6000 12804
rect 6052 12832 6058 12844
rect 6822 12832 6828 12844
rect 6052 12804 6828 12832
rect 6052 12792 6058 12804
rect 6822 12792 6828 12804
rect 6880 12792 6886 12844
rect 7282 12832 7288 12844
rect 7243 12804 7288 12832
rect 7282 12792 7288 12804
rect 7340 12832 7346 12844
rect 7340 12804 7880 12832
rect 7340 12792 7346 12804
rect 5718 12764 5724 12776
rect 5776 12773 5782 12776
rect 5776 12767 5799 12773
rect 4908 12736 5580 12764
rect 5651 12736 5724 12764
rect 2682 12696 2688 12708
rect 1964 12668 2688 12696
rect 2682 12656 2688 12668
rect 2740 12656 2746 12708
rect 4096 12699 4154 12705
rect 4096 12665 4108 12699
rect 4142 12696 4154 12699
rect 4890 12696 4896 12708
rect 4142 12668 4896 12696
rect 4142 12665 4154 12668
rect 4096 12659 4154 12665
rect 4890 12656 4896 12668
rect 4948 12656 4954 12708
rect 5552 12696 5580 12736
rect 5718 12724 5724 12736
rect 5787 12764 5799 12767
rect 5902 12764 5908 12776
rect 5787 12736 5908 12764
rect 5787 12733 5799 12736
rect 5776 12727 5799 12733
rect 5776 12724 5782 12727
rect 5902 12724 5908 12736
rect 5960 12724 5966 12776
rect 7466 12764 7472 12776
rect 6012 12736 7472 12764
rect 6012 12696 6040 12736
rect 7466 12724 7472 12736
rect 7524 12724 7530 12776
rect 7742 12764 7748 12776
rect 7703 12736 7748 12764
rect 7742 12724 7748 12736
rect 7800 12724 7806 12776
rect 7852 12764 7880 12804
rect 8001 12767 8059 12773
rect 8001 12764 8013 12767
rect 7852 12736 8013 12764
rect 8001 12733 8013 12736
rect 8047 12733 8059 12767
rect 8001 12727 8059 12733
rect 5552 12668 6040 12696
rect 7101 12699 7159 12705
rect 7101 12665 7113 12699
rect 7147 12696 7159 12699
rect 7558 12696 7564 12708
rect 7147 12668 7564 12696
rect 7147 12665 7159 12668
rect 7101 12659 7159 12665
rect 7558 12656 7564 12668
rect 7616 12656 7622 12708
rect 8772 12696 8800 12940
rect 9122 12928 9128 12940
rect 9180 12928 9186 12980
rect 12526 12968 12532 12980
rect 9600 12940 12532 12968
rect 9600 12773 9628 12940
rect 12526 12928 12532 12940
rect 12584 12928 12590 12980
rect 13541 12971 13599 12977
rect 13541 12937 13553 12971
rect 13587 12968 13599 12971
rect 13630 12968 13636 12980
rect 13587 12940 13636 12968
rect 13587 12937 13599 12940
rect 13541 12931 13599 12937
rect 13630 12928 13636 12940
rect 13688 12928 13694 12980
rect 15013 12971 15071 12977
rect 15013 12937 15025 12971
rect 15059 12968 15071 12971
rect 15654 12968 15660 12980
rect 15059 12940 15660 12968
rect 15059 12937 15071 12940
rect 15013 12931 15071 12937
rect 15654 12928 15660 12940
rect 15712 12928 15718 12980
rect 18601 12971 18659 12977
rect 18601 12937 18613 12971
rect 18647 12968 18659 12971
rect 18782 12968 18788 12980
rect 18647 12940 18788 12968
rect 18647 12937 18659 12940
rect 18601 12931 18659 12937
rect 18782 12928 18788 12940
rect 18840 12928 18846 12980
rect 9766 12860 9772 12912
rect 9824 12900 9830 12912
rect 9861 12903 9919 12909
rect 9861 12900 9873 12903
rect 9824 12872 9873 12900
rect 9824 12860 9830 12872
rect 9861 12869 9873 12872
rect 9907 12900 9919 12903
rect 10042 12900 10048 12912
rect 9907 12872 10048 12900
rect 9907 12869 9919 12872
rect 9861 12863 9919 12869
rect 10042 12860 10048 12872
rect 10100 12860 10106 12912
rect 10594 12900 10600 12912
rect 10555 12872 10600 12900
rect 10594 12860 10600 12872
rect 10652 12860 10658 12912
rect 10965 12903 11023 12909
rect 10965 12869 10977 12903
rect 11011 12900 11023 12903
rect 12250 12900 12256 12912
rect 11011 12872 12256 12900
rect 11011 12869 11023 12872
rect 10965 12863 11023 12869
rect 12250 12860 12256 12872
rect 12308 12860 12314 12912
rect 14366 12900 14372 12912
rect 14200 12872 14372 12900
rect 13262 12832 13268 12844
rect 13223 12804 13268 12832
rect 13262 12792 13268 12804
rect 13320 12792 13326 12844
rect 13998 12832 14004 12844
rect 13959 12804 14004 12832
rect 13998 12792 14004 12804
rect 14056 12792 14062 12844
rect 14200 12841 14228 12872
rect 14366 12860 14372 12872
rect 14424 12900 14430 12912
rect 14734 12900 14740 12912
rect 14424 12872 14740 12900
rect 14424 12860 14430 12872
rect 14734 12860 14740 12872
rect 14792 12860 14798 12912
rect 14185 12835 14243 12841
rect 14185 12801 14197 12835
rect 14231 12801 14243 12835
rect 14185 12795 14243 12801
rect 16393 12835 16451 12841
rect 16393 12801 16405 12835
rect 16439 12832 16451 12835
rect 17310 12832 17316 12844
rect 16439 12804 17316 12832
rect 16439 12801 16451 12804
rect 16393 12795 16451 12801
rect 17310 12792 17316 12804
rect 17368 12792 17374 12844
rect 17770 12832 17776 12844
rect 17731 12804 17776 12832
rect 17770 12792 17776 12804
rect 17828 12792 17834 12844
rect 17865 12835 17923 12841
rect 17865 12801 17877 12835
rect 17911 12832 17923 12835
rect 18046 12832 18052 12844
rect 17911 12804 18052 12832
rect 17911 12801 17923 12804
rect 17865 12795 17923 12801
rect 18046 12792 18052 12804
rect 18104 12792 18110 12844
rect 19150 12832 19156 12844
rect 19111 12804 19156 12832
rect 19150 12792 19156 12804
rect 19208 12792 19214 12844
rect 9585 12767 9643 12773
rect 9585 12733 9597 12767
rect 9631 12733 9643 12767
rect 11698 12764 11704 12776
rect 9585 12727 9643 12733
rect 9692 12736 11704 12764
rect 9692 12696 9720 12736
rect 11698 12724 11704 12736
rect 11756 12724 11762 12776
rect 11974 12724 11980 12776
rect 12032 12764 12038 12776
rect 12998 12767 13056 12773
rect 12998 12764 13010 12767
rect 12032 12736 13010 12764
rect 12032 12724 12038 12736
rect 12998 12733 13010 12736
rect 13044 12733 13056 12767
rect 12998 12727 13056 12733
rect 13814 12724 13820 12776
rect 13872 12764 13878 12776
rect 13872 12736 14596 12764
rect 13872 12724 13878 12736
rect 13909 12699 13967 12705
rect 13909 12696 13921 12699
rect 8772 12668 9720 12696
rect 11256 12668 13921 12696
rect 2958 12628 2964 12640
rect 2919 12600 2964 12628
rect 2958 12588 2964 12600
rect 3016 12588 3022 12640
rect 4617 12631 4675 12637
rect 4617 12597 4629 12631
rect 4663 12628 4675 12631
rect 5534 12628 5540 12640
rect 4663 12600 5540 12628
rect 4663 12597 4675 12600
rect 4617 12591 4675 12597
rect 5534 12588 5540 12600
rect 5592 12588 5598 12640
rect 7190 12628 7196 12640
rect 7151 12600 7196 12628
rect 7190 12588 7196 12600
rect 7248 12588 7254 12640
rect 8754 12588 8760 12640
rect 8812 12628 8818 12640
rect 9401 12631 9459 12637
rect 9401 12628 9413 12631
rect 8812 12600 9413 12628
rect 8812 12588 8818 12600
rect 9401 12597 9413 12600
rect 9447 12597 9459 12631
rect 9401 12591 9459 12597
rect 11146 12588 11152 12640
rect 11204 12628 11210 12640
rect 11256 12637 11284 12668
rect 13909 12665 13921 12668
rect 13955 12665 13967 12699
rect 13909 12659 13967 12665
rect 11241 12631 11299 12637
rect 11241 12628 11253 12631
rect 11204 12600 11253 12628
rect 11204 12588 11210 12600
rect 11241 12597 11253 12600
rect 11287 12597 11299 12631
rect 11241 12591 11299 12597
rect 11790 12588 11796 12640
rect 11848 12628 11854 12640
rect 14568 12637 14596 12736
rect 14642 12724 14648 12776
rect 14700 12764 14706 12776
rect 14737 12767 14795 12773
rect 14737 12764 14749 12767
rect 14700 12736 14749 12764
rect 14700 12724 14706 12736
rect 14737 12733 14749 12736
rect 14783 12733 14795 12767
rect 14737 12727 14795 12733
rect 17129 12767 17187 12773
rect 17129 12733 17141 12767
rect 17175 12733 17187 12767
rect 17129 12727 17187 12733
rect 16114 12696 16120 12708
rect 16172 12705 16178 12708
rect 16084 12668 16120 12696
rect 16114 12656 16120 12668
rect 16172 12659 16184 12705
rect 16172 12656 16178 12659
rect 11885 12631 11943 12637
rect 11885 12628 11897 12631
rect 11848 12600 11897 12628
rect 11848 12588 11854 12600
rect 11885 12597 11897 12600
rect 11931 12597 11943 12631
rect 11885 12591 11943 12597
rect 14553 12631 14611 12637
rect 14553 12597 14565 12631
rect 14599 12628 14611 12631
rect 17144 12628 17172 12727
rect 17586 12724 17592 12776
rect 17644 12764 17650 12776
rect 17957 12767 18015 12773
rect 17957 12764 17969 12767
rect 17644 12736 17969 12764
rect 17644 12724 17650 12736
rect 17957 12733 17969 12736
rect 18003 12733 18015 12767
rect 18966 12764 18972 12776
rect 18927 12736 18972 12764
rect 17957 12727 18015 12733
rect 18966 12724 18972 12736
rect 19024 12724 19030 12776
rect 19061 12699 19119 12705
rect 19061 12696 19073 12699
rect 18340 12668 19073 12696
rect 17310 12628 17316 12640
rect 14599 12600 17172 12628
rect 17271 12600 17316 12628
rect 14599 12597 14611 12600
rect 14553 12591 14611 12597
rect 17310 12588 17316 12600
rect 17368 12588 17374 12640
rect 18340 12637 18368 12668
rect 19061 12665 19073 12668
rect 19107 12665 19119 12699
rect 19061 12659 19119 12665
rect 18325 12631 18383 12637
rect 18325 12597 18337 12631
rect 18371 12597 18383 12631
rect 18325 12591 18383 12597
rect 1104 12538 21896 12560
rect 1104 12486 7912 12538
rect 7964 12486 7976 12538
rect 8028 12486 8040 12538
rect 8092 12486 8104 12538
rect 8156 12486 14843 12538
rect 14895 12486 14907 12538
rect 14959 12486 14971 12538
rect 15023 12486 15035 12538
rect 15087 12486 21896 12538
rect 1104 12464 21896 12486
rect 1762 12424 1768 12436
rect 1723 12396 1768 12424
rect 1762 12384 1768 12396
rect 1820 12384 1826 12436
rect 2406 12424 2412 12436
rect 2367 12396 2412 12424
rect 2406 12384 2412 12396
rect 2464 12384 2470 12436
rect 2682 12424 2688 12436
rect 2643 12396 2688 12424
rect 2682 12384 2688 12396
rect 2740 12384 2746 12436
rect 3329 12427 3387 12433
rect 3329 12393 3341 12427
rect 3375 12424 3387 12427
rect 5445 12427 5503 12433
rect 3375 12396 5396 12424
rect 3375 12393 3387 12396
rect 3329 12387 3387 12393
rect 4706 12356 4712 12368
rect 2884 12328 4712 12356
rect 1949 12291 2007 12297
rect 1949 12257 1961 12291
rect 1995 12288 2007 12291
rect 2038 12288 2044 12300
rect 1995 12260 2044 12288
rect 1995 12257 2007 12260
rect 1949 12251 2007 12257
rect 2038 12248 2044 12260
rect 2096 12248 2102 12300
rect 2225 12291 2283 12297
rect 2225 12257 2237 12291
rect 2271 12288 2283 12291
rect 2498 12288 2504 12300
rect 2271 12260 2504 12288
rect 2271 12257 2283 12260
rect 2225 12251 2283 12257
rect 2498 12248 2504 12260
rect 2556 12248 2562 12300
rect 2884 12297 2912 12328
rect 4706 12316 4712 12328
rect 4764 12316 4770 12368
rect 5368 12356 5396 12396
rect 5445 12393 5457 12427
rect 5491 12424 5503 12427
rect 5718 12424 5724 12436
rect 5491 12396 5724 12424
rect 5491 12393 5503 12396
rect 5445 12387 5503 12393
rect 5718 12384 5724 12396
rect 5776 12384 5782 12436
rect 7558 12424 7564 12436
rect 6748 12396 7236 12424
rect 7519 12396 7564 12424
rect 6748 12356 6776 12396
rect 5368 12328 6776 12356
rect 6822 12316 6828 12368
rect 6880 12316 6886 12368
rect 7006 12316 7012 12368
rect 7064 12365 7070 12368
rect 7064 12356 7076 12365
rect 7208 12356 7236 12396
rect 7558 12384 7564 12396
rect 7616 12384 7622 12436
rect 9214 12424 9220 12436
rect 9175 12396 9220 12424
rect 9214 12384 9220 12396
rect 9272 12384 9278 12436
rect 10505 12427 10563 12433
rect 10505 12393 10517 12427
rect 10551 12424 10563 12427
rect 12618 12424 12624 12436
rect 10551 12396 12434 12424
rect 12579 12396 12624 12424
rect 10551 12393 10563 12396
rect 10505 12387 10563 12393
rect 10045 12359 10103 12365
rect 10045 12356 10057 12359
rect 7064 12328 7109 12356
rect 7208 12328 10057 12356
rect 7064 12319 7076 12328
rect 10045 12325 10057 12328
rect 10091 12325 10103 12359
rect 12406 12356 12434 12396
rect 12618 12384 12624 12396
rect 12676 12384 12682 12436
rect 16209 12427 16267 12433
rect 16209 12393 16221 12427
rect 16255 12424 16267 12427
rect 16482 12424 16488 12436
rect 16255 12396 16488 12424
rect 16255 12393 16267 12396
rect 16209 12387 16267 12393
rect 16482 12384 16488 12396
rect 16540 12384 16546 12436
rect 17954 12384 17960 12436
rect 18012 12424 18018 12436
rect 18969 12427 19027 12433
rect 18969 12424 18981 12427
rect 18012 12396 18981 12424
rect 18012 12384 18018 12396
rect 18969 12393 18981 12396
rect 19015 12393 19027 12427
rect 18969 12387 19027 12393
rect 12989 12359 13047 12365
rect 12989 12356 13001 12359
rect 12406 12328 13001 12356
rect 10045 12319 10103 12325
rect 12989 12325 13001 12328
rect 13035 12325 13047 12359
rect 13998 12356 14004 12368
rect 12989 12319 13047 12325
rect 13188 12328 14004 12356
rect 7064 12316 7070 12319
rect 2869 12291 2927 12297
rect 2869 12257 2881 12291
rect 2915 12257 2927 12291
rect 3142 12288 3148 12300
rect 3103 12260 3148 12288
rect 2869 12251 2927 12257
rect 3142 12248 3148 12260
rect 3200 12248 3206 12300
rect 3878 12288 3884 12300
rect 3791 12260 3884 12288
rect 1489 12223 1547 12229
rect 1489 12189 1501 12223
rect 1535 12220 1547 12223
rect 1535 12192 2774 12220
rect 1535 12189 1547 12192
rect 1489 12183 1547 12189
rect 2746 12152 2774 12192
rect 2958 12180 2964 12232
rect 3016 12220 3022 12232
rect 3804 12220 3832 12260
rect 3878 12248 3884 12260
rect 3936 12288 3942 12300
rect 4321 12291 4379 12297
rect 4321 12288 4333 12291
rect 3936 12260 4333 12288
rect 3936 12248 3942 12260
rect 4321 12257 4333 12260
rect 4367 12257 4379 12291
rect 4321 12251 4379 12257
rect 4798 12248 4804 12300
rect 4856 12288 4862 12300
rect 5994 12288 6000 12300
rect 4856 12260 6000 12288
rect 4856 12248 4862 12260
rect 5994 12248 6000 12260
rect 6052 12248 6058 12300
rect 6840 12288 6868 12316
rect 7285 12291 7343 12297
rect 7285 12288 7297 12291
rect 6840 12260 7297 12288
rect 7285 12257 7297 12260
rect 7331 12257 7343 12291
rect 7285 12251 7343 12257
rect 7929 12291 7987 12297
rect 7929 12257 7941 12291
rect 7975 12288 7987 12291
rect 8662 12288 8668 12300
rect 7975 12260 8668 12288
rect 7975 12257 7987 12260
rect 7929 12251 7987 12257
rect 8662 12248 8668 12260
rect 8720 12248 8726 12300
rect 8754 12248 8760 12300
rect 8812 12288 8818 12300
rect 10137 12291 10195 12297
rect 8812 12260 8857 12288
rect 8812 12248 8818 12260
rect 10137 12257 10149 12291
rect 10183 12288 10195 12291
rect 10781 12291 10839 12297
rect 10781 12288 10793 12291
rect 10183 12260 10793 12288
rect 10183 12257 10195 12260
rect 10137 12251 10195 12257
rect 10781 12257 10793 12260
rect 10827 12257 10839 12291
rect 10781 12251 10839 12257
rect 11333 12291 11391 12297
rect 11333 12257 11345 12291
rect 11379 12288 11391 12291
rect 11885 12291 11943 12297
rect 11885 12288 11897 12291
rect 11379 12260 11897 12288
rect 11379 12257 11391 12260
rect 11333 12251 11391 12257
rect 11885 12257 11897 12260
rect 11931 12257 11943 12291
rect 11885 12251 11943 12257
rect 11977 12291 12035 12297
rect 11977 12257 11989 12291
rect 12023 12288 12035 12291
rect 13188 12288 13216 12328
rect 13998 12316 14004 12328
rect 14056 12316 14062 12368
rect 17580 12359 17638 12365
rect 17580 12325 17592 12359
rect 17626 12356 17638 12359
rect 17770 12356 17776 12368
rect 17626 12328 17776 12356
rect 17626 12325 17638 12328
rect 17580 12319 17638 12325
rect 17770 12316 17776 12328
rect 17828 12316 17834 12368
rect 19242 12316 19248 12368
rect 19300 12356 19306 12368
rect 19300 12328 21404 12356
rect 19300 12316 19306 12328
rect 13814 12288 13820 12300
rect 12023 12260 13216 12288
rect 13775 12260 13820 12288
rect 12023 12257 12035 12260
rect 11977 12251 12035 12257
rect 3016 12192 3832 12220
rect 4065 12223 4123 12229
rect 3016 12180 3022 12192
rect 4065 12189 4077 12223
rect 4111 12189 4123 12223
rect 4065 12183 4123 12189
rect 3326 12152 3332 12164
rect 2746 12124 3332 12152
rect 3326 12112 3332 12124
rect 3384 12112 3390 12164
rect 4080 12084 4108 12183
rect 7558 12180 7564 12232
rect 7616 12220 7622 12232
rect 8021 12223 8079 12229
rect 8021 12220 8033 12223
rect 7616 12192 8033 12220
rect 7616 12180 7622 12192
rect 8021 12189 8033 12192
rect 8067 12189 8079 12223
rect 8202 12220 8208 12232
rect 8163 12192 8208 12220
rect 8021 12183 8079 12189
rect 8202 12180 8208 12192
rect 8260 12180 8266 12232
rect 9950 12220 9956 12232
rect 9863 12192 9956 12220
rect 9950 12180 9956 12192
rect 10008 12220 10014 12232
rect 11790 12220 11796 12232
rect 10008 12192 11796 12220
rect 10008 12180 10014 12192
rect 11790 12180 11796 12192
rect 11848 12180 11854 12232
rect 8478 12152 8484 12164
rect 7300 12124 8484 12152
rect 4246 12084 4252 12096
rect 4080 12056 4252 12084
rect 4246 12044 4252 12056
rect 4304 12084 4310 12096
rect 4798 12084 4804 12096
rect 4304 12056 4804 12084
rect 4304 12044 4310 12056
rect 4798 12044 4804 12056
rect 4856 12044 4862 12096
rect 4982 12044 4988 12096
rect 5040 12084 5046 12096
rect 5902 12084 5908 12096
rect 5040 12056 5908 12084
rect 5040 12044 5046 12056
rect 5902 12044 5908 12056
rect 5960 12044 5966 12096
rect 5994 12044 6000 12096
rect 6052 12084 6058 12096
rect 7300 12084 7328 12124
rect 8478 12112 8484 12124
rect 8536 12112 8542 12164
rect 8570 12084 8576 12096
rect 6052 12056 7328 12084
rect 8531 12056 8576 12084
rect 6052 12044 6058 12056
rect 8570 12044 8576 12056
rect 8628 12044 8634 12096
rect 11900 12084 11928 12251
rect 13814 12248 13820 12260
rect 13872 12248 13878 12300
rect 14820 12291 14878 12297
rect 14820 12257 14832 12291
rect 14866 12288 14878 12291
rect 15286 12288 15292 12300
rect 14866 12260 15292 12288
rect 14866 12257 14878 12260
rect 14820 12251 14878 12257
rect 15286 12248 15292 12260
rect 15344 12248 15350 12300
rect 16298 12248 16304 12300
rect 16356 12288 16362 12300
rect 16577 12291 16635 12297
rect 16577 12288 16589 12291
rect 16356 12260 16589 12288
rect 16356 12248 16362 12260
rect 16577 12257 16589 12260
rect 16623 12257 16635 12291
rect 17310 12288 17316 12300
rect 17223 12260 17316 12288
rect 16577 12251 16635 12257
rect 17310 12248 17316 12260
rect 17368 12288 17374 12300
rect 19260 12288 19288 12316
rect 21082 12288 21088 12300
rect 21140 12297 21146 12300
rect 21376 12297 21404 12328
rect 17368 12260 19288 12288
rect 21052 12260 21088 12288
rect 17368 12248 17374 12260
rect 21082 12248 21088 12260
rect 21140 12251 21152 12297
rect 21361 12291 21419 12297
rect 21361 12257 21373 12291
rect 21407 12257 21419 12291
rect 21361 12251 21419 12257
rect 21140 12248 21146 12251
rect 13081 12223 13139 12229
rect 13081 12220 13093 12223
rect 12360 12192 13093 12220
rect 12360 12161 12388 12192
rect 13081 12189 13093 12192
rect 13127 12189 13139 12223
rect 13081 12183 13139 12189
rect 13173 12223 13231 12229
rect 13173 12189 13185 12223
rect 13219 12189 13231 12223
rect 14553 12223 14611 12229
rect 14553 12220 14565 12223
rect 13173 12183 13231 12189
rect 14016 12192 14565 12220
rect 12345 12155 12403 12161
rect 12345 12121 12357 12155
rect 12391 12121 12403 12155
rect 12345 12115 12403 12121
rect 12710 12112 12716 12164
rect 12768 12152 12774 12164
rect 13188 12152 13216 12183
rect 13906 12152 13912 12164
rect 12768 12124 13216 12152
rect 13280 12124 13912 12152
rect 12768 12112 12774 12124
rect 13280 12084 13308 12124
rect 13906 12112 13912 12124
rect 13964 12112 13970 12164
rect 11900 12056 13308 12084
rect 13354 12044 13360 12096
rect 13412 12084 13418 12096
rect 13630 12084 13636 12096
rect 13412 12056 13636 12084
rect 13412 12044 13418 12056
rect 13630 12044 13636 12056
rect 13688 12084 13694 12096
rect 14016 12084 14044 12192
rect 14553 12189 14565 12192
rect 14599 12189 14611 12223
rect 14553 12183 14611 12189
rect 15838 12180 15844 12232
rect 15896 12220 15902 12232
rect 16669 12223 16727 12229
rect 16669 12220 16681 12223
rect 15896 12192 16681 12220
rect 15896 12180 15902 12192
rect 16669 12189 16681 12192
rect 16715 12189 16727 12223
rect 16669 12183 16727 12189
rect 16761 12223 16819 12229
rect 16761 12189 16773 12223
rect 16807 12189 16819 12223
rect 16761 12183 16819 12189
rect 15933 12155 15991 12161
rect 15933 12121 15945 12155
rect 15979 12152 15991 12155
rect 16114 12152 16120 12164
rect 15979 12124 16120 12152
rect 15979 12121 15991 12124
rect 15933 12115 15991 12121
rect 16114 12112 16120 12124
rect 16172 12152 16178 12164
rect 16776 12152 16804 12183
rect 16172 12124 16804 12152
rect 18693 12155 18751 12161
rect 16172 12112 16178 12124
rect 18693 12121 18705 12155
rect 18739 12152 18751 12155
rect 18782 12152 18788 12164
rect 18739 12124 18788 12152
rect 18739 12121 18751 12124
rect 18693 12115 18751 12121
rect 18782 12112 18788 12124
rect 18840 12152 18846 12164
rect 19150 12152 19156 12164
rect 18840 12124 19156 12152
rect 18840 12112 18846 12124
rect 19150 12112 19156 12124
rect 19208 12112 19214 12164
rect 13688 12056 14044 12084
rect 13688 12044 13694 12056
rect 14366 12044 14372 12096
rect 14424 12084 14430 12096
rect 19981 12087 20039 12093
rect 19981 12084 19993 12087
rect 14424 12056 19993 12084
rect 14424 12044 14430 12056
rect 19981 12053 19993 12056
rect 20027 12053 20039 12087
rect 19981 12047 20039 12053
rect 1104 11994 21896 12016
rect 1104 11942 4447 11994
rect 4499 11942 4511 11994
rect 4563 11942 4575 11994
rect 4627 11942 4639 11994
rect 4691 11942 11378 11994
rect 11430 11942 11442 11994
rect 11494 11942 11506 11994
rect 11558 11942 11570 11994
rect 11622 11942 18308 11994
rect 18360 11942 18372 11994
rect 18424 11942 18436 11994
rect 18488 11942 18500 11994
rect 18552 11942 21896 11994
rect 1104 11920 21896 11942
rect 1670 11840 1676 11892
rect 1728 11880 1734 11892
rect 1765 11883 1823 11889
rect 1765 11880 1777 11883
rect 1728 11852 1777 11880
rect 1728 11840 1734 11852
rect 1765 11849 1777 11852
rect 1811 11849 1823 11883
rect 1765 11843 1823 11849
rect 2038 11840 2044 11892
rect 2096 11880 2102 11892
rect 2225 11883 2283 11889
rect 2225 11880 2237 11883
rect 2096 11852 2237 11880
rect 2096 11840 2102 11852
rect 2225 11849 2237 11852
rect 2271 11849 2283 11883
rect 2225 11843 2283 11849
rect 2498 11840 2504 11892
rect 2556 11880 2562 11892
rect 3329 11883 3387 11889
rect 3329 11880 3341 11883
rect 2556 11852 3341 11880
rect 2556 11840 2562 11852
rect 3329 11849 3341 11852
rect 3375 11849 3387 11883
rect 3329 11843 3387 11849
rect 4062 11840 4068 11892
rect 4120 11880 4126 11892
rect 5353 11883 5411 11889
rect 5353 11880 5365 11883
rect 4120 11852 5365 11880
rect 4120 11840 4126 11852
rect 5353 11849 5365 11852
rect 5399 11849 5411 11883
rect 5353 11843 5411 11849
rect 5905 11883 5963 11889
rect 5905 11849 5917 11883
rect 5951 11880 5963 11883
rect 6086 11880 6092 11892
rect 5951 11852 6092 11880
rect 5951 11849 5963 11852
rect 5905 11843 5963 11849
rect 6086 11840 6092 11852
rect 6144 11840 6150 11892
rect 7190 11840 7196 11892
rect 7248 11880 7254 11892
rect 7929 11883 7987 11889
rect 7929 11880 7941 11883
rect 7248 11852 7941 11880
rect 7248 11840 7254 11852
rect 7929 11849 7941 11852
rect 7975 11849 7987 11883
rect 7929 11843 7987 11849
rect 8294 11840 8300 11892
rect 8352 11880 8358 11892
rect 11054 11880 11060 11892
rect 8352 11852 10640 11880
rect 10967 11852 11060 11880
rect 8352 11840 8358 11852
rect 4157 11815 4215 11821
rect 4157 11781 4169 11815
rect 4203 11812 4215 11815
rect 6641 11815 6699 11821
rect 6641 11812 6653 11815
rect 4203 11784 6653 11812
rect 4203 11781 4215 11784
rect 4157 11775 4215 11781
rect 6641 11781 6653 11784
rect 6687 11781 6699 11815
rect 8570 11812 8576 11824
rect 6641 11775 6699 11781
rect 7033 11784 8576 11812
rect 3878 11744 3884 11756
rect 3839 11716 3884 11744
rect 3878 11704 3884 11716
rect 3936 11704 3942 11756
rect 4890 11744 4896 11756
rect 4851 11716 4896 11744
rect 4890 11704 4896 11716
rect 4948 11704 4954 11756
rect 1854 11636 1860 11688
rect 1912 11676 1918 11688
rect 1949 11679 2007 11685
rect 1949 11676 1961 11679
rect 1912 11648 1961 11676
rect 1912 11636 1918 11648
rect 1949 11645 1961 11648
rect 1995 11645 2007 11679
rect 1949 11639 2007 11645
rect 2409 11679 2467 11685
rect 2409 11645 2421 11679
rect 2455 11676 2467 11679
rect 2498 11676 2504 11688
rect 2455 11648 2504 11676
rect 2455 11645 2467 11648
rect 2409 11639 2467 11645
rect 2498 11636 2504 11648
rect 2556 11636 2562 11688
rect 2685 11679 2743 11685
rect 2685 11645 2697 11679
rect 2731 11676 2743 11679
rect 3418 11676 3424 11688
rect 2731 11648 3424 11676
rect 2731 11645 2743 11648
rect 2685 11639 2743 11645
rect 3418 11636 3424 11648
rect 3476 11636 3482 11688
rect 6089 11679 6147 11685
rect 6089 11645 6101 11679
rect 6135 11676 6147 11679
rect 7033 11676 7061 11784
rect 8570 11772 8576 11784
rect 8628 11772 8634 11824
rect 10612 11812 10640 11852
rect 11054 11840 11060 11852
rect 11112 11880 11118 11892
rect 12710 11880 12716 11892
rect 11112 11852 12716 11880
rect 11112 11840 11118 11852
rect 12710 11840 12716 11852
rect 12768 11840 12774 11892
rect 12805 11883 12863 11889
rect 12805 11849 12817 11883
rect 12851 11880 12863 11883
rect 12986 11880 12992 11892
rect 12851 11852 12992 11880
rect 12851 11849 12863 11852
rect 12805 11843 12863 11849
rect 12986 11840 12992 11852
rect 13044 11840 13050 11892
rect 14182 11840 14188 11892
rect 14240 11880 14246 11892
rect 14829 11883 14887 11889
rect 14829 11880 14841 11883
rect 14240 11852 14841 11880
rect 14240 11840 14246 11852
rect 14829 11849 14841 11852
rect 14875 11849 14887 11883
rect 15838 11880 15844 11892
rect 15799 11852 15844 11880
rect 14829 11843 14887 11849
rect 15838 11840 15844 11852
rect 15896 11840 15902 11892
rect 21082 11840 21088 11892
rect 21140 11880 21146 11892
rect 21177 11883 21235 11889
rect 21177 11880 21189 11883
rect 21140 11852 21189 11880
rect 21140 11840 21146 11852
rect 21177 11849 21189 11852
rect 21223 11849 21235 11883
rect 21177 11843 21235 11849
rect 10612 11784 13952 11812
rect 7098 11704 7104 11756
rect 7156 11744 7162 11756
rect 7285 11747 7343 11753
rect 7156 11716 7201 11744
rect 7156 11704 7162 11716
rect 7285 11713 7297 11747
rect 7331 11744 7343 11747
rect 7466 11744 7472 11756
rect 7331 11716 7472 11744
rect 7331 11713 7343 11716
rect 7285 11707 7343 11713
rect 7466 11704 7472 11716
rect 7524 11704 7530 11756
rect 8202 11704 8208 11756
rect 8260 11744 8266 11756
rect 8481 11747 8539 11753
rect 8481 11744 8493 11747
rect 8260 11716 8493 11744
rect 8260 11704 8266 11716
rect 8481 11713 8493 11716
rect 8527 11713 8539 11747
rect 8481 11707 8539 11713
rect 12066 11704 12072 11756
rect 12124 11744 12130 11756
rect 12161 11747 12219 11753
rect 12161 11744 12173 11747
rect 12124 11716 12173 11744
rect 12124 11704 12130 11716
rect 12161 11713 12173 11716
rect 12207 11713 12219 11747
rect 13265 11747 13323 11753
rect 12161 11707 12219 11713
rect 12268 11716 12756 11744
rect 6135 11648 7061 11676
rect 8389 11679 8447 11685
rect 6135 11645 6147 11648
rect 6089 11639 6147 11645
rect 8389 11645 8401 11679
rect 8435 11676 8447 11679
rect 9674 11676 9680 11688
rect 8435 11648 9076 11676
rect 9635 11648 9680 11676
rect 8435 11645 8447 11648
rect 8389 11639 8447 11645
rect 3697 11611 3755 11617
rect 3697 11577 3709 11611
rect 3743 11608 3755 11611
rect 3743 11580 4384 11608
rect 3743 11577 3755 11580
rect 3697 11571 3755 11577
rect 1394 11540 1400 11552
rect 1355 11512 1400 11540
rect 1394 11500 1400 11512
rect 1452 11500 1458 11552
rect 2866 11540 2872 11552
rect 2827 11512 2872 11540
rect 2866 11500 2872 11512
rect 2924 11500 2930 11552
rect 4356 11549 4384 11580
rect 4430 11568 4436 11620
rect 4488 11608 4494 11620
rect 7009 11611 7067 11617
rect 7009 11608 7021 11611
rect 4488 11580 7021 11608
rect 4488 11568 4494 11580
rect 7009 11577 7021 11580
rect 7055 11608 7067 11611
rect 7742 11608 7748 11620
rect 7055 11580 7748 11608
rect 7055 11577 7067 11580
rect 7009 11571 7067 11577
rect 7742 11568 7748 11580
rect 7800 11608 7806 11620
rect 8297 11611 8355 11617
rect 8297 11608 8309 11611
rect 7800 11580 8309 11608
rect 7800 11568 7806 11580
rect 8297 11577 8309 11580
rect 8343 11577 8355 11611
rect 9048 11608 9076 11648
rect 9674 11636 9680 11648
rect 9732 11636 9738 11688
rect 9950 11685 9956 11688
rect 9944 11676 9956 11685
rect 9911 11648 9956 11676
rect 9944 11639 9956 11648
rect 9950 11636 9956 11639
rect 10008 11636 10014 11688
rect 12268 11676 12296 11716
rect 11532 11648 12296 11676
rect 12728 11676 12756 11716
rect 13265 11713 13277 11747
rect 13311 11744 13323 11747
rect 13814 11744 13820 11756
rect 13311 11716 13820 11744
rect 13311 11713 13323 11716
rect 13265 11707 13323 11713
rect 13814 11704 13820 11716
rect 13872 11704 13878 11756
rect 13449 11679 13507 11685
rect 13449 11676 13461 11679
rect 12728 11648 13461 11676
rect 10502 11608 10508 11620
rect 9048 11580 10508 11608
rect 8297 11571 8355 11577
rect 10502 11568 10508 11580
rect 10560 11568 10566 11620
rect 3789 11543 3847 11549
rect 3789 11509 3801 11543
rect 3835 11540 3847 11543
rect 4157 11543 4215 11549
rect 4157 11540 4169 11543
rect 3835 11512 4169 11540
rect 3835 11509 3847 11512
rect 3789 11503 3847 11509
rect 4157 11509 4169 11512
rect 4203 11509 4215 11543
rect 4157 11503 4215 11509
rect 4341 11543 4399 11549
rect 4341 11509 4353 11543
rect 4387 11509 4399 11543
rect 4706 11540 4712 11552
rect 4667 11512 4712 11540
rect 4341 11503 4399 11509
rect 4706 11500 4712 11512
rect 4764 11500 4770 11552
rect 4801 11543 4859 11549
rect 4801 11509 4813 11543
rect 4847 11540 4859 11543
rect 4982 11540 4988 11552
rect 4847 11512 4988 11540
rect 4847 11509 4859 11512
rect 4801 11503 4859 11509
rect 4982 11500 4988 11512
rect 5040 11500 5046 11552
rect 9122 11500 9128 11552
rect 9180 11540 9186 11552
rect 11532 11540 11560 11648
rect 13449 11645 13461 11648
rect 13495 11645 13507 11679
rect 13449 11639 13507 11645
rect 12342 11608 12348 11620
rect 12303 11580 12348 11608
rect 12342 11568 12348 11580
rect 12400 11568 12406 11620
rect 12437 11611 12495 11617
rect 12437 11577 12449 11611
rect 12483 11608 12495 11611
rect 12894 11608 12900 11620
rect 12483 11580 12900 11608
rect 12483 11577 12495 11580
rect 12437 11571 12495 11577
rect 12894 11568 12900 11580
rect 12952 11568 12958 11620
rect 13924 11608 13952 11784
rect 16482 11772 16488 11824
rect 16540 11812 16546 11824
rect 17681 11815 17739 11821
rect 17681 11812 17693 11815
rect 16540 11784 17693 11812
rect 16540 11772 16546 11784
rect 17681 11781 17693 11784
rect 17727 11781 17739 11815
rect 17681 11775 17739 11781
rect 14274 11744 14280 11756
rect 14235 11716 14280 11744
rect 14274 11704 14280 11716
rect 14332 11704 14338 11756
rect 15286 11744 15292 11756
rect 15247 11716 15292 11744
rect 15286 11704 15292 11716
rect 15344 11704 15350 11756
rect 16298 11744 16304 11756
rect 16259 11716 16304 11744
rect 16298 11704 16304 11716
rect 16356 11704 16362 11756
rect 19061 11747 19119 11753
rect 19061 11713 19073 11747
rect 19107 11744 19119 11747
rect 19242 11744 19248 11756
rect 19107 11716 19248 11744
rect 19107 11713 19119 11716
rect 19061 11707 19119 11713
rect 19242 11704 19248 11716
rect 19300 11704 19306 11756
rect 15194 11636 15200 11688
rect 15252 11676 15258 11688
rect 15381 11679 15439 11685
rect 15381 11676 15393 11679
rect 15252 11648 15393 11676
rect 15252 11636 15258 11648
rect 15381 11645 15393 11648
rect 15427 11676 15439 11679
rect 16945 11679 17003 11685
rect 16945 11676 16957 11679
rect 15427 11648 16957 11676
rect 15427 11645 15439 11648
rect 15381 11639 15439 11645
rect 16945 11645 16957 11648
rect 16991 11645 17003 11679
rect 16945 11639 17003 11645
rect 18782 11636 18788 11688
rect 18840 11685 18846 11688
rect 18840 11676 18852 11685
rect 20901 11679 20959 11685
rect 18840 11648 18885 11676
rect 18840 11639 18852 11648
rect 20901 11645 20913 11679
rect 20947 11676 20959 11679
rect 21358 11676 21364 11688
rect 20947 11648 21364 11676
rect 20947 11645 20959 11648
rect 20901 11639 20959 11645
rect 18840 11636 18846 11639
rect 21358 11636 21364 11648
rect 21416 11636 21422 11688
rect 15473 11611 15531 11617
rect 15473 11608 15485 11611
rect 13924 11580 15485 11608
rect 15473 11577 15485 11580
rect 15519 11577 15531 11611
rect 15473 11571 15531 11577
rect 9180 11512 11560 11540
rect 11793 11543 11851 11549
rect 9180 11500 9186 11512
rect 11793 11509 11805 11543
rect 11839 11540 11851 11543
rect 13357 11543 13415 11549
rect 13357 11540 13369 11543
rect 11839 11512 13369 11540
rect 11839 11509 11851 11512
rect 11793 11503 11851 11509
rect 13357 11509 13369 11512
rect 13403 11540 13415 11543
rect 13446 11540 13452 11552
rect 13403 11512 13452 11540
rect 13403 11509 13415 11512
rect 13357 11503 13415 11509
rect 13446 11500 13452 11512
rect 13504 11500 13510 11552
rect 13817 11543 13875 11549
rect 13817 11509 13829 11543
rect 13863 11540 13875 11543
rect 14369 11543 14427 11549
rect 14369 11540 14381 11543
rect 13863 11512 14381 11540
rect 13863 11509 13875 11512
rect 13817 11503 13875 11509
rect 14369 11509 14381 11512
rect 14415 11509 14427 11543
rect 14369 11503 14427 11509
rect 14458 11500 14464 11552
rect 14516 11540 14522 11552
rect 14516 11512 14561 11540
rect 14516 11500 14522 11512
rect 1104 11450 21896 11472
rect 1104 11398 7912 11450
rect 7964 11398 7976 11450
rect 8028 11398 8040 11450
rect 8092 11398 8104 11450
rect 8156 11398 14843 11450
rect 14895 11398 14907 11450
rect 14959 11398 14971 11450
rect 15023 11398 15035 11450
rect 15087 11398 21896 11450
rect 1104 11376 21896 11398
rect 1581 11339 1639 11345
rect 1581 11305 1593 11339
rect 1627 11305 1639 11339
rect 1854 11336 1860 11348
rect 1815 11308 1860 11336
rect 1581 11299 1639 11305
rect 1596 11268 1624 11299
rect 1854 11296 1860 11308
rect 1912 11296 1918 11348
rect 3418 11336 3424 11348
rect 3379 11308 3424 11336
rect 3418 11296 3424 11308
rect 3476 11296 3482 11348
rect 4154 11296 4160 11348
rect 4212 11336 4218 11348
rect 4430 11336 4436 11348
rect 4212 11308 4436 11336
rect 4212 11296 4218 11308
rect 4430 11296 4436 11308
rect 4488 11296 4494 11348
rect 4706 11296 4712 11348
rect 4764 11336 4770 11348
rect 5077 11339 5135 11345
rect 5077 11336 5089 11339
rect 4764 11308 5089 11336
rect 4764 11296 4770 11308
rect 5077 11305 5089 11308
rect 5123 11305 5135 11339
rect 5077 11299 5135 11305
rect 5166 11296 5172 11348
rect 5224 11336 5230 11348
rect 7101 11339 7159 11345
rect 7101 11336 7113 11339
rect 5224 11308 7113 11336
rect 5224 11296 5230 11308
rect 7101 11305 7113 11308
rect 7147 11305 7159 11339
rect 7101 11299 7159 11305
rect 7193 11339 7251 11345
rect 7193 11305 7205 11339
rect 7239 11336 7251 11339
rect 7282 11336 7288 11348
rect 7239 11308 7288 11336
rect 7239 11305 7251 11308
rect 7193 11299 7251 11305
rect 7282 11296 7288 11308
rect 7340 11296 7346 11348
rect 8294 11336 8300 11348
rect 7392 11308 8300 11336
rect 6273 11271 6331 11277
rect 1596 11240 6132 11268
rect 1394 11200 1400 11212
rect 1355 11172 1400 11200
rect 1394 11160 1400 11172
rect 1452 11160 1458 11212
rect 2041 11203 2099 11209
rect 2041 11169 2053 11203
rect 2087 11169 2099 11203
rect 2041 11163 2099 11169
rect 2056 11064 2084 11163
rect 2774 11160 2780 11212
rect 2832 11200 2838 11212
rect 2832 11172 2877 11200
rect 2832 11160 2838 11172
rect 2866 11132 2872 11144
rect 2827 11104 2872 11132
rect 2866 11092 2872 11104
rect 2924 11092 2930 11144
rect 3050 11132 3056 11144
rect 3011 11104 3056 11132
rect 3050 11092 3056 11104
rect 3108 11092 3114 11144
rect 4062 11092 4068 11144
rect 4120 11132 4126 11144
rect 4157 11135 4215 11141
rect 4157 11132 4169 11135
rect 4120 11104 4169 11132
rect 4120 11092 4126 11104
rect 4157 11101 4169 11104
rect 4203 11101 4215 11135
rect 4157 11095 4215 11101
rect 4341 11135 4399 11141
rect 4341 11101 4353 11135
rect 4387 11132 4399 11135
rect 5994 11132 6000 11144
rect 4387 11104 6000 11132
rect 4387 11101 4399 11104
rect 4341 11095 4399 11101
rect 5994 11092 6000 11104
rect 6052 11092 6058 11144
rect 5813 11067 5871 11073
rect 5813 11064 5825 11067
rect 2056 11036 5825 11064
rect 5813 11033 5825 11036
rect 5859 11033 5871 11067
rect 6104 11064 6132 11240
rect 6273 11237 6285 11271
rect 6319 11268 6331 11271
rect 7006 11268 7012 11280
rect 6319 11240 7012 11268
rect 6319 11237 6331 11240
rect 6273 11231 6331 11237
rect 7006 11228 7012 11240
rect 7064 11228 7070 11280
rect 6181 11203 6239 11209
rect 6181 11169 6193 11203
rect 6227 11200 6239 11203
rect 6638 11200 6644 11212
rect 6227 11172 6644 11200
rect 6227 11169 6239 11172
rect 6181 11163 6239 11169
rect 6638 11160 6644 11172
rect 6696 11160 6702 11212
rect 7392 11200 7420 11308
rect 8294 11296 8300 11308
rect 8352 11296 8358 11348
rect 8662 11296 8668 11348
rect 8720 11336 8726 11348
rect 9309 11339 9367 11345
rect 9309 11336 9321 11339
rect 8720 11308 9321 11336
rect 8720 11296 8726 11308
rect 9309 11305 9321 11308
rect 9355 11305 9367 11339
rect 12250 11336 12256 11348
rect 9309 11299 9367 11305
rect 9416 11308 12256 11336
rect 9416 11268 9444 11308
rect 12250 11296 12256 11308
rect 12308 11296 12314 11348
rect 13541 11339 13599 11345
rect 13541 11305 13553 11339
rect 13587 11336 13599 11339
rect 13814 11336 13820 11348
rect 13587 11308 13820 11336
rect 13587 11305 13599 11308
rect 13541 11299 13599 11305
rect 13814 11296 13820 11308
rect 13872 11296 13878 11348
rect 14001 11339 14059 11345
rect 14001 11305 14013 11339
rect 14047 11336 14059 11339
rect 14458 11336 14464 11348
rect 14047 11308 14464 11336
rect 14047 11305 14059 11308
rect 14001 11299 14059 11305
rect 14458 11296 14464 11308
rect 14516 11296 14522 11348
rect 15286 11296 15292 11348
rect 15344 11336 15350 11348
rect 15933 11339 15991 11345
rect 15933 11336 15945 11339
rect 15344 11308 15945 11336
rect 15344 11296 15350 11308
rect 15933 11305 15945 11308
rect 15979 11305 15991 11339
rect 15933 11299 15991 11305
rect 7944 11240 9444 11268
rect 10496 11271 10554 11277
rect 7944 11200 7972 11240
rect 10496 11237 10508 11271
rect 10542 11268 10554 11271
rect 11054 11268 11060 11280
rect 10542 11240 11060 11268
rect 10542 11237 10554 11240
rect 10496 11231 10554 11237
rect 11054 11228 11060 11240
rect 11112 11228 11118 11280
rect 12710 11268 12716 11280
rect 12176 11240 12716 11268
rect 6840 11172 7420 11200
rect 7576 11172 7972 11200
rect 6457 11135 6515 11141
rect 6457 11101 6469 11135
rect 6503 11132 6515 11135
rect 6730 11132 6736 11144
rect 6503 11104 6736 11132
rect 6503 11101 6515 11104
rect 6457 11095 6515 11101
rect 6730 11092 6736 11104
rect 6788 11092 6794 11144
rect 6840 11064 6868 11172
rect 6917 11135 6975 11141
rect 6917 11101 6929 11135
rect 6963 11132 6975 11135
rect 7374 11132 7380 11144
rect 6963 11104 7380 11132
rect 6963 11101 6975 11104
rect 6917 11095 6975 11101
rect 7374 11092 7380 11104
rect 7432 11132 7438 11144
rect 7576 11132 7604 11172
rect 8018 11160 8024 11212
rect 8076 11200 8082 11212
rect 12176 11209 12204 11240
rect 12710 11228 12716 11240
rect 12768 11228 12774 11280
rect 14274 11228 14280 11280
rect 14332 11268 14338 11280
rect 14798 11271 14856 11277
rect 14798 11268 14810 11271
rect 14332 11240 14810 11268
rect 14332 11228 14338 11240
rect 14798 11237 14810 11240
rect 14844 11268 14856 11271
rect 14918 11268 14924 11280
rect 14844 11240 14924 11268
rect 14844 11237 14856 11240
rect 14798 11231 14856 11237
rect 14918 11228 14924 11240
rect 14976 11228 14982 11280
rect 16482 11277 16488 11280
rect 16476 11268 16488 11277
rect 16443 11240 16488 11268
rect 16476 11231 16488 11240
rect 16482 11228 16488 11231
rect 16540 11228 16546 11280
rect 8306 11203 8364 11209
rect 8306 11200 8318 11203
rect 8076 11172 8318 11200
rect 8076 11160 8082 11172
rect 8306 11169 8318 11172
rect 8352 11169 8364 11203
rect 8306 11163 8364 11169
rect 12161 11203 12219 11209
rect 12161 11169 12173 11203
rect 12207 11169 12219 11203
rect 12428 11203 12486 11209
rect 12428 11200 12440 11203
rect 12161 11163 12219 11169
rect 12268 11172 12440 11200
rect 7432 11104 7604 11132
rect 8573 11135 8631 11141
rect 7432 11092 7438 11104
rect 8573 11101 8585 11135
rect 8619 11132 8631 11135
rect 9674 11132 9680 11144
rect 8619 11104 9680 11132
rect 8619 11101 8631 11104
rect 8573 11095 8631 11101
rect 6104 11036 6868 11064
rect 7101 11067 7159 11073
rect 5813 11027 5871 11033
rect 7101 11033 7113 11067
rect 7147 11064 7159 11067
rect 7558 11064 7564 11076
rect 7147 11036 7564 11064
rect 7147 11033 7159 11036
rect 7101 11027 7159 11033
rect 7558 11024 7564 11036
rect 7616 11024 7622 11076
rect 2406 10996 2412 11008
rect 2367 10968 2412 10996
rect 2406 10956 2412 10968
rect 2464 10956 2470 11008
rect 4798 10996 4804 11008
rect 4759 10968 4804 10996
rect 4798 10956 4804 10968
rect 4856 10956 4862 11008
rect 7650 10956 7656 11008
rect 7708 10996 7714 11008
rect 8588 10996 8616 11095
rect 9674 11092 9680 11104
rect 9732 11132 9738 11144
rect 10229 11135 10287 11141
rect 10229 11132 10241 11135
rect 9732 11104 10241 11132
rect 9732 11092 9738 11104
rect 10229 11101 10241 11104
rect 10275 11101 10287 11135
rect 10229 11095 10287 11101
rect 12066 11092 12072 11144
rect 12124 11132 12130 11144
rect 12268 11132 12296 11172
rect 12428 11169 12440 11172
rect 12474 11200 12486 11203
rect 13262 11200 13268 11212
rect 12474 11172 13268 11200
rect 12474 11169 12486 11172
rect 12428 11163 12486 11169
rect 13262 11160 13268 11172
rect 13320 11160 13326 11212
rect 13630 11160 13636 11212
rect 13688 11200 13694 11212
rect 14553 11203 14611 11209
rect 14553 11200 14565 11203
rect 13688 11172 14565 11200
rect 13688 11160 13694 11172
rect 14553 11169 14565 11172
rect 14599 11169 14611 11203
rect 14553 11163 14611 11169
rect 16209 11203 16267 11209
rect 16209 11169 16221 11203
rect 16255 11200 16267 11203
rect 17310 11200 17316 11212
rect 16255 11172 17316 11200
rect 16255 11169 16267 11172
rect 16209 11163 16267 11169
rect 17310 11160 17316 11172
rect 17368 11160 17374 11212
rect 12124 11104 12296 11132
rect 12124 11092 12130 11104
rect 7708 10968 8616 10996
rect 7708 10956 7714 10968
rect 11238 10956 11244 11008
rect 11296 10996 11302 11008
rect 11609 10999 11667 11005
rect 11609 10996 11621 10999
rect 11296 10968 11621 10996
rect 11296 10956 11302 10968
rect 11609 10965 11621 10968
rect 11655 10965 11667 10999
rect 17586 10996 17592 11008
rect 17547 10968 17592 10996
rect 11609 10959 11667 10965
rect 17586 10956 17592 10968
rect 17644 10956 17650 11008
rect 1104 10906 21896 10928
rect 1104 10854 4447 10906
rect 4499 10854 4511 10906
rect 4563 10854 4575 10906
rect 4627 10854 4639 10906
rect 4691 10854 11378 10906
rect 11430 10854 11442 10906
rect 11494 10854 11506 10906
rect 11558 10854 11570 10906
rect 11622 10854 18308 10906
rect 18360 10854 18372 10906
rect 18424 10854 18436 10906
rect 18488 10854 18500 10906
rect 18552 10854 21896 10906
rect 1104 10832 21896 10854
rect 2498 10792 2504 10804
rect 2459 10764 2504 10792
rect 2498 10752 2504 10764
rect 2556 10752 2562 10804
rect 2777 10795 2835 10801
rect 2777 10761 2789 10795
rect 2823 10792 2835 10795
rect 3050 10792 3056 10804
rect 2823 10764 3056 10792
rect 2823 10761 2835 10764
rect 2777 10755 2835 10761
rect 3050 10752 3056 10764
rect 3108 10792 3114 10804
rect 7650 10792 7656 10804
rect 3108 10764 5028 10792
rect 3108 10752 3114 10764
rect 1949 10659 2007 10665
rect 1949 10625 1961 10659
rect 1995 10656 2007 10659
rect 2038 10656 2044 10668
rect 1995 10628 2044 10656
rect 1995 10625 2007 10628
rect 1949 10619 2007 10625
rect 2038 10616 2044 10628
rect 2096 10616 2102 10668
rect 4157 10659 4215 10665
rect 4157 10625 4169 10659
rect 4203 10656 4215 10659
rect 4246 10656 4252 10668
rect 4203 10628 4252 10656
rect 4203 10625 4215 10628
rect 4157 10619 4215 10625
rect 4246 10616 4252 10628
rect 4304 10616 4310 10668
rect 4798 10616 4804 10668
rect 4856 10656 4862 10668
rect 5000 10665 5028 10764
rect 6656 10764 7656 10792
rect 6656 10665 6684 10764
rect 7650 10752 7656 10764
rect 7708 10752 7714 10804
rect 8018 10792 8024 10804
rect 7979 10764 8024 10792
rect 8018 10752 8024 10764
rect 8076 10752 8082 10804
rect 9674 10752 9680 10804
rect 9732 10792 9738 10804
rect 9769 10795 9827 10801
rect 9769 10792 9781 10795
rect 9732 10764 9781 10792
rect 9732 10752 9738 10764
rect 9769 10761 9781 10764
rect 9815 10792 9827 10795
rect 10686 10792 10692 10804
rect 9815 10764 10692 10792
rect 9815 10761 9827 10764
rect 9769 10755 9827 10761
rect 10686 10752 10692 10764
rect 10744 10752 10750 10804
rect 11333 10795 11391 10801
rect 11333 10761 11345 10795
rect 11379 10792 11391 10795
rect 11790 10792 11796 10804
rect 11379 10764 11796 10792
rect 11379 10761 11391 10764
rect 11333 10755 11391 10761
rect 11790 10752 11796 10764
rect 11848 10752 11854 10804
rect 13262 10792 13268 10804
rect 11900 10764 13124 10792
rect 13223 10764 13268 10792
rect 11900 10724 11928 10764
rect 7668 10696 11928 10724
rect 13096 10724 13124 10764
rect 13262 10752 13268 10764
rect 13320 10752 13326 10804
rect 14918 10792 14924 10804
rect 13556 10764 14780 10792
rect 14879 10764 14924 10792
rect 13556 10724 13584 10764
rect 13096 10696 13584 10724
rect 14752 10724 14780 10764
rect 14918 10752 14924 10764
rect 14976 10752 14982 10804
rect 17129 10727 17187 10733
rect 17129 10724 17141 10727
rect 14752 10696 17141 10724
rect 4893 10659 4951 10665
rect 4893 10656 4905 10659
rect 4856 10628 4905 10656
rect 4856 10616 4862 10628
rect 4893 10625 4905 10628
rect 4939 10625 4951 10659
rect 4893 10619 4951 10625
rect 4985 10659 5043 10665
rect 4985 10625 4997 10659
rect 5031 10625 5043 10659
rect 4985 10619 5043 10625
rect 6641 10659 6699 10665
rect 6641 10625 6653 10659
rect 6687 10625 6699 10659
rect 6641 10619 6699 10625
rect 2133 10591 2191 10597
rect 2133 10557 2145 10591
rect 2179 10588 2191 10591
rect 2406 10588 2412 10600
rect 2179 10560 2412 10588
rect 2179 10557 2191 10560
rect 2133 10551 2191 10557
rect 2406 10548 2412 10560
rect 2464 10548 2470 10600
rect 6730 10548 6736 10600
rect 6788 10588 6794 10600
rect 6897 10591 6955 10597
rect 6897 10588 6909 10591
rect 6788 10560 6909 10588
rect 6788 10548 6794 10560
rect 6897 10557 6909 10560
rect 6943 10557 6955 10591
rect 6897 10551 6955 10557
rect 2041 10523 2099 10529
rect 2041 10489 2053 10523
rect 2087 10520 2099 10523
rect 3912 10523 3970 10529
rect 2087 10492 3648 10520
rect 2087 10489 2099 10492
rect 2041 10483 2099 10489
rect 1394 10452 1400 10464
rect 1355 10424 1400 10452
rect 1394 10412 1400 10424
rect 1452 10412 1458 10464
rect 3620 10452 3648 10492
rect 3912 10489 3924 10523
rect 3958 10520 3970 10523
rect 4062 10520 4068 10532
rect 3958 10492 4068 10520
rect 3958 10489 3970 10492
rect 3912 10483 3970 10489
rect 4062 10480 4068 10492
rect 4120 10520 4126 10532
rect 7668 10520 7696 10696
rect 17129 10693 17141 10696
rect 17175 10693 17187 10727
rect 17129 10687 17187 10693
rect 7742 10616 7748 10668
rect 7800 10656 7806 10668
rect 8294 10656 8300 10668
rect 7800 10628 8300 10656
rect 7800 10616 7806 10628
rect 8294 10616 8300 10628
rect 8352 10616 8358 10668
rect 9030 10656 9036 10668
rect 8991 10628 9036 10656
rect 9030 10616 9036 10628
rect 9088 10616 9094 10668
rect 9217 10659 9275 10665
rect 9217 10625 9229 10659
rect 9263 10656 9275 10659
rect 9674 10656 9680 10668
rect 9263 10628 9680 10656
rect 9263 10625 9275 10628
rect 9217 10619 9275 10625
rect 9674 10616 9680 10628
rect 9732 10616 9738 10668
rect 15565 10659 15623 10665
rect 15565 10625 15577 10659
rect 15611 10656 15623 10659
rect 16482 10656 16488 10668
rect 15611 10628 16488 10656
rect 15611 10625 15623 10628
rect 15565 10619 15623 10625
rect 16482 10616 16488 10628
rect 16540 10616 16546 10668
rect 18509 10659 18567 10665
rect 18509 10625 18521 10659
rect 18555 10656 18567 10659
rect 19242 10656 19248 10668
rect 18555 10628 19248 10656
rect 18555 10625 18567 10628
rect 18509 10619 18567 10625
rect 19242 10616 19248 10628
rect 19300 10616 19306 10668
rect 8570 10548 8576 10600
rect 8628 10588 8634 10600
rect 9585 10591 9643 10597
rect 9585 10588 9597 10591
rect 8628 10560 9597 10588
rect 8628 10548 8634 10560
rect 9585 10557 9597 10560
rect 9631 10557 9643 10591
rect 9585 10551 9643 10557
rect 11238 10548 11244 10600
rect 11296 10548 11302 10600
rect 11885 10591 11943 10597
rect 11885 10557 11897 10591
rect 11931 10588 11943 10591
rect 12710 10588 12716 10600
rect 11931 10560 12716 10588
rect 11931 10557 11943 10560
rect 11885 10551 11943 10557
rect 12710 10548 12716 10560
rect 12768 10588 12774 10600
rect 13541 10591 13599 10597
rect 13541 10588 13553 10591
rect 12768 10560 13553 10588
rect 12768 10548 12774 10560
rect 13541 10557 13553 10560
rect 13587 10588 13599 10591
rect 13630 10588 13636 10600
rect 13587 10560 13636 10588
rect 13587 10557 13599 10560
rect 13541 10551 13599 10557
rect 13630 10548 13636 10560
rect 13688 10548 13694 10600
rect 13814 10597 13820 10600
rect 13808 10588 13820 10597
rect 13775 10560 13820 10588
rect 13808 10551 13820 10560
rect 13814 10548 13820 10551
rect 13872 10548 13878 10600
rect 9766 10520 9772 10532
rect 4120 10492 7696 10520
rect 8128 10492 9772 10520
rect 4120 10480 4126 10492
rect 4433 10455 4491 10461
rect 4433 10452 4445 10455
rect 3620 10424 4445 10452
rect 4433 10421 4445 10424
rect 4479 10421 4491 10455
rect 4798 10452 4804 10464
rect 4759 10424 4804 10452
rect 4433 10415 4491 10421
rect 4798 10412 4804 10424
rect 4856 10412 4862 10464
rect 5350 10412 5356 10464
rect 5408 10452 5414 10464
rect 5445 10455 5503 10461
rect 5445 10452 5457 10455
rect 5408 10424 5457 10452
rect 5408 10412 5414 10424
rect 5445 10421 5457 10424
rect 5491 10421 5503 10455
rect 5445 10415 5503 10421
rect 5718 10412 5724 10464
rect 5776 10452 5782 10464
rect 5813 10455 5871 10461
rect 5813 10452 5825 10455
rect 5776 10424 5825 10452
rect 5776 10412 5782 10424
rect 5813 10421 5825 10424
rect 5859 10452 5871 10455
rect 6362 10452 6368 10464
rect 5859 10424 6368 10452
rect 5859 10421 5871 10424
rect 5813 10415 5871 10421
rect 6362 10412 6368 10424
rect 6420 10452 6426 10464
rect 8128 10452 8156 10492
rect 9766 10480 9772 10492
rect 9824 10520 9830 10532
rect 10042 10520 10048 10532
rect 9824 10492 10048 10520
rect 9824 10480 9830 10492
rect 10042 10480 10048 10492
rect 10100 10480 10106 10532
rect 11256 10520 11284 10548
rect 12130 10523 12188 10529
rect 12130 10520 12142 10523
rect 11256 10492 12142 10520
rect 12130 10489 12142 10492
rect 12176 10489 12188 10523
rect 12130 10483 12188 10489
rect 12526 10480 12532 10532
rect 12584 10520 12590 10532
rect 15194 10520 15200 10532
rect 12584 10492 15200 10520
rect 12584 10480 12590 10492
rect 15194 10480 15200 10492
rect 15252 10520 15258 10532
rect 15657 10523 15715 10529
rect 15657 10520 15669 10523
rect 15252 10492 15669 10520
rect 15252 10480 15258 10492
rect 15657 10489 15669 10492
rect 15703 10489 15715 10523
rect 15657 10483 15715 10489
rect 17586 10480 17592 10532
rect 17644 10520 17650 10532
rect 18242 10523 18300 10529
rect 18242 10520 18254 10523
rect 17644 10492 18254 10520
rect 17644 10480 17650 10492
rect 18242 10489 18254 10492
rect 18288 10489 18300 10523
rect 18242 10483 18300 10489
rect 6420 10424 8156 10452
rect 6420 10412 6426 10424
rect 8202 10412 8208 10464
rect 8260 10452 8266 10464
rect 8573 10455 8631 10461
rect 8573 10452 8585 10455
rect 8260 10424 8585 10452
rect 8260 10412 8266 10424
rect 8573 10421 8585 10424
rect 8619 10421 8631 10455
rect 8938 10452 8944 10464
rect 8899 10424 8944 10452
rect 8573 10415 8631 10421
rect 8938 10412 8944 10424
rect 8996 10412 9002 10464
rect 15746 10412 15752 10464
rect 15804 10452 15810 10464
rect 16114 10452 16120 10464
rect 15804 10424 15849 10452
rect 16075 10424 16120 10452
rect 15804 10412 15810 10424
rect 16114 10412 16120 10424
rect 16172 10412 16178 10464
rect 16577 10455 16635 10461
rect 16577 10421 16589 10455
rect 16623 10452 16635 10455
rect 16942 10452 16948 10464
rect 16623 10424 16948 10452
rect 16623 10421 16635 10424
rect 16577 10415 16635 10421
rect 16942 10412 16948 10424
rect 17000 10412 17006 10464
rect 1104 10362 21896 10384
rect 1104 10310 7912 10362
rect 7964 10310 7976 10362
rect 8028 10310 8040 10362
rect 8092 10310 8104 10362
rect 8156 10310 14843 10362
rect 14895 10310 14907 10362
rect 14959 10310 14971 10362
rect 15023 10310 15035 10362
rect 15087 10310 21896 10362
rect 1104 10288 21896 10310
rect 1581 10251 1639 10257
rect 1581 10217 1593 10251
rect 1627 10248 1639 10251
rect 2590 10248 2596 10260
rect 1627 10220 2596 10248
rect 1627 10217 1639 10220
rect 1581 10211 1639 10217
rect 2590 10208 2596 10220
rect 2648 10208 2654 10260
rect 4798 10248 4804 10260
rect 4759 10220 4804 10248
rect 4798 10208 4804 10220
rect 4856 10208 4862 10260
rect 5074 10208 5080 10260
rect 5132 10248 5138 10260
rect 5810 10248 5816 10260
rect 5132 10220 5816 10248
rect 5132 10208 5138 10220
rect 5810 10208 5816 10220
rect 5868 10208 5874 10260
rect 6641 10251 6699 10257
rect 6641 10217 6653 10251
rect 6687 10248 6699 10251
rect 6730 10248 6736 10260
rect 6687 10220 6736 10248
rect 6687 10217 6699 10220
rect 6641 10211 6699 10217
rect 6730 10208 6736 10220
rect 6788 10208 6794 10260
rect 7006 10208 7012 10260
rect 7064 10248 7070 10260
rect 7745 10251 7803 10257
rect 7745 10248 7757 10251
rect 7064 10220 7757 10248
rect 7064 10208 7070 10220
rect 7745 10217 7757 10220
rect 7791 10217 7803 10251
rect 8202 10248 8208 10260
rect 8163 10220 8208 10248
rect 7745 10211 7803 10217
rect 8202 10208 8208 10220
rect 8260 10208 8266 10260
rect 11517 10251 11575 10257
rect 11517 10217 11529 10251
rect 11563 10248 11575 10251
rect 11698 10248 11704 10260
rect 11563 10220 11704 10248
rect 11563 10217 11575 10220
rect 11517 10211 11575 10217
rect 11698 10208 11704 10220
rect 11756 10208 11762 10260
rect 11885 10251 11943 10257
rect 11885 10217 11897 10251
rect 11931 10248 11943 10251
rect 12342 10248 12348 10260
rect 11931 10220 12348 10248
rect 11931 10217 11943 10220
rect 11885 10211 11943 10217
rect 12342 10208 12348 10220
rect 12400 10208 12406 10260
rect 12437 10251 12495 10257
rect 12437 10217 12449 10251
rect 12483 10248 12495 10251
rect 12894 10248 12900 10260
rect 12483 10220 12900 10248
rect 12483 10217 12495 10220
rect 12437 10211 12495 10217
rect 12894 10208 12900 10220
rect 12952 10208 12958 10260
rect 15194 10248 15200 10260
rect 15155 10220 15200 10248
rect 15194 10208 15200 10220
rect 15252 10208 15258 10260
rect 16942 10248 16948 10260
rect 16903 10220 16948 10248
rect 16942 10208 16948 10220
rect 17000 10208 17006 10260
rect 17313 10251 17371 10257
rect 17313 10217 17325 10251
rect 17359 10248 17371 10251
rect 18690 10248 18696 10260
rect 17359 10220 18696 10248
rect 17359 10217 17371 10220
rect 17313 10211 17371 10217
rect 18690 10208 18696 10220
rect 18748 10208 18754 10260
rect 15746 10180 15752 10192
rect 2746 10152 15752 10180
rect 1394 10112 1400 10124
rect 1355 10084 1400 10112
rect 1394 10072 1400 10084
rect 1452 10072 1458 10124
rect 1578 10072 1584 10124
rect 1636 10112 1642 10124
rect 2746 10112 2774 10152
rect 15746 10140 15752 10152
rect 15804 10140 15810 10192
rect 16114 10140 16120 10192
rect 16172 10180 16178 10192
rect 16853 10183 16911 10189
rect 16853 10180 16865 10183
rect 16172 10152 16865 10180
rect 16172 10140 16178 10152
rect 16853 10149 16865 10152
rect 16899 10149 16911 10183
rect 16853 10143 16911 10149
rect 1636 10084 2774 10112
rect 1636 10072 1642 10084
rect 2958 10072 2964 10124
rect 3016 10121 3022 10124
rect 3016 10112 3028 10121
rect 4433 10115 4491 10121
rect 3016 10084 3061 10112
rect 3016 10075 3028 10084
rect 4433 10081 4445 10115
rect 4479 10112 4491 10115
rect 5074 10112 5080 10124
rect 4479 10084 5080 10112
rect 4479 10081 4491 10084
rect 4433 10075 4491 10081
rect 3016 10072 3022 10075
rect 5074 10072 5080 10084
rect 5132 10072 5138 10124
rect 5528 10115 5586 10121
rect 5528 10081 5540 10115
rect 5574 10112 5586 10115
rect 6822 10112 6828 10124
rect 5574 10084 6828 10112
rect 5574 10081 5586 10084
rect 5528 10075 5586 10081
rect 6822 10072 6828 10084
rect 6880 10112 6886 10124
rect 8113 10115 8171 10121
rect 6880 10084 7604 10112
rect 6880 10072 6886 10084
rect 3237 10047 3295 10053
rect 3237 10013 3249 10047
rect 3283 10013 3295 10047
rect 3237 10007 3295 10013
rect 3252 9976 3280 10007
rect 4062 10004 4068 10056
rect 4120 10044 4126 10056
rect 4157 10047 4215 10053
rect 4157 10044 4169 10047
rect 4120 10016 4169 10044
rect 4120 10004 4126 10016
rect 4157 10013 4169 10016
rect 4203 10013 4215 10047
rect 4338 10044 4344 10056
rect 4299 10016 4344 10044
rect 4157 10007 4215 10013
rect 4338 10004 4344 10016
rect 4396 10004 4402 10056
rect 5261 10047 5319 10053
rect 5261 10013 5273 10047
rect 5307 10013 5319 10047
rect 7098 10044 7104 10056
rect 7059 10016 7104 10044
rect 5261 10007 5319 10013
rect 4246 9976 4252 9988
rect 3252 9948 4252 9976
rect 4246 9936 4252 9948
rect 4304 9976 4310 9988
rect 4890 9976 4896 9988
rect 4304 9948 4896 9976
rect 4304 9936 4310 9948
rect 4890 9936 4896 9948
rect 4948 9976 4954 9988
rect 5276 9976 5304 10007
rect 7098 10004 7104 10016
rect 7156 10004 7162 10056
rect 7576 10044 7604 10084
rect 8113 10081 8125 10115
rect 8159 10112 8171 10115
rect 9582 10112 9588 10124
rect 8159 10084 9588 10112
rect 8159 10081 8171 10084
rect 8113 10075 8171 10081
rect 9582 10072 9588 10084
rect 9640 10072 9646 10124
rect 9674 10072 9680 10124
rect 9732 10112 9738 10124
rect 10422 10115 10480 10121
rect 10422 10112 10434 10115
rect 9732 10084 10434 10112
rect 9732 10072 9738 10084
rect 10422 10081 10434 10084
rect 10468 10081 10480 10115
rect 10686 10112 10692 10124
rect 10647 10084 10692 10112
rect 10422 10075 10480 10081
rect 10686 10072 10692 10084
rect 10744 10072 10750 10124
rect 11054 10072 11060 10124
rect 11112 10112 11118 10124
rect 11425 10115 11483 10121
rect 11425 10112 11437 10115
rect 11112 10084 11437 10112
rect 11112 10072 11118 10084
rect 11425 10081 11437 10084
rect 11471 10112 11483 10115
rect 12526 10112 12532 10124
rect 11471 10084 12532 10112
rect 11471 10081 11483 10084
rect 11425 10075 11483 10081
rect 12526 10072 12532 10084
rect 12584 10072 12590 10124
rect 8297 10047 8355 10053
rect 8297 10044 8309 10047
rect 7576 10016 8309 10044
rect 8297 10013 8309 10016
rect 8343 10013 8355 10047
rect 11238 10044 11244 10056
rect 11199 10016 11244 10044
rect 8297 10007 8355 10013
rect 4948 9948 5304 9976
rect 8312 9976 8340 10007
rect 11238 10004 11244 10016
rect 11296 10004 11302 10056
rect 16761 10047 16819 10053
rect 16761 10013 16773 10047
rect 16807 10044 16819 10047
rect 17586 10044 17592 10056
rect 16807 10016 17592 10044
rect 16807 10013 16819 10016
rect 16761 10007 16819 10013
rect 17586 10004 17592 10016
rect 17644 10004 17650 10056
rect 9309 9979 9367 9985
rect 9309 9976 9321 9979
rect 8312 9948 9321 9976
rect 4948 9936 4954 9948
rect 9309 9945 9321 9948
rect 9355 9945 9367 9979
rect 9309 9939 9367 9945
rect 1857 9911 1915 9917
rect 1857 9877 1869 9911
rect 1903 9908 1915 9911
rect 2038 9908 2044 9920
rect 1903 9880 2044 9908
rect 1903 9877 1915 9880
rect 1857 9871 1915 9877
rect 2038 9868 2044 9880
rect 2096 9868 2102 9920
rect 1104 9818 21896 9840
rect 1104 9766 4447 9818
rect 4499 9766 4511 9818
rect 4563 9766 4575 9818
rect 4627 9766 4639 9818
rect 4691 9766 11378 9818
rect 11430 9766 11442 9818
rect 11494 9766 11506 9818
rect 11558 9766 11570 9818
rect 11622 9766 18308 9818
rect 18360 9766 18372 9818
rect 18424 9766 18436 9818
rect 18488 9766 18500 9818
rect 18552 9766 21896 9818
rect 1104 9744 21896 9766
rect 9309 9707 9367 9713
rect 9309 9673 9321 9707
rect 9355 9704 9367 9707
rect 9674 9704 9680 9716
rect 9355 9676 9680 9704
rect 9355 9673 9367 9676
rect 9309 9667 9367 9673
rect 9674 9664 9680 9676
rect 9732 9664 9738 9716
rect 11054 9704 11060 9716
rect 11015 9676 11060 9704
rect 11054 9664 11060 9676
rect 11112 9664 11118 9716
rect 1581 9639 1639 9645
rect 1581 9605 1593 9639
rect 1627 9636 1639 9639
rect 2314 9636 2320 9648
rect 1627 9608 2320 9636
rect 1627 9605 1639 9608
rect 1581 9599 1639 9605
rect 2314 9596 2320 9608
rect 2372 9596 2378 9648
rect 2866 9596 2872 9648
rect 2924 9636 2930 9648
rect 2961 9639 3019 9645
rect 2961 9636 2973 9639
rect 2924 9608 2973 9636
rect 2924 9596 2930 9608
rect 2961 9605 2973 9608
rect 3007 9605 3019 9639
rect 2961 9599 3019 9605
rect 3878 9596 3884 9648
rect 3936 9636 3942 9648
rect 4709 9639 4767 9645
rect 4709 9636 4721 9639
rect 3936 9608 4721 9636
rect 3936 9596 3942 9608
rect 4709 9605 4721 9608
rect 4755 9636 4767 9639
rect 5074 9636 5080 9648
rect 4755 9608 5080 9636
rect 4755 9605 4767 9608
rect 4709 9599 4767 9605
rect 5074 9596 5080 9608
rect 5132 9596 5138 9648
rect 6638 9636 6644 9648
rect 6599 9608 6644 9636
rect 6638 9596 6644 9608
rect 6696 9596 6702 9648
rect 9582 9636 9588 9648
rect 9543 9608 9588 9636
rect 9582 9596 9588 9608
rect 9640 9596 9646 9648
rect 2685 9571 2743 9577
rect 2685 9537 2697 9571
rect 2731 9568 2743 9571
rect 2774 9568 2780 9580
rect 2731 9540 2780 9568
rect 2731 9537 2743 9540
rect 2685 9531 2743 9537
rect 2774 9528 2780 9540
rect 2832 9528 2838 9580
rect 3605 9571 3663 9577
rect 3605 9537 3617 9571
rect 3651 9568 3663 9571
rect 4062 9568 4068 9580
rect 3651 9540 4068 9568
rect 3651 9537 3663 9540
rect 3605 9531 3663 9537
rect 4062 9528 4068 9540
rect 4120 9528 4126 9580
rect 4982 9568 4988 9580
rect 4264 9540 4988 9568
rect 1394 9500 1400 9512
rect 1355 9472 1400 9500
rect 1394 9460 1400 9472
rect 1452 9460 1458 9512
rect 1854 9500 1860 9512
rect 1815 9472 1860 9500
rect 1854 9460 1860 9472
rect 1912 9460 1918 9512
rect 3329 9503 3387 9509
rect 3329 9469 3341 9503
rect 3375 9500 3387 9503
rect 4264 9500 4292 9540
rect 4982 9528 4988 9540
rect 5040 9528 5046 9580
rect 6822 9528 6828 9580
rect 6880 9568 6886 9580
rect 7193 9571 7251 9577
rect 7193 9568 7205 9571
rect 6880 9540 7205 9568
rect 6880 9528 6886 9540
rect 7193 9537 7205 9540
rect 7239 9537 7251 9571
rect 7193 9531 7251 9537
rect 7650 9528 7656 9580
rect 7708 9568 7714 9580
rect 7929 9571 7987 9577
rect 7929 9568 7941 9571
rect 7708 9540 7941 9568
rect 7708 9528 7714 9540
rect 7929 9537 7941 9540
rect 7975 9537 7987 9571
rect 9692 9568 9720 9664
rect 10137 9571 10195 9577
rect 10137 9568 10149 9571
rect 9692 9540 10149 9568
rect 7929 9531 7987 9537
rect 10137 9537 10149 9540
rect 10183 9537 10195 9571
rect 10137 9531 10195 9537
rect 3375 9472 4292 9500
rect 3375 9469 3387 9472
rect 3329 9463 3387 9469
rect 4338 9460 4344 9512
rect 4396 9500 4402 9512
rect 4433 9503 4491 9509
rect 4433 9500 4445 9503
rect 4396 9472 4445 9500
rect 4396 9460 4402 9472
rect 4433 9469 4445 9472
rect 4479 9500 4491 9503
rect 5350 9500 5356 9512
rect 4479 9472 5356 9500
rect 4479 9469 4491 9472
rect 4433 9463 4491 9469
rect 5350 9460 5356 9472
rect 5408 9460 5414 9512
rect 7009 9503 7067 9509
rect 7009 9469 7021 9503
rect 7055 9500 7067 9503
rect 7098 9500 7104 9512
rect 7055 9472 7104 9500
rect 7055 9469 7067 9472
rect 7009 9463 7067 9469
rect 7098 9460 7104 9472
rect 7156 9460 7162 9512
rect 9766 9460 9772 9512
rect 9824 9500 9830 9512
rect 10045 9503 10103 9509
rect 10045 9500 10057 9503
rect 9824 9472 10057 9500
rect 9824 9460 9830 9472
rect 10045 9469 10057 9472
rect 10091 9469 10103 9503
rect 10045 9463 10103 9469
rect 2746 9404 7236 9432
rect 2041 9367 2099 9373
rect 2041 9333 2053 9367
rect 2087 9364 2099 9367
rect 2746 9364 2774 9404
rect 3418 9364 3424 9376
rect 2087 9336 2774 9364
rect 3379 9336 3424 9364
rect 2087 9333 2099 9336
rect 2041 9327 2099 9333
rect 3418 9324 3424 9336
rect 3476 9364 3482 9376
rect 3973 9367 4031 9373
rect 3973 9364 3985 9367
rect 3476 9336 3985 9364
rect 3476 9324 3482 9336
rect 3973 9333 3985 9336
rect 4019 9333 4031 9367
rect 3973 9327 4031 9333
rect 4062 9324 4068 9376
rect 4120 9364 4126 9376
rect 6546 9364 6552 9376
rect 4120 9336 6552 9364
rect 4120 9324 4126 9336
rect 6546 9324 6552 9336
rect 6604 9364 6610 9376
rect 7101 9367 7159 9373
rect 7101 9364 7113 9367
rect 6604 9336 7113 9364
rect 6604 9324 6610 9336
rect 7101 9333 7113 9336
rect 7147 9333 7159 9367
rect 7208 9364 7236 9404
rect 7650 9392 7656 9444
rect 7708 9432 7714 9444
rect 8174 9435 8232 9441
rect 8174 9432 8186 9435
rect 7708 9404 8186 9432
rect 7708 9392 7714 9404
rect 8174 9401 8186 9404
rect 8220 9401 8232 9435
rect 8174 9395 8232 9401
rect 8312 9404 12434 9432
rect 8312 9364 8340 9404
rect 7208 9336 8340 9364
rect 7101 9327 7159 9333
rect 8846 9324 8852 9376
rect 8904 9364 8910 9376
rect 9398 9364 9404 9376
rect 8904 9336 9404 9364
rect 8904 9324 8910 9336
rect 9398 9324 9404 9336
rect 9456 9364 9462 9376
rect 9953 9367 10011 9373
rect 9953 9364 9965 9367
rect 9456 9336 9965 9364
rect 9456 9324 9462 9336
rect 9953 9333 9965 9336
rect 9999 9333 10011 9367
rect 12406 9364 12434 9404
rect 14090 9364 14096 9376
rect 12406 9336 14096 9364
rect 9953 9327 10011 9333
rect 14090 9324 14096 9336
rect 14148 9324 14154 9376
rect 1104 9274 21896 9296
rect 1104 9222 7912 9274
rect 7964 9222 7976 9274
rect 8028 9222 8040 9274
rect 8092 9222 8104 9274
rect 8156 9222 14843 9274
rect 14895 9222 14907 9274
rect 14959 9222 14971 9274
rect 15023 9222 15035 9274
rect 15087 9222 21896 9274
rect 1104 9200 21896 9222
rect 1854 9120 1860 9172
rect 1912 9160 1918 9172
rect 3145 9163 3203 9169
rect 3145 9160 3157 9163
rect 1912 9132 3157 9160
rect 1912 9120 1918 9132
rect 3145 9129 3157 9132
rect 3191 9129 3203 9163
rect 3145 9123 3203 9129
rect 5353 9163 5411 9169
rect 5353 9129 5365 9163
rect 5399 9160 5411 9163
rect 5442 9160 5448 9172
rect 5399 9132 5448 9160
rect 5399 9129 5411 9132
rect 5353 9123 5411 9129
rect 5442 9120 5448 9132
rect 5500 9120 5506 9172
rect 7101 9163 7159 9169
rect 7101 9129 7113 9163
rect 7147 9129 7159 9163
rect 9766 9160 9772 9172
rect 9727 9132 9772 9160
rect 7101 9123 7159 9129
rect 1394 9092 1400 9104
rect 1355 9064 1400 9092
rect 1394 9052 1400 9064
rect 1452 9052 1458 9104
rect 7116 9092 7144 9123
rect 9766 9120 9772 9132
rect 9824 9120 9830 9172
rect 8938 9092 8944 9104
rect 2424 9064 7144 9092
rect 7208 9064 8944 9092
rect 2424 9033 2452 9064
rect 1765 9027 1823 9033
rect 1765 8993 1777 9027
rect 1811 9024 1823 9027
rect 2409 9027 2467 9033
rect 1811 8996 2268 9024
rect 1811 8993 1823 8996
rect 1765 8987 1823 8993
rect 1949 8891 2007 8897
rect 1949 8857 1961 8891
rect 1995 8888 2007 8891
rect 2130 8888 2136 8900
rect 1995 8860 2136 8888
rect 1995 8857 2007 8860
rect 1949 8851 2007 8857
rect 2130 8848 2136 8860
rect 2188 8848 2194 8900
rect 2240 8897 2268 8996
rect 2409 8993 2421 9027
rect 2455 8993 2467 9027
rect 2409 8987 2467 8993
rect 2685 9027 2743 9033
rect 2685 8993 2697 9027
rect 2731 9024 2743 9027
rect 2774 9024 2780 9036
rect 2731 8996 2780 9024
rect 2731 8993 2743 8996
rect 2685 8987 2743 8993
rect 2774 8984 2780 8996
rect 2832 9024 2838 9036
rect 3881 9027 3939 9033
rect 3881 9024 3893 9027
rect 2832 8996 3893 9024
rect 2832 8984 2838 8996
rect 3881 8993 3893 8996
rect 3927 8993 3939 9027
rect 5261 9027 5319 9033
rect 5261 9024 5273 9027
rect 3881 8987 3939 8993
rect 5092 8996 5273 9024
rect 2590 8916 2596 8968
rect 2648 8956 2654 8968
rect 5092 8956 5120 8996
rect 5261 8993 5273 8996
rect 5307 9024 5319 9027
rect 7208 9024 7236 9064
rect 8938 9052 8944 9064
rect 8996 9052 9002 9104
rect 5307 8996 7236 9024
rect 5307 8993 5319 8996
rect 5261 8987 5319 8993
rect 7282 8984 7288 9036
rect 7340 9024 7346 9036
rect 7469 9027 7527 9033
rect 7469 9024 7481 9027
rect 7340 8996 7481 9024
rect 7340 8984 7346 8996
rect 7469 8993 7481 8996
rect 7515 8993 7527 9027
rect 7469 8987 7527 8993
rect 7561 9027 7619 9033
rect 7561 8993 7573 9027
rect 7607 9024 7619 9027
rect 9306 9024 9312 9036
rect 7607 8996 9312 9024
rect 7607 8993 7619 8996
rect 7561 8987 7619 8993
rect 9306 8984 9312 8996
rect 9364 8984 9370 9036
rect 2648 8928 5120 8956
rect 2648 8916 2654 8928
rect 5166 8916 5172 8968
rect 5224 8956 5230 8968
rect 5445 8959 5503 8965
rect 5445 8956 5457 8959
rect 5224 8928 5457 8956
rect 5224 8916 5230 8928
rect 5445 8925 5457 8928
rect 5491 8925 5503 8959
rect 5445 8919 5503 8925
rect 7650 8916 7656 8968
rect 7708 8956 7714 8968
rect 7708 8928 7753 8956
rect 7708 8916 7714 8928
rect 2225 8891 2283 8897
rect 2225 8857 2237 8891
rect 2271 8857 2283 8891
rect 2225 8851 2283 8857
rect 2869 8891 2927 8897
rect 2869 8857 2881 8891
rect 2915 8888 2927 8891
rect 17494 8888 17500 8900
rect 2915 8860 17500 8888
rect 2915 8857 2927 8860
rect 2869 8851 2927 8857
rect 17494 8848 17500 8860
rect 17552 8848 17558 8900
rect 4798 8780 4804 8832
rect 4856 8820 4862 8832
rect 4893 8823 4951 8829
rect 4893 8820 4905 8823
rect 4856 8792 4905 8820
rect 4856 8780 4862 8792
rect 4893 8789 4905 8792
rect 4939 8789 4951 8823
rect 9398 8820 9404 8832
rect 9359 8792 9404 8820
rect 4893 8783 4951 8789
rect 9398 8780 9404 8792
rect 9456 8780 9462 8832
rect 1104 8730 21896 8752
rect 1104 8678 4447 8730
rect 4499 8678 4511 8730
rect 4563 8678 4575 8730
rect 4627 8678 4639 8730
rect 4691 8678 11378 8730
rect 11430 8678 11442 8730
rect 11494 8678 11506 8730
rect 11558 8678 11570 8730
rect 11622 8678 18308 8730
rect 18360 8678 18372 8730
rect 18424 8678 18436 8730
rect 18488 8678 18500 8730
rect 18552 8678 21896 8730
rect 1104 8656 21896 8678
rect 1765 8619 1823 8625
rect 1765 8585 1777 8619
rect 1811 8616 1823 8619
rect 1946 8616 1952 8628
rect 1811 8588 1952 8616
rect 1811 8585 1823 8588
rect 1765 8579 1823 8585
rect 1946 8576 1952 8588
rect 2004 8576 2010 8628
rect 3697 8619 3755 8625
rect 3697 8585 3709 8619
rect 3743 8616 3755 8619
rect 5166 8616 5172 8628
rect 3743 8588 5172 8616
rect 3743 8585 3755 8588
rect 3697 8579 3755 8585
rect 5166 8576 5172 8588
rect 5224 8576 5230 8628
rect 9033 8551 9091 8557
rect 9033 8517 9045 8551
rect 9079 8548 9091 8551
rect 9766 8548 9772 8560
rect 9079 8520 9772 8548
rect 9079 8517 9091 8520
rect 9033 8511 9091 8517
rect 9766 8508 9772 8520
rect 9824 8508 9830 8560
rect 8386 8480 8392 8492
rect 8347 8452 8392 8480
rect 8386 8440 8392 8452
rect 8444 8440 8450 8492
rect 8573 8483 8631 8489
rect 8573 8449 8585 8483
rect 8619 8480 8631 8483
rect 13078 8480 13084 8492
rect 8619 8452 13084 8480
rect 8619 8449 8631 8452
rect 8573 8443 8631 8449
rect 13078 8440 13084 8452
rect 13136 8440 13142 8492
rect 1946 8412 1952 8424
rect 1907 8384 1952 8412
rect 1946 8372 1952 8384
rect 2004 8372 2010 8424
rect 2317 8415 2375 8421
rect 2317 8381 2329 8415
rect 2363 8412 2375 8415
rect 4065 8415 4123 8421
rect 4065 8412 4077 8415
rect 2363 8384 4077 8412
rect 2363 8381 2375 8384
rect 2317 8375 2375 8381
rect 4065 8381 4077 8384
rect 4111 8412 4123 8415
rect 4890 8412 4896 8424
rect 4111 8384 4896 8412
rect 4111 8381 4123 8384
rect 4065 8375 4123 8381
rect 4890 8372 4896 8384
rect 4948 8412 4954 8424
rect 6641 8415 6699 8421
rect 6641 8412 6653 8415
rect 4948 8384 6653 8412
rect 4948 8372 4954 8384
rect 6641 8381 6653 8384
rect 6687 8381 6699 8415
rect 6641 8375 6699 8381
rect 6908 8415 6966 8421
rect 6908 8381 6920 8415
rect 6954 8412 6966 8415
rect 8404 8412 8432 8440
rect 6954 8384 8432 8412
rect 6954 8381 6966 8384
rect 6908 8375 6966 8381
rect 2038 8304 2044 8356
rect 2096 8344 2102 8356
rect 2562 8347 2620 8353
rect 2562 8344 2574 8347
rect 2096 8316 2574 8344
rect 2096 8304 2102 8316
rect 2562 8313 2574 8316
rect 2608 8313 2620 8347
rect 2562 8307 2620 8313
rect 4246 8304 4252 8356
rect 4304 8353 4310 8356
rect 4304 8347 4368 8353
rect 4304 8313 4322 8347
rect 4356 8313 4368 8347
rect 4304 8307 4368 8313
rect 4304 8304 4310 8307
rect 8294 8304 8300 8356
rect 8352 8344 8358 8356
rect 8665 8347 8723 8353
rect 8665 8344 8677 8347
rect 8352 8316 8677 8344
rect 8352 8304 8358 8316
rect 8665 8313 8677 8316
rect 8711 8313 8723 8347
rect 8665 8307 8723 8313
rect 1394 8276 1400 8288
rect 1355 8248 1400 8276
rect 1394 8236 1400 8248
rect 1452 8236 1458 8288
rect 4430 8236 4436 8288
rect 4488 8276 4494 8288
rect 5442 8276 5448 8288
rect 4488 8248 5448 8276
rect 4488 8236 4494 8248
rect 5442 8236 5448 8248
rect 5500 8236 5506 8288
rect 8021 8279 8079 8285
rect 8021 8245 8033 8279
rect 8067 8276 8079 8279
rect 8202 8276 8208 8288
rect 8067 8248 8208 8276
rect 8067 8245 8079 8248
rect 8021 8239 8079 8245
rect 8202 8236 8208 8248
rect 8260 8236 8266 8288
rect 1104 8186 21896 8208
rect 1104 8134 7912 8186
rect 7964 8134 7976 8186
rect 8028 8134 8040 8186
rect 8092 8134 8104 8186
rect 8156 8134 14843 8186
rect 14895 8134 14907 8186
rect 14959 8134 14971 8186
rect 15023 8134 15035 8186
rect 15087 8134 21896 8186
rect 1104 8112 21896 8134
rect 1578 8072 1584 8084
rect 1539 8044 1584 8072
rect 1578 8032 1584 8044
rect 1636 8032 1642 8084
rect 1946 8032 1952 8084
rect 2004 8072 2010 8084
rect 2041 8075 2099 8081
rect 2041 8072 2053 8075
rect 2004 8044 2053 8072
rect 2004 8032 2010 8044
rect 2041 8041 2053 8044
rect 2087 8041 2099 8075
rect 2041 8035 2099 8041
rect 2777 8075 2835 8081
rect 2777 8041 2789 8075
rect 2823 8041 2835 8075
rect 2777 8035 2835 8041
rect 7377 8075 7435 8081
rect 7377 8041 7389 8075
rect 7423 8072 7435 8075
rect 7650 8072 7656 8084
rect 7423 8044 7656 8072
rect 7423 8041 7435 8044
rect 7377 8035 7435 8041
rect 1394 7936 1400 7948
rect 1355 7908 1400 7936
rect 1394 7896 1400 7908
rect 1452 7896 1458 7948
rect 2225 7939 2283 7945
rect 2225 7905 2237 7939
rect 2271 7936 2283 7939
rect 2792 7936 2820 8035
rect 7650 8032 7656 8044
rect 7708 8032 7714 8084
rect 9306 8072 9312 8084
rect 9267 8044 9312 8072
rect 9306 8032 9312 8044
rect 9364 8032 9370 8084
rect 9766 8072 9772 8084
rect 9727 8044 9772 8072
rect 9766 8032 9772 8044
rect 9824 8032 9830 8084
rect 3237 8007 3295 8013
rect 3237 7973 3249 8007
rect 3283 8004 3295 8007
rect 4338 8004 4344 8016
rect 3283 7976 4344 8004
rect 3283 7973 3295 7976
rect 3237 7967 3295 7973
rect 4338 7964 4344 7976
rect 4396 7964 4402 8016
rect 5166 7964 5172 8016
rect 5224 8013 5230 8016
rect 5224 8004 5236 8013
rect 5224 7976 5269 8004
rect 5224 7967 5236 7976
rect 5224 7964 5230 7967
rect 5442 7964 5448 8016
rect 5500 8004 5506 8016
rect 5966 8007 6024 8013
rect 5966 8004 5978 8007
rect 5500 7976 5978 8004
rect 5500 7964 5506 7976
rect 5966 7973 5978 7976
rect 6012 7973 6024 8007
rect 5966 7967 6024 7973
rect 7742 7964 7748 8016
rect 7800 8004 7806 8016
rect 7800 7976 8800 8004
rect 7800 7964 7806 7976
rect 2271 7908 2820 7936
rect 3145 7939 3203 7945
rect 2271 7905 2283 7908
rect 2225 7899 2283 7905
rect 3145 7905 3157 7939
rect 3191 7936 3203 7939
rect 3602 7936 3608 7948
rect 3191 7908 3608 7936
rect 3191 7905 3203 7908
rect 3145 7899 3203 7905
rect 3602 7896 3608 7908
rect 3660 7896 3666 7948
rect 4890 7896 4896 7948
rect 4948 7936 4954 7948
rect 5721 7939 5779 7945
rect 5721 7936 5733 7939
rect 4948 7908 5733 7936
rect 4948 7896 4954 7908
rect 3421 7871 3479 7877
rect 3421 7837 3433 7871
rect 3467 7868 3479 7871
rect 4430 7868 4436 7880
rect 3467 7840 4436 7868
rect 3467 7837 3479 7840
rect 3421 7831 3479 7837
rect 4430 7828 4436 7840
rect 4488 7828 4494 7880
rect 5460 7877 5488 7908
rect 5721 7905 5733 7908
rect 5767 7905 5779 7939
rect 5721 7899 5779 7905
rect 8202 7896 8208 7948
rect 8260 7936 8266 7948
rect 8772 7945 8800 7976
rect 8490 7939 8548 7945
rect 8490 7936 8502 7939
rect 8260 7908 8502 7936
rect 8260 7896 8266 7908
rect 8490 7905 8502 7908
rect 8536 7936 8548 7939
rect 8757 7939 8815 7945
rect 8536 7908 8708 7936
rect 8536 7905 8548 7908
rect 8490 7899 8548 7905
rect 5445 7871 5503 7877
rect 5445 7837 5457 7871
rect 5491 7837 5503 7871
rect 8680 7868 8708 7908
rect 8757 7905 8769 7939
rect 8803 7905 8815 7939
rect 8757 7899 8815 7905
rect 8846 7896 8852 7948
rect 8904 7936 8910 7948
rect 9677 7939 9735 7945
rect 9677 7936 9689 7939
rect 8904 7908 9689 7936
rect 8904 7896 8910 7908
rect 9677 7905 9689 7908
rect 9723 7905 9735 7939
rect 9677 7899 9735 7905
rect 9861 7871 9919 7877
rect 9861 7868 9873 7871
rect 8680 7840 9873 7868
rect 5445 7831 5503 7837
rect 9861 7837 9873 7840
rect 9907 7837 9919 7871
rect 9861 7831 9919 7837
rect 4065 7735 4123 7741
rect 4065 7701 4077 7735
rect 4111 7732 4123 7735
rect 4246 7732 4252 7744
rect 4111 7704 4252 7732
rect 4111 7701 4123 7704
rect 4065 7695 4123 7701
rect 4246 7692 4252 7704
rect 4304 7692 4310 7744
rect 7101 7735 7159 7741
rect 7101 7701 7113 7735
rect 7147 7732 7159 7735
rect 8386 7732 8392 7744
rect 7147 7704 8392 7732
rect 7147 7701 7159 7704
rect 7101 7695 7159 7701
rect 8386 7692 8392 7704
rect 8444 7692 8450 7744
rect 1104 7642 21896 7664
rect 1104 7590 4447 7642
rect 4499 7590 4511 7642
rect 4563 7590 4575 7642
rect 4627 7590 4639 7642
rect 4691 7590 11378 7642
rect 11430 7590 11442 7642
rect 11494 7590 11506 7642
rect 11558 7590 11570 7642
rect 11622 7590 18308 7642
rect 18360 7590 18372 7642
rect 18424 7590 18436 7642
rect 18488 7590 18500 7642
rect 18552 7590 21896 7642
rect 1104 7568 21896 7590
rect 3602 7528 3608 7540
rect 3563 7500 3608 7528
rect 3602 7488 3608 7500
rect 3660 7488 3666 7540
rect 3694 7488 3700 7540
rect 3752 7528 3758 7540
rect 6733 7531 6791 7537
rect 6733 7528 6745 7531
rect 3752 7500 6745 7528
rect 3752 7488 3758 7500
rect 6733 7497 6745 7500
rect 6779 7528 6791 7531
rect 7009 7531 7067 7537
rect 7009 7528 7021 7531
rect 6779 7500 7021 7528
rect 6779 7497 6791 7500
rect 6733 7491 6791 7497
rect 7009 7497 7021 7500
rect 7055 7497 7067 7531
rect 8846 7528 8852 7540
rect 8807 7500 8852 7528
rect 7009 7491 7067 7497
rect 8846 7488 8852 7500
rect 8904 7488 8910 7540
rect 18601 7531 18659 7537
rect 18601 7497 18613 7531
rect 18647 7528 18659 7531
rect 18874 7528 18880 7540
rect 18647 7500 18880 7528
rect 18647 7497 18659 7500
rect 18601 7491 18659 7497
rect 18874 7488 18880 7500
rect 18932 7488 18938 7540
rect 19245 7531 19303 7537
rect 19245 7497 19257 7531
rect 19291 7528 19303 7531
rect 19702 7528 19708 7540
rect 19291 7500 19708 7528
rect 19291 7497 19303 7500
rect 19245 7491 19303 7497
rect 19702 7488 19708 7500
rect 19760 7488 19766 7540
rect 2041 7463 2099 7469
rect 2041 7429 2053 7463
rect 2087 7460 2099 7463
rect 6914 7460 6920 7472
rect 2087 7432 6920 7460
rect 2087 7429 2099 7432
rect 2041 7423 2099 7429
rect 6914 7420 6920 7432
rect 6972 7420 6978 7472
rect 7190 7420 7196 7472
rect 7248 7460 7254 7472
rect 17218 7460 17224 7472
rect 7248 7432 17224 7460
rect 7248 7420 7254 7432
rect 17218 7420 17224 7432
rect 17276 7420 17282 7472
rect 4246 7392 4252 7404
rect 4207 7364 4252 7392
rect 4246 7352 4252 7364
rect 4304 7352 4310 7404
rect 5166 7392 5172 7404
rect 5127 7364 5172 7392
rect 5166 7352 5172 7364
rect 5224 7352 5230 7404
rect 7285 7395 7343 7401
rect 7285 7361 7297 7395
rect 7331 7392 7343 7395
rect 8297 7395 8355 7401
rect 8297 7392 8309 7395
rect 7331 7364 8309 7392
rect 7331 7361 7343 7364
rect 7285 7355 7343 7361
rect 8297 7361 8309 7364
rect 8343 7392 8355 7395
rect 8386 7392 8392 7404
rect 8343 7364 8392 7392
rect 8343 7361 8355 7364
rect 8297 7355 8355 7361
rect 8386 7352 8392 7364
rect 8444 7352 8450 7404
rect 1394 7324 1400 7336
rect 1355 7296 1400 7324
rect 1394 7284 1400 7296
rect 1452 7284 1458 7336
rect 1854 7324 1860 7336
rect 1815 7296 1860 7324
rect 1854 7284 1860 7296
rect 1912 7324 1918 7336
rect 2685 7327 2743 7333
rect 2685 7324 2697 7327
rect 1912 7296 2697 7324
rect 1912 7284 1918 7296
rect 2685 7293 2697 7296
rect 2731 7293 2743 7327
rect 2685 7287 2743 7293
rect 4982 7284 4988 7336
rect 5040 7324 5046 7336
rect 7469 7327 7527 7333
rect 7469 7324 7481 7327
rect 5040 7296 7481 7324
rect 5040 7284 5046 7296
rect 7469 7293 7481 7296
rect 7515 7293 7527 7327
rect 7469 7287 7527 7293
rect 7558 7284 7564 7336
rect 7616 7324 7622 7336
rect 9398 7324 9404 7336
rect 7616 7296 9404 7324
rect 7616 7284 7622 7296
rect 9398 7284 9404 7296
rect 9456 7284 9462 7336
rect 18782 7324 18788 7336
rect 18743 7296 18788 7324
rect 18782 7284 18788 7296
rect 18840 7284 18846 7336
rect 19058 7324 19064 7336
rect 19019 7296 19064 7324
rect 19058 7284 19064 7296
rect 19116 7284 19122 7336
rect 1412 7256 1440 7284
rect 2317 7259 2375 7265
rect 2317 7256 2329 7259
rect 1412 7228 2329 7256
rect 2317 7225 2329 7228
rect 2363 7225 2375 7259
rect 2317 7219 2375 7225
rect 3973 7259 4031 7265
rect 3973 7225 3985 7259
rect 4019 7256 4031 7259
rect 5629 7259 5687 7265
rect 5629 7256 5641 7259
rect 4019 7228 5641 7256
rect 4019 7225 4031 7228
rect 3973 7219 4031 7225
rect 5629 7225 5641 7228
rect 5675 7225 5687 7259
rect 8389 7259 8447 7265
rect 8389 7256 8401 7259
rect 5629 7219 5687 7225
rect 6104 7228 8401 7256
rect 1578 7188 1584 7200
rect 1539 7160 1584 7188
rect 1578 7148 1584 7160
rect 1636 7148 1642 7200
rect 3234 7188 3240 7200
rect 3195 7160 3240 7188
rect 3234 7148 3240 7160
rect 3292 7148 3298 7200
rect 4062 7188 4068 7200
rect 4023 7160 4068 7188
rect 4062 7148 4068 7160
rect 4120 7148 4126 7200
rect 4617 7191 4675 7197
rect 4617 7157 4629 7191
rect 4663 7188 4675 7191
rect 4706 7188 4712 7200
rect 4663 7160 4712 7188
rect 4663 7157 4675 7160
rect 4617 7151 4675 7157
rect 4706 7148 4712 7160
rect 4764 7148 4770 7200
rect 4890 7148 4896 7200
rect 4948 7188 4954 7200
rect 4985 7191 5043 7197
rect 4985 7188 4997 7191
rect 4948 7160 4997 7188
rect 4948 7148 4954 7160
rect 4985 7157 4997 7160
rect 5031 7157 5043 7191
rect 4985 7151 5043 7157
rect 5077 7191 5135 7197
rect 5077 7157 5089 7191
rect 5123 7188 5135 7191
rect 5166 7188 5172 7200
rect 5123 7160 5172 7188
rect 5123 7157 5135 7160
rect 5077 7151 5135 7157
rect 5166 7148 5172 7160
rect 5224 7148 5230 7200
rect 5442 7148 5448 7200
rect 5500 7188 5506 7200
rect 6104 7188 6132 7228
rect 8389 7225 8401 7228
rect 8435 7256 8447 7259
rect 9125 7259 9183 7265
rect 9125 7256 9137 7259
rect 8435 7228 9137 7256
rect 8435 7225 8447 7228
rect 8389 7219 8447 7225
rect 9125 7225 9137 7228
rect 9171 7225 9183 7259
rect 9125 7219 9183 7225
rect 5500 7160 6132 7188
rect 7009 7191 7067 7197
rect 5500 7148 5506 7160
rect 7009 7157 7021 7191
rect 7055 7188 7067 7191
rect 7377 7191 7435 7197
rect 7377 7188 7389 7191
rect 7055 7160 7389 7188
rect 7055 7157 7067 7160
rect 7009 7151 7067 7157
rect 7377 7157 7389 7160
rect 7423 7157 7435 7191
rect 7377 7151 7435 7157
rect 7742 7148 7748 7200
rect 7800 7188 7806 7200
rect 7837 7191 7895 7197
rect 7837 7188 7849 7191
rect 7800 7160 7849 7188
rect 7800 7148 7806 7160
rect 7837 7157 7849 7160
rect 7883 7157 7895 7191
rect 8478 7188 8484 7200
rect 8439 7160 8484 7188
rect 7837 7151 7895 7157
rect 8478 7148 8484 7160
rect 8536 7188 8542 7200
rect 9493 7191 9551 7197
rect 9493 7188 9505 7191
rect 8536 7160 9505 7188
rect 8536 7148 8542 7160
rect 9493 7157 9505 7160
rect 9539 7157 9551 7191
rect 9493 7151 9551 7157
rect 1104 7098 21896 7120
rect 1104 7046 7912 7098
rect 7964 7046 7976 7098
rect 8028 7046 8040 7098
rect 8092 7046 8104 7098
rect 8156 7046 14843 7098
rect 14895 7046 14907 7098
rect 14959 7046 14971 7098
rect 15023 7046 15035 7098
rect 15087 7046 21896 7098
rect 1104 7024 21896 7046
rect 4338 6984 4344 6996
rect 4299 6956 4344 6984
rect 4338 6944 4344 6956
rect 4396 6944 4402 6996
rect 4706 6984 4712 6996
rect 4667 6956 4712 6984
rect 4706 6944 4712 6956
rect 4764 6944 4770 6996
rect 4890 6944 4896 6996
rect 4948 6984 4954 6996
rect 7558 6984 7564 6996
rect 4948 6956 7564 6984
rect 4948 6944 4954 6956
rect 7558 6944 7564 6956
rect 7616 6944 7622 6996
rect 7742 6984 7748 6996
rect 7703 6956 7748 6984
rect 7742 6944 7748 6956
rect 7800 6944 7806 6996
rect 3234 6876 3240 6928
rect 3292 6916 3298 6928
rect 5166 6916 5172 6928
rect 3292 6888 5172 6916
rect 3292 6876 3298 6888
rect 5166 6876 5172 6888
rect 5224 6916 5230 6928
rect 5718 6916 5724 6928
rect 5224 6888 5724 6916
rect 5224 6876 5230 6888
rect 5718 6876 5724 6888
rect 5776 6876 5782 6928
rect 7653 6919 7711 6925
rect 7653 6885 7665 6919
rect 7699 6916 7711 6919
rect 7699 6888 8340 6916
rect 7699 6885 7711 6888
rect 7653 6879 7711 6885
rect 1394 6848 1400 6860
rect 1355 6820 1400 6848
rect 1394 6808 1400 6820
rect 1452 6848 1458 6860
rect 1857 6851 1915 6857
rect 1857 6848 1869 6851
rect 1452 6820 1869 6848
rect 1452 6808 1458 6820
rect 1857 6817 1869 6820
rect 1903 6817 1915 6851
rect 4798 6848 4804 6860
rect 4759 6820 4804 6848
rect 1857 6811 1915 6817
rect 4798 6808 4804 6820
rect 4856 6808 4862 6860
rect 8312 6857 8340 6888
rect 8297 6851 8355 6857
rect 8297 6817 8309 6851
rect 8343 6817 8355 6851
rect 19794 6848 19800 6860
rect 19755 6820 19800 6848
rect 8297 6811 8355 6817
rect 19794 6808 19800 6820
rect 19852 6848 19858 6860
rect 20257 6851 20315 6857
rect 20257 6848 20269 6851
rect 19852 6820 20269 6848
rect 19852 6808 19858 6820
rect 20257 6817 20269 6820
rect 20303 6817 20315 6851
rect 20257 6811 20315 6817
rect 4246 6740 4252 6792
rect 4304 6780 4310 6792
rect 4893 6783 4951 6789
rect 4893 6780 4905 6783
rect 4304 6752 4905 6780
rect 4304 6740 4310 6752
rect 4893 6749 4905 6752
rect 4939 6749 4951 6783
rect 4893 6743 4951 6749
rect 7929 6783 7987 6789
rect 7929 6749 7941 6783
rect 7975 6780 7987 6783
rect 8202 6780 8208 6792
rect 7975 6752 8208 6780
rect 7975 6749 7987 6752
rect 7929 6743 7987 6749
rect 8202 6740 8208 6752
rect 8260 6740 8266 6792
rect 1581 6715 1639 6721
rect 1581 6681 1593 6715
rect 1627 6712 1639 6715
rect 7282 6712 7288 6724
rect 1627 6684 5212 6712
rect 7243 6684 7288 6712
rect 1627 6681 1639 6684
rect 1581 6675 1639 6681
rect 3970 6644 3976 6656
rect 3931 6616 3976 6644
rect 3970 6604 3976 6616
rect 4028 6644 4034 6656
rect 4890 6644 4896 6656
rect 4028 6616 4896 6644
rect 4028 6604 4034 6616
rect 4890 6604 4896 6616
rect 4948 6604 4954 6656
rect 5184 6644 5212 6684
rect 7282 6672 7288 6684
rect 7340 6672 7346 6724
rect 19978 6712 19984 6724
rect 19939 6684 19984 6712
rect 19978 6672 19984 6684
rect 20036 6672 20042 6724
rect 19058 6644 19064 6656
rect 5184 6616 19064 6644
rect 19058 6604 19064 6616
rect 19116 6604 19122 6656
rect 1104 6554 21896 6576
rect 1104 6502 4447 6554
rect 4499 6502 4511 6554
rect 4563 6502 4575 6554
rect 4627 6502 4639 6554
rect 4691 6502 11378 6554
rect 11430 6502 11442 6554
rect 11494 6502 11506 6554
rect 11558 6502 11570 6554
rect 11622 6502 18308 6554
rect 18360 6502 18372 6554
rect 18424 6502 18436 6554
rect 18488 6502 18500 6554
rect 18552 6502 21896 6554
rect 1104 6480 21896 6502
rect 19886 6400 19892 6452
rect 19944 6440 19950 6452
rect 20257 6443 20315 6449
rect 20257 6440 20269 6443
rect 19944 6412 20269 6440
rect 19944 6400 19950 6412
rect 20257 6409 20269 6412
rect 20303 6409 20315 6443
rect 20257 6403 20315 6409
rect 1394 6236 1400 6248
rect 1355 6208 1400 6236
rect 1394 6196 1400 6208
rect 1452 6236 1458 6248
rect 1857 6239 1915 6245
rect 1857 6236 1869 6239
rect 1452 6208 1869 6236
rect 1452 6196 1458 6208
rect 1857 6205 1869 6208
rect 1903 6205 1915 6239
rect 20070 6236 20076 6248
rect 20031 6208 20076 6236
rect 1857 6199 1915 6205
rect 20070 6196 20076 6208
rect 20128 6236 20134 6248
rect 20533 6239 20591 6245
rect 20533 6236 20545 6239
rect 20128 6208 20545 6236
rect 20128 6196 20134 6208
rect 20533 6205 20545 6208
rect 20579 6205 20591 6239
rect 20533 6199 20591 6205
rect 1578 6100 1584 6112
rect 1539 6072 1584 6100
rect 1578 6060 1584 6072
rect 1636 6060 1642 6112
rect 1104 6010 21896 6032
rect 1104 5958 7912 6010
rect 7964 5958 7976 6010
rect 8028 5958 8040 6010
rect 8092 5958 8104 6010
rect 8156 5958 14843 6010
rect 14895 5958 14907 6010
rect 14959 5958 14971 6010
rect 15023 5958 15035 6010
rect 15087 5958 21896 6010
rect 1104 5936 21896 5958
rect 1578 5856 1584 5908
rect 1636 5896 1642 5908
rect 19794 5896 19800 5908
rect 1636 5868 19800 5896
rect 1636 5856 1642 5868
rect 19794 5856 19800 5868
rect 19852 5856 19858 5908
rect 20530 5896 20536 5908
rect 20491 5868 20536 5896
rect 20530 5856 20536 5868
rect 20588 5856 20594 5908
rect 1394 5760 1400 5772
rect 1355 5732 1400 5760
rect 1394 5720 1400 5732
rect 1452 5760 1458 5772
rect 1857 5763 1915 5769
rect 1857 5760 1869 5763
rect 1452 5732 1869 5760
rect 1452 5720 1458 5732
rect 1857 5729 1869 5732
rect 1903 5729 1915 5763
rect 1857 5723 1915 5729
rect 20717 5763 20775 5769
rect 20717 5729 20729 5763
rect 20763 5729 20775 5763
rect 20717 5723 20775 5729
rect 1670 5652 1676 5704
rect 1728 5692 1734 5704
rect 20732 5692 20760 5723
rect 20993 5695 21051 5701
rect 20993 5692 21005 5695
rect 1728 5664 21005 5692
rect 1728 5652 1734 5664
rect 20993 5661 21005 5664
rect 21039 5661 21051 5695
rect 20993 5655 21051 5661
rect 1581 5627 1639 5633
rect 1581 5593 1593 5627
rect 1627 5624 1639 5627
rect 20070 5624 20076 5636
rect 1627 5596 20076 5624
rect 1627 5593 1639 5596
rect 1581 5587 1639 5593
rect 20070 5584 20076 5596
rect 20128 5584 20134 5636
rect 1104 5466 21896 5488
rect 1104 5414 4447 5466
rect 4499 5414 4511 5466
rect 4563 5414 4575 5466
rect 4627 5414 4639 5466
rect 4691 5414 11378 5466
rect 11430 5414 11442 5466
rect 11494 5414 11506 5466
rect 11558 5414 11570 5466
rect 11622 5414 18308 5466
rect 18360 5414 18372 5466
rect 18424 5414 18436 5466
rect 18488 5414 18500 5466
rect 18552 5414 21896 5466
rect 1104 5392 21896 5414
rect 1581 5355 1639 5361
rect 1581 5321 1593 5355
rect 1627 5352 1639 5355
rect 1670 5352 1676 5364
rect 1627 5324 1676 5352
rect 1627 5321 1639 5324
rect 1581 5315 1639 5321
rect 1670 5312 1676 5324
rect 1728 5312 1734 5364
rect 20806 5352 20812 5364
rect 20767 5324 20812 5352
rect 20806 5312 20812 5324
rect 20864 5312 20870 5364
rect 1394 5148 1400 5160
rect 1355 5120 1400 5148
rect 1394 5108 1400 5120
rect 1452 5148 1458 5160
rect 2225 5151 2283 5157
rect 2225 5148 2237 5151
rect 1452 5120 2237 5148
rect 1452 5108 1458 5120
rect 2225 5117 2237 5120
rect 2271 5117 2283 5151
rect 20990 5148 20996 5160
rect 20951 5120 20996 5148
rect 2225 5111 2283 5117
rect 20990 5108 20996 5120
rect 21048 5148 21054 5160
rect 21269 5151 21327 5157
rect 21269 5148 21281 5151
rect 21048 5120 21281 5148
rect 21048 5108 21054 5120
rect 21269 5117 21281 5120
rect 21315 5117 21327 5151
rect 21269 5111 21327 5117
rect 1854 5012 1860 5024
rect 1815 4984 1860 5012
rect 1854 4972 1860 4984
rect 1912 4972 1918 5024
rect 1104 4922 21896 4944
rect 1104 4870 7912 4922
rect 7964 4870 7976 4922
rect 8028 4870 8040 4922
rect 8092 4870 8104 4922
rect 8156 4870 14843 4922
rect 14895 4870 14907 4922
rect 14959 4870 14971 4922
rect 15023 4870 15035 4922
rect 15087 4870 21896 4922
rect 1104 4848 21896 4870
rect 2317 4743 2375 4749
rect 2317 4740 2329 4743
rect 1412 4712 2329 4740
rect 1412 4684 1440 4712
rect 2317 4709 2329 4712
rect 2363 4709 2375 4743
rect 2317 4703 2375 4709
rect 1394 4672 1400 4684
rect 1355 4644 1400 4672
rect 1394 4632 1400 4644
rect 1452 4632 1458 4684
rect 1854 4672 1860 4684
rect 1815 4644 1860 4672
rect 1854 4632 1860 4644
rect 1912 4632 1918 4684
rect 11146 4604 11152 4616
rect 1596 4576 11152 4604
rect 1596 4545 1624 4576
rect 11146 4564 11152 4576
rect 11204 4564 11210 4616
rect 1581 4539 1639 4545
rect 1581 4505 1593 4539
rect 1627 4505 1639 4539
rect 1581 4499 1639 4505
rect 2041 4539 2099 4545
rect 2041 4505 2053 4539
rect 2087 4536 2099 4539
rect 2087 4508 2774 4536
rect 2087 4505 2099 4508
rect 2041 4499 2099 4505
rect 2746 4468 2774 4508
rect 20990 4468 20996 4480
rect 2746 4440 20996 4468
rect 20990 4428 20996 4440
rect 21048 4428 21054 4480
rect 1104 4378 21896 4400
rect 1104 4326 4447 4378
rect 4499 4326 4511 4378
rect 4563 4326 4575 4378
rect 4627 4326 4639 4378
rect 4691 4326 11378 4378
rect 11430 4326 11442 4378
rect 11494 4326 11506 4378
rect 11558 4326 11570 4378
rect 11622 4326 18308 4378
rect 18360 4326 18372 4378
rect 18424 4326 18436 4378
rect 18488 4326 18500 4378
rect 18552 4326 21896 4378
rect 1104 4304 21896 4326
rect 1857 4131 1915 4137
rect 1857 4097 1869 4131
rect 1903 4128 1915 4131
rect 4982 4128 4988 4140
rect 1903 4100 4988 4128
rect 1903 4097 1915 4100
rect 1857 4091 1915 4097
rect 4982 4088 4988 4100
rect 5040 4088 5046 4140
rect 1670 3992 1676 4004
rect 1631 3964 1676 3992
rect 1670 3952 1676 3964
rect 1728 3992 1734 4004
rect 2501 3995 2559 4001
rect 2501 3992 2513 3995
rect 1728 3964 2513 3992
rect 1728 3952 1734 3964
rect 2501 3961 2513 3964
rect 2547 3961 2559 3995
rect 2501 3955 2559 3961
rect 1762 3884 1768 3936
rect 1820 3924 1826 3936
rect 2133 3927 2191 3933
rect 2133 3924 2145 3927
rect 1820 3896 2145 3924
rect 1820 3884 1826 3896
rect 2133 3893 2145 3896
rect 2179 3893 2191 3927
rect 2133 3887 2191 3893
rect 1104 3834 21896 3856
rect 1104 3782 7912 3834
rect 7964 3782 7976 3834
rect 8028 3782 8040 3834
rect 8092 3782 8104 3834
rect 8156 3782 14843 3834
rect 14895 3782 14907 3834
rect 14959 3782 14971 3834
rect 15023 3782 15035 3834
rect 15087 3782 21896 3834
rect 1104 3760 21896 3782
rect 1765 3723 1823 3729
rect 1765 3689 1777 3723
rect 1811 3720 1823 3723
rect 4062 3720 4068 3732
rect 1811 3692 4068 3720
rect 1811 3689 1823 3692
rect 1765 3683 1823 3689
rect 4062 3680 4068 3692
rect 4120 3680 4126 3732
rect 2409 3655 2467 3661
rect 2409 3621 2421 3655
rect 2455 3652 2467 3655
rect 3234 3652 3240 3664
rect 2455 3624 3240 3652
rect 2455 3621 2467 3624
rect 2409 3615 2467 3621
rect 3234 3612 3240 3624
rect 3292 3612 3298 3664
rect 1670 3584 1676 3596
rect 1631 3556 1676 3584
rect 1670 3544 1676 3556
rect 1728 3544 1734 3596
rect 2225 3587 2283 3593
rect 2225 3553 2237 3587
rect 2271 3584 2283 3587
rect 3142 3584 3148 3596
rect 2271 3556 3148 3584
rect 2271 3553 2283 3556
rect 2225 3547 2283 3553
rect 3142 3544 3148 3556
rect 3200 3544 3206 3596
rect 1688 3516 1716 3544
rect 2685 3519 2743 3525
rect 2685 3516 2697 3519
rect 1688 3488 2697 3516
rect 2685 3485 2697 3488
rect 2731 3485 2743 3519
rect 2685 3479 2743 3485
rect 3142 3380 3148 3392
rect 3103 3352 3148 3380
rect 3142 3340 3148 3352
rect 3200 3340 3206 3392
rect 1104 3290 21896 3312
rect 1104 3238 4447 3290
rect 4499 3238 4511 3290
rect 4563 3238 4575 3290
rect 4627 3238 4639 3290
rect 4691 3238 11378 3290
rect 11430 3238 11442 3290
rect 11494 3238 11506 3290
rect 11558 3238 11570 3290
rect 11622 3238 18308 3290
rect 18360 3238 18372 3290
rect 18424 3238 18436 3290
rect 18488 3238 18500 3290
rect 18552 3238 21896 3290
rect 1104 3216 21896 3238
rect 1673 3179 1731 3185
rect 1673 3145 1685 3179
rect 1719 3176 1731 3179
rect 3418 3176 3424 3188
rect 1719 3148 3424 3176
rect 1719 3145 1731 3148
rect 1673 3139 1731 3145
rect 3418 3136 3424 3148
rect 3476 3136 3482 3188
rect 2409 3111 2467 3117
rect 2409 3077 2421 3111
rect 2455 3108 2467 3111
rect 2590 3108 2596 3120
rect 2455 3080 2596 3108
rect 2455 3077 2467 3080
rect 2409 3071 2467 3077
rect 2590 3068 2596 3080
rect 2648 3068 2654 3120
rect 2961 3111 3019 3117
rect 2700 3080 2912 3108
rect 2130 3000 2136 3052
rect 2188 3040 2194 3052
rect 2700 3040 2728 3080
rect 2188 3012 2728 3040
rect 2884 3040 2912 3080
rect 2961 3077 2973 3111
rect 3007 3108 3019 3111
rect 3878 3108 3884 3120
rect 3007 3080 3884 3108
rect 3007 3077 3019 3080
rect 2961 3071 3019 3077
rect 3878 3068 3884 3080
rect 3936 3068 3942 3120
rect 3237 3043 3295 3049
rect 3237 3040 3249 3043
rect 2884 3012 3249 3040
rect 2188 3000 2194 3012
rect 3237 3009 3249 3012
rect 3283 3009 3295 3043
rect 3237 3003 3295 3009
rect 1762 2972 1768 2984
rect 1723 2944 1768 2972
rect 1762 2932 1768 2944
rect 1820 2932 1826 2984
rect 2777 2975 2835 2981
rect 2777 2941 2789 2975
rect 2823 2972 2835 2975
rect 2823 2944 2912 2972
rect 2823 2941 2835 2944
rect 2777 2935 2835 2941
rect 2222 2904 2228 2916
rect 2183 2876 2228 2904
rect 2222 2864 2228 2876
rect 2280 2864 2286 2916
rect 2884 2904 2912 2944
rect 3878 2904 3884 2916
rect 2884 2876 3884 2904
rect 3878 2864 3884 2876
rect 3936 2904 3942 2916
rect 3973 2907 4031 2913
rect 3973 2904 3985 2907
rect 3936 2876 3985 2904
rect 3936 2864 3942 2876
rect 3973 2873 3985 2876
rect 4019 2873 4031 2907
rect 3973 2867 4031 2873
rect 2240 2836 2268 2864
rect 3605 2839 3663 2845
rect 3605 2836 3617 2839
rect 2240 2808 3617 2836
rect 3605 2805 3617 2808
rect 3651 2805 3663 2839
rect 3605 2799 3663 2805
rect 1104 2746 21896 2768
rect 1104 2694 7912 2746
rect 7964 2694 7976 2746
rect 8028 2694 8040 2746
rect 8092 2694 8104 2746
rect 8156 2694 14843 2746
rect 14895 2694 14907 2746
rect 14959 2694 14971 2746
rect 15023 2694 15035 2746
rect 15087 2694 21896 2746
rect 1104 2672 21896 2694
rect 2317 2635 2375 2641
rect 2317 2601 2329 2635
rect 2363 2632 2375 2635
rect 4338 2632 4344 2644
rect 2363 2604 4344 2632
rect 2363 2601 2375 2604
rect 2317 2595 2375 2601
rect 4338 2592 4344 2604
rect 4396 2592 4402 2644
rect 2961 2567 3019 2573
rect 2961 2533 2973 2567
rect 3007 2564 3019 2567
rect 5442 2564 5448 2576
rect 3007 2536 5448 2564
rect 3007 2533 3019 2536
rect 2961 2527 3019 2533
rect 5442 2524 5448 2536
rect 5500 2524 5506 2576
rect 12250 2564 12256 2576
rect 12211 2536 12256 2564
rect 12250 2524 12256 2536
rect 12308 2564 12314 2576
rect 12621 2567 12679 2573
rect 12621 2564 12633 2567
rect 12308 2536 12633 2564
rect 12308 2524 12314 2536
rect 12621 2533 12633 2536
rect 12667 2533 12679 2567
rect 12621 2527 12679 2533
rect 1670 2496 1676 2508
rect 1631 2468 1676 2496
rect 1670 2456 1676 2468
rect 1728 2456 1734 2508
rect 2130 2456 2136 2508
rect 2188 2496 2194 2508
rect 2225 2499 2283 2505
rect 2225 2496 2237 2499
rect 2188 2468 2237 2496
rect 2188 2456 2194 2468
rect 2225 2465 2237 2468
rect 2271 2465 2283 2499
rect 2774 2496 2780 2508
rect 2735 2468 2780 2496
rect 2225 2459 2283 2465
rect 2774 2456 2780 2468
rect 2832 2496 2838 2508
rect 3881 2499 3939 2505
rect 3881 2496 3893 2499
rect 2832 2468 3893 2496
rect 2832 2456 2838 2468
rect 3881 2465 3893 2468
rect 3927 2465 3939 2499
rect 3881 2459 3939 2465
rect 1688 2428 1716 2456
rect 3237 2431 3295 2437
rect 3237 2428 3249 2431
rect 1688 2400 3249 2428
rect 3237 2397 3249 2400
rect 3283 2397 3295 2431
rect 3237 2391 3295 2397
rect 1857 2363 1915 2369
rect 1857 2329 1869 2363
rect 1903 2360 1915 2363
rect 3970 2360 3976 2372
rect 1903 2332 3976 2360
rect 1903 2329 1915 2332
rect 1857 2323 1915 2329
rect 3970 2320 3976 2332
rect 4028 2320 4034 2372
rect 11698 2320 11704 2372
rect 11756 2360 11762 2372
rect 12069 2363 12127 2369
rect 12069 2360 12081 2363
rect 11756 2332 12081 2360
rect 11756 2320 11762 2332
rect 12069 2329 12081 2332
rect 12115 2329 12127 2363
rect 12069 2323 12127 2329
rect 1104 2202 21896 2224
rect 1104 2150 4447 2202
rect 4499 2150 4511 2202
rect 4563 2150 4575 2202
rect 4627 2150 4639 2202
rect 4691 2150 11378 2202
rect 11430 2150 11442 2202
rect 11494 2150 11506 2202
rect 11558 2150 11570 2202
rect 11622 2150 18308 2202
rect 18360 2150 18372 2202
rect 18424 2150 18436 2202
rect 18488 2150 18500 2202
rect 18552 2150 21896 2202
rect 1104 2128 21896 2150
<< via1 >>
rect 3976 20816 4028 20868
rect 7840 20816 7892 20868
rect 9404 20816 9456 20868
rect 10140 20816 10192 20868
rect 4068 20748 4120 20800
rect 7288 20748 7340 20800
rect 8944 20748 8996 20800
rect 10048 20748 10100 20800
rect 4447 20646 4499 20698
rect 4511 20646 4563 20698
rect 4575 20646 4627 20698
rect 4639 20646 4691 20698
rect 11378 20646 11430 20698
rect 11442 20646 11494 20698
rect 11506 20646 11558 20698
rect 11570 20646 11622 20698
rect 18308 20646 18360 20698
rect 18372 20646 18424 20698
rect 18436 20646 18488 20698
rect 18500 20646 18552 20698
rect 7564 20544 7616 20596
rect 7656 20544 7708 20596
rect 2780 20476 2832 20528
rect 7104 20476 7156 20528
rect 7288 20519 7340 20528
rect 7288 20485 7297 20519
rect 7297 20485 7331 20519
rect 7331 20485 7340 20519
rect 7288 20476 7340 20485
rect 7840 20519 7892 20528
rect 7840 20485 7849 20519
rect 7849 20485 7883 20519
rect 7883 20485 7892 20519
rect 7840 20476 7892 20485
rect 8484 20544 8536 20596
rect 14464 20544 14516 20596
rect 19524 20544 19576 20596
rect 1584 20408 1636 20460
rect 204 20340 256 20392
rect 1308 20340 1360 20392
rect 4160 20408 4212 20460
rect 3608 20340 3660 20392
rect 4252 20340 4304 20392
rect 6092 20451 6144 20460
rect 6092 20417 6101 20451
rect 6101 20417 6135 20451
rect 6135 20417 6144 20451
rect 6092 20408 6144 20417
rect 6552 20408 6604 20460
rect 9680 20408 9732 20460
rect 4988 20340 5040 20392
rect 6736 20340 6788 20392
rect 7656 20340 7708 20392
rect 664 20272 716 20324
rect 2228 20315 2280 20324
rect 2228 20281 2237 20315
rect 2237 20281 2271 20315
rect 2271 20281 2280 20315
rect 2228 20272 2280 20281
rect 1124 20204 1176 20256
rect 3700 20272 3752 20324
rect 6828 20315 6880 20324
rect 6828 20281 6837 20315
rect 6837 20281 6871 20315
rect 6871 20281 6880 20315
rect 6828 20272 6880 20281
rect 7012 20272 7064 20324
rect 3424 20204 3476 20256
rect 4068 20247 4120 20256
rect 4068 20213 4077 20247
rect 4077 20213 4111 20247
rect 4111 20213 4120 20247
rect 4068 20204 4120 20213
rect 4620 20204 4672 20256
rect 5080 20247 5132 20256
rect 5080 20213 5089 20247
rect 5089 20213 5123 20247
rect 5123 20213 5132 20247
rect 5080 20204 5132 20213
rect 5448 20247 5500 20256
rect 5448 20213 5457 20247
rect 5457 20213 5491 20247
rect 5491 20213 5500 20247
rect 5448 20204 5500 20213
rect 5816 20247 5868 20256
rect 5816 20213 5825 20247
rect 5825 20213 5859 20247
rect 5859 20213 5868 20247
rect 5816 20204 5868 20213
rect 6552 20204 6604 20256
rect 9312 20272 9364 20324
rect 8484 20204 8536 20256
rect 9680 20204 9732 20256
rect 11336 20476 11388 20528
rect 11612 20476 11664 20528
rect 13084 20519 13136 20528
rect 13084 20485 13093 20519
rect 13093 20485 13127 20519
rect 13127 20485 13136 20519
rect 13084 20476 13136 20485
rect 13544 20476 13596 20528
rect 14004 20476 14056 20528
rect 17684 20519 17736 20528
rect 9956 20451 10008 20460
rect 9956 20417 9965 20451
rect 9965 20417 9999 20451
rect 9999 20417 10008 20451
rect 9956 20408 10008 20417
rect 14924 20408 14976 20460
rect 16580 20408 16632 20460
rect 17684 20485 17693 20519
rect 17693 20485 17727 20519
rect 17727 20485 17736 20519
rect 17684 20476 17736 20485
rect 18144 20476 18196 20528
rect 18604 20476 18656 20528
rect 19064 20476 19116 20528
rect 21364 20408 21416 20460
rect 10048 20340 10100 20392
rect 10968 20340 11020 20392
rect 10140 20272 10192 20324
rect 12808 20340 12860 20392
rect 10048 20204 10100 20256
rect 10416 20247 10468 20256
rect 10416 20213 10425 20247
rect 10425 20213 10459 20247
rect 10459 20213 10468 20247
rect 10416 20204 10468 20213
rect 10508 20204 10560 20256
rect 12256 20204 12308 20256
rect 14280 20340 14332 20392
rect 13268 20315 13320 20324
rect 13268 20281 13277 20315
rect 13277 20281 13311 20315
rect 13311 20281 13320 20315
rect 13268 20272 13320 20281
rect 13820 20315 13872 20324
rect 13820 20281 13829 20315
rect 13829 20281 13863 20315
rect 13863 20281 13872 20315
rect 13820 20272 13872 20281
rect 13912 20272 13964 20324
rect 15568 20315 15620 20324
rect 15568 20281 15577 20315
rect 15577 20281 15611 20315
rect 15611 20281 15620 20315
rect 15568 20272 15620 20281
rect 16120 20315 16172 20324
rect 16120 20281 16129 20315
rect 16129 20281 16163 20315
rect 16163 20281 16172 20315
rect 16120 20272 16172 20281
rect 13636 20204 13688 20256
rect 18052 20272 18104 20324
rect 18604 20272 18656 20324
rect 18972 20315 19024 20324
rect 18972 20281 18981 20315
rect 18981 20281 19015 20315
rect 19015 20281 19024 20315
rect 18972 20272 19024 20281
rect 19340 20340 19392 20392
rect 22744 20340 22796 20392
rect 21824 20272 21876 20324
rect 18880 20204 18932 20256
rect 19248 20204 19300 20256
rect 21180 20247 21232 20256
rect 21180 20213 21189 20247
rect 21189 20213 21223 20247
rect 21223 20213 21232 20247
rect 21180 20204 21232 20213
rect 7912 20102 7964 20154
rect 7976 20102 8028 20154
rect 8040 20102 8092 20154
rect 8104 20102 8156 20154
rect 14843 20102 14895 20154
rect 14907 20102 14959 20154
rect 14971 20102 15023 20154
rect 15035 20102 15087 20154
rect 4068 20000 4120 20052
rect 5448 20000 5500 20052
rect 6000 20000 6052 20052
rect 7288 20000 7340 20052
rect 8392 20043 8444 20052
rect 8392 20009 8401 20043
rect 8401 20009 8435 20043
rect 8435 20009 8444 20043
rect 8392 20000 8444 20009
rect 10416 20000 10468 20052
rect 10508 20000 10560 20052
rect 12808 20043 12860 20052
rect 12808 20009 12817 20043
rect 12817 20009 12851 20043
rect 12851 20009 12860 20043
rect 12808 20000 12860 20009
rect 13912 20000 13964 20052
rect 16120 20000 16172 20052
rect 1308 19932 1360 19984
rect 5080 19932 5132 19984
rect 6092 19932 6144 19984
rect 7564 19932 7616 19984
rect 10876 19932 10928 19984
rect 11060 19932 11112 19984
rect 15384 19975 15436 19984
rect 15384 19941 15393 19975
rect 15393 19941 15427 19975
rect 15427 19941 15436 19975
rect 15384 19932 15436 19941
rect 15844 19932 15896 19984
rect 16304 19932 16356 19984
rect 16764 19932 16816 19984
rect 17224 20000 17276 20052
rect 18972 20000 19024 20052
rect 19156 19932 19208 19984
rect 19984 19975 20036 19984
rect 19984 19941 19993 19975
rect 19993 19941 20027 19975
rect 20027 19941 20036 19975
rect 19984 19932 20036 19941
rect 20444 19932 20496 19984
rect 20904 19932 20956 19984
rect 2044 19864 2096 19916
rect 2504 19864 2556 19916
rect 6368 19864 6420 19916
rect 6828 19864 6880 19916
rect 1584 19771 1636 19780
rect 1584 19737 1593 19771
rect 1593 19737 1627 19771
rect 1627 19737 1636 19771
rect 1584 19728 1636 19737
rect 3148 19728 3200 19780
rect 5356 19728 5408 19780
rect 5540 19771 5592 19780
rect 5540 19737 5549 19771
rect 5549 19737 5583 19771
rect 5583 19737 5592 19771
rect 5540 19728 5592 19737
rect 5172 19660 5224 19712
rect 8668 19864 8720 19916
rect 9588 19864 9640 19916
rect 10692 19864 10744 19916
rect 11336 19864 11388 19916
rect 12348 19907 12400 19916
rect 8852 19796 8904 19848
rect 8760 19728 8812 19780
rect 7288 19660 7340 19712
rect 7656 19703 7708 19712
rect 7656 19669 7665 19703
rect 7665 19669 7699 19703
rect 7699 19669 7708 19703
rect 7656 19660 7708 19669
rect 7748 19660 7800 19712
rect 8208 19660 8260 19712
rect 11796 19660 11848 19712
rect 12348 19873 12357 19907
rect 12357 19873 12391 19907
rect 12391 19873 12400 19907
rect 12348 19864 12400 19873
rect 14188 19864 14240 19916
rect 15200 19864 15252 19916
rect 16120 19907 16172 19916
rect 16120 19873 16129 19907
rect 16129 19873 16163 19907
rect 16163 19873 16172 19907
rect 16120 19864 16172 19873
rect 16672 19907 16724 19916
rect 16672 19873 16681 19907
rect 16681 19873 16715 19907
rect 16715 19873 16724 19907
rect 16672 19864 16724 19873
rect 17224 19907 17276 19916
rect 17224 19873 17233 19907
rect 17233 19873 17267 19907
rect 17267 19873 17276 19907
rect 17224 19864 17276 19873
rect 17776 19907 17828 19916
rect 17776 19873 17785 19907
rect 17785 19873 17819 19907
rect 17819 19873 17828 19907
rect 17776 19864 17828 19873
rect 18144 19907 18196 19916
rect 18144 19873 18153 19907
rect 18153 19873 18187 19907
rect 18187 19873 18196 19907
rect 18144 19864 18196 19873
rect 18696 19864 18748 19916
rect 19708 19864 19760 19916
rect 14004 19796 14056 19848
rect 19432 19796 19484 19848
rect 19984 19796 20036 19848
rect 13636 19771 13688 19780
rect 13176 19660 13228 19712
rect 13636 19737 13645 19771
rect 13645 19737 13679 19771
rect 13679 19737 13688 19771
rect 13636 19728 13688 19737
rect 19248 19728 19300 19780
rect 19800 19728 19852 19780
rect 15292 19660 15344 19712
rect 18972 19660 19024 19712
rect 4447 19558 4499 19610
rect 4511 19558 4563 19610
rect 4575 19558 4627 19610
rect 4639 19558 4691 19610
rect 11378 19558 11430 19610
rect 11442 19558 11494 19610
rect 11506 19558 11558 19610
rect 11570 19558 11622 19610
rect 18308 19558 18360 19610
rect 18372 19558 18424 19610
rect 18436 19558 18488 19610
rect 18500 19558 18552 19610
rect 3424 19456 3476 19508
rect 4252 19499 4304 19508
rect 2228 19388 2280 19440
rect 4252 19465 4261 19499
rect 4261 19465 4295 19499
rect 4295 19465 4304 19499
rect 4252 19456 4304 19465
rect 5172 19456 5224 19508
rect 6460 19456 6512 19508
rect 6828 19456 6880 19508
rect 7104 19456 7156 19508
rect 1584 19295 1636 19304
rect 1584 19261 1593 19295
rect 1593 19261 1627 19295
rect 1627 19261 1636 19295
rect 1584 19252 1636 19261
rect 2780 19252 2832 19304
rect 4068 19295 4120 19304
rect 4068 19261 4077 19295
rect 4077 19261 4111 19295
rect 4111 19261 4120 19295
rect 4068 19252 4120 19261
rect 6644 19388 6696 19440
rect 10876 19456 10928 19508
rect 13084 19456 13136 19508
rect 13268 19456 13320 19508
rect 13820 19499 13872 19508
rect 13820 19465 13829 19499
rect 13829 19465 13863 19499
rect 13863 19465 13872 19499
rect 13820 19456 13872 19465
rect 14280 19499 14332 19508
rect 14280 19465 14289 19499
rect 14289 19465 14323 19499
rect 14323 19465 14332 19499
rect 14280 19456 14332 19465
rect 16120 19456 16172 19508
rect 17224 19456 17276 19508
rect 17776 19499 17828 19508
rect 17776 19465 17785 19499
rect 17785 19465 17819 19499
rect 17819 19465 17828 19499
rect 17776 19456 17828 19465
rect 18052 19499 18104 19508
rect 18052 19465 18061 19499
rect 18061 19465 18095 19499
rect 18095 19465 18104 19499
rect 18052 19456 18104 19465
rect 18604 19456 18656 19508
rect 19432 19499 19484 19508
rect 19432 19465 19441 19499
rect 19441 19465 19475 19499
rect 19475 19465 19484 19499
rect 19432 19456 19484 19465
rect 11152 19388 11204 19440
rect 11336 19388 11388 19440
rect 12532 19388 12584 19440
rect 2228 19184 2280 19236
rect 2412 19116 2464 19168
rect 3148 19116 3200 19168
rect 5540 19252 5592 19304
rect 6276 19252 6328 19304
rect 6368 19252 6420 19304
rect 4436 19116 4488 19168
rect 7288 19116 7340 19168
rect 7472 19159 7524 19168
rect 7472 19125 7481 19159
rect 7481 19125 7515 19159
rect 7515 19125 7524 19159
rect 7472 19116 7524 19125
rect 8760 19252 8812 19304
rect 9220 19252 9272 19304
rect 9956 19295 10008 19304
rect 9956 19261 9990 19295
rect 9990 19261 10008 19295
rect 9956 19252 10008 19261
rect 10968 19252 11020 19304
rect 12072 19295 12124 19304
rect 12072 19261 12081 19295
rect 12081 19261 12115 19295
rect 12115 19261 12124 19295
rect 12072 19252 12124 19261
rect 12532 19295 12584 19304
rect 12532 19261 12541 19295
rect 12541 19261 12575 19295
rect 12575 19261 12584 19295
rect 12532 19252 12584 19261
rect 12808 19388 12860 19440
rect 13452 19388 13504 19440
rect 16672 19388 16724 19440
rect 15568 19320 15620 19372
rect 14004 19295 14056 19304
rect 8116 19184 8168 19236
rect 10416 19184 10468 19236
rect 9312 19116 9364 19168
rect 9680 19116 9732 19168
rect 11060 19159 11112 19168
rect 11060 19125 11069 19159
rect 11069 19125 11103 19159
rect 11103 19125 11112 19159
rect 11060 19116 11112 19125
rect 13360 19184 13412 19236
rect 14004 19261 14013 19295
rect 14013 19261 14047 19295
rect 14047 19261 14056 19295
rect 14004 19252 14056 19261
rect 15292 19295 15344 19304
rect 13268 19116 13320 19168
rect 15292 19261 15301 19295
rect 15301 19261 15335 19295
rect 15335 19261 15344 19295
rect 15292 19252 15344 19261
rect 16488 19295 16540 19304
rect 15200 19116 15252 19168
rect 16488 19261 16497 19295
rect 16497 19261 16531 19295
rect 16531 19261 16540 19295
rect 16488 19252 16540 19261
rect 17316 19295 17368 19304
rect 17316 19261 17325 19295
rect 17325 19261 17359 19295
rect 17359 19261 17368 19295
rect 17316 19252 17368 19261
rect 17868 19252 17920 19304
rect 17960 19252 18012 19304
rect 18328 19252 18380 19304
rect 18972 19295 19024 19304
rect 18972 19261 18981 19295
rect 18981 19261 19015 19295
rect 19015 19261 19024 19295
rect 18972 19252 19024 19261
rect 19340 19116 19392 19168
rect 21364 19295 21416 19304
rect 21364 19261 21373 19295
rect 21373 19261 21407 19295
rect 21407 19261 21416 19295
rect 21364 19252 21416 19261
rect 22284 19252 22336 19304
rect 20720 19184 20772 19236
rect 20812 19116 20864 19168
rect 7912 19014 7964 19066
rect 7976 19014 8028 19066
rect 8040 19014 8092 19066
rect 8104 19014 8156 19066
rect 14843 19014 14895 19066
rect 14907 19014 14959 19066
rect 14971 19014 15023 19066
rect 15035 19014 15087 19066
rect 2872 18912 2924 18964
rect 4528 18912 4580 18964
rect 5908 18912 5960 18964
rect 6092 18912 6144 18964
rect 6736 18912 6788 18964
rect 7748 18955 7800 18964
rect 7748 18921 7757 18955
rect 7757 18921 7791 18955
rect 7791 18921 7800 18955
rect 7748 18912 7800 18921
rect 9956 18912 10008 18964
rect 1584 18819 1636 18828
rect 1584 18785 1593 18819
rect 1593 18785 1627 18819
rect 1627 18785 1636 18819
rect 1584 18776 1636 18785
rect 2136 18776 2188 18828
rect 4068 18776 4120 18828
rect 4252 18819 4304 18828
rect 4252 18785 4261 18819
rect 4261 18785 4295 18819
rect 4295 18785 4304 18819
rect 4252 18776 4304 18785
rect 6000 18844 6052 18896
rect 7104 18887 7156 18896
rect 5080 18776 5132 18828
rect 5264 18819 5316 18828
rect 5264 18785 5298 18819
rect 5298 18785 5316 18819
rect 5264 18776 5316 18785
rect 5724 18776 5776 18828
rect 7104 18853 7113 18887
rect 7113 18853 7147 18887
rect 7147 18853 7156 18887
rect 7104 18844 7156 18853
rect 7564 18844 7616 18896
rect 11152 18912 11204 18964
rect 12164 18912 12216 18964
rect 12440 18912 12492 18964
rect 13268 18912 13320 18964
rect 14004 18955 14056 18964
rect 14004 18921 14013 18955
rect 14013 18921 14047 18955
rect 14047 18921 14056 18955
rect 14004 18912 14056 18921
rect 14280 18912 14332 18964
rect 17868 18955 17920 18964
rect 17868 18921 17877 18955
rect 17877 18921 17911 18955
rect 17911 18921 17920 18955
rect 17868 18912 17920 18921
rect 18328 18955 18380 18964
rect 18328 18921 18337 18955
rect 18337 18921 18371 18955
rect 18371 18921 18380 18955
rect 18328 18912 18380 18921
rect 21364 18955 21416 18964
rect 21364 18921 21373 18955
rect 21373 18921 21407 18955
rect 21407 18921 21416 18955
rect 21364 18912 21416 18921
rect 10324 18844 10376 18896
rect 6644 18819 6696 18828
rect 6644 18785 6653 18819
rect 6653 18785 6687 18819
rect 6687 18785 6696 18819
rect 6644 18776 6696 18785
rect 2320 18640 2372 18692
rect 2688 18615 2740 18624
rect 2688 18581 2697 18615
rect 2697 18581 2731 18615
rect 2731 18581 2740 18615
rect 2688 18572 2740 18581
rect 2964 18572 3016 18624
rect 6184 18708 6236 18760
rect 7472 18708 7524 18760
rect 9312 18776 9364 18828
rect 10140 18776 10192 18828
rect 10600 18776 10652 18828
rect 13544 18844 13596 18896
rect 12164 18819 12216 18828
rect 12164 18785 12173 18819
rect 12173 18785 12207 18819
rect 12207 18785 12216 18819
rect 12164 18776 12216 18785
rect 12992 18819 13044 18828
rect 12992 18785 13001 18819
rect 13001 18785 13035 18819
rect 13035 18785 13044 18819
rect 12992 18776 13044 18785
rect 13820 18819 13872 18828
rect 13820 18785 13829 18819
rect 13829 18785 13863 18819
rect 13863 18785 13872 18819
rect 13820 18776 13872 18785
rect 8668 18708 8720 18760
rect 8852 18640 8904 18692
rect 8024 18572 8076 18624
rect 9220 18572 9272 18624
rect 11336 18708 11388 18760
rect 11980 18751 12032 18760
rect 11980 18717 11989 18751
rect 11989 18717 12023 18751
rect 12023 18717 12032 18751
rect 11980 18708 12032 18717
rect 12716 18708 12768 18760
rect 14372 18751 14424 18760
rect 14372 18717 14381 18751
rect 14381 18717 14415 18751
rect 14415 18717 14424 18751
rect 14372 18708 14424 18717
rect 16304 18844 16356 18896
rect 16396 18776 16448 18828
rect 16764 18776 16816 18828
rect 17684 18819 17736 18828
rect 17684 18785 17693 18819
rect 17693 18785 17727 18819
rect 17727 18785 17736 18819
rect 17684 18776 17736 18785
rect 18604 18776 18656 18828
rect 18788 18819 18840 18828
rect 18788 18785 18797 18819
rect 18797 18785 18831 18819
rect 18831 18785 18840 18819
rect 18788 18776 18840 18785
rect 17500 18708 17552 18760
rect 21180 18708 21232 18760
rect 12256 18640 12308 18692
rect 14740 18640 14792 18692
rect 18144 18640 18196 18692
rect 10968 18615 11020 18624
rect 10968 18581 10977 18615
rect 10977 18581 11011 18615
rect 11011 18581 11020 18615
rect 10968 18572 11020 18581
rect 11704 18572 11756 18624
rect 13360 18572 13412 18624
rect 15844 18572 15896 18624
rect 16028 18615 16080 18624
rect 16028 18581 16037 18615
rect 16037 18581 16071 18615
rect 16071 18581 16080 18615
rect 16028 18572 16080 18581
rect 19156 18615 19208 18624
rect 19156 18581 19165 18615
rect 19165 18581 19199 18615
rect 19199 18581 19208 18615
rect 19156 18572 19208 18581
rect 20536 18572 20588 18624
rect 4447 18470 4499 18522
rect 4511 18470 4563 18522
rect 4575 18470 4627 18522
rect 4639 18470 4691 18522
rect 11378 18470 11430 18522
rect 11442 18470 11494 18522
rect 11506 18470 11558 18522
rect 11570 18470 11622 18522
rect 18308 18470 18360 18522
rect 18372 18470 18424 18522
rect 18436 18470 18488 18522
rect 18500 18470 18552 18522
rect 1676 18411 1728 18420
rect 1676 18377 1685 18411
rect 1685 18377 1719 18411
rect 1719 18377 1728 18411
rect 1676 18368 1728 18377
rect 3056 18368 3108 18420
rect 4896 18368 4948 18420
rect 6368 18368 6420 18420
rect 6644 18368 6696 18420
rect 8852 18411 8904 18420
rect 8852 18377 8861 18411
rect 8861 18377 8895 18411
rect 8895 18377 8904 18411
rect 8852 18368 8904 18377
rect 4068 18300 4120 18352
rect 4804 18232 4856 18284
rect 5264 18232 5316 18284
rect 5448 18232 5500 18284
rect 6828 18232 6880 18284
rect 7380 18275 7432 18284
rect 7380 18241 7389 18275
rect 7389 18241 7423 18275
rect 7423 18241 7432 18275
rect 7380 18232 7432 18241
rect 11704 18368 11756 18420
rect 12716 18368 12768 18420
rect 13820 18368 13872 18420
rect 17316 18411 17368 18420
rect 17316 18377 17325 18411
rect 17325 18377 17359 18411
rect 17359 18377 17368 18411
rect 17316 18368 17368 18377
rect 17960 18411 18012 18420
rect 17960 18377 17969 18411
rect 17969 18377 18003 18411
rect 18003 18377 18012 18411
rect 17960 18368 18012 18377
rect 9772 18275 9824 18284
rect 2320 18207 2372 18216
rect 2320 18173 2329 18207
rect 2329 18173 2363 18207
rect 2363 18173 2372 18207
rect 2320 18164 2372 18173
rect 3148 18207 3200 18216
rect 3148 18173 3182 18207
rect 3182 18173 3200 18207
rect 2504 18096 2556 18148
rect 3148 18164 3200 18173
rect 3608 18164 3660 18216
rect 9772 18241 9781 18275
rect 9781 18241 9815 18275
rect 9815 18241 9824 18275
rect 9772 18232 9824 18241
rect 11060 18232 11112 18284
rect 12808 18300 12860 18352
rect 17500 18300 17552 18352
rect 18052 18300 18104 18352
rect 12716 18232 12768 18284
rect 8024 18207 8076 18216
rect 8024 18173 8033 18207
rect 8033 18173 8067 18207
rect 8067 18173 8076 18207
rect 8024 18164 8076 18173
rect 9680 18207 9732 18216
rect 3884 18096 3936 18148
rect 1952 18028 2004 18080
rect 4896 18096 4948 18148
rect 4160 18028 4212 18080
rect 4988 18028 5040 18080
rect 5264 18071 5316 18080
rect 5264 18037 5273 18071
rect 5273 18037 5307 18071
rect 5307 18037 5316 18071
rect 5264 18028 5316 18037
rect 5540 18028 5592 18080
rect 6276 18028 6328 18080
rect 7196 18071 7248 18080
rect 7196 18037 7205 18071
rect 7205 18037 7239 18071
rect 7239 18037 7248 18071
rect 7196 18028 7248 18037
rect 7288 18071 7340 18080
rect 7288 18037 7297 18071
rect 7297 18037 7331 18071
rect 7331 18037 7340 18071
rect 9680 18173 9689 18207
rect 9689 18173 9723 18207
rect 9723 18173 9732 18207
rect 9680 18164 9732 18173
rect 9864 18164 9916 18216
rect 10784 18164 10836 18216
rect 11704 18164 11756 18216
rect 12900 18164 12952 18216
rect 14004 18164 14056 18216
rect 16028 18232 16080 18284
rect 16672 18232 16724 18284
rect 15844 18164 15896 18216
rect 17132 18207 17184 18216
rect 17132 18173 17141 18207
rect 17141 18173 17175 18207
rect 17175 18173 17184 18207
rect 17132 18164 17184 18173
rect 18144 18164 18196 18216
rect 7288 18028 7340 18037
rect 10324 18071 10376 18080
rect 10324 18037 10333 18071
rect 10333 18037 10367 18071
rect 10367 18037 10376 18071
rect 10324 18028 10376 18037
rect 10784 18071 10836 18080
rect 10784 18037 10793 18071
rect 10793 18037 10827 18071
rect 10827 18037 10836 18071
rect 10784 18028 10836 18037
rect 11060 18028 11112 18080
rect 12440 18028 12492 18080
rect 13268 18071 13320 18080
rect 13268 18037 13277 18071
rect 13277 18037 13311 18071
rect 13311 18037 13320 18071
rect 13268 18028 13320 18037
rect 13360 18071 13412 18080
rect 13360 18037 13369 18071
rect 13369 18037 13403 18071
rect 13403 18037 13412 18071
rect 16764 18096 16816 18148
rect 13360 18028 13412 18037
rect 16212 18071 16264 18080
rect 16212 18037 16221 18071
rect 16221 18037 16255 18071
rect 16255 18037 16264 18071
rect 16212 18028 16264 18037
rect 7912 17926 7964 17978
rect 7976 17926 8028 17978
rect 8040 17926 8092 17978
rect 8104 17926 8156 17978
rect 14843 17926 14895 17978
rect 14907 17926 14959 17978
rect 14971 17926 15023 17978
rect 15035 17926 15087 17978
rect 4804 17867 4856 17876
rect 4804 17833 4813 17867
rect 4813 17833 4847 17867
rect 4847 17833 4856 17867
rect 4804 17824 4856 17833
rect 4896 17824 4948 17876
rect 7564 17824 7616 17876
rect 10324 17824 10376 17876
rect 10508 17824 10560 17876
rect 14740 17824 14792 17876
rect 15384 17824 15436 17876
rect 16396 17824 16448 17876
rect 2688 17756 2740 17808
rect 2872 17756 2924 17808
rect 5540 17756 5592 17808
rect 5632 17756 5684 17808
rect 6000 17756 6052 17808
rect 6460 17756 6512 17808
rect 7472 17799 7524 17808
rect 3148 17731 3200 17740
rect 3148 17697 3157 17731
rect 3157 17697 3191 17731
rect 3191 17697 3200 17731
rect 3148 17688 3200 17697
rect 7472 17765 7506 17799
rect 7506 17765 7524 17799
rect 7472 17756 7524 17765
rect 9864 17688 9916 17740
rect 10140 17688 10192 17740
rect 10324 17688 10376 17740
rect 2872 17663 2924 17672
rect 2872 17629 2881 17663
rect 2881 17629 2915 17663
rect 2915 17629 2924 17663
rect 2872 17620 2924 17629
rect 4344 17620 4396 17672
rect 6184 17663 6236 17672
rect 6184 17629 6193 17663
rect 6193 17629 6227 17663
rect 6227 17629 6236 17663
rect 6184 17620 6236 17629
rect 10048 17620 10100 17672
rect 11244 17688 11296 17740
rect 12808 17731 12860 17740
rect 12808 17697 12826 17731
rect 12826 17697 12860 17731
rect 13544 17731 13596 17740
rect 12808 17688 12860 17697
rect 13544 17697 13553 17731
rect 13553 17697 13587 17731
rect 13587 17697 13596 17731
rect 13544 17688 13596 17697
rect 14004 17731 14056 17740
rect 14004 17697 14013 17731
rect 14013 17697 14047 17731
rect 14047 17697 14056 17731
rect 14004 17688 14056 17697
rect 15292 17688 15344 17740
rect 15752 17688 15804 17740
rect 11336 17620 11388 17672
rect 14372 17620 14424 17672
rect 2688 17552 2740 17604
rect 2228 17527 2280 17536
rect 2228 17493 2237 17527
rect 2237 17493 2271 17527
rect 2271 17493 2280 17527
rect 2228 17484 2280 17493
rect 9036 17552 9088 17604
rect 8116 17484 8168 17536
rect 9772 17484 9824 17536
rect 10140 17484 10192 17536
rect 10508 17552 10560 17604
rect 16304 17620 16356 17672
rect 15200 17552 15252 17604
rect 16212 17552 16264 17604
rect 12716 17484 12768 17536
rect 13544 17484 13596 17536
rect 13636 17484 13688 17536
rect 14464 17484 14516 17536
rect 19892 17620 19944 17672
rect 17960 17552 18012 17604
rect 18972 17484 19024 17536
rect 4447 17382 4499 17434
rect 4511 17382 4563 17434
rect 4575 17382 4627 17434
rect 4639 17382 4691 17434
rect 11378 17382 11430 17434
rect 11442 17382 11494 17434
rect 11506 17382 11558 17434
rect 11570 17382 11622 17434
rect 18308 17382 18360 17434
rect 18372 17382 18424 17434
rect 18436 17382 18488 17434
rect 18500 17382 18552 17434
rect 2780 17280 2832 17332
rect 4344 17323 4396 17332
rect 4344 17289 4353 17323
rect 4353 17289 4387 17323
rect 4387 17289 4396 17323
rect 4344 17280 4396 17289
rect 5264 17280 5316 17332
rect 6368 17280 6420 17332
rect 7380 17280 7432 17332
rect 5448 17212 5500 17264
rect 8576 17280 8628 17332
rect 10600 17323 10652 17332
rect 9128 17212 9180 17264
rect 10600 17289 10609 17323
rect 10609 17289 10643 17323
rect 10643 17289 10652 17323
rect 10600 17280 10652 17289
rect 11704 17323 11756 17332
rect 11704 17289 11713 17323
rect 11713 17289 11747 17323
rect 11747 17289 11756 17323
rect 11704 17280 11756 17289
rect 12256 17280 12308 17332
rect 12440 17280 12492 17332
rect 12624 17280 12676 17332
rect 13176 17280 13228 17332
rect 13360 17280 13412 17332
rect 14004 17280 14056 17332
rect 16304 17280 16356 17332
rect 18144 17280 18196 17332
rect 11244 17212 11296 17264
rect 19340 17212 19392 17264
rect 4160 17144 4212 17196
rect 5632 17144 5684 17196
rect 11888 17144 11940 17196
rect 12440 17144 12492 17196
rect 12808 17144 12860 17196
rect 13084 17187 13136 17196
rect 13084 17153 13093 17187
rect 13093 17153 13127 17187
rect 13127 17153 13136 17187
rect 13084 17144 13136 17153
rect 18972 17144 19024 17196
rect 2964 17076 3016 17128
rect 4068 17119 4120 17128
rect 4068 17085 4077 17119
rect 4077 17085 4111 17119
rect 4111 17085 4120 17119
rect 4068 17076 4120 17085
rect 7748 17076 7800 17128
rect 8116 17119 8168 17128
rect 8116 17085 8134 17119
rect 8134 17085 8168 17119
rect 8116 17076 8168 17085
rect 9220 17119 9272 17128
rect 9220 17085 9229 17119
rect 9229 17085 9263 17119
rect 9263 17085 9272 17119
rect 9220 17076 9272 17085
rect 1584 17051 1636 17060
rect 1584 17017 1593 17051
rect 1593 17017 1627 17051
rect 1627 17017 1636 17051
rect 1584 17008 1636 17017
rect 1768 17051 1820 17060
rect 1768 17017 1777 17051
rect 1777 17017 1811 17051
rect 1811 17017 1820 17051
rect 1768 17008 1820 17017
rect 4160 17008 4212 17060
rect 6184 17008 6236 17060
rect 10048 17008 10100 17060
rect 2872 16940 2924 16992
rect 3332 16940 3384 16992
rect 5632 16940 5684 16992
rect 6368 16940 6420 16992
rect 9680 16940 9732 16992
rect 11152 17076 11204 17128
rect 14372 17076 14424 17128
rect 15384 17076 15436 17128
rect 17776 17076 17828 17128
rect 19892 17119 19944 17128
rect 19892 17085 19901 17119
rect 19901 17085 19935 17119
rect 19935 17085 19944 17119
rect 19892 17076 19944 17085
rect 10416 17008 10468 17060
rect 11888 16940 11940 16992
rect 12348 16983 12400 16992
rect 12348 16949 12357 16983
rect 12357 16949 12391 16983
rect 12391 16949 12400 16983
rect 12348 16940 12400 16949
rect 13912 17008 13964 17060
rect 15200 17008 15252 17060
rect 15292 17008 15344 17060
rect 15476 17008 15528 17060
rect 13452 16940 13504 16992
rect 17316 16983 17368 16992
rect 17316 16949 17325 16983
rect 17325 16949 17359 16983
rect 17359 16949 17368 16983
rect 17316 16940 17368 16949
rect 17960 17008 18012 17060
rect 19156 17008 19208 17060
rect 18052 16940 18104 16992
rect 7912 16838 7964 16890
rect 7976 16838 8028 16890
rect 8040 16838 8092 16890
rect 8104 16838 8156 16890
rect 14843 16838 14895 16890
rect 14907 16838 14959 16890
rect 14971 16838 15023 16890
rect 15035 16838 15087 16890
rect 1768 16736 1820 16788
rect 2504 16736 2556 16788
rect 3148 16779 3200 16788
rect 3148 16745 3157 16779
rect 3157 16745 3191 16779
rect 3191 16745 3200 16779
rect 3148 16736 3200 16745
rect 4252 16779 4304 16788
rect 4252 16745 4261 16779
rect 4261 16745 4295 16779
rect 4295 16745 4304 16779
rect 4252 16736 4304 16745
rect 4896 16736 4948 16788
rect 1584 16643 1636 16652
rect 1584 16609 1593 16643
rect 1593 16609 1627 16643
rect 1627 16609 1636 16643
rect 1584 16600 1636 16609
rect 1768 16643 1820 16652
rect 1768 16609 1777 16643
rect 1777 16609 1811 16643
rect 1811 16609 1820 16643
rect 1768 16600 1820 16609
rect 3056 16668 3108 16720
rect 5540 16668 5592 16720
rect 3516 16600 3568 16652
rect 4988 16600 5040 16652
rect 5172 16643 5224 16652
rect 5172 16609 5181 16643
rect 5181 16609 5215 16643
rect 5215 16609 5224 16643
rect 5172 16600 5224 16609
rect 5908 16736 5960 16788
rect 7196 16779 7248 16788
rect 7196 16745 7205 16779
rect 7205 16745 7239 16779
rect 7239 16745 7248 16779
rect 7196 16736 7248 16745
rect 7288 16736 7340 16788
rect 7748 16736 7800 16788
rect 9680 16779 9732 16788
rect 9680 16745 9689 16779
rect 9689 16745 9723 16779
rect 9723 16745 9732 16779
rect 9680 16736 9732 16745
rect 9772 16779 9824 16788
rect 9772 16745 9781 16779
rect 9781 16745 9815 16779
rect 9815 16745 9824 16779
rect 9772 16736 9824 16745
rect 5264 16575 5316 16584
rect 5264 16541 5273 16575
rect 5273 16541 5307 16575
rect 5307 16541 5316 16575
rect 5264 16532 5316 16541
rect 5356 16532 5408 16584
rect 6460 16600 6512 16652
rect 6644 16600 6696 16652
rect 2780 16464 2832 16516
rect 7012 16464 7064 16516
rect 8300 16600 8352 16652
rect 8668 16643 8720 16652
rect 8668 16609 8677 16643
rect 8677 16609 8711 16643
rect 8711 16609 8720 16643
rect 8668 16600 8720 16609
rect 10232 16668 10284 16720
rect 8208 16532 8260 16584
rect 10416 16600 10468 16652
rect 10692 16600 10744 16652
rect 11244 16668 11296 16720
rect 13268 16736 13320 16788
rect 13912 16779 13964 16788
rect 13912 16745 13921 16779
rect 13921 16745 13955 16779
rect 13955 16745 13964 16779
rect 13912 16736 13964 16745
rect 15752 16779 15804 16788
rect 15752 16745 15761 16779
rect 15761 16745 15795 16779
rect 15795 16745 15804 16779
rect 15752 16736 15804 16745
rect 19156 16779 19208 16788
rect 13176 16643 13228 16652
rect 13176 16609 13185 16643
rect 13185 16609 13219 16643
rect 13219 16609 13228 16643
rect 13176 16600 13228 16609
rect 10600 16532 10652 16584
rect 12808 16532 12860 16584
rect 13360 16600 13412 16652
rect 15936 16600 15988 16652
rect 17224 16668 17276 16720
rect 19156 16745 19165 16779
rect 19165 16745 19199 16779
rect 19199 16745 19208 16779
rect 19156 16736 19208 16745
rect 18144 16668 18196 16720
rect 14464 16532 14516 16584
rect 15200 16575 15252 16584
rect 15200 16541 15209 16575
rect 15209 16541 15243 16575
rect 15243 16541 15252 16575
rect 15200 16532 15252 16541
rect 15292 16575 15344 16584
rect 15292 16541 15301 16575
rect 15301 16541 15335 16575
rect 15335 16541 15344 16575
rect 15292 16532 15344 16541
rect 17776 16575 17828 16584
rect 11980 16464 12032 16516
rect 4160 16396 4212 16448
rect 6184 16439 6236 16448
rect 6184 16405 6193 16439
rect 6193 16405 6227 16439
rect 6227 16405 6236 16439
rect 6184 16396 6236 16405
rect 10324 16439 10376 16448
rect 10324 16405 10333 16439
rect 10333 16405 10367 16439
rect 10367 16405 10376 16439
rect 10324 16396 10376 16405
rect 11888 16396 11940 16448
rect 12808 16396 12860 16448
rect 15384 16396 15436 16448
rect 16764 16396 16816 16448
rect 17776 16541 17785 16575
rect 17785 16541 17819 16575
rect 17819 16541 17828 16575
rect 17776 16532 17828 16541
rect 17592 16396 17644 16448
rect 19892 16396 19944 16448
rect 4447 16294 4499 16346
rect 4511 16294 4563 16346
rect 4575 16294 4627 16346
rect 4639 16294 4691 16346
rect 11378 16294 11430 16346
rect 11442 16294 11494 16346
rect 11506 16294 11558 16346
rect 11570 16294 11622 16346
rect 18308 16294 18360 16346
rect 18372 16294 18424 16346
rect 18436 16294 18488 16346
rect 18500 16294 18552 16346
rect 1768 16192 1820 16244
rect 2320 16192 2372 16244
rect 3056 16235 3108 16244
rect 3056 16201 3065 16235
rect 3065 16201 3099 16235
rect 3099 16201 3108 16235
rect 3056 16192 3108 16201
rect 3516 16235 3568 16244
rect 3516 16201 3525 16235
rect 3525 16201 3559 16235
rect 3559 16201 3568 16235
rect 3516 16192 3568 16201
rect 4988 16192 5040 16244
rect 6000 16235 6052 16244
rect 6000 16201 6009 16235
rect 6009 16201 6043 16235
rect 6043 16201 6052 16235
rect 6000 16192 6052 16201
rect 6552 16192 6604 16244
rect 10048 16235 10100 16244
rect 10048 16201 10057 16235
rect 10057 16201 10091 16235
rect 10091 16201 10100 16235
rect 10048 16192 10100 16201
rect 11152 16192 11204 16244
rect 12164 16192 12216 16244
rect 15200 16235 15252 16244
rect 1584 16099 1636 16108
rect 1584 16065 1593 16099
rect 1593 16065 1627 16099
rect 1627 16065 1636 16099
rect 1584 16056 1636 16065
rect 8300 16099 8352 16108
rect 2320 16031 2372 16040
rect 2320 15997 2329 16031
rect 2329 15997 2363 16031
rect 2363 15997 2372 16031
rect 2320 15988 2372 15997
rect 8300 16065 8309 16099
rect 8309 16065 8343 16099
rect 8343 16065 8352 16099
rect 8300 16056 8352 16065
rect 4160 16031 4212 16040
rect 1768 15963 1820 15972
rect 1768 15929 1777 15963
rect 1777 15929 1811 15963
rect 1811 15929 1820 15963
rect 1768 15920 1820 15929
rect 4160 15997 4169 16031
rect 4169 15997 4203 16031
rect 4203 15997 4212 16031
rect 4160 15988 4212 15997
rect 4620 16031 4672 16040
rect 4620 15997 4629 16031
rect 4629 15997 4663 16031
rect 4663 15997 4672 16031
rect 4620 15988 4672 15997
rect 5264 15988 5316 16040
rect 6828 16031 6880 16040
rect 6828 15997 6837 16031
rect 6837 15997 6871 16031
rect 6871 15997 6880 16031
rect 6828 15988 6880 15997
rect 7104 15988 7156 16040
rect 10876 16056 10928 16108
rect 11244 16056 11296 16108
rect 12716 16056 12768 16108
rect 5356 15920 5408 15972
rect 8208 15920 8260 15972
rect 10416 15988 10468 16040
rect 11704 15988 11756 16040
rect 12348 15988 12400 16040
rect 15200 16201 15209 16235
rect 15209 16201 15243 16235
rect 15243 16201 15252 16235
rect 15200 16192 15252 16201
rect 17684 16192 17736 16244
rect 19892 16235 19944 16244
rect 19892 16201 19901 16235
rect 19901 16201 19935 16235
rect 19935 16201 19944 16235
rect 19892 16192 19944 16201
rect 16672 16124 16724 16176
rect 15936 16099 15988 16108
rect 15936 16065 15945 16099
rect 15945 16065 15979 16099
rect 15979 16065 15988 16099
rect 15936 16056 15988 16065
rect 17224 16099 17276 16108
rect 17224 16065 17233 16099
rect 17233 16065 17267 16099
rect 17267 16065 17276 16099
rect 17224 16056 17276 16065
rect 9220 15920 9272 15972
rect 11888 15920 11940 15972
rect 6276 15852 6328 15904
rect 7656 15895 7708 15904
rect 7656 15861 7665 15895
rect 7665 15861 7699 15895
rect 7699 15861 7708 15895
rect 7656 15852 7708 15861
rect 9312 15852 9364 15904
rect 10600 15895 10652 15904
rect 10600 15861 10609 15895
rect 10609 15861 10643 15895
rect 10643 15861 10652 15895
rect 10600 15852 10652 15861
rect 11060 15895 11112 15904
rect 11060 15861 11069 15895
rect 11069 15861 11103 15895
rect 11103 15861 11112 15895
rect 11060 15852 11112 15861
rect 12256 15852 12308 15904
rect 12900 15895 12952 15904
rect 12900 15861 12909 15895
rect 12909 15861 12943 15895
rect 12943 15861 12952 15895
rect 14372 15988 14424 16040
rect 17316 15988 17368 16040
rect 19340 16031 19392 16040
rect 19340 15997 19358 16031
rect 19358 15997 19392 16031
rect 19340 15988 19392 15997
rect 14096 15963 14148 15972
rect 14096 15929 14130 15963
rect 14130 15929 14148 15963
rect 14096 15920 14148 15929
rect 14556 15920 14608 15972
rect 12900 15852 12952 15861
rect 15292 15852 15344 15904
rect 16580 15920 16632 15972
rect 17592 15920 17644 15972
rect 17776 15920 17828 15972
rect 18236 15895 18288 15904
rect 18236 15861 18245 15895
rect 18245 15861 18279 15895
rect 18279 15861 18288 15895
rect 18236 15852 18288 15861
rect 7912 15750 7964 15802
rect 7976 15750 8028 15802
rect 8040 15750 8092 15802
rect 8104 15750 8156 15802
rect 14843 15750 14895 15802
rect 14907 15750 14959 15802
rect 14971 15750 15023 15802
rect 15035 15750 15087 15802
rect 2136 15691 2188 15700
rect 2136 15657 2145 15691
rect 2145 15657 2179 15691
rect 2179 15657 2188 15691
rect 2136 15648 2188 15657
rect 1584 15555 1636 15564
rect 1584 15521 1593 15555
rect 1593 15521 1627 15555
rect 1627 15521 1636 15555
rect 1584 15512 1636 15521
rect 1860 15512 1912 15564
rect 5264 15648 5316 15700
rect 5540 15648 5592 15700
rect 7656 15648 7708 15700
rect 9312 15691 9364 15700
rect 9312 15657 9321 15691
rect 9321 15657 9355 15691
rect 9355 15657 9364 15691
rect 9312 15648 9364 15657
rect 10968 15648 11020 15700
rect 2596 15555 2648 15564
rect 2596 15521 2605 15555
rect 2605 15521 2639 15555
rect 2639 15521 2648 15555
rect 2596 15512 2648 15521
rect 7380 15580 7432 15632
rect 11980 15623 12032 15632
rect 11980 15589 11998 15623
rect 11998 15589 12032 15623
rect 12900 15648 12952 15700
rect 11980 15580 12032 15589
rect 2320 15376 2372 15428
rect 2780 15351 2832 15360
rect 2780 15317 2789 15351
rect 2789 15317 2823 15351
rect 2823 15317 2832 15351
rect 2780 15308 2832 15317
rect 5816 15512 5868 15564
rect 7196 15512 7248 15564
rect 9680 15555 9732 15564
rect 6000 15444 6052 15496
rect 6460 15444 6512 15496
rect 9680 15521 9689 15555
rect 9689 15521 9723 15555
rect 9723 15521 9732 15555
rect 9680 15512 9732 15521
rect 10048 15512 10100 15564
rect 9864 15487 9916 15496
rect 9864 15453 9873 15487
rect 9873 15453 9907 15487
rect 9907 15453 9916 15487
rect 9864 15444 9916 15453
rect 8760 15376 8812 15428
rect 10692 15512 10744 15564
rect 12440 15580 12492 15632
rect 15292 15648 15344 15700
rect 15936 15648 15988 15700
rect 14740 15580 14792 15632
rect 13084 15512 13136 15564
rect 12256 15376 12308 15428
rect 13084 15376 13136 15428
rect 13544 15376 13596 15428
rect 14004 15512 14056 15564
rect 14648 15512 14700 15564
rect 16764 15580 16816 15632
rect 17960 15580 18012 15632
rect 18144 15580 18196 15632
rect 16028 15555 16080 15564
rect 16028 15521 16062 15555
rect 16062 15521 16080 15555
rect 16028 15512 16080 15521
rect 13728 15376 13780 15428
rect 13912 15376 13964 15428
rect 14556 15376 14608 15428
rect 18144 15444 18196 15496
rect 18052 15376 18104 15428
rect 18236 15376 18288 15428
rect 6644 15308 6696 15360
rect 6920 15308 6972 15360
rect 8392 15308 8444 15360
rect 9312 15308 9364 15360
rect 9956 15308 10008 15360
rect 10232 15308 10284 15360
rect 10968 15308 11020 15360
rect 13268 15351 13320 15360
rect 13268 15317 13277 15351
rect 13277 15317 13311 15351
rect 13311 15317 13320 15351
rect 13268 15308 13320 15317
rect 13636 15308 13688 15360
rect 13820 15308 13872 15360
rect 15108 15308 15160 15360
rect 16672 15308 16724 15360
rect 17960 15308 18012 15360
rect 4447 15206 4499 15258
rect 4511 15206 4563 15258
rect 4575 15206 4627 15258
rect 4639 15206 4691 15258
rect 11378 15206 11430 15258
rect 11442 15206 11494 15258
rect 11506 15206 11558 15258
rect 11570 15206 11622 15258
rect 18308 15206 18360 15258
rect 18372 15206 18424 15258
rect 18436 15206 18488 15258
rect 18500 15206 18552 15258
rect 1676 15147 1728 15156
rect 1676 15113 1685 15147
rect 1685 15113 1719 15147
rect 1719 15113 1728 15147
rect 1676 15104 1728 15113
rect 1768 15104 1820 15156
rect 5172 15104 5224 15156
rect 5264 15036 5316 15088
rect 8300 15147 8352 15156
rect 8300 15113 8309 15147
rect 8309 15113 8343 15147
rect 8343 15113 8352 15147
rect 8300 15104 8352 15113
rect 10140 15104 10192 15156
rect 10416 15104 10468 15156
rect 12072 15104 12124 15156
rect 12532 15104 12584 15156
rect 11704 15079 11756 15088
rect 4344 14968 4396 15020
rect 5908 15011 5960 15020
rect 5908 14977 5917 15011
rect 5917 14977 5951 15011
rect 5951 14977 5960 15011
rect 5908 14968 5960 14977
rect 2320 14943 2372 14952
rect 2320 14909 2329 14943
rect 2329 14909 2363 14943
rect 2363 14909 2372 14943
rect 2320 14900 2372 14909
rect 2872 14943 2924 14952
rect 2872 14909 2906 14943
rect 2906 14909 2924 14943
rect 1768 14875 1820 14884
rect 1768 14841 1777 14875
rect 1777 14841 1811 14875
rect 1811 14841 1820 14875
rect 1768 14832 1820 14841
rect 2872 14900 2924 14909
rect 4896 14900 4948 14952
rect 11704 15045 11713 15079
rect 11713 15045 11747 15079
rect 11747 15045 11756 15079
rect 11704 15036 11756 15045
rect 14096 15104 14148 15156
rect 14740 15147 14792 15156
rect 14740 15113 14749 15147
rect 14749 15113 14783 15147
rect 14783 15113 14792 15147
rect 14740 15104 14792 15113
rect 17132 15104 17184 15156
rect 6920 14968 6972 15020
rect 8208 14968 8260 15020
rect 10324 14968 10376 15020
rect 13268 14968 13320 15020
rect 14740 14968 14792 15020
rect 15384 14968 15436 15020
rect 16028 14968 16080 15020
rect 17776 14968 17828 15020
rect 4068 14832 4120 14884
rect 9956 14900 10008 14952
rect 11336 14943 11388 14952
rect 11336 14909 11345 14943
rect 11345 14909 11379 14943
rect 11379 14909 11388 14943
rect 11336 14900 11388 14909
rect 12440 14943 12492 14952
rect 12440 14909 12449 14943
rect 12449 14909 12483 14943
rect 12483 14909 12492 14943
rect 12440 14900 12492 14909
rect 13728 14900 13780 14952
rect 14372 14900 14424 14952
rect 18052 14900 18104 14952
rect 4252 14807 4304 14816
rect 4252 14773 4261 14807
rect 4261 14773 4295 14807
rect 4295 14773 4304 14807
rect 4252 14764 4304 14773
rect 5264 14764 5316 14816
rect 7196 14832 7248 14884
rect 8576 14832 8628 14884
rect 9864 14832 9916 14884
rect 6552 14764 6604 14816
rect 7104 14764 7156 14816
rect 9680 14764 9732 14816
rect 10876 14832 10928 14884
rect 10968 14832 11020 14884
rect 11244 14832 11296 14884
rect 10048 14764 10100 14816
rect 12532 14832 12584 14884
rect 13176 14832 13228 14884
rect 14464 14764 14516 14816
rect 15844 14764 15896 14816
rect 16120 14807 16172 14816
rect 16120 14773 16129 14807
rect 16129 14773 16163 14807
rect 16163 14773 16172 14807
rect 16120 14764 16172 14773
rect 16212 14807 16264 14816
rect 16212 14773 16221 14807
rect 16221 14773 16255 14807
rect 16255 14773 16264 14807
rect 16948 14807 17000 14816
rect 16212 14764 16264 14773
rect 16948 14773 16957 14807
rect 16957 14773 16991 14807
rect 16991 14773 17000 14807
rect 16948 14764 17000 14773
rect 17500 14807 17552 14816
rect 17500 14773 17509 14807
rect 17509 14773 17543 14807
rect 17543 14773 17552 14807
rect 17500 14764 17552 14773
rect 17868 14764 17920 14816
rect 19064 14764 19116 14816
rect 7912 14662 7964 14714
rect 7976 14662 8028 14714
rect 8040 14662 8092 14714
rect 8104 14662 8156 14714
rect 14843 14662 14895 14714
rect 14907 14662 14959 14714
rect 14971 14662 15023 14714
rect 15035 14662 15087 14714
rect 2228 14603 2280 14612
rect 2228 14569 2237 14603
rect 2237 14569 2271 14603
rect 2271 14569 2280 14603
rect 2228 14560 2280 14569
rect 4252 14560 4304 14612
rect 4344 14535 4396 14544
rect 4344 14501 4378 14535
rect 4378 14501 4396 14535
rect 4344 14492 4396 14501
rect 1952 14424 2004 14476
rect 2228 14424 2280 14476
rect 3148 14467 3200 14476
rect 3148 14433 3157 14467
rect 3157 14433 3191 14467
rect 3191 14433 3200 14467
rect 3148 14424 3200 14433
rect 7380 14560 7432 14612
rect 7012 14492 7064 14544
rect 8668 14560 8720 14612
rect 10600 14560 10652 14612
rect 11060 14560 11112 14612
rect 12164 14492 12216 14544
rect 12808 14560 12860 14612
rect 13452 14560 13504 14612
rect 14004 14603 14056 14612
rect 14004 14569 14013 14603
rect 14013 14569 14047 14603
rect 14047 14569 14056 14603
rect 14004 14560 14056 14569
rect 14648 14560 14700 14612
rect 15200 14560 15252 14612
rect 15384 14603 15436 14612
rect 15384 14569 15393 14603
rect 15393 14569 15427 14603
rect 15427 14569 15436 14603
rect 15384 14560 15436 14569
rect 13544 14535 13596 14544
rect 13544 14501 13553 14535
rect 13553 14501 13587 14535
rect 13587 14501 13596 14535
rect 13544 14492 13596 14501
rect 17408 14560 17460 14612
rect 17960 14603 18012 14612
rect 17960 14569 17969 14603
rect 17969 14569 18003 14603
rect 18003 14569 18012 14603
rect 17960 14560 18012 14569
rect 18144 14560 18196 14612
rect 18604 14560 18656 14612
rect 6460 14424 6512 14476
rect 6920 14424 6972 14476
rect 7564 14424 7616 14476
rect 4068 14399 4120 14408
rect 4068 14365 4077 14399
rect 4077 14365 4111 14399
rect 4111 14365 4120 14399
rect 4068 14356 4120 14365
rect 1676 14263 1728 14272
rect 1676 14229 1685 14263
rect 1685 14229 1719 14263
rect 1719 14229 1728 14263
rect 1676 14220 1728 14229
rect 2780 14263 2832 14272
rect 2780 14229 2789 14263
rect 2789 14229 2823 14263
rect 2823 14229 2832 14263
rect 2780 14220 2832 14229
rect 3608 14220 3660 14272
rect 6736 14220 6788 14272
rect 7748 14263 7800 14272
rect 7748 14229 7757 14263
rect 7757 14229 7791 14263
rect 7791 14229 7800 14263
rect 7748 14220 7800 14229
rect 8852 14424 8904 14476
rect 9220 14424 9272 14476
rect 9956 14467 10008 14476
rect 9956 14433 9965 14467
rect 9965 14433 9999 14467
rect 9999 14433 10008 14467
rect 9956 14424 10008 14433
rect 10692 14424 10744 14476
rect 10876 14467 10928 14476
rect 10876 14433 10910 14467
rect 10910 14433 10928 14467
rect 10876 14424 10928 14433
rect 11244 14424 11296 14476
rect 12256 14424 12308 14476
rect 12716 14424 12768 14476
rect 10048 14288 10100 14340
rect 10416 14288 10468 14340
rect 10140 14220 10192 14272
rect 12164 14356 12216 14408
rect 14740 14424 14792 14476
rect 13544 14356 13596 14408
rect 16948 14492 17000 14544
rect 15660 14424 15712 14476
rect 16764 14467 16816 14476
rect 16764 14433 16773 14467
rect 16773 14433 16807 14467
rect 16807 14433 16816 14467
rect 16764 14424 16816 14433
rect 19064 14356 19116 14408
rect 13176 14288 13228 14340
rect 11980 14263 12032 14272
rect 11980 14229 11989 14263
rect 11989 14229 12023 14263
rect 12023 14229 12032 14263
rect 11980 14220 12032 14229
rect 12072 14220 12124 14272
rect 14280 14220 14332 14272
rect 14372 14220 14424 14272
rect 15200 14220 15252 14272
rect 15476 14220 15528 14272
rect 4447 14118 4499 14170
rect 4511 14118 4563 14170
rect 4575 14118 4627 14170
rect 4639 14118 4691 14170
rect 11378 14118 11430 14170
rect 11442 14118 11494 14170
rect 11506 14118 11558 14170
rect 11570 14118 11622 14170
rect 18308 14118 18360 14170
rect 18372 14118 18424 14170
rect 18436 14118 18488 14170
rect 18500 14118 18552 14170
rect 2044 14016 2096 14068
rect 2320 14016 2372 14068
rect 4344 14016 4396 14068
rect 5908 14016 5960 14068
rect 6644 14059 6696 14068
rect 6644 14025 6653 14059
rect 6653 14025 6687 14059
rect 6687 14025 6696 14059
rect 6644 14016 6696 14025
rect 6736 14016 6788 14068
rect 5080 13948 5132 14000
rect 6092 13948 6144 14000
rect 9680 14016 9732 14068
rect 9864 14016 9916 14068
rect 8208 13948 8260 14000
rect 9496 13948 9548 14000
rect 3148 13923 3200 13932
rect 3148 13889 3157 13923
rect 3157 13889 3191 13923
rect 3191 13889 3200 13923
rect 3148 13880 3200 13889
rect 1584 13855 1636 13864
rect 1584 13821 1593 13855
rect 1593 13821 1627 13855
rect 1627 13821 1636 13855
rect 1584 13812 1636 13821
rect 1768 13855 1820 13864
rect 1768 13821 1777 13855
rect 1777 13821 1811 13855
rect 1811 13821 1820 13855
rect 1768 13812 1820 13821
rect 2320 13855 2372 13864
rect 2320 13821 2329 13855
rect 2329 13821 2363 13855
rect 2363 13821 2372 13855
rect 2320 13812 2372 13821
rect 3608 13855 3660 13864
rect 3608 13821 3617 13855
rect 3617 13821 3651 13855
rect 3651 13821 3660 13855
rect 4068 13855 4120 13864
rect 3608 13812 3660 13821
rect 4068 13821 4077 13855
rect 4077 13821 4111 13855
rect 4111 13821 4120 13855
rect 4068 13812 4120 13821
rect 6920 13880 6972 13932
rect 7748 13880 7800 13932
rect 12072 14016 12124 14068
rect 13728 14016 13780 14068
rect 13268 13948 13320 14000
rect 6000 13812 6052 13864
rect 9404 13812 9456 13864
rect 12716 13880 12768 13932
rect 14280 13880 14332 13932
rect 16120 14016 16172 14068
rect 15660 13923 15712 13932
rect 15660 13889 15669 13923
rect 15669 13889 15703 13923
rect 15703 13889 15712 13923
rect 15660 13880 15712 13889
rect 15844 13923 15896 13932
rect 15844 13889 15853 13923
rect 15853 13889 15887 13923
rect 15887 13889 15896 13923
rect 15844 13880 15896 13889
rect 5540 13744 5592 13796
rect 7012 13787 7064 13796
rect 7012 13753 7021 13787
rect 7021 13753 7055 13787
rect 7055 13753 7064 13787
rect 7012 13744 7064 13753
rect 7104 13787 7156 13796
rect 7104 13753 7113 13787
rect 7113 13753 7147 13787
rect 7147 13753 7156 13787
rect 7104 13744 7156 13753
rect 9128 13744 9180 13796
rect 9634 13744 9686 13796
rect 10600 13744 10652 13796
rect 13268 13812 13320 13864
rect 14740 13812 14792 13864
rect 20720 14016 20772 14068
rect 17408 13991 17460 14000
rect 17408 13957 17417 13991
rect 17417 13957 17451 13991
rect 17451 13957 17460 13991
rect 17408 13948 17460 13957
rect 18052 13948 18104 14000
rect 19064 13812 19116 13864
rect 19248 13812 19300 13864
rect 6828 13676 6880 13728
rect 7472 13676 7524 13728
rect 12532 13676 12584 13728
rect 13176 13676 13228 13728
rect 15476 13676 15528 13728
rect 17776 13719 17828 13728
rect 17776 13685 17785 13719
rect 17785 13685 17819 13719
rect 17819 13685 17828 13719
rect 17776 13676 17828 13685
rect 7912 13574 7964 13626
rect 7976 13574 8028 13626
rect 8040 13574 8092 13626
rect 8104 13574 8156 13626
rect 14843 13574 14895 13626
rect 14907 13574 14959 13626
rect 14971 13574 15023 13626
rect 15035 13574 15087 13626
rect 2320 13472 2372 13524
rect 2596 13472 2648 13524
rect 8392 13472 8444 13524
rect 9956 13472 10008 13524
rect 11888 13515 11940 13524
rect 11888 13481 11897 13515
rect 11897 13481 11931 13515
rect 11931 13481 11940 13515
rect 11888 13472 11940 13481
rect 12348 13515 12400 13524
rect 12348 13481 12357 13515
rect 12357 13481 12391 13515
rect 12391 13481 12400 13515
rect 12348 13472 12400 13481
rect 12440 13472 12492 13524
rect 15476 13515 15528 13524
rect 15476 13481 15485 13515
rect 15485 13481 15519 13515
rect 15519 13481 15528 13515
rect 15476 13472 15528 13481
rect 16212 13472 16264 13524
rect 16580 13515 16632 13524
rect 16580 13481 16589 13515
rect 16589 13481 16623 13515
rect 16623 13481 16632 13515
rect 16580 13472 16632 13481
rect 1492 13336 1544 13388
rect 3148 13404 3200 13456
rect 2780 13336 2832 13388
rect 2872 13336 2924 13388
rect 8944 13404 8996 13456
rect 10784 13404 10836 13456
rect 17224 13404 17276 13456
rect 5540 13268 5592 13320
rect 5908 13311 5960 13320
rect 5908 13277 5917 13311
rect 5917 13277 5951 13311
rect 5951 13277 5960 13311
rect 5908 13268 5960 13277
rect 6460 13268 6512 13320
rect 10232 13336 10284 13388
rect 10876 13336 10928 13388
rect 6644 13200 6696 13252
rect 8208 13200 8260 13252
rect 9496 13268 9548 13320
rect 11796 13336 11848 13388
rect 17960 13379 18012 13388
rect 17960 13345 17969 13379
rect 17969 13345 18003 13379
rect 18003 13345 18012 13379
rect 17960 13336 18012 13345
rect 9128 13200 9180 13252
rect 10140 13200 10192 13252
rect 6736 13132 6788 13184
rect 6920 13132 6972 13184
rect 8116 13132 8168 13184
rect 12164 13268 12216 13320
rect 13636 13311 13688 13320
rect 13636 13277 13645 13311
rect 13645 13277 13679 13311
rect 13679 13277 13688 13311
rect 13636 13268 13688 13277
rect 13728 13311 13780 13320
rect 13728 13277 13737 13311
rect 13737 13277 13771 13311
rect 13771 13277 13780 13311
rect 17776 13311 17828 13320
rect 13728 13268 13780 13277
rect 17776 13277 17785 13311
rect 17785 13277 17819 13311
rect 17819 13277 17828 13311
rect 17776 13268 17828 13277
rect 14004 13132 14056 13184
rect 17592 13132 17644 13184
rect 18972 13132 19024 13184
rect 4447 13030 4499 13082
rect 4511 13030 4563 13082
rect 4575 13030 4627 13082
rect 4639 13030 4691 13082
rect 11378 13030 11430 13082
rect 11442 13030 11494 13082
rect 11506 13030 11558 13082
rect 11570 13030 11622 13082
rect 18308 13030 18360 13082
rect 18372 13030 18424 13082
rect 18436 13030 18488 13082
rect 18500 13030 18552 13082
rect 1492 12971 1544 12980
rect 1492 12937 1501 12971
rect 1501 12937 1535 12971
rect 1535 12937 1544 12971
rect 1492 12928 1544 12937
rect 1860 12928 1912 12980
rect 2412 12928 2464 12980
rect 6828 12928 6880 12980
rect 9128 12971 9180 12980
rect 4712 12860 4764 12912
rect 6000 12835 6052 12844
rect 2412 12767 2464 12776
rect 2412 12733 2421 12767
rect 2421 12733 2455 12767
rect 2455 12733 2464 12767
rect 2412 12724 2464 12733
rect 2596 12724 2648 12776
rect 4804 12724 4856 12776
rect 6000 12801 6009 12835
rect 6009 12801 6043 12835
rect 6043 12801 6052 12835
rect 6000 12792 6052 12801
rect 6828 12792 6880 12844
rect 7288 12835 7340 12844
rect 7288 12801 7297 12835
rect 7297 12801 7331 12835
rect 7331 12801 7340 12835
rect 7288 12792 7340 12801
rect 5724 12767 5776 12776
rect 2688 12656 2740 12708
rect 4896 12656 4948 12708
rect 5724 12733 5753 12767
rect 5753 12733 5776 12767
rect 5724 12724 5776 12733
rect 5908 12724 5960 12776
rect 7472 12724 7524 12776
rect 7748 12767 7800 12776
rect 7748 12733 7757 12767
rect 7757 12733 7791 12767
rect 7791 12733 7800 12767
rect 7748 12724 7800 12733
rect 7564 12656 7616 12708
rect 9128 12937 9137 12971
rect 9137 12937 9171 12971
rect 9171 12937 9180 12971
rect 9128 12928 9180 12937
rect 12532 12928 12584 12980
rect 13636 12928 13688 12980
rect 15660 12928 15712 12980
rect 18788 12928 18840 12980
rect 9772 12860 9824 12912
rect 10048 12860 10100 12912
rect 10600 12903 10652 12912
rect 10600 12869 10609 12903
rect 10609 12869 10643 12903
rect 10643 12869 10652 12903
rect 10600 12860 10652 12869
rect 12256 12860 12308 12912
rect 13268 12835 13320 12844
rect 13268 12801 13277 12835
rect 13277 12801 13311 12835
rect 13311 12801 13320 12835
rect 13268 12792 13320 12801
rect 14004 12835 14056 12844
rect 14004 12801 14013 12835
rect 14013 12801 14047 12835
rect 14047 12801 14056 12835
rect 14004 12792 14056 12801
rect 14372 12860 14424 12912
rect 14740 12860 14792 12912
rect 17316 12792 17368 12844
rect 17776 12835 17828 12844
rect 17776 12801 17785 12835
rect 17785 12801 17819 12835
rect 17819 12801 17828 12835
rect 17776 12792 17828 12801
rect 18052 12792 18104 12844
rect 19156 12835 19208 12844
rect 19156 12801 19165 12835
rect 19165 12801 19199 12835
rect 19199 12801 19208 12835
rect 19156 12792 19208 12801
rect 11704 12724 11756 12776
rect 11980 12724 12032 12776
rect 13820 12724 13872 12776
rect 2964 12631 3016 12640
rect 2964 12597 2973 12631
rect 2973 12597 3007 12631
rect 3007 12597 3016 12631
rect 2964 12588 3016 12597
rect 5540 12588 5592 12640
rect 7196 12631 7248 12640
rect 7196 12597 7205 12631
rect 7205 12597 7239 12631
rect 7239 12597 7248 12631
rect 7196 12588 7248 12597
rect 8760 12588 8812 12640
rect 11152 12588 11204 12640
rect 11796 12588 11848 12640
rect 14648 12724 14700 12776
rect 16120 12699 16172 12708
rect 16120 12665 16138 12699
rect 16138 12665 16172 12699
rect 16120 12656 16172 12665
rect 17592 12724 17644 12776
rect 18972 12767 19024 12776
rect 18972 12733 18981 12767
rect 18981 12733 19015 12767
rect 19015 12733 19024 12767
rect 18972 12724 19024 12733
rect 17316 12631 17368 12640
rect 17316 12597 17325 12631
rect 17325 12597 17359 12631
rect 17359 12597 17368 12631
rect 17316 12588 17368 12597
rect 7912 12486 7964 12538
rect 7976 12486 8028 12538
rect 8040 12486 8092 12538
rect 8104 12486 8156 12538
rect 14843 12486 14895 12538
rect 14907 12486 14959 12538
rect 14971 12486 15023 12538
rect 15035 12486 15087 12538
rect 1768 12427 1820 12436
rect 1768 12393 1777 12427
rect 1777 12393 1811 12427
rect 1811 12393 1820 12427
rect 1768 12384 1820 12393
rect 2412 12427 2464 12436
rect 2412 12393 2421 12427
rect 2421 12393 2455 12427
rect 2455 12393 2464 12427
rect 2412 12384 2464 12393
rect 2688 12427 2740 12436
rect 2688 12393 2697 12427
rect 2697 12393 2731 12427
rect 2731 12393 2740 12427
rect 2688 12384 2740 12393
rect 2044 12248 2096 12300
rect 2504 12248 2556 12300
rect 4712 12316 4764 12368
rect 5724 12384 5776 12436
rect 7564 12427 7616 12436
rect 6828 12316 6880 12368
rect 7012 12359 7064 12368
rect 7012 12325 7030 12359
rect 7030 12325 7064 12359
rect 7564 12393 7573 12427
rect 7573 12393 7607 12427
rect 7607 12393 7616 12427
rect 7564 12384 7616 12393
rect 9220 12427 9272 12436
rect 9220 12393 9229 12427
rect 9229 12393 9263 12427
rect 9263 12393 9272 12427
rect 9220 12384 9272 12393
rect 12624 12427 12676 12436
rect 7012 12316 7064 12325
rect 12624 12393 12633 12427
rect 12633 12393 12667 12427
rect 12667 12393 12676 12427
rect 12624 12384 12676 12393
rect 16488 12384 16540 12436
rect 17960 12384 18012 12436
rect 3148 12291 3200 12300
rect 3148 12257 3157 12291
rect 3157 12257 3191 12291
rect 3191 12257 3200 12291
rect 3148 12248 3200 12257
rect 2964 12180 3016 12232
rect 3884 12248 3936 12300
rect 4804 12248 4856 12300
rect 6000 12248 6052 12300
rect 8668 12248 8720 12300
rect 8760 12291 8812 12300
rect 8760 12257 8769 12291
rect 8769 12257 8803 12291
rect 8803 12257 8812 12291
rect 8760 12248 8812 12257
rect 14004 12316 14056 12368
rect 17776 12316 17828 12368
rect 19248 12316 19300 12368
rect 13820 12291 13872 12300
rect 3332 12112 3384 12164
rect 7564 12180 7616 12232
rect 8208 12223 8260 12232
rect 8208 12189 8217 12223
rect 8217 12189 8251 12223
rect 8251 12189 8260 12223
rect 8208 12180 8260 12189
rect 9956 12223 10008 12232
rect 9956 12189 9965 12223
rect 9965 12189 9999 12223
rect 9999 12189 10008 12223
rect 11796 12223 11848 12232
rect 9956 12180 10008 12189
rect 11796 12189 11805 12223
rect 11805 12189 11839 12223
rect 11839 12189 11848 12223
rect 11796 12180 11848 12189
rect 4252 12044 4304 12096
rect 4804 12044 4856 12096
rect 4988 12044 5040 12096
rect 5908 12087 5960 12096
rect 5908 12053 5917 12087
rect 5917 12053 5951 12087
rect 5951 12053 5960 12087
rect 5908 12044 5960 12053
rect 6000 12044 6052 12096
rect 8484 12112 8536 12164
rect 8576 12087 8628 12096
rect 8576 12053 8585 12087
rect 8585 12053 8619 12087
rect 8619 12053 8628 12087
rect 8576 12044 8628 12053
rect 13820 12257 13829 12291
rect 13829 12257 13863 12291
rect 13863 12257 13872 12291
rect 13820 12248 13872 12257
rect 15292 12248 15344 12300
rect 16304 12248 16356 12300
rect 17316 12291 17368 12300
rect 17316 12257 17325 12291
rect 17325 12257 17359 12291
rect 17359 12257 17368 12291
rect 21088 12291 21140 12300
rect 17316 12248 17368 12257
rect 21088 12257 21106 12291
rect 21106 12257 21140 12291
rect 21088 12248 21140 12257
rect 12716 12112 12768 12164
rect 13912 12112 13964 12164
rect 13360 12044 13412 12096
rect 13636 12087 13688 12096
rect 13636 12053 13645 12087
rect 13645 12053 13679 12087
rect 13679 12053 13688 12087
rect 15844 12180 15896 12232
rect 16120 12112 16172 12164
rect 18788 12112 18840 12164
rect 19156 12112 19208 12164
rect 13636 12044 13688 12053
rect 14372 12044 14424 12096
rect 4447 11942 4499 11994
rect 4511 11942 4563 11994
rect 4575 11942 4627 11994
rect 4639 11942 4691 11994
rect 11378 11942 11430 11994
rect 11442 11942 11494 11994
rect 11506 11942 11558 11994
rect 11570 11942 11622 11994
rect 18308 11942 18360 11994
rect 18372 11942 18424 11994
rect 18436 11942 18488 11994
rect 18500 11942 18552 11994
rect 1676 11840 1728 11892
rect 2044 11840 2096 11892
rect 2504 11840 2556 11892
rect 4068 11840 4120 11892
rect 6092 11840 6144 11892
rect 7196 11840 7248 11892
rect 8300 11840 8352 11892
rect 11060 11883 11112 11892
rect 3884 11747 3936 11756
rect 3884 11713 3893 11747
rect 3893 11713 3927 11747
rect 3927 11713 3936 11747
rect 3884 11704 3936 11713
rect 4896 11747 4948 11756
rect 4896 11713 4905 11747
rect 4905 11713 4939 11747
rect 4939 11713 4948 11747
rect 4896 11704 4948 11713
rect 1860 11636 1912 11688
rect 2504 11636 2556 11688
rect 3424 11636 3476 11688
rect 8576 11772 8628 11824
rect 11060 11849 11069 11883
rect 11069 11849 11103 11883
rect 11103 11849 11112 11883
rect 11060 11840 11112 11849
rect 12716 11840 12768 11892
rect 12992 11840 13044 11892
rect 14188 11840 14240 11892
rect 15844 11883 15896 11892
rect 15844 11849 15853 11883
rect 15853 11849 15887 11883
rect 15887 11849 15896 11883
rect 15844 11840 15896 11849
rect 21088 11840 21140 11892
rect 7104 11747 7156 11756
rect 7104 11713 7113 11747
rect 7113 11713 7147 11747
rect 7147 11713 7156 11747
rect 7104 11704 7156 11713
rect 7472 11704 7524 11756
rect 8208 11704 8260 11756
rect 12072 11704 12124 11756
rect 9680 11679 9732 11688
rect 1400 11543 1452 11552
rect 1400 11509 1409 11543
rect 1409 11509 1443 11543
rect 1443 11509 1452 11543
rect 1400 11500 1452 11509
rect 2872 11543 2924 11552
rect 2872 11509 2881 11543
rect 2881 11509 2915 11543
rect 2915 11509 2924 11543
rect 2872 11500 2924 11509
rect 4436 11568 4488 11620
rect 7748 11568 7800 11620
rect 9680 11645 9689 11679
rect 9689 11645 9723 11679
rect 9723 11645 9732 11679
rect 9680 11636 9732 11645
rect 9956 11679 10008 11688
rect 9956 11645 9990 11679
rect 9990 11645 10008 11679
rect 9956 11636 10008 11645
rect 13820 11704 13872 11756
rect 10508 11568 10560 11620
rect 4712 11543 4764 11552
rect 4712 11509 4721 11543
rect 4721 11509 4755 11543
rect 4755 11509 4764 11543
rect 4712 11500 4764 11509
rect 4988 11500 5040 11552
rect 9128 11500 9180 11552
rect 12348 11611 12400 11620
rect 12348 11577 12357 11611
rect 12357 11577 12391 11611
rect 12391 11577 12400 11611
rect 12348 11568 12400 11577
rect 12900 11568 12952 11620
rect 16488 11772 16540 11824
rect 14280 11747 14332 11756
rect 14280 11713 14289 11747
rect 14289 11713 14323 11747
rect 14323 11713 14332 11747
rect 14280 11704 14332 11713
rect 15292 11747 15344 11756
rect 15292 11713 15301 11747
rect 15301 11713 15335 11747
rect 15335 11713 15344 11747
rect 15292 11704 15344 11713
rect 16304 11747 16356 11756
rect 16304 11713 16313 11747
rect 16313 11713 16347 11747
rect 16347 11713 16356 11747
rect 16304 11704 16356 11713
rect 19248 11704 19300 11756
rect 15200 11636 15252 11688
rect 18788 11679 18840 11688
rect 18788 11645 18806 11679
rect 18806 11645 18840 11679
rect 18788 11636 18840 11645
rect 21364 11679 21416 11688
rect 21364 11645 21373 11679
rect 21373 11645 21407 11679
rect 21407 11645 21416 11679
rect 21364 11636 21416 11645
rect 13452 11500 13504 11552
rect 14464 11543 14516 11552
rect 14464 11509 14473 11543
rect 14473 11509 14507 11543
rect 14507 11509 14516 11543
rect 14464 11500 14516 11509
rect 7912 11398 7964 11450
rect 7976 11398 8028 11450
rect 8040 11398 8092 11450
rect 8104 11398 8156 11450
rect 14843 11398 14895 11450
rect 14907 11398 14959 11450
rect 14971 11398 15023 11450
rect 15035 11398 15087 11450
rect 1860 11339 1912 11348
rect 1860 11305 1869 11339
rect 1869 11305 1903 11339
rect 1903 11305 1912 11339
rect 1860 11296 1912 11305
rect 3424 11339 3476 11348
rect 3424 11305 3433 11339
rect 3433 11305 3467 11339
rect 3467 11305 3476 11339
rect 3424 11296 3476 11305
rect 4160 11296 4212 11348
rect 4436 11339 4488 11348
rect 4436 11305 4445 11339
rect 4445 11305 4479 11339
rect 4479 11305 4488 11339
rect 4436 11296 4488 11305
rect 4712 11296 4764 11348
rect 5172 11296 5224 11348
rect 7288 11296 7340 11348
rect 1400 11203 1452 11212
rect 1400 11169 1409 11203
rect 1409 11169 1443 11203
rect 1443 11169 1452 11203
rect 1400 11160 1452 11169
rect 2780 11203 2832 11212
rect 2780 11169 2789 11203
rect 2789 11169 2823 11203
rect 2823 11169 2832 11203
rect 2780 11160 2832 11169
rect 2872 11135 2924 11144
rect 2872 11101 2881 11135
rect 2881 11101 2915 11135
rect 2915 11101 2924 11135
rect 2872 11092 2924 11101
rect 3056 11135 3108 11144
rect 3056 11101 3065 11135
rect 3065 11101 3099 11135
rect 3099 11101 3108 11135
rect 3056 11092 3108 11101
rect 4068 11092 4120 11144
rect 6000 11092 6052 11144
rect 7012 11228 7064 11280
rect 6644 11160 6696 11212
rect 8300 11296 8352 11348
rect 8668 11296 8720 11348
rect 12256 11296 12308 11348
rect 13820 11296 13872 11348
rect 14464 11296 14516 11348
rect 15292 11296 15344 11348
rect 11060 11228 11112 11280
rect 6736 11092 6788 11144
rect 7380 11092 7432 11144
rect 8024 11160 8076 11212
rect 12716 11228 12768 11280
rect 14280 11228 14332 11280
rect 14924 11228 14976 11280
rect 16488 11271 16540 11280
rect 16488 11237 16522 11271
rect 16522 11237 16540 11271
rect 16488 11228 16540 11237
rect 7564 11024 7616 11076
rect 2412 10999 2464 11008
rect 2412 10965 2421 10999
rect 2421 10965 2455 10999
rect 2455 10965 2464 10999
rect 2412 10956 2464 10965
rect 4804 10999 4856 11008
rect 4804 10965 4813 10999
rect 4813 10965 4847 10999
rect 4847 10965 4856 10999
rect 4804 10956 4856 10965
rect 7656 10956 7708 11008
rect 9680 11092 9732 11144
rect 12072 11092 12124 11144
rect 13268 11160 13320 11212
rect 13636 11160 13688 11212
rect 17316 11160 17368 11212
rect 11244 10956 11296 11008
rect 17592 10999 17644 11008
rect 17592 10965 17601 10999
rect 17601 10965 17635 10999
rect 17635 10965 17644 10999
rect 17592 10956 17644 10965
rect 4447 10854 4499 10906
rect 4511 10854 4563 10906
rect 4575 10854 4627 10906
rect 4639 10854 4691 10906
rect 11378 10854 11430 10906
rect 11442 10854 11494 10906
rect 11506 10854 11558 10906
rect 11570 10854 11622 10906
rect 18308 10854 18360 10906
rect 18372 10854 18424 10906
rect 18436 10854 18488 10906
rect 18500 10854 18552 10906
rect 2504 10795 2556 10804
rect 2504 10761 2513 10795
rect 2513 10761 2547 10795
rect 2547 10761 2556 10795
rect 2504 10752 2556 10761
rect 3056 10752 3108 10804
rect 2044 10616 2096 10668
rect 4252 10616 4304 10668
rect 4804 10616 4856 10668
rect 7656 10752 7708 10804
rect 8024 10795 8076 10804
rect 8024 10761 8033 10795
rect 8033 10761 8067 10795
rect 8067 10761 8076 10795
rect 8024 10752 8076 10761
rect 9680 10752 9732 10804
rect 10692 10752 10744 10804
rect 11796 10752 11848 10804
rect 13268 10795 13320 10804
rect 13268 10761 13277 10795
rect 13277 10761 13311 10795
rect 13311 10761 13320 10795
rect 13268 10752 13320 10761
rect 14924 10795 14976 10804
rect 14924 10761 14933 10795
rect 14933 10761 14967 10795
rect 14967 10761 14976 10795
rect 14924 10752 14976 10761
rect 2412 10548 2464 10600
rect 6736 10548 6788 10600
rect 1400 10455 1452 10464
rect 1400 10421 1409 10455
rect 1409 10421 1443 10455
rect 1443 10421 1452 10455
rect 1400 10412 1452 10421
rect 4068 10480 4120 10532
rect 7748 10616 7800 10668
rect 8300 10616 8352 10668
rect 9036 10659 9088 10668
rect 9036 10625 9045 10659
rect 9045 10625 9079 10659
rect 9079 10625 9088 10659
rect 9036 10616 9088 10625
rect 9680 10616 9732 10668
rect 16488 10616 16540 10668
rect 19248 10616 19300 10668
rect 8576 10548 8628 10600
rect 11244 10548 11296 10600
rect 12716 10548 12768 10600
rect 13636 10548 13688 10600
rect 13820 10591 13872 10600
rect 13820 10557 13854 10591
rect 13854 10557 13872 10591
rect 13820 10548 13872 10557
rect 4804 10455 4856 10464
rect 4804 10421 4813 10455
rect 4813 10421 4847 10455
rect 4847 10421 4856 10455
rect 4804 10412 4856 10421
rect 5356 10412 5408 10464
rect 5724 10412 5776 10464
rect 6368 10412 6420 10464
rect 9772 10480 9824 10532
rect 10048 10480 10100 10532
rect 12532 10480 12584 10532
rect 15200 10480 15252 10532
rect 17592 10480 17644 10532
rect 8208 10412 8260 10464
rect 8944 10455 8996 10464
rect 8944 10421 8953 10455
rect 8953 10421 8987 10455
rect 8987 10421 8996 10455
rect 8944 10412 8996 10421
rect 15752 10455 15804 10464
rect 15752 10421 15761 10455
rect 15761 10421 15795 10455
rect 15795 10421 15804 10455
rect 16120 10455 16172 10464
rect 15752 10412 15804 10421
rect 16120 10421 16129 10455
rect 16129 10421 16163 10455
rect 16163 10421 16172 10455
rect 16120 10412 16172 10421
rect 16948 10412 17000 10464
rect 7912 10310 7964 10362
rect 7976 10310 8028 10362
rect 8040 10310 8092 10362
rect 8104 10310 8156 10362
rect 14843 10310 14895 10362
rect 14907 10310 14959 10362
rect 14971 10310 15023 10362
rect 15035 10310 15087 10362
rect 2596 10208 2648 10260
rect 4804 10251 4856 10260
rect 4804 10217 4813 10251
rect 4813 10217 4847 10251
rect 4847 10217 4856 10251
rect 4804 10208 4856 10217
rect 5080 10208 5132 10260
rect 5816 10208 5868 10260
rect 6736 10208 6788 10260
rect 7012 10208 7064 10260
rect 8208 10251 8260 10260
rect 8208 10217 8217 10251
rect 8217 10217 8251 10251
rect 8251 10217 8260 10251
rect 8208 10208 8260 10217
rect 11704 10208 11756 10260
rect 12348 10208 12400 10260
rect 12900 10208 12952 10260
rect 15200 10251 15252 10260
rect 15200 10217 15209 10251
rect 15209 10217 15243 10251
rect 15243 10217 15252 10251
rect 15200 10208 15252 10217
rect 16948 10251 17000 10260
rect 16948 10217 16957 10251
rect 16957 10217 16991 10251
rect 16991 10217 17000 10251
rect 16948 10208 17000 10217
rect 18696 10208 18748 10260
rect 1400 10115 1452 10124
rect 1400 10081 1409 10115
rect 1409 10081 1443 10115
rect 1443 10081 1452 10115
rect 1400 10072 1452 10081
rect 1584 10072 1636 10124
rect 15752 10140 15804 10192
rect 16120 10140 16172 10192
rect 2964 10115 3016 10124
rect 2964 10081 2982 10115
rect 2982 10081 3016 10115
rect 2964 10072 3016 10081
rect 5080 10072 5132 10124
rect 6828 10072 6880 10124
rect 4068 10004 4120 10056
rect 4344 10047 4396 10056
rect 4344 10013 4353 10047
rect 4353 10013 4387 10047
rect 4387 10013 4396 10047
rect 4344 10004 4396 10013
rect 7104 10047 7156 10056
rect 4252 9936 4304 9988
rect 4896 9936 4948 9988
rect 7104 10013 7113 10047
rect 7113 10013 7147 10047
rect 7147 10013 7156 10047
rect 7104 10004 7156 10013
rect 9588 10072 9640 10124
rect 9680 10072 9732 10124
rect 10692 10115 10744 10124
rect 10692 10081 10701 10115
rect 10701 10081 10735 10115
rect 10735 10081 10744 10115
rect 10692 10072 10744 10081
rect 11060 10072 11112 10124
rect 12532 10072 12584 10124
rect 11244 10047 11296 10056
rect 11244 10013 11253 10047
rect 11253 10013 11287 10047
rect 11287 10013 11296 10047
rect 11244 10004 11296 10013
rect 17592 10004 17644 10056
rect 2044 9868 2096 9920
rect 4447 9766 4499 9818
rect 4511 9766 4563 9818
rect 4575 9766 4627 9818
rect 4639 9766 4691 9818
rect 11378 9766 11430 9818
rect 11442 9766 11494 9818
rect 11506 9766 11558 9818
rect 11570 9766 11622 9818
rect 18308 9766 18360 9818
rect 18372 9766 18424 9818
rect 18436 9766 18488 9818
rect 18500 9766 18552 9818
rect 9680 9664 9732 9716
rect 11060 9707 11112 9716
rect 11060 9673 11069 9707
rect 11069 9673 11103 9707
rect 11103 9673 11112 9707
rect 11060 9664 11112 9673
rect 2320 9596 2372 9648
rect 2872 9596 2924 9648
rect 3884 9596 3936 9648
rect 5080 9596 5132 9648
rect 6644 9639 6696 9648
rect 6644 9605 6653 9639
rect 6653 9605 6687 9639
rect 6687 9605 6696 9639
rect 6644 9596 6696 9605
rect 9588 9639 9640 9648
rect 9588 9605 9597 9639
rect 9597 9605 9631 9639
rect 9631 9605 9640 9639
rect 9588 9596 9640 9605
rect 2780 9528 2832 9580
rect 4068 9528 4120 9580
rect 1400 9503 1452 9512
rect 1400 9469 1409 9503
rect 1409 9469 1443 9503
rect 1443 9469 1452 9503
rect 1400 9460 1452 9469
rect 1860 9503 1912 9512
rect 1860 9469 1869 9503
rect 1869 9469 1903 9503
rect 1903 9469 1912 9503
rect 1860 9460 1912 9469
rect 4988 9528 5040 9580
rect 6828 9528 6880 9580
rect 7656 9528 7708 9580
rect 4344 9460 4396 9512
rect 5356 9460 5408 9512
rect 7104 9460 7156 9512
rect 9772 9460 9824 9512
rect 3424 9367 3476 9376
rect 3424 9333 3433 9367
rect 3433 9333 3467 9367
rect 3467 9333 3476 9367
rect 3424 9324 3476 9333
rect 4068 9324 4120 9376
rect 6552 9324 6604 9376
rect 7656 9392 7708 9444
rect 8852 9324 8904 9376
rect 9404 9324 9456 9376
rect 14096 9324 14148 9376
rect 7912 9222 7964 9274
rect 7976 9222 8028 9274
rect 8040 9222 8092 9274
rect 8104 9222 8156 9274
rect 14843 9222 14895 9274
rect 14907 9222 14959 9274
rect 14971 9222 15023 9274
rect 15035 9222 15087 9274
rect 1860 9120 1912 9172
rect 5448 9120 5500 9172
rect 9772 9163 9824 9172
rect 1400 9095 1452 9104
rect 1400 9061 1409 9095
rect 1409 9061 1443 9095
rect 1443 9061 1452 9095
rect 1400 9052 1452 9061
rect 9772 9129 9781 9163
rect 9781 9129 9815 9163
rect 9815 9129 9824 9163
rect 9772 9120 9824 9129
rect 2136 8848 2188 8900
rect 2780 8984 2832 9036
rect 2596 8916 2648 8968
rect 8944 9052 8996 9104
rect 7288 8984 7340 9036
rect 9312 8984 9364 9036
rect 5172 8916 5224 8968
rect 7656 8959 7708 8968
rect 7656 8925 7665 8959
rect 7665 8925 7699 8959
rect 7699 8925 7708 8959
rect 7656 8916 7708 8925
rect 17500 8848 17552 8900
rect 4804 8780 4856 8832
rect 9404 8823 9456 8832
rect 9404 8789 9413 8823
rect 9413 8789 9447 8823
rect 9447 8789 9456 8823
rect 9404 8780 9456 8789
rect 4447 8678 4499 8730
rect 4511 8678 4563 8730
rect 4575 8678 4627 8730
rect 4639 8678 4691 8730
rect 11378 8678 11430 8730
rect 11442 8678 11494 8730
rect 11506 8678 11558 8730
rect 11570 8678 11622 8730
rect 18308 8678 18360 8730
rect 18372 8678 18424 8730
rect 18436 8678 18488 8730
rect 18500 8678 18552 8730
rect 1952 8576 2004 8628
rect 5172 8576 5224 8628
rect 9772 8508 9824 8560
rect 8392 8483 8444 8492
rect 8392 8449 8401 8483
rect 8401 8449 8435 8483
rect 8435 8449 8444 8483
rect 8392 8440 8444 8449
rect 13084 8440 13136 8492
rect 1952 8415 2004 8424
rect 1952 8381 1961 8415
rect 1961 8381 1995 8415
rect 1995 8381 2004 8415
rect 1952 8372 2004 8381
rect 4896 8372 4948 8424
rect 2044 8304 2096 8356
rect 4252 8304 4304 8356
rect 8300 8304 8352 8356
rect 1400 8279 1452 8288
rect 1400 8245 1409 8279
rect 1409 8245 1443 8279
rect 1443 8245 1452 8279
rect 1400 8236 1452 8245
rect 4436 8236 4488 8288
rect 5448 8279 5500 8288
rect 5448 8245 5457 8279
rect 5457 8245 5491 8279
rect 5491 8245 5500 8279
rect 5448 8236 5500 8245
rect 8208 8236 8260 8288
rect 7912 8134 7964 8186
rect 7976 8134 8028 8186
rect 8040 8134 8092 8186
rect 8104 8134 8156 8186
rect 14843 8134 14895 8186
rect 14907 8134 14959 8186
rect 14971 8134 15023 8186
rect 15035 8134 15087 8186
rect 1584 8075 1636 8084
rect 1584 8041 1593 8075
rect 1593 8041 1627 8075
rect 1627 8041 1636 8075
rect 1584 8032 1636 8041
rect 1952 8032 2004 8084
rect 1400 7939 1452 7948
rect 1400 7905 1409 7939
rect 1409 7905 1443 7939
rect 1443 7905 1452 7939
rect 1400 7896 1452 7905
rect 7656 8032 7708 8084
rect 9312 8075 9364 8084
rect 9312 8041 9321 8075
rect 9321 8041 9355 8075
rect 9355 8041 9364 8075
rect 9312 8032 9364 8041
rect 9772 8075 9824 8084
rect 9772 8041 9781 8075
rect 9781 8041 9815 8075
rect 9815 8041 9824 8075
rect 9772 8032 9824 8041
rect 4344 7964 4396 8016
rect 5172 8007 5224 8016
rect 5172 7973 5190 8007
rect 5190 7973 5224 8007
rect 5172 7964 5224 7973
rect 5448 7964 5500 8016
rect 7748 7964 7800 8016
rect 3608 7896 3660 7948
rect 4896 7896 4948 7948
rect 4436 7828 4488 7880
rect 8208 7896 8260 7948
rect 8852 7896 8904 7948
rect 4252 7692 4304 7744
rect 8392 7692 8444 7744
rect 4447 7590 4499 7642
rect 4511 7590 4563 7642
rect 4575 7590 4627 7642
rect 4639 7590 4691 7642
rect 11378 7590 11430 7642
rect 11442 7590 11494 7642
rect 11506 7590 11558 7642
rect 11570 7590 11622 7642
rect 18308 7590 18360 7642
rect 18372 7590 18424 7642
rect 18436 7590 18488 7642
rect 18500 7590 18552 7642
rect 3608 7531 3660 7540
rect 3608 7497 3617 7531
rect 3617 7497 3651 7531
rect 3651 7497 3660 7531
rect 3608 7488 3660 7497
rect 3700 7488 3752 7540
rect 8852 7531 8904 7540
rect 8852 7497 8861 7531
rect 8861 7497 8895 7531
rect 8895 7497 8904 7531
rect 8852 7488 8904 7497
rect 18880 7488 18932 7540
rect 19708 7488 19760 7540
rect 6920 7420 6972 7472
rect 7196 7420 7248 7472
rect 17224 7420 17276 7472
rect 4252 7395 4304 7404
rect 4252 7361 4261 7395
rect 4261 7361 4295 7395
rect 4295 7361 4304 7395
rect 4252 7352 4304 7361
rect 5172 7395 5224 7404
rect 5172 7361 5181 7395
rect 5181 7361 5215 7395
rect 5215 7361 5224 7395
rect 5172 7352 5224 7361
rect 8392 7352 8444 7404
rect 1400 7327 1452 7336
rect 1400 7293 1409 7327
rect 1409 7293 1443 7327
rect 1443 7293 1452 7327
rect 1400 7284 1452 7293
rect 1860 7327 1912 7336
rect 1860 7293 1869 7327
rect 1869 7293 1903 7327
rect 1903 7293 1912 7327
rect 1860 7284 1912 7293
rect 4988 7284 5040 7336
rect 7564 7284 7616 7336
rect 9404 7284 9456 7336
rect 18788 7327 18840 7336
rect 18788 7293 18797 7327
rect 18797 7293 18831 7327
rect 18831 7293 18840 7327
rect 18788 7284 18840 7293
rect 19064 7327 19116 7336
rect 19064 7293 19073 7327
rect 19073 7293 19107 7327
rect 19107 7293 19116 7327
rect 19064 7284 19116 7293
rect 1584 7191 1636 7200
rect 1584 7157 1593 7191
rect 1593 7157 1627 7191
rect 1627 7157 1636 7191
rect 1584 7148 1636 7157
rect 3240 7191 3292 7200
rect 3240 7157 3249 7191
rect 3249 7157 3283 7191
rect 3283 7157 3292 7191
rect 3240 7148 3292 7157
rect 4068 7191 4120 7200
rect 4068 7157 4077 7191
rect 4077 7157 4111 7191
rect 4111 7157 4120 7191
rect 4068 7148 4120 7157
rect 4712 7148 4764 7200
rect 4896 7148 4948 7200
rect 5172 7148 5224 7200
rect 5448 7148 5500 7200
rect 7748 7148 7800 7200
rect 8484 7191 8536 7200
rect 8484 7157 8493 7191
rect 8493 7157 8527 7191
rect 8527 7157 8536 7191
rect 8484 7148 8536 7157
rect 7912 7046 7964 7098
rect 7976 7046 8028 7098
rect 8040 7046 8092 7098
rect 8104 7046 8156 7098
rect 14843 7046 14895 7098
rect 14907 7046 14959 7098
rect 14971 7046 15023 7098
rect 15035 7046 15087 7098
rect 4344 6987 4396 6996
rect 4344 6953 4353 6987
rect 4353 6953 4387 6987
rect 4387 6953 4396 6987
rect 4344 6944 4396 6953
rect 4712 6987 4764 6996
rect 4712 6953 4721 6987
rect 4721 6953 4755 6987
rect 4755 6953 4764 6987
rect 4712 6944 4764 6953
rect 4896 6944 4948 6996
rect 7564 6944 7616 6996
rect 7748 6987 7800 6996
rect 7748 6953 7757 6987
rect 7757 6953 7791 6987
rect 7791 6953 7800 6987
rect 7748 6944 7800 6953
rect 3240 6876 3292 6928
rect 5172 6876 5224 6928
rect 5724 6876 5776 6928
rect 1400 6851 1452 6860
rect 1400 6817 1409 6851
rect 1409 6817 1443 6851
rect 1443 6817 1452 6851
rect 1400 6808 1452 6817
rect 4804 6851 4856 6860
rect 4804 6817 4813 6851
rect 4813 6817 4847 6851
rect 4847 6817 4856 6851
rect 4804 6808 4856 6817
rect 19800 6851 19852 6860
rect 19800 6817 19809 6851
rect 19809 6817 19843 6851
rect 19843 6817 19852 6851
rect 19800 6808 19852 6817
rect 4252 6740 4304 6792
rect 8208 6740 8260 6792
rect 7288 6715 7340 6724
rect 3976 6647 4028 6656
rect 3976 6613 3985 6647
rect 3985 6613 4019 6647
rect 4019 6613 4028 6647
rect 3976 6604 4028 6613
rect 4896 6604 4948 6656
rect 7288 6681 7297 6715
rect 7297 6681 7331 6715
rect 7331 6681 7340 6715
rect 7288 6672 7340 6681
rect 19984 6715 20036 6724
rect 19984 6681 19993 6715
rect 19993 6681 20027 6715
rect 20027 6681 20036 6715
rect 19984 6672 20036 6681
rect 19064 6604 19116 6656
rect 4447 6502 4499 6554
rect 4511 6502 4563 6554
rect 4575 6502 4627 6554
rect 4639 6502 4691 6554
rect 11378 6502 11430 6554
rect 11442 6502 11494 6554
rect 11506 6502 11558 6554
rect 11570 6502 11622 6554
rect 18308 6502 18360 6554
rect 18372 6502 18424 6554
rect 18436 6502 18488 6554
rect 18500 6502 18552 6554
rect 19892 6400 19944 6452
rect 1400 6239 1452 6248
rect 1400 6205 1409 6239
rect 1409 6205 1443 6239
rect 1443 6205 1452 6239
rect 1400 6196 1452 6205
rect 20076 6239 20128 6248
rect 20076 6205 20085 6239
rect 20085 6205 20119 6239
rect 20119 6205 20128 6239
rect 20076 6196 20128 6205
rect 1584 6103 1636 6112
rect 1584 6069 1593 6103
rect 1593 6069 1627 6103
rect 1627 6069 1636 6103
rect 1584 6060 1636 6069
rect 7912 5958 7964 6010
rect 7976 5958 8028 6010
rect 8040 5958 8092 6010
rect 8104 5958 8156 6010
rect 14843 5958 14895 6010
rect 14907 5958 14959 6010
rect 14971 5958 15023 6010
rect 15035 5958 15087 6010
rect 1584 5856 1636 5908
rect 19800 5856 19852 5908
rect 20536 5899 20588 5908
rect 20536 5865 20545 5899
rect 20545 5865 20579 5899
rect 20579 5865 20588 5899
rect 20536 5856 20588 5865
rect 1400 5763 1452 5772
rect 1400 5729 1409 5763
rect 1409 5729 1443 5763
rect 1443 5729 1452 5763
rect 1400 5720 1452 5729
rect 1676 5652 1728 5704
rect 20076 5584 20128 5636
rect 4447 5414 4499 5466
rect 4511 5414 4563 5466
rect 4575 5414 4627 5466
rect 4639 5414 4691 5466
rect 11378 5414 11430 5466
rect 11442 5414 11494 5466
rect 11506 5414 11558 5466
rect 11570 5414 11622 5466
rect 18308 5414 18360 5466
rect 18372 5414 18424 5466
rect 18436 5414 18488 5466
rect 18500 5414 18552 5466
rect 1676 5312 1728 5364
rect 20812 5355 20864 5364
rect 20812 5321 20821 5355
rect 20821 5321 20855 5355
rect 20855 5321 20864 5355
rect 20812 5312 20864 5321
rect 1400 5151 1452 5160
rect 1400 5117 1409 5151
rect 1409 5117 1443 5151
rect 1443 5117 1452 5151
rect 1400 5108 1452 5117
rect 20996 5151 21048 5160
rect 20996 5117 21005 5151
rect 21005 5117 21039 5151
rect 21039 5117 21048 5151
rect 20996 5108 21048 5117
rect 1860 5015 1912 5024
rect 1860 4981 1869 5015
rect 1869 4981 1903 5015
rect 1903 4981 1912 5015
rect 1860 4972 1912 4981
rect 7912 4870 7964 4922
rect 7976 4870 8028 4922
rect 8040 4870 8092 4922
rect 8104 4870 8156 4922
rect 14843 4870 14895 4922
rect 14907 4870 14959 4922
rect 14971 4870 15023 4922
rect 15035 4870 15087 4922
rect 1400 4675 1452 4684
rect 1400 4641 1409 4675
rect 1409 4641 1443 4675
rect 1443 4641 1452 4675
rect 1400 4632 1452 4641
rect 1860 4675 1912 4684
rect 1860 4641 1869 4675
rect 1869 4641 1903 4675
rect 1903 4641 1912 4675
rect 1860 4632 1912 4641
rect 11152 4564 11204 4616
rect 20996 4428 21048 4480
rect 4447 4326 4499 4378
rect 4511 4326 4563 4378
rect 4575 4326 4627 4378
rect 4639 4326 4691 4378
rect 11378 4326 11430 4378
rect 11442 4326 11494 4378
rect 11506 4326 11558 4378
rect 11570 4326 11622 4378
rect 18308 4326 18360 4378
rect 18372 4326 18424 4378
rect 18436 4326 18488 4378
rect 18500 4326 18552 4378
rect 4988 4088 5040 4140
rect 1676 3995 1728 4004
rect 1676 3961 1685 3995
rect 1685 3961 1719 3995
rect 1719 3961 1728 3995
rect 1676 3952 1728 3961
rect 1768 3884 1820 3936
rect 7912 3782 7964 3834
rect 7976 3782 8028 3834
rect 8040 3782 8092 3834
rect 8104 3782 8156 3834
rect 14843 3782 14895 3834
rect 14907 3782 14959 3834
rect 14971 3782 15023 3834
rect 15035 3782 15087 3834
rect 4068 3680 4120 3732
rect 3240 3612 3292 3664
rect 1676 3587 1728 3596
rect 1676 3553 1685 3587
rect 1685 3553 1719 3587
rect 1719 3553 1728 3587
rect 1676 3544 1728 3553
rect 3148 3544 3200 3596
rect 3148 3383 3200 3392
rect 3148 3349 3157 3383
rect 3157 3349 3191 3383
rect 3191 3349 3200 3383
rect 3148 3340 3200 3349
rect 4447 3238 4499 3290
rect 4511 3238 4563 3290
rect 4575 3238 4627 3290
rect 4639 3238 4691 3290
rect 11378 3238 11430 3290
rect 11442 3238 11494 3290
rect 11506 3238 11558 3290
rect 11570 3238 11622 3290
rect 18308 3238 18360 3290
rect 18372 3238 18424 3290
rect 18436 3238 18488 3290
rect 18500 3238 18552 3290
rect 3424 3136 3476 3188
rect 2596 3068 2648 3120
rect 2136 3000 2188 3052
rect 3884 3068 3936 3120
rect 1768 2975 1820 2984
rect 1768 2941 1777 2975
rect 1777 2941 1811 2975
rect 1811 2941 1820 2975
rect 1768 2932 1820 2941
rect 2228 2907 2280 2916
rect 2228 2873 2237 2907
rect 2237 2873 2271 2907
rect 2271 2873 2280 2907
rect 2228 2864 2280 2873
rect 3884 2864 3936 2916
rect 7912 2694 7964 2746
rect 7976 2694 8028 2746
rect 8040 2694 8092 2746
rect 8104 2694 8156 2746
rect 14843 2694 14895 2746
rect 14907 2694 14959 2746
rect 14971 2694 15023 2746
rect 15035 2694 15087 2746
rect 4344 2592 4396 2644
rect 5448 2524 5500 2576
rect 12256 2567 12308 2576
rect 12256 2533 12265 2567
rect 12265 2533 12299 2567
rect 12299 2533 12308 2567
rect 12256 2524 12308 2533
rect 1676 2499 1728 2508
rect 1676 2465 1685 2499
rect 1685 2465 1719 2499
rect 1719 2465 1728 2499
rect 1676 2456 1728 2465
rect 2136 2456 2188 2508
rect 2780 2499 2832 2508
rect 2780 2465 2789 2499
rect 2789 2465 2823 2499
rect 2823 2465 2832 2499
rect 2780 2456 2832 2465
rect 3976 2320 4028 2372
rect 11704 2320 11756 2372
rect 4447 2150 4499 2202
rect 4511 2150 4563 2202
rect 4575 2150 4627 2202
rect 4639 2150 4691 2202
rect 11378 2150 11430 2202
rect 11442 2150 11494 2202
rect 11506 2150 11558 2202
rect 11570 2150 11622 2202
rect 18308 2150 18360 2202
rect 18372 2150 18424 2202
rect 18436 2150 18488 2202
rect 18500 2150 18552 2202
<< metal2 >>
rect 202 22200 258 23000
rect 662 22200 718 23000
rect 1122 22200 1178 23000
rect 1582 22200 1638 23000
rect 2042 22200 2098 23000
rect 2502 22200 2558 23000
rect 2962 22200 3018 23000
rect 3422 22200 3478 23000
rect 3882 22200 3938 23000
rect 3974 22672 4030 22681
rect 3974 22607 4030 22616
rect 216 20398 244 22200
rect 204 20392 256 20398
rect 204 20334 256 20340
rect 676 20330 704 22200
rect 664 20324 716 20330
rect 664 20266 716 20272
rect 1136 20262 1164 22200
rect 1596 20466 1624 22200
rect 1584 20460 1636 20466
rect 1584 20402 1636 20408
rect 1308 20392 1360 20398
rect 1308 20334 1360 20340
rect 1124 20256 1176 20262
rect 1124 20198 1176 20204
rect 1320 19990 1348 20334
rect 2056 20074 2084 22200
rect 2228 20324 2280 20330
rect 2228 20266 2280 20272
rect 1964 20046 2084 20074
rect 1308 19984 1360 19990
rect 1308 19926 1360 19932
rect 1582 19816 1638 19825
rect 1582 19751 1584 19760
rect 1636 19751 1638 19760
rect 1584 19722 1636 19728
rect 1582 19408 1638 19417
rect 1582 19343 1638 19352
rect 1596 19310 1624 19343
rect 1584 19304 1636 19310
rect 1584 19246 1636 19252
rect 1582 18864 1638 18873
rect 1582 18799 1584 18808
rect 1636 18799 1638 18808
rect 1584 18770 1636 18776
rect 1674 18456 1730 18465
rect 1674 18391 1676 18400
rect 1728 18391 1730 18400
rect 1676 18362 1728 18368
rect 1964 18086 1992 20046
rect 2044 19916 2096 19922
rect 2044 19858 2096 19864
rect 1952 18080 2004 18086
rect 1952 18022 2004 18028
rect 1582 17096 1638 17105
rect 1582 17031 1584 17040
rect 1636 17031 1638 17040
rect 1768 17060 1820 17066
rect 1584 17002 1636 17008
rect 1768 17002 1820 17008
rect 1780 16794 1808 17002
rect 1768 16788 1820 16794
rect 1768 16730 1820 16736
rect 1584 16652 1636 16658
rect 1584 16594 1636 16600
rect 1768 16652 1820 16658
rect 1768 16594 1820 16600
rect 1596 16561 1624 16594
rect 1582 16552 1638 16561
rect 1582 16487 1638 16496
rect 1780 16250 1808 16594
rect 1768 16244 1820 16250
rect 1768 16186 1820 16192
rect 1582 16144 1638 16153
rect 1582 16079 1584 16088
rect 1636 16079 1638 16088
rect 1584 16050 1636 16056
rect 1768 15972 1820 15978
rect 1768 15914 1820 15920
rect 1582 15600 1638 15609
rect 1582 15535 1584 15544
rect 1636 15535 1638 15544
rect 1584 15506 1636 15512
rect 1674 15192 1730 15201
rect 1780 15162 1808 15914
rect 1860 15564 1912 15570
rect 1860 15506 1912 15512
rect 1674 15127 1676 15136
rect 1728 15127 1730 15136
rect 1768 15156 1820 15162
rect 1676 15098 1728 15104
rect 1768 15098 1820 15104
rect 1768 14884 1820 14890
rect 1768 14826 1820 14832
rect 1676 14272 1728 14278
rect 1674 14240 1676 14249
rect 1728 14240 1730 14249
rect 1674 14175 1730 14184
rect 1780 13954 1808 14826
rect 1688 13926 1808 13954
rect 1584 13864 1636 13870
rect 1582 13832 1584 13841
rect 1636 13832 1638 13841
rect 1582 13767 1638 13776
rect 1492 13388 1544 13394
rect 1492 13330 1544 13336
rect 1504 12986 1532 13330
rect 1492 12980 1544 12986
rect 1492 12922 1544 12928
rect 1400 11552 1452 11558
rect 1400 11494 1452 11500
rect 1412 11218 1440 11494
rect 1504 11393 1532 12922
rect 1688 11898 1716 13926
rect 1768 13864 1820 13870
rect 1768 13806 1820 13812
rect 1780 12442 1808 13806
rect 1872 12986 1900 15506
rect 1952 14476 2004 14482
rect 1952 14418 2004 14424
rect 1860 12980 1912 12986
rect 1860 12922 1912 12928
rect 1768 12436 1820 12442
rect 1768 12378 1820 12384
rect 1676 11892 1728 11898
rect 1676 11834 1728 11840
rect 1860 11688 1912 11694
rect 1860 11630 1912 11636
rect 1490 11384 1546 11393
rect 1872 11354 1900 11630
rect 1490 11319 1546 11328
rect 1860 11348 1912 11354
rect 1860 11290 1912 11296
rect 1400 11212 1452 11218
rect 1400 11154 1452 11160
rect 1412 10577 1440 11154
rect 1398 10568 1454 10577
rect 1398 10503 1454 10512
rect 1400 10464 1452 10470
rect 1400 10406 1452 10412
rect 1412 10130 1440 10406
rect 1400 10124 1452 10130
rect 1400 10066 1452 10072
rect 1584 10124 1636 10130
rect 1584 10066 1636 10072
rect 1412 10033 1440 10066
rect 1398 10024 1454 10033
rect 1398 9959 1454 9968
rect 1400 9512 1452 9518
rect 1400 9454 1452 9460
rect 1412 9110 1440 9454
rect 1400 9104 1452 9110
rect 1398 9072 1400 9081
rect 1452 9072 1454 9081
rect 1398 9007 1454 9016
rect 1400 8288 1452 8294
rect 1400 8230 1452 8236
rect 1412 7954 1440 8230
rect 1596 8090 1624 10066
rect 1860 9512 1912 9518
rect 1858 9480 1860 9489
rect 1912 9480 1914 9489
rect 1858 9415 1914 9424
rect 1872 9178 1900 9415
rect 1860 9172 1912 9178
rect 1860 9114 1912 9120
rect 1964 8634 1992 14418
rect 2056 14074 2084 19858
rect 2240 19446 2268 20266
rect 2516 19922 2544 22200
rect 2976 21842 3004 22200
rect 2976 21814 3372 21842
rect 2962 21720 3018 21729
rect 2962 21655 3018 21664
rect 2870 20768 2926 20777
rect 2870 20703 2926 20712
rect 2780 20528 2832 20534
rect 2778 20496 2780 20505
rect 2832 20496 2834 20505
rect 2778 20431 2834 20440
rect 2778 20360 2834 20369
rect 2778 20295 2834 20304
rect 2504 19916 2556 19922
rect 2504 19858 2556 19864
rect 2228 19440 2280 19446
rect 2228 19382 2280 19388
rect 2228 19236 2280 19242
rect 2228 19178 2280 19184
rect 2136 18828 2188 18834
rect 2136 18770 2188 18776
rect 2148 15706 2176 18770
rect 2240 17626 2268 19178
rect 2412 19168 2464 19174
rect 2412 19110 2464 19116
rect 2320 18692 2372 18698
rect 2320 18634 2372 18640
rect 2332 18222 2360 18634
rect 2320 18216 2372 18222
rect 2320 18158 2372 18164
rect 2240 17598 2360 17626
rect 2228 17536 2280 17542
rect 2226 17504 2228 17513
rect 2280 17504 2282 17513
rect 2226 17439 2282 17448
rect 2332 16250 2360 17598
rect 2320 16244 2372 16250
rect 2320 16186 2372 16192
rect 2320 16040 2372 16046
rect 2320 15982 2372 15988
rect 2136 15700 2188 15706
rect 2136 15642 2188 15648
rect 2332 15434 2360 15982
rect 2320 15428 2372 15434
rect 2320 15370 2372 15376
rect 2320 14952 2372 14958
rect 2320 14894 2372 14900
rect 2226 14648 2282 14657
rect 2226 14583 2228 14592
rect 2280 14583 2282 14592
rect 2228 14554 2280 14560
rect 2228 14476 2280 14482
rect 2228 14418 2280 14424
rect 2044 14068 2096 14074
rect 2044 14010 2096 14016
rect 2240 12434 2268 14418
rect 2332 14074 2360 14894
rect 2320 14068 2372 14074
rect 2320 14010 2372 14016
rect 2320 13864 2372 13870
rect 2320 13806 2372 13812
rect 2332 13530 2360 13806
rect 2320 13524 2372 13530
rect 2320 13466 2372 13472
rect 2424 12986 2452 19110
rect 2516 18737 2544 19858
rect 2792 19310 2820 20295
rect 2780 19304 2832 19310
rect 2780 19246 2832 19252
rect 2884 18970 2912 20703
rect 2872 18964 2924 18970
rect 2872 18906 2924 18912
rect 2502 18728 2558 18737
rect 2976 18714 3004 21655
rect 3054 21312 3110 21321
rect 3054 21247 3110 21256
rect 2502 18663 2558 18672
rect 2884 18686 3004 18714
rect 2688 18624 2740 18630
rect 2688 18566 2740 18572
rect 2504 18148 2556 18154
rect 2504 18090 2556 18096
rect 2516 16794 2544 18090
rect 2700 17814 2728 18566
rect 2778 18048 2834 18057
rect 2778 17983 2834 17992
rect 2688 17808 2740 17814
rect 2688 17750 2740 17756
rect 2688 17604 2740 17610
rect 2688 17546 2740 17552
rect 2504 16788 2556 16794
rect 2504 16730 2556 16736
rect 2596 15564 2648 15570
rect 2596 15506 2648 15512
rect 2608 13530 2636 15506
rect 2596 13524 2648 13530
rect 2596 13466 2648 13472
rect 2700 13172 2728 17546
rect 2792 17338 2820 17983
rect 2884 17814 2912 18686
rect 2964 18624 3016 18630
rect 2964 18566 3016 18572
rect 2872 17808 2924 17814
rect 2872 17750 2924 17756
rect 2872 17672 2924 17678
rect 2872 17614 2924 17620
rect 2780 17332 2832 17338
rect 2780 17274 2832 17280
rect 2884 16998 2912 17614
rect 2976 17134 3004 18566
rect 3068 18426 3096 21247
rect 3148 19780 3200 19786
rect 3148 19722 3200 19728
rect 3160 19174 3188 19722
rect 3148 19168 3200 19174
rect 3148 19110 3200 19116
rect 3056 18420 3108 18426
rect 3056 18362 3108 18368
rect 3160 18222 3188 19110
rect 3148 18216 3200 18222
rect 3344 18193 3372 21814
rect 3436 20482 3464 22200
rect 3436 20454 3740 20482
rect 3608 20392 3660 20398
rect 3608 20334 3660 20340
rect 3424 20256 3476 20262
rect 3424 20198 3476 20204
rect 3436 19514 3464 20198
rect 3424 19508 3476 19514
rect 3424 19450 3476 19456
rect 3620 18222 3648 20334
rect 3712 20330 3740 20454
rect 3700 20324 3752 20330
rect 3700 20266 3752 20272
rect 3896 19394 3924 22200
rect 3988 20874 4016 22607
rect 4066 22264 4122 22273
rect 4066 22199 4122 22208
rect 4342 22200 4398 23000
rect 4802 22200 4858 23000
rect 5262 22200 5318 23000
rect 5722 22200 5778 23000
rect 6182 22200 6238 23000
rect 6642 22200 6698 23000
rect 7102 22200 7158 23000
rect 7562 22200 7618 23000
rect 8022 22200 8078 23000
rect 8482 22200 8538 23000
rect 8942 22200 8998 23000
rect 9402 22200 9458 23000
rect 9862 22200 9918 23000
rect 10322 22200 10378 23000
rect 10782 22200 10838 23000
rect 11242 22200 11298 23000
rect 11702 22200 11758 23000
rect 12162 22200 12218 23000
rect 12622 22200 12678 23000
rect 13082 22200 13138 23000
rect 13542 22200 13598 23000
rect 14002 22200 14058 23000
rect 14462 22200 14518 23000
rect 14922 22200 14978 23000
rect 15382 22200 15438 23000
rect 15842 22200 15898 23000
rect 16302 22200 16358 23000
rect 16762 22200 16818 23000
rect 17222 22200 17278 23000
rect 17682 22200 17738 23000
rect 18142 22200 18198 23000
rect 18602 22200 18658 23000
rect 19062 22200 19118 23000
rect 19522 22200 19578 23000
rect 19982 22200 20038 23000
rect 20442 22200 20498 23000
rect 20902 22200 20958 23000
rect 21362 22200 21418 23000
rect 21822 22200 21878 23000
rect 22282 22200 22338 23000
rect 22742 22200 22798 23000
rect 3976 20868 4028 20874
rect 3976 20810 4028 20816
rect 4080 20806 4108 22199
rect 4068 20800 4120 20806
rect 4068 20742 4120 20748
rect 4356 20584 4384 22200
rect 4421 20700 4717 20720
rect 4477 20698 4501 20700
rect 4557 20698 4581 20700
rect 4637 20698 4661 20700
rect 4499 20646 4501 20698
rect 4563 20646 4575 20698
rect 4637 20646 4639 20698
rect 4477 20644 4501 20646
rect 4557 20644 4581 20646
rect 4637 20644 4661 20646
rect 4421 20624 4717 20644
rect 4816 20618 4844 22200
rect 4816 20590 4936 20618
rect 4356 20556 4476 20584
rect 4158 20496 4214 20505
rect 4158 20431 4160 20440
rect 4212 20431 4214 20440
rect 4160 20402 4212 20408
rect 4252 20392 4304 20398
rect 4448 20380 4476 20556
rect 4252 20334 4304 20340
rect 4356 20352 4476 20380
rect 4068 20256 4120 20262
rect 4068 20198 4120 20204
rect 4080 20058 4108 20198
rect 4068 20052 4120 20058
rect 4068 19994 4120 20000
rect 4264 19514 4292 20334
rect 4252 19508 4304 19514
rect 4252 19450 4304 19456
rect 3896 19366 4200 19394
rect 4068 19304 4120 19310
rect 4066 19272 4068 19281
rect 4120 19272 4122 19281
rect 4066 19207 4122 19216
rect 4172 19156 4200 19366
rect 4356 19258 4384 20352
rect 4620 20256 4672 20262
rect 4620 20198 4672 20204
rect 4632 20097 4660 20198
rect 4618 20088 4674 20097
rect 4618 20023 4674 20032
rect 4421 19612 4717 19632
rect 4477 19610 4501 19612
rect 4557 19610 4581 19612
rect 4637 19610 4661 19612
rect 4499 19558 4501 19610
rect 4563 19558 4575 19610
rect 4637 19558 4639 19610
rect 4477 19556 4501 19558
rect 4557 19556 4581 19558
rect 4637 19556 4661 19558
rect 4421 19536 4717 19556
rect 4356 19230 4568 19258
rect 4436 19168 4488 19174
rect 4172 19128 4436 19156
rect 4436 19110 4488 19116
rect 4540 18970 4568 19230
rect 4528 18964 4580 18970
rect 4528 18906 4580 18912
rect 4068 18828 4120 18834
rect 4068 18770 4120 18776
rect 4252 18828 4304 18834
rect 4252 18770 4304 18776
rect 4080 18358 4108 18770
rect 4068 18352 4120 18358
rect 4068 18294 4120 18300
rect 3608 18216 3660 18222
rect 3148 18158 3200 18164
rect 3330 18184 3386 18193
rect 3608 18158 3660 18164
rect 3330 18119 3386 18128
rect 3884 18148 3936 18154
rect 3884 18090 3936 18096
rect 3148 17740 3200 17746
rect 3148 17682 3200 17688
rect 2964 17128 3016 17134
rect 2964 17070 3016 17076
rect 2872 16992 2924 16998
rect 2872 16934 2924 16940
rect 2780 16516 2832 16522
rect 2780 16458 2832 16464
rect 2792 15366 2820 16458
rect 2780 15360 2832 15366
rect 2780 15302 2832 15308
rect 2884 14958 2912 16934
rect 3160 16794 3188 17682
rect 3896 17116 3924 18090
rect 4160 18080 4212 18086
rect 4160 18022 4212 18028
rect 4172 17202 4200 18022
rect 4160 17196 4212 17202
rect 4160 17138 4212 17144
rect 4068 17128 4120 17134
rect 3896 17088 4068 17116
rect 4068 17070 4120 17076
rect 3332 16992 3384 16998
rect 3332 16934 3384 16940
rect 3148 16788 3200 16794
rect 3148 16730 3200 16736
rect 3056 16720 3108 16726
rect 3056 16662 3108 16668
rect 3068 16250 3096 16662
rect 3056 16244 3108 16250
rect 3056 16186 3108 16192
rect 2872 14952 2924 14958
rect 2872 14894 2924 14900
rect 3148 14476 3200 14482
rect 3148 14418 3200 14424
rect 2780 14272 2832 14278
rect 2780 14214 2832 14220
rect 2792 13394 2820 14214
rect 3160 13938 3188 14418
rect 3148 13932 3200 13938
rect 3148 13874 3200 13880
rect 3148 13456 3200 13462
rect 3148 13398 3200 13404
rect 2780 13388 2832 13394
rect 2780 13330 2832 13336
rect 2872 13388 2924 13394
rect 2872 13330 2924 13336
rect 2516 13144 2728 13172
rect 2412 12980 2464 12986
rect 2412 12922 2464 12928
rect 2516 12866 2544 13144
rect 2148 12406 2268 12434
rect 2332 12838 2544 12866
rect 2044 12300 2096 12306
rect 2044 12242 2096 12248
rect 2056 11898 2084 12242
rect 2044 11892 2096 11898
rect 2044 11834 2096 11840
rect 2044 10668 2096 10674
rect 2044 10610 2096 10616
rect 2056 9926 2084 10610
rect 2044 9920 2096 9926
rect 2044 9862 2096 9868
rect 1952 8628 2004 8634
rect 1952 8570 2004 8576
rect 1952 8424 2004 8430
rect 1952 8366 2004 8372
rect 1858 8120 1914 8129
rect 1584 8084 1636 8090
rect 1964 8090 1992 8366
rect 2056 8362 2084 9862
rect 2148 8906 2176 12406
rect 2332 9654 2360 12838
rect 2412 12776 2464 12782
rect 2412 12718 2464 12724
rect 2596 12776 2648 12782
rect 2596 12718 2648 12724
rect 2424 12442 2452 12718
rect 2412 12436 2464 12442
rect 2412 12378 2464 12384
rect 2504 12300 2556 12306
rect 2504 12242 2556 12248
rect 2516 11898 2544 12242
rect 2504 11892 2556 11898
rect 2504 11834 2556 11840
rect 2504 11688 2556 11694
rect 2504 11630 2556 11636
rect 2412 11008 2464 11014
rect 2412 10950 2464 10956
rect 2424 10606 2452 10950
rect 2516 10810 2544 11630
rect 2504 10804 2556 10810
rect 2504 10746 2556 10752
rect 2412 10600 2464 10606
rect 2412 10542 2464 10548
rect 2608 10266 2636 12718
rect 2688 12708 2740 12714
rect 2688 12650 2740 12656
rect 2700 12442 2728 12650
rect 2688 12436 2740 12442
rect 2688 12378 2740 12384
rect 2884 12345 2912 13330
rect 2964 12640 3016 12646
rect 2964 12582 3016 12588
rect 2870 12336 2926 12345
rect 2870 12271 2926 12280
rect 2976 12238 3004 12582
rect 3160 12306 3188 13398
rect 3148 12300 3200 12306
rect 3148 12242 3200 12248
rect 2964 12232 3016 12238
rect 2964 12174 3016 12180
rect 3160 11937 3188 12242
rect 3344 12170 3372 16934
rect 3516 16652 3568 16658
rect 3516 16594 3568 16600
rect 3528 16250 3556 16594
rect 3516 16244 3568 16250
rect 3516 16186 3568 16192
rect 4080 16017 4108 17070
rect 4172 17066 4200 17138
rect 4160 17060 4212 17066
rect 4160 17002 4212 17008
rect 4264 16794 4292 18770
rect 4421 18524 4717 18544
rect 4477 18522 4501 18524
rect 4557 18522 4581 18524
rect 4637 18522 4661 18524
rect 4499 18470 4501 18522
rect 4563 18470 4575 18522
rect 4637 18470 4639 18522
rect 4477 18468 4501 18470
rect 4557 18468 4581 18470
rect 4637 18468 4661 18470
rect 4421 18448 4717 18468
rect 4908 18426 4936 20590
rect 4988 20392 5040 20398
rect 4988 20334 5040 20340
rect 4896 18420 4948 18426
rect 4896 18362 4948 18368
rect 4804 18284 4856 18290
rect 4804 18226 4856 18232
rect 4816 17882 4844 18226
rect 5000 18170 5028 20334
rect 5080 20256 5132 20262
rect 5080 20198 5132 20204
rect 5092 19990 5120 20198
rect 5080 19984 5132 19990
rect 5080 19926 5132 19932
rect 5172 19712 5224 19718
rect 5172 19654 5224 19660
rect 5184 19514 5212 19654
rect 5172 19508 5224 19514
rect 5172 19450 5224 19456
rect 5078 19272 5134 19281
rect 5078 19207 5134 19216
rect 5092 18834 5120 19207
rect 5276 18952 5304 22200
rect 5448 20256 5500 20262
rect 5448 20198 5500 20204
rect 5460 20058 5488 20198
rect 5448 20052 5500 20058
rect 5448 19994 5500 20000
rect 5354 19816 5410 19825
rect 5354 19751 5356 19760
rect 5408 19751 5410 19760
rect 5540 19780 5592 19786
rect 5356 19722 5408 19728
rect 5540 19722 5592 19728
rect 5552 19310 5580 19722
rect 5540 19304 5592 19310
rect 5540 19246 5592 19252
rect 5276 18924 5488 18952
rect 5080 18828 5132 18834
rect 5080 18770 5132 18776
rect 5264 18828 5316 18834
rect 5264 18770 5316 18776
rect 5092 18601 5120 18770
rect 5078 18592 5134 18601
rect 5078 18527 5134 18536
rect 5276 18290 5304 18770
rect 5460 18290 5488 18924
rect 5736 18834 5764 22200
rect 5814 20632 5870 20641
rect 5814 20567 5870 20576
rect 5828 20262 5856 20567
rect 6092 20460 6144 20466
rect 6092 20402 6144 20408
rect 5816 20256 5868 20262
rect 5816 20198 5868 20204
rect 5724 18828 5776 18834
rect 5724 18770 5776 18776
rect 5828 18306 5856 20198
rect 6000 20052 6052 20058
rect 6000 19994 6052 20000
rect 5908 18964 5960 18970
rect 5908 18906 5960 18912
rect 5264 18284 5316 18290
rect 5264 18226 5316 18232
rect 5448 18284 5500 18290
rect 5448 18226 5500 18232
rect 5736 18278 5856 18306
rect 4896 18148 4948 18154
rect 5000 18142 5120 18170
rect 4896 18090 4948 18096
rect 4908 17882 4936 18090
rect 4988 18080 5040 18086
rect 4988 18022 5040 18028
rect 4804 17876 4856 17882
rect 4804 17818 4856 17824
rect 4896 17876 4948 17882
rect 4896 17818 4948 17824
rect 4344 17672 4396 17678
rect 4344 17614 4396 17620
rect 4356 17338 4384 17614
rect 4421 17436 4717 17456
rect 4477 17434 4501 17436
rect 4557 17434 4581 17436
rect 4637 17434 4661 17436
rect 4499 17382 4501 17434
rect 4563 17382 4575 17434
rect 4637 17382 4639 17434
rect 4477 17380 4501 17382
rect 4557 17380 4581 17382
rect 4637 17380 4661 17382
rect 4421 17360 4717 17380
rect 4344 17332 4396 17338
rect 4344 17274 4396 17280
rect 4252 16788 4304 16794
rect 4252 16730 4304 16736
rect 4896 16788 4948 16794
rect 4896 16730 4948 16736
rect 4160 16448 4212 16454
rect 4160 16390 4212 16396
rect 4172 16046 4200 16390
rect 4421 16348 4717 16368
rect 4477 16346 4501 16348
rect 4557 16346 4581 16348
rect 4637 16346 4661 16348
rect 4499 16294 4501 16346
rect 4563 16294 4575 16346
rect 4637 16294 4639 16346
rect 4477 16292 4501 16294
rect 4557 16292 4581 16294
rect 4637 16292 4661 16294
rect 4421 16272 4717 16292
rect 4160 16040 4212 16046
rect 4066 16008 4122 16017
rect 4620 16040 4672 16046
rect 4160 15982 4212 15988
rect 4618 16008 4620 16017
rect 4672 16008 4674 16017
rect 4066 15943 4122 15952
rect 4618 15943 4674 15952
rect 4080 14890 4108 15943
rect 4421 15260 4717 15280
rect 4477 15258 4501 15260
rect 4557 15258 4581 15260
rect 4637 15258 4661 15260
rect 4499 15206 4501 15258
rect 4563 15206 4575 15258
rect 4637 15206 4639 15258
rect 4477 15204 4501 15206
rect 4557 15204 4581 15206
rect 4637 15204 4661 15206
rect 4421 15184 4717 15204
rect 4344 15020 4396 15026
rect 4344 14962 4396 14968
rect 4068 14884 4120 14890
rect 4068 14826 4120 14832
rect 4080 14414 4108 14826
rect 4252 14816 4304 14822
rect 4252 14758 4304 14764
rect 4264 14618 4292 14758
rect 4252 14612 4304 14618
rect 4252 14554 4304 14560
rect 4356 14550 4384 14962
rect 4908 14958 4936 16730
rect 5000 16658 5028 18022
rect 4988 16652 5040 16658
rect 4988 16594 5040 16600
rect 4988 16244 5040 16250
rect 5092 16232 5120 18142
rect 5264 18080 5316 18086
rect 5264 18022 5316 18028
rect 5540 18080 5592 18086
rect 5540 18022 5592 18028
rect 5276 17338 5304 18022
rect 5552 17814 5580 18022
rect 5540 17808 5592 17814
rect 5540 17750 5592 17756
rect 5632 17808 5684 17814
rect 5632 17750 5684 17756
rect 5264 17332 5316 17338
rect 5264 17274 5316 17280
rect 5448 17264 5500 17270
rect 5448 17206 5500 17212
rect 5172 16652 5224 16658
rect 5172 16594 5224 16600
rect 5040 16204 5120 16232
rect 4988 16186 5040 16192
rect 5184 15162 5212 16594
rect 5264 16584 5316 16590
rect 5264 16526 5316 16532
rect 5356 16584 5408 16590
rect 5356 16526 5408 16532
rect 5276 16046 5304 16526
rect 5264 16040 5316 16046
rect 5264 15982 5316 15988
rect 5276 15706 5304 15982
rect 5368 15978 5396 16526
rect 5356 15972 5408 15978
rect 5356 15914 5408 15920
rect 5264 15700 5316 15706
rect 5264 15642 5316 15648
rect 5172 15156 5224 15162
rect 5172 15098 5224 15104
rect 5264 15088 5316 15094
rect 5264 15030 5316 15036
rect 4896 14952 4948 14958
rect 4896 14894 4948 14900
rect 5276 14822 5304 15030
rect 5264 14816 5316 14822
rect 5264 14758 5316 14764
rect 4344 14544 4396 14550
rect 4344 14486 4396 14492
rect 4068 14408 4120 14414
rect 4068 14350 4120 14356
rect 3608 14272 3660 14278
rect 3608 14214 3660 14220
rect 3620 13870 3648 14214
rect 4421 14172 4717 14192
rect 4477 14170 4501 14172
rect 4557 14170 4581 14172
rect 4637 14170 4661 14172
rect 4499 14118 4501 14170
rect 4563 14118 4575 14170
rect 4637 14118 4639 14170
rect 4477 14116 4501 14118
rect 4557 14116 4581 14118
rect 4637 14116 4661 14118
rect 4421 14096 4717 14116
rect 5078 14104 5134 14113
rect 4344 14068 4396 14074
rect 5078 14039 5134 14048
rect 4344 14010 4396 14016
rect 4356 13977 4384 14010
rect 5092 14006 5120 14039
rect 5080 14000 5132 14006
rect 4342 13968 4398 13977
rect 5080 13942 5132 13948
rect 4342 13903 4398 13912
rect 3608 13864 3660 13870
rect 3608 13806 3660 13812
rect 4068 13864 4120 13870
rect 4068 13806 4120 13812
rect 3620 12889 3648 13806
rect 4080 13297 4108 13806
rect 4066 13288 4122 13297
rect 4066 13223 4122 13232
rect 3606 12880 3662 12889
rect 3606 12815 3662 12824
rect 3884 12300 3936 12306
rect 3884 12242 3936 12248
rect 3332 12164 3384 12170
rect 3332 12106 3384 12112
rect 3146 11928 3202 11937
rect 3146 11863 3202 11872
rect 2870 11656 2926 11665
rect 2870 11591 2926 11600
rect 2884 11558 2912 11591
rect 2872 11552 2924 11558
rect 2872 11494 2924 11500
rect 2780 11212 2832 11218
rect 2780 11154 2832 11160
rect 2596 10260 2648 10266
rect 2596 10202 2648 10208
rect 2320 9648 2372 9654
rect 2320 9590 2372 9596
rect 2792 9586 2820 11154
rect 2872 11144 2924 11150
rect 2872 11086 2924 11092
rect 3056 11144 3108 11150
rect 3056 11086 3108 11092
rect 2884 9654 2912 11086
rect 3068 10810 3096 11086
rect 3344 10826 3372 12106
rect 3896 11762 3924 12242
rect 4080 11898 4108 13223
rect 4421 13084 4717 13104
rect 4477 13082 4501 13084
rect 4557 13082 4581 13084
rect 4637 13082 4661 13084
rect 4499 13030 4501 13082
rect 4563 13030 4575 13082
rect 4637 13030 4639 13082
rect 4477 13028 4501 13030
rect 4557 13028 4581 13030
rect 4637 13028 4661 13030
rect 4421 13008 4717 13028
rect 4712 12912 4764 12918
rect 4712 12854 4764 12860
rect 4724 12374 4752 12854
rect 4804 12776 4856 12782
rect 4804 12718 4856 12724
rect 4712 12368 4764 12374
rect 4712 12310 4764 12316
rect 4816 12306 4844 12718
rect 4896 12708 4948 12714
rect 4896 12650 4948 12656
rect 4804 12300 4856 12306
rect 4804 12242 4856 12248
rect 4816 12102 4844 12242
rect 4252 12096 4304 12102
rect 4252 12038 4304 12044
rect 4804 12096 4856 12102
rect 4804 12038 4856 12044
rect 4908 12084 4936 12650
rect 5276 12434 5304 14758
rect 5276 12406 5396 12434
rect 4988 12096 5040 12102
rect 4908 12056 4988 12084
rect 4068 11892 4120 11898
rect 4068 11834 4120 11840
rect 3884 11756 3936 11762
rect 3884 11698 3936 11704
rect 3424 11688 3476 11694
rect 3424 11630 3476 11636
rect 3436 11354 3464 11630
rect 3424 11348 3476 11354
rect 3424 11290 3476 11296
rect 4160 11348 4212 11354
rect 4160 11290 4212 11296
rect 3436 10985 3464 11290
rect 4068 11144 4120 11150
rect 4068 11086 4120 11092
rect 3422 10976 3478 10985
rect 3422 10911 3478 10920
rect 3056 10804 3108 10810
rect 2976 10764 3056 10792
rect 2976 10130 3004 10764
rect 3344 10798 3464 10826
rect 3056 10746 3108 10752
rect 2964 10124 3016 10130
rect 2964 10066 3016 10072
rect 2872 9648 2924 9654
rect 2872 9590 2924 9596
rect 2780 9580 2832 9586
rect 2780 9522 2832 9528
rect 3436 9382 3464 10798
rect 4080 10538 4108 11086
rect 4068 10532 4120 10538
rect 4068 10474 4120 10480
rect 4080 10062 4108 10474
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 3884 9648 3936 9654
rect 3884 9590 3936 9596
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 2780 9036 2832 9042
rect 2780 8978 2832 8984
rect 2596 8968 2648 8974
rect 2596 8910 2648 8916
rect 2136 8900 2188 8906
rect 2136 8842 2188 8848
rect 2044 8356 2096 8362
rect 2044 8298 2096 8304
rect 1858 8055 1914 8064
rect 1952 8084 2004 8090
rect 1584 8026 1636 8032
rect 1400 7948 1452 7954
rect 1400 7890 1452 7896
rect 1412 7721 1440 7890
rect 1398 7712 1454 7721
rect 1398 7647 1454 7656
rect 1872 7342 1900 8055
rect 1952 8026 2004 8032
rect 1400 7336 1452 7342
rect 1860 7336 1912 7342
rect 1400 7278 1452 7284
rect 1582 7304 1638 7313
rect 1412 7177 1440 7278
rect 1860 7278 1912 7284
rect 1582 7239 1638 7248
rect 1596 7206 1624 7239
rect 1584 7200 1636 7206
rect 1398 7168 1454 7177
rect 1584 7142 1636 7148
rect 1398 7103 1454 7112
rect 1400 6860 1452 6866
rect 1400 6802 1452 6808
rect 1412 6769 1440 6802
rect 1398 6760 1454 6769
rect 1398 6695 1454 6704
rect 1400 6248 1452 6254
rect 1398 6216 1400 6225
rect 1452 6216 1454 6225
rect 1398 6151 1454 6160
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 1596 5914 1624 6054
rect 1584 5908 1636 5914
rect 1584 5850 1636 5856
rect 1398 5808 1454 5817
rect 1398 5743 1400 5752
rect 1452 5743 1454 5752
rect 1400 5714 1452 5720
rect 1676 5704 1728 5710
rect 1676 5646 1728 5652
rect 1688 5370 1716 5646
rect 1676 5364 1728 5370
rect 1676 5306 1728 5312
rect 1398 5264 1454 5273
rect 1398 5199 1454 5208
rect 1412 5166 1440 5199
rect 1400 5160 1452 5166
rect 1400 5102 1452 5108
rect 1860 5024 1912 5030
rect 1860 4966 1912 4972
rect 1872 4865 1900 4966
rect 1858 4856 1914 4865
rect 1858 4791 1914 4800
rect 1872 4690 1900 4791
rect 1400 4684 1452 4690
rect 1400 4626 1452 4632
rect 1860 4684 1912 4690
rect 1860 4626 1912 4632
rect 1412 4457 1440 4626
rect 1398 4448 1454 4457
rect 1398 4383 1454 4392
rect 1676 4004 1728 4010
rect 1676 3946 1728 3952
rect 1688 3913 1716 3946
rect 1768 3936 1820 3942
rect 1674 3904 1730 3913
rect 1768 3878 1820 3884
rect 1674 3839 1730 3848
rect 1676 3596 1728 3602
rect 1676 3538 1728 3544
rect 1688 3505 1716 3538
rect 1674 3496 1730 3505
rect 1674 3431 1730 3440
rect 1780 2990 1808 3878
rect 2608 3126 2636 8910
rect 2792 8673 2820 8978
rect 2778 8664 2834 8673
rect 2778 8599 2834 8608
rect 3436 7426 3464 9318
rect 3608 7948 3660 7954
rect 3608 7890 3660 7896
rect 3620 7546 3648 7890
rect 3608 7540 3660 7546
rect 3608 7482 3660 7488
rect 3700 7540 3752 7546
rect 3700 7482 3752 7488
rect 3712 7426 3740 7482
rect 3896 7449 3924 9590
rect 4080 9586 4108 9998
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 3436 7398 3740 7426
rect 3882 7440 3938 7449
rect 3240 7200 3292 7206
rect 3240 7142 3292 7148
rect 3252 6934 3280 7142
rect 3240 6928 3292 6934
rect 3240 6870 3292 6876
rect 3252 3670 3280 6870
rect 3240 3664 3292 3670
rect 3240 3606 3292 3612
rect 3148 3596 3200 3602
rect 3148 3538 3200 3544
rect 3160 3398 3188 3538
rect 3148 3392 3200 3398
rect 3148 3334 3200 3340
rect 2596 3120 2648 3126
rect 2596 3062 2648 3068
rect 2136 3052 2188 3058
rect 2136 2994 2188 3000
rect 1768 2984 1820 2990
rect 1766 2952 1768 2961
rect 1820 2952 1822 2961
rect 1766 2887 1822 2896
rect 1674 2544 1730 2553
rect 2148 2514 2176 2994
rect 2228 2916 2280 2922
rect 2228 2858 2280 2864
rect 1674 2479 1676 2488
rect 1728 2479 1730 2488
rect 2136 2508 2188 2514
rect 1676 2450 1728 2456
rect 2136 2450 2188 2456
rect 2148 241 2176 2450
rect 2240 649 2268 2858
rect 2780 2508 2832 2514
rect 2780 2450 2832 2456
rect 2792 1057 2820 2450
rect 3160 1601 3188 3334
rect 3436 3194 3464 7398
rect 3882 7375 3938 7384
rect 3424 3188 3476 3194
rect 3424 3130 3476 3136
rect 3896 3126 3924 7375
rect 4080 7206 4108 9318
rect 4068 7200 4120 7206
rect 4068 7142 4120 7148
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 3884 3120 3936 3126
rect 3884 3062 3936 3068
rect 3884 2916 3936 2922
rect 3884 2858 3936 2864
rect 3896 2009 3924 2858
rect 3988 2378 4016 6598
rect 4080 3738 4108 7142
rect 4068 3732 4120 3738
rect 4068 3674 4120 3680
rect 4172 2774 4200 11290
rect 4264 10674 4292 12038
rect 4421 11996 4717 12016
rect 4477 11994 4501 11996
rect 4557 11994 4581 11996
rect 4637 11994 4661 11996
rect 4499 11942 4501 11994
rect 4563 11942 4575 11994
rect 4637 11942 4639 11994
rect 4477 11940 4501 11942
rect 4557 11940 4581 11942
rect 4637 11940 4661 11942
rect 4421 11920 4717 11940
rect 4908 11762 4936 12056
rect 4988 12038 5040 12044
rect 4896 11756 4948 11762
rect 4896 11698 4948 11704
rect 4436 11620 4488 11626
rect 4436 11562 4488 11568
rect 4448 11354 4476 11562
rect 4712 11552 4764 11558
rect 4712 11494 4764 11500
rect 4988 11552 5040 11558
rect 4988 11494 5040 11500
rect 4724 11354 4752 11494
rect 5000 11370 5028 11494
rect 5000 11354 5212 11370
rect 4436 11348 4488 11354
rect 4436 11290 4488 11296
rect 4712 11348 4764 11354
rect 4712 11290 4764 11296
rect 5000 11348 5224 11354
rect 5000 11342 5172 11348
rect 4804 11008 4856 11014
rect 4804 10950 4856 10956
rect 4421 10908 4717 10928
rect 4477 10906 4501 10908
rect 4557 10906 4581 10908
rect 4637 10906 4661 10908
rect 4499 10854 4501 10906
rect 4563 10854 4575 10906
rect 4637 10854 4639 10906
rect 4477 10852 4501 10854
rect 4557 10852 4581 10854
rect 4637 10852 4661 10854
rect 4421 10832 4717 10852
rect 4816 10674 4844 10950
rect 4252 10668 4304 10674
rect 4252 10610 4304 10616
rect 4804 10668 4856 10674
rect 4804 10610 4856 10616
rect 4264 9994 4292 10610
rect 4804 10464 4856 10470
rect 4804 10406 4856 10412
rect 4816 10266 4844 10406
rect 4804 10260 4856 10266
rect 4804 10202 4856 10208
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 4252 9988 4304 9994
rect 4252 9930 4304 9936
rect 4356 9518 4384 9998
rect 4896 9988 4948 9994
rect 4896 9930 4948 9936
rect 4421 9820 4717 9840
rect 4477 9818 4501 9820
rect 4557 9818 4581 9820
rect 4637 9818 4661 9820
rect 4499 9766 4501 9818
rect 4563 9766 4575 9818
rect 4637 9766 4639 9818
rect 4477 9764 4501 9766
rect 4557 9764 4581 9766
rect 4637 9764 4661 9766
rect 4421 9744 4717 9764
rect 4344 9512 4396 9518
rect 4344 9454 4396 9460
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 4421 8732 4717 8752
rect 4477 8730 4501 8732
rect 4557 8730 4581 8732
rect 4637 8730 4661 8732
rect 4499 8678 4501 8730
rect 4563 8678 4575 8730
rect 4637 8678 4639 8730
rect 4477 8676 4501 8678
rect 4557 8676 4581 8678
rect 4637 8676 4661 8678
rect 4421 8656 4717 8676
rect 4252 8356 4304 8362
rect 4252 8298 4304 8304
rect 4264 7750 4292 8298
rect 4436 8288 4488 8294
rect 4436 8230 4488 8236
rect 4344 8016 4396 8022
rect 4344 7958 4396 7964
rect 4252 7744 4304 7750
rect 4252 7686 4304 7692
rect 4264 7410 4292 7686
rect 4252 7404 4304 7410
rect 4252 7346 4304 7352
rect 4264 6798 4292 7346
rect 4356 7002 4384 7958
rect 4448 7886 4476 8230
rect 4436 7880 4488 7886
rect 4436 7822 4488 7828
rect 4421 7644 4717 7664
rect 4477 7642 4501 7644
rect 4557 7642 4581 7644
rect 4637 7642 4661 7644
rect 4499 7590 4501 7642
rect 4563 7590 4575 7642
rect 4637 7590 4639 7642
rect 4477 7588 4501 7590
rect 4557 7588 4581 7590
rect 4637 7588 4661 7590
rect 4421 7568 4717 7588
rect 4712 7200 4764 7206
rect 4712 7142 4764 7148
rect 4724 7002 4752 7142
rect 4344 6996 4396 7002
rect 4344 6938 4396 6944
rect 4712 6996 4764 7002
rect 4712 6938 4764 6944
rect 4816 6866 4844 8774
rect 4908 8430 4936 9930
rect 5000 9586 5028 11342
rect 5172 11290 5224 11296
rect 5368 10470 5396 12406
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 5080 10260 5132 10266
rect 5080 10202 5132 10208
rect 5092 10130 5120 10202
rect 5080 10124 5132 10130
rect 5080 10066 5132 10072
rect 5092 9654 5120 10066
rect 5080 9648 5132 9654
rect 5080 9590 5132 9596
rect 4988 9580 5040 9586
rect 4988 9522 5040 9528
rect 4896 8424 4948 8430
rect 4896 8366 4948 8372
rect 4908 7954 4936 8366
rect 4896 7948 4948 7954
rect 4896 7890 4948 7896
rect 5000 7342 5028 9522
rect 5368 9518 5396 10406
rect 5356 9512 5408 9518
rect 5356 9454 5408 9460
rect 5172 8968 5224 8974
rect 5172 8910 5224 8916
rect 5184 8634 5212 8910
rect 5172 8628 5224 8634
rect 5172 8570 5224 8576
rect 5184 8022 5212 8570
rect 5172 8016 5224 8022
rect 5172 7958 5224 7964
rect 5184 7410 5212 7958
rect 5368 7834 5396 9454
rect 5460 9178 5488 17206
rect 5644 17202 5672 17750
rect 5632 17196 5684 17202
rect 5632 17138 5684 17144
rect 5632 16992 5684 16998
rect 5632 16934 5684 16940
rect 5540 16720 5592 16726
rect 5644 16697 5672 16934
rect 5540 16662 5592 16668
rect 5630 16688 5686 16697
rect 5552 15706 5580 16662
rect 5630 16623 5686 16632
rect 5540 15700 5592 15706
rect 5540 15642 5592 15648
rect 5736 15450 5764 18278
rect 5920 16794 5948 18906
rect 6012 18902 6040 19994
rect 6104 19990 6132 20402
rect 6092 19984 6144 19990
rect 6092 19926 6144 19932
rect 6104 18970 6132 19926
rect 6092 18964 6144 18970
rect 6092 18906 6144 18912
rect 6000 18896 6052 18902
rect 6000 18838 6052 18844
rect 6196 18766 6224 22200
rect 6550 20496 6606 20505
rect 6550 20431 6552 20440
rect 6604 20431 6606 20440
rect 6552 20402 6604 20408
rect 6552 20256 6604 20262
rect 6552 20198 6604 20204
rect 6368 19916 6420 19922
rect 6368 19858 6420 19864
rect 6380 19310 6408 19858
rect 6460 19508 6512 19514
rect 6460 19450 6512 19456
rect 6276 19304 6328 19310
rect 6276 19246 6328 19252
rect 6368 19304 6420 19310
rect 6368 19246 6420 19252
rect 6184 18760 6236 18766
rect 6184 18702 6236 18708
rect 6090 18592 6146 18601
rect 6288 18578 6316 19246
rect 6146 18550 6316 18578
rect 6090 18527 6146 18536
rect 6000 17808 6052 17814
rect 6000 17750 6052 17756
rect 5908 16788 5960 16794
rect 5908 16730 5960 16736
rect 6012 16250 6040 17750
rect 6104 17660 6132 18527
rect 6368 18420 6420 18426
rect 6368 18362 6420 18368
rect 6276 18080 6328 18086
rect 6276 18022 6328 18028
rect 6184 17672 6236 17678
rect 6104 17632 6184 17660
rect 6000 16244 6052 16250
rect 6000 16186 6052 16192
rect 5998 16008 6054 16017
rect 6104 15994 6132 17632
rect 6184 17614 6236 17620
rect 6184 17060 6236 17066
rect 6184 17002 6236 17008
rect 6196 16454 6224 17002
rect 6184 16448 6236 16454
rect 6184 16390 6236 16396
rect 6054 15966 6132 15994
rect 5998 15943 6054 15952
rect 5816 15564 5868 15570
rect 5868 15524 5948 15552
rect 5816 15506 5868 15512
rect 5736 15422 5856 15450
rect 5540 13796 5592 13802
rect 5540 13738 5592 13744
rect 5552 13326 5580 13738
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 5552 12646 5580 13262
rect 5724 12776 5776 12782
rect 5724 12718 5776 12724
rect 5540 12640 5592 12646
rect 5540 12582 5592 12588
rect 5736 12442 5764 12718
rect 5724 12436 5776 12442
rect 5724 12378 5776 12384
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 5460 8022 5488 8230
rect 5448 8016 5500 8022
rect 5448 7958 5500 7964
rect 5368 7806 5488 7834
rect 5172 7404 5224 7410
rect 5172 7346 5224 7352
rect 4988 7336 5040 7342
rect 4988 7278 5040 7284
rect 4896 7200 4948 7206
rect 4896 7142 4948 7148
rect 4908 7002 4936 7142
rect 4896 6996 4948 7002
rect 4896 6938 4948 6944
rect 4804 6860 4856 6866
rect 4804 6802 4856 6808
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 4908 6662 4936 6938
rect 4896 6656 4948 6662
rect 4896 6598 4948 6604
rect 4421 6556 4717 6576
rect 4477 6554 4501 6556
rect 4557 6554 4581 6556
rect 4637 6554 4661 6556
rect 4499 6502 4501 6554
rect 4563 6502 4575 6554
rect 4637 6502 4639 6554
rect 4477 6500 4501 6502
rect 4557 6500 4581 6502
rect 4637 6500 4661 6502
rect 4421 6480 4717 6500
rect 4421 5468 4717 5488
rect 4477 5466 4501 5468
rect 4557 5466 4581 5468
rect 4637 5466 4661 5468
rect 4499 5414 4501 5466
rect 4563 5414 4575 5466
rect 4637 5414 4639 5466
rect 4477 5412 4501 5414
rect 4557 5412 4581 5414
rect 4637 5412 4661 5414
rect 4421 5392 4717 5412
rect 4421 4380 4717 4400
rect 4477 4378 4501 4380
rect 4557 4378 4581 4380
rect 4637 4378 4661 4380
rect 4499 4326 4501 4378
rect 4563 4326 4575 4378
rect 4637 4326 4639 4378
rect 4477 4324 4501 4326
rect 4557 4324 4581 4326
rect 4637 4324 4661 4326
rect 4421 4304 4717 4324
rect 5000 4146 5028 7278
rect 5460 7206 5488 7806
rect 5172 7200 5224 7206
rect 5172 7142 5224 7148
rect 5448 7200 5500 7206
rect 5448 7142 5500 7148
rect 5184 6934 5212 7142
rect 5172 6928 5224 6934
rect 5172 6870 5224 6876
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 4421 3292 4717 3312
rect 4477 3290 4501 3292
rect 4557 3290 4581 3292
rect 4637 3290 4661 3292
rect 4499 3238 4501 3290
rect 4563 3238 4575 3290
rect 4637 3238 4639 3290
rect 4477 3236 4501 3238
rect 4557 3236 4581 3238
rect 4637 3236 4661 3238
rect 4421 3216 4717 3236
rect 4172 2746 4384 2774
rect 4356 2650 4384 2746
rect 4344 2644 4396 2650
rect 4344 2586 4396 2592
rect 5460 2582 5488 7142
rect 5736 6934 5764 10406
rect 5828 10266 5856 15422
rect 5920 15026 5948 15524
rect 6012 15502 6040 15943
rect 6288 15910 6316 18022
rect 6380 17338 6408 18362
rect 6472 17814 6500 19450
rect 6460 17808 6512 17814
rect 6460 17750 6512 17756
rect 6368 17332 6420 17338
rect 6420 17292 6500 17320
rect 6368 17274 6420 17280
rect 6368 16992 6420 16998
rect 6368 16934 6420 16940
rect 6276 15904 6328 15910
rect 6276 15846 6328 15852
rect 6000 15496 6052 15502
rect 6000 15438 6052 15444
rect 5908 15020 5960 15026
rect 5908 14962 5960 14968
rect 5920 14074 5948 14962
rect 5908 14068 5960 14074
rect 5908 14010 5960 14016
rect 6092 14000 6144 14006
rect 6090 13968 6092 13977
rect 6144 13968 6146 13977
rect 6090 13903 6146 13912
rect 6000 13864 6052 13870
rect 6000 13806 6052 13812
rect 5908 13320 5960 13326
rect 5908 13262 5960 13268
rect 5920 12782 5948 13262
rect 6012 12850 6040 13806
rect 6000 12844 6052 12850
rect 6000 12786 6052 12792
rect 5908 12776 5960 12782
rect 5908 12718 5960 12724
rect 6012 12306 6040 12786
rect 6000 12300 6052 12306
rect 6052 12260 6132 12288
rect 6000 12242 6052 12248
rect 5908 12096 5960 12102
rect 5908 12038 5960 12044
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 5920 11801 5948 12038
rect 5906 11792 5962 11801
rect 5906 11727 5962 11736
rect 6012 11150 6040 12038
rect 6104 11898 6132 12260
rect 6092 11892 6144 11898
rect 6092 11834 6144 11840
rect 6000 11144 6052 11150
rect 6000 11086 6052 11092
rect 6380 10470 6408 16934
rect 6472 16658 6500 17292
rect 6460 16652 6512 16658
rect 6460 16594 6512 16600
rect 6564 16250 6592 20198
rect 6656 19446 6684 22200
rect 7116 20618 7144 22200
rect 7288 20800 7340 20806
rect 7576 20754 7604 22200
rect 7840 20868 7892 20874
rect 7840 20810 7892 20816
rect 7288 20742 7340 20748
rect 6932 20590 7144 20618
rect 6826 20496 6882 20505
rect 6826 20431 6882 20440
rect 6736 20392 6788 20398
rect 6736 20334 6788 20340
rect 6644 19440 6696 19446
rect 6644 19382 6696 19388
rect 6748 18970 6776 20334
rect 6840 20330 6868 20431
rect 6828 20324 6880 20330
rect 6828 20266 6880 20272
rect 6828 19916 6880 19922
rect 6828 19858 6880 19864
rect 6840 19514 6868 19858
rect 6828 19508 6880 19514
rect 6828 19450 6880 19456
rect 6736 18964 6788 18970
rect 6736 18906 6788 18912
rect 6644 18828 6696 18834
rect 6644 18770 6696 18776
rect 6656 18426 6684 18770
rect 6644 18420 6696 18426
rect 6644 18362 6696 18368
rect 6828 18284 6880 18290
rect 6828 18226 6880 18232
rect 6642 16688 6698 16697
rect 6642 16623 6644 16632
rect 6696 16623 6698 16632
rect 6644 16594 6696 16600
rect 6552 16244 6604 16250
rect 6552 16186 6604 16192
rect 6840 16046 6868 18226
rect 6828 16040 6880 16046
rect 6828 15982 6880 15988
rect 6932 15586 6960 20590
rect 7300 20534 7328 20742
rect 7484 20726 7604 20754
rect 7104 20528 7156 20534
rect 7104 20470 7156 20476
rect 7288 20528 7340 20534
rect 7288 20470 7340 20476
rect 7012 20324 7064 20330
rect 7012 20266 7064 20272
rect 7024 16522 7052 20266
rect 7116 19514 7144 20470
rect 7286 20088 7342 20097
rect 7286 20023 7288 20032
rect 7340 20023 7342 20032
rect 7288 19994 7340 20000
rect 7288 19712 7340 19718
rect 7288 19654 7340 19660
rect 7104 19508 7156 19514
rect 7104 19450 7156 19456
rect 7300 19174 7328 19654
rect 7484 19258 7512 20726
rect 7654 20632 7710 20641
rect 7564 20596 7616 20602
rect 7654 20567 7656 20576
rect 7564 20538 7616 20544
rect 7708 20567 7710 20576
rect 7656 20538 7708 20544
rect 7576 19990 7604 20538
rect 7852 20534 7880 20810
rect 7840 20528 7892 20534
rect 7840 20470 7892 20476
rect 7656 20392 7708 20398
rect 7656 20334 7708 20340
rect 7564 19984 7616 19990
rect 7564 19926 7616 19932
rect 7668 19718 7696 20334
rect 8036 20244 8064 22200
rect 8496 20602 8524 22200
rect 8956 20806 8984 22200
rect 9416 20874 9444 22200
rect 9404 20868 9456 20874
rect 9404 20810 9456 20816
rect 8944 20800 8996 20806
rect 8944 20742 8996 20748
rect 8484 20596 8536 20602
rect 8484 20538 8536 20544
rect 8496 20346 8524 20538
rect 9680 20460 9732 20466
rect 9680 20402 9732 20408
rect 9692 20346 9720 20402
rect 8496 20318 8708 20346
rect 8484 20256 8536 20262
rect 8036 20216 8248 20244
rect 7886 20156 8182 20176
rect 7942 20154 7966 20156
rect 8022 20154 8046 20156
rect 8102 20154 8126 20156
rect 7964 20102 7966 20154
rect 8028 20102 8040 20154
rect 8102 20102 8104 20154
rect 7942 20100 7966 20102
rect 8022 20100 8046 20102
rect 8102 20100 8126 20102
rect 7886 20080 8182 20100
rect 8220 19802 8248 20216
rect 8484 20198 8536 20204
rect 8390 20088 8446 20097
rect 8390 20023 8392 20032
rect 8444 20023 8446 20032
rect 8392 19994 8444 20000
rect 8128 19774 8248 19802
rect 7656 19712 7708 19718
rect 7656 19654 7708 19660
rect 7748 19712 7800 19718
rect 7748 19654 7800 19660
rect 7484 19230 7604 19258
rect 7288 19168 7340 19174
rect 7288 19110 7340 19116
rect 7472 19168 7524 19174
rect 7472 19110 7524 19116
rect 7104 18896 7156 18902
rect 7104 18838 7156 18844
rect 7012 16516 7064 16522
rect 7012 16458 7064 16464
rect 7116 16046 7144 18838
rect 7484 18766 7512 19110
rect 7576 18902 7604 19230
rect 7760 18970 7788 19654
rect 8128 19242 8156 19774
rect 8208 19712 8260 19718
rect 8208 19654 8260 19660
rect 8116 19236 8168 19242
rect 8116 19178 8168 19184
rect 7886 19068 8182 19088
rect 7942 19066 7966 19068
rect 8022 19066 8046 19068
rect 8102 19066 8126 19068
rect 7964 19014 7966 19066
rect 8028 19014 8040 19066
rect 8102 19014 8104 19066
rect 7942 19012 7966 19014
rect 8022 19012 8046 19014
rect 8102 19012 8126 19014
rect 7886 18992 8182 19012
rect 7748 18964 7800 18970
rect 7748 18906 7800 18912
rect 7564 18896 7616 18902
rect 7564 18838 7616 18844
rect 7472 18760 7524 18766
rect 7472 18702 7524 18708
rect 7380 18284 7432 18290
rect 7380 18226 7432 18232
rect 7196 18080 7248 18086
rect 7196 18022 7248 18028
rect 7288 18080 7340 18086
rect 7288 18022 7340 18028
rect 7208 16794 7236 18022
rect 7300 16794 7328 18022
rect 7392 17338 7420 18226
rect 7484 17814 7512 18702
rect 8024 18624 8076 18630
rect 8024 18566 8076 18572
rect 8036 18222 8064 18566
rect 8024 18216 8076 18222
rect 8024 18158 8076 18164
rect 7886 17980 8182 18000
rect 7942 17978 7966 17980
rect 8022 17978 8046 17980
rect 8102 17978 8126 17980
rect 7964 17926 7966 17978
rect 8028 17926 8040 17978
rect 8102 17926 8104 17978
rect 7942 17924 7966 17926
rect 8022 17924 8046 17926
rect 8102 17924 8126 17926
rect 7886 17904 8182 17924
rect 7564 17876 7616 17882
rect 7564 17818 7616 17824
rect 7472 17808 7524 17814
rect 7472 17750 7524 17756
rect 7380 17332 7432 17338
rect 7380 17274 7432 17280
rect 7196 16788 7248 16794
rect 7196 16730 7248 16736
rect 7288 16788 7340 16794
rect 7288 16730 7340 16736
rect 7104 16040 7156 16046
rect 7104 15982 7156 15988
rect 7392 15638 7420 17274
rect 7380 15632 7432 15638
rect 6932 15570 7236 15586
rect 7380 15574 7432 15580
rect 6932 15564 7248 15570
rect 6932 15558 7196 15564
rect 7196 15506 7248 15512
rect 6460 15496 6512 15502
rect 6460 15438 6512 15444
rect 6472 14482 6500 15438
rect 6644 15360 6696 15366
rect 6644 15302 6696 15308
rect 6920 15360 6972 15366
rect 6920 15302 6972 15308
rect 6552 14816 6604 14822
rect 6552 14758 6604 14764
rect 6460 14476 6512 14482
rect 6460 14418 6512 14424
rect 6472 13326 6500 14418
rect 6460 13320 6512 13326
rect 6460 13262 6512 13268
rect 6368 10464 6420 10470
rect 6368 10406 6420 10412
rect 5816 10260 5868 10266
rect 5816 10202 5868 10208
rect 6564 9382 6592 14758
rect 6656 14074 6684 15302
rect 6932 15026 6960 15302
rect 6920 15020 6972 15026
rect 6920 14962 6972 14968
rect 6932 14482 6960 14962
rect 7196 14884 7248 14890
rect 7196 14826 7248 14832
rect 7104 14816 7156 14822
rect 7104 14758 7156 14764
rect 7012 14544 7064 14550
rect 7012 14486 7064 14492
rect 6920 14476 6972 14482
rect 6920 14418 6972 14424
rect 6736 14272 6788 14278
rect 6736 14214 6788 14220
rect 6748 14074 6776 14214
rect 6644 14068 6696 14074
rect 6644 14010 6696 14016
rect 6736 14068 6788 14074
rect 6736 14010 6788 14016
rect 6920 13932 6972 13938
rect 6920 13874 6972 13880
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 6932 13682 6960 13874
rect 7024 13802 7052 14486
rect 7116 13802 7144 14758
rect 7012 13796 7064 13802
rect 7012 13738 7064 13744
rect 7104 13796 7156 13802
rect 7104 13738 7156 13744
rect 6644 13252 6696 13258
rect 6644 13194 6696 13200
rect 6656 13161 6684 13194
rect 6736 13184 6788 13190
rect 6642 13152 6698 13161
rect 6840 13172 6868 13670
rect 6932 13654 7052 13682
rect 6920 13184 6972 13190
rect 6840 13144 6920 13172
rect 6736 13126 6788 13132
rect 6920 13126 6972 13132
rect 6642 13087 6698 13096
rect 6748 12968 6776 13126
rect 6828 12980 6880 12986
rect 6748 12940 6828 12968
rect 6828 12922 6880 12928
rect 6828 12844 6880 12850
rect 6828 12786 6880 12792
rect 6840 12374 6868 12786
rect 7024 12374 7052 13654
rect 7208 12832 7236 14826
rect 7380 14612 7432 14618
rect 7380 14554 7432 14560
rect 7116 12804 7236 12832
rect 7288 12844 7340 12850
rect 6828 12368 6880 12374
rect 6828 12310 6880 12316
rect 7012 12368 7064 12374
rect 7012 12310 7064 12316
rect 7116 11762 7144 12804
rect 7288 12786 7340 12792
rect 7196 12640 7248 12646
rect 7196 12582 7248 12588
rect 7208 11898 7236 12582
rect 7196 11892 7248 11898
rect 7196 11834 7248 11840
rect 7104 11756 7156 11762
rect 7104 11698 7156 11704
rect 7300 11354 7328 12786
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 7012 11280 7064 11286
rect 7012 11222 7064 11228
rect 6644 11212 6696 11218
rect 6644 11154 6696 11160
rect 6656 9654 6684 11154
rect 6736 11144 6788 11150
rect 6736 11086 6788 11092
rect 6748 10606 6776 11086
rect 6736 10600 6788 10606
rect 6736 10542 6788 10548
rect 6748 10266 6776 10542
rect 7024 10266 7052 11222
rect 7392 11150 7420 14554
rect 7576 14482 7604 17818
rect 8116 17536 8168 17542
rect 8116 17478 8168 17484
rect 8128 17134 8156 17478
rect 8220 17184 8248 19654
rect 8220 17156 8340 17184
rect 7748 17128 7800 17134
rect 7748 17070 7800 17076
rect 8116 17128 8168 17134
rect 8168 17076 8248 17082
rect 8116 17070 8248 17076
rect 7760 16794 7788 17070
rect 8128 17054 8248 17070
rect 7886 16892 8182 16912
rect 7942 16890 7966 16892
rect 8022 16890 8046 16892
rect 8102 16890 8126 16892
rect 7964 16838 7966 16890
rect 8028 16838 8040 16890
rect 8102 16838 8104 16890
rect 7942 16836 7966 16838
rect 8022 16836 8046 16838
rect 8102 16836 8126 16838
rect 7886 16816 8182 16836
rect 7748 16788 7800 16794
rect 7748 16730 7800 16736
rect 8220 16590 8248 17054
rect 8312 16658 8340 17156
rect 8300 16652 8352 16658
rect 8300 16594 8352 16600
rect 8208 16584 8260 16590
rect 8208 16526 8260 16532
rect 8300 16108 8352 16114
rect 8300 16050 8352 16056
rect 8208 15972 8260 15978
rect 8208 15914 8260 15920
rect 7656 15904 7708 15910
rect 7656 15846 7708 15852
rect 7668 15706 7696 15846
rect 7886 15804 8182 15824
rect 7942 15802 7966 15804
rect 8022 15802 8046 15804
rect 8102 15802 8126 15804
rect 7964 15750 7966 15802
rect 8028 15750 8040 15802
rect 8102 15750 8104 15802
rect 7942 15748 7966 15750
rect 8022 15748 8046 15750
rect 8102 15748 8126 15750
rect 7886 15728 8182 15748
rect 7656 15700 7708 15706
rect 7656 15642 7708 15648
rect 8220 15026 8248 15914
rect 8312 15162 8340 16050
rect 8392 15360 8444 15366
rect 8392 15302 8444 15308
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 8208 15020 8260 15026
rect 8208 14962 8260 14968
rect 7886 14716 8182 14736
rect 7942 14714 7966 14716
rect 8022 14714 8046 14716
rect 8102 14714 8126 14716
rect 7964 14662 7966 14714
rect 8028 14662 8040 14714
rect 8102 14662 8104 14714
rect 7942 14660 7966 14662
rect 8022 14660 8046 14662
rect 8102 14660 8126 14662
rect 7886 14640 8182 14660
rect 7564 14476 7616 14482
rect 7564 14418 7616 14424
rect 7748 14272 7800 14278
rect 7748 14214 7800 14220
rect 7760 13938 7788 14214
rect 8208 14000 8260 14006
rect 8208 13942 8260 13948
rect 7748 13932 7800 13938
rect 7748 13874 7800 13880
rect 7472 13728 7524 13734
rect 7472 13670 7524 13676
rect 7484 12782 7512 13670
rect 7886 13628 8182 13648
rect 7942 13626 7966 13628
rect 8022 13626 8046 13628
rect 8102 13626 8126 13628
rect 7964 13574 7966 13626
rect 8028 13574 8040 13626
rect 8102 13574 8104 13626
rect 7942 13572 7966 13574
rect 8022 13572 8046 13574
rect 8102 13572 8126 13574
rect 7886 13552 8182 13572
rect 8220 13258 8248 13942
rect 8404 13530 8432 15302
rect 8392 13524 8444 13530
rect 8392 13466 8444 13472
rect 8208 13252 8260 13258
rect 8208 13194 8260 13200
rect 8116 13184 8168 13190
rect 8114 13152 8116 13161
rect 8168 13152 8170 13161
rect 8114 13087 8170 13096
rect 7472 12776 7524 12782
rect 7472 12718 7524 12724
rect 7748 12776 7800 12782
rect 7748 12718 7800 12724
rect 7564 12708 7616 12714
rect 7564 12650 7616 12656
rect 7576 12442 7604 12650
rect 7564 12436 7616 12442
rect 7760 12434 7788 12718
rect 7886 12540 8182 12560
rect 7942 12538 7966 12540
rect 8022 12538 8046 12540
rect 8102 12538 8126 12540
rect 7964 12486 7966 12538
rect 8028 12486 8040 12538
rect 8102 12486 8104 12538
rect 7942 12484 7966 12486
rect 8022 12484 8046 12486
rect 8102 12484 8126 12486
rect 7886 12464 8182 12484
rect 7564 12378 7616 12384
rect 7668 12406 7788 12434
rect 7564 12232 7616 12238
rect 7564 12174 7616 12180
rect 7470 11792 7526 11801
rect 7470 11727 7472 11736
rect 7524 11727 7526 11736
rect 7472 11698 7524 11704
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 7576 11082 7604 12174
rect 7564 11076 7616 11082
rect 7564 11018 7616 11024
rect 7668 11014 7696 12406
rect 8208 12232 8260 12238
rect 8208 12174 8260 12180
rect 8220 11762 8248 12174
rect 8496 12170 8524 20198
rect 8680 19922 8708 20318
rect 9312 20324 9364 20330
rect 9312 20266 9364 20272
rect 9600 20318 9720 20346
rect 8942 20088 8998 20097
rect 8942 20023 8998 20032
rect 8668 19916 8720 19922
rect 8668 19858 8720 19864
rect 8852 19848 8904 19854
rect 8850 19816 8852 19825
rect 8904 19816 8906 19825
rect 8760 19780 8812 19786
rect 8850 19751 8906 19760
rect 8760 19722 8812 19728
rect 8772 19310 8800 19722
rect 8760 19304 8812 19310
rect 8760 19246 8812 19252
rect 8668 18760 8720 18766
rect 8668 18702 8720 18708
rect 8576 17332 8628 17338
rect 8576 17274 8628 17280
rect 8588 14890 8616 17274
rect 8680 16658 8708 18702
rect 8852 18692 8904 18698
rect 8852 18634 8904 18640
rect 8864 18426 8892 18634
rect 8852 18420 8904 18426
rect 8852 18362 8904 18368
rect 8850 18184 8906 18193
rect 8850 18119 8906 18128
rect 8668 16652 8720 16658
rect 8668 16594 8720 16600
rect 8576 14884 8628 14890
rect 8576 14826 8628 14832
rect 8680 14618 8708 16594
rect 8760 15428 8812 15434
rect 8760 15370 8812 15376
rect 8668 14612 8720 14618
rect 8668 14554 8720 14560
rect 8772 12646 8800 15370
rect 8864 14482 8892 18119
rect 8852 14476 8904 14482
rect 8852 14418 8904 14424
rect 8956 14362 8984 20023
rect 9220 19304 9272 19310
rect 9220 19246 9272 19252
rect 9324 19258 9352 20266
rect 9600 19922 9628 20318
rect 9680 20256 9732 20262
rect 9732 20216 9812 20244
rect 9680 20198 9732 20204
rect 9588 19916 9640 19922
rect 9588 19858 9640 19864
rect 9232 18630 9260 19246
rect 9324 19230 9444 19258
rect 9312 19168 9364 19174
rect 9312 19110 9364 19116
rect 9324 18834 9352 19110
rect 9312 18828 9364 18834
rect 9312 18770 9364 18776
rect 9220 18624 9272 18630
rect 9220 18566 9272 18572
rect 9126 17776 9182 17785
rect 9126 17711 9182 17720
rect 9036 17604 9088 17610
rect 9036 17546 9088 17552
rect 8864 14334 8984 14362
rect 8760 12640 8812 12646
rect 8760 12582 8812 12588
rect 8772 12306 8800 12582
rect 8668 12300 8720 12306
rect 8668 12242 8720 12248
rect 8760 12300 8812 12306
rect 8760 12242 8812 12248
rect 8484 12164 8536 12170
rect 8484 12106 8536 12112
rect 8576 12096 8628 12102
rect 8576 12038 8628 12044
rect 8300 11892 8352 11898
rect 8300 11834 8352 11840
rect 8208 11756 8260 11762
rect 8208 11698 8260 11704
rect 7748 11620 7800 11626
rect 7748 11562 7800 11568
rect 7656 11008 7708 11014
rect 7656 10950 7708 10956
rect 7668 10810 7696 10950
rect 7656 10804 7708 10810
rect 7656 10746 7708 10752
rect 6736 10260 6788 10266
rect 6736 10202 6788 10208
rect 7012 10260 7064 10266
rect 7012 10202 7064 10208
rect 6828 10124 6880 10130
rect 6828 10066 6880 10072
rect 6644 9648 6696 9654
rect 6644 9590 6696 9596
rect 6840 9586 6868 10066
rect 7104 10056 7156 10062
rect 7104 9998 7156 10004
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 7116 9518 7144 9998
rect 7668 9602 7696 10746
rect 7760 10674 7788 11562
rect 7886 11452 8182 11472
rect 7942 11450 7966 11452
rect 8022 11450 8046 11452
rect 8102 11450 8126 11452
rect 7964 11398 7966 11450
rect 8028 11398 8040 11450
rect 8102 11398 8104 11450
rect 7942 11396 7966 11398
rect 8022 11396 8046 11398
rect 8102 11396 8126 11398
rect 7886 11376 8182 11396
rect 8024 11212 8076 11218
rect 8220 11200 8248 11698
rect 8312 11354 8340 11834
rect 8588 11830 8616 12038
rect 8576 11824 8628 11830
rect 8576 11766 8628 11772
rect 8300 11348 8352 11354
rect 8300 11290 8352 11296
rect 8076 11172 8248 11200
rect 8024 11154 8076 11160
rect 8036 10810 8064 11154
rect 8024 10804 8076 10810
rect 8024 10746 8076 10752
rect 7748 10668 7800 10674
rect 7748 10610 7800 10616
rect 8300 10668 8352 10674
rect 8300 10610 8352 10616
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 7886 10364 8182 10384
rect 7942 10362 7966 10364
rect 8022 10362 8046 10364
rect 8102 10362 8126 10364
rect 7964 10310 7966 10362
rect 8028 10310 8040 10362
rect 8102 10310 8104 10362
rect 7942 10308 7966 10310
rect 8022 10308 8046 10310
rect 8102 10308 8126 10310
rect 7886 10288 8182 10308
rect 8220 10266 8248 10406
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 7668 9586 7788 9602
rect 7656 9580 7788 9586
rect 7708 9574 7788 9580
rect 7656 9522 7708 9528
rect 7104 9512 7156 9518
rect 7104 9454 7156 9460
rect 7656 9444 7708 9450
rect 7656 9386 7708 9392
rect 6552 9376 6604 9382
rect 6552 9318 6604 9324
rect 7288 9036 7340 9042
rect 7288 8978 7340 8984
rect 6920 7472 6972 7478
rect 7196 7472 7248 7478
rect 6972 7420 7196 7426
rect 6920 7414 7248 7420
rect 6932 7398 7236 7414
rect 5724 6928 5776 6934
rect 5724 6870 5776 6876
rect 7300 6730 7328 8978
rect 7668 8974 7696 9386
rect 7656 8968 7708 8974
rect 7656 8910 7708 8916
rect 7668 8090 7696 8910
rect 7656 8084 7708 8090
rect 7656 8026 7708 8032
rect 7760 8022 7788 9574
rect 7886 9276 8182 9296
rect 7942 9274 7966 9276
rect 8022 9274 8046 9276
rect 8102 9274 8126 9276
rect 7964 9222 7966 9274
rect 8028 9222 8040 9274
rect 8102 9222 8104 9274
rect 7942 9220 7966 9222
rect 8022 9220 8046 9222
rect 8102 9220 8126 9222
rect 7886 9200 8182 9220
rect 8312 8362 8340 10610
rect 8588 10606 8616 11766
rect 8680 11354 8708 12242
rect 8668 11348 8720 11354
rect 8668 11290 8720 11296
rect 8576 10600 8628 10606
rect 8576 10542 8628 10548
rect 8864 9382 8892 14334
rect 8944 13456 8996 13462
rect 8944 13398 8996 13404
rect 8956 10470 8984 13398
rect 9048 10674 9076 17546
rect 9140 17270 9168 17711
rect 9128 17264 9180 17270
rect 9128 17206 9180 17212
rect 9232 17134 9260 18566
rect 9220 17128 9272 17134
rect 9220 17070 9272 17076
rect 9232 15978 9260 17070
rect 9416 16697 9444 19230
rect 9680 19168 9732 19174
rect 9680 19110 9732 19116
rect 9692 18222 9720 19110
rect 9784 18290 9812 20216
rect 9772 18284 9824 18290
rect 9772 18226 9824 18232
rect 9876 18222 9904 22200
rect 10140 20868 10192 20874
rect 10140 20810 10192 20816
rect 10048 20800 10100 20806
rect 10048 20742 10100 20748
rect 9956 20460 10008 20466
rect 9956 20402 10008 20408
rect 9968 19310 9996 20402
rect 10060 20398 10088 20742
rect 10048 20392 10100 20398
rect 10048 20334 10100 20340
rect 10152 20330 10180 20810
rect 10140 20324 10192 20330
rect 10140 20266 10192 20272
rect 10048 20256 10100 20262
rect 10046 20224 10048 20233
rect 10100 20224 10102 20233
rect 10046 20159 10102 20168
rect 9956 19304 10008 19310
rect 9956 19246 10008 19252
rect 9968 18970 9996 19246
rect 9956 18964 10008 18970
rect 9956 18906 10008 18912
rect 10336 18902 10364 22200
rect 10506 20360 10562 20369
rect 10506 20295 10562 20304
rect 10520 20262 10548 20295
rect 10416 20256 10468 20262
rect 10416 20198 10468 20204
rect 10508 20256 10560 20262
rect 10508 20198 10560 20204
rect 10428 20058 10456 20198
rect 10506 20088 10562 20097
rect 10416 20052 10468 20058
rect 10506 20023 10508 20032
rect 10416 19994 10468 20000
rect 10560 20023 10562 20032
rect 10508 19994 10560 20000
rect 10692 19916 10744 19922
rect 10692 19858 10744 19864
rect 10416 19236 10468 19242
rect 10416 19178 10468 19184
rect 10324 18896 10376 18902
rect 10324 18838 10376 18844
rect 10140 18828 10192 18834
rect 10140 18770 10192 18776
rect 9680 18216 9732 18222
rect 9680 18158 9732 18164
rect 9864 18216 9916 18222
rect 9864 18158 9916 18164
rect 10152 17746 10180 18770
rect 10324 18080 10376 18086
rect 10324 18022 10376 18028
rect 10336 17882 10364 18022
rect 10324 17876 10376 17882
rect 10324 17818 10376 17824
rect 9864 17740 9916 17746
rect 9864 17682 9916 17688
rect 10140 17740 10192 17746
rect 10140 17682 10192 17688
rect 10324 17740 10376 17746
rect 10324 17682 10376 17688
rect 9772 17536 9824 17542
rect 9772 17478 9824 17484
rect 9680 16992 9732 16998
rect 9680 16934 9732 16940
rect 9692 16794 9720 16934
rect 9784 16794 9812 17478
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 9772 16788 9824 16794
rect 9772 16730 9824 16736
rect 9402 16688 9458 16697
rect 9402 16623 9458 16632
rect 9220 15972 9272 15978
rect 9220 15914 9272 15920
rect 9232 15348 9260 15914
rect 9312 15904 9364 15910
rect 9312 15846 9364 15852
rect 9324 15706 9352 15846
rect 9312 15700 9364 15706
rect 9312 15642 9364 15648
rect 9876 15586 9904 17682
rect 10048 17672 10100 17678
rect 10048 17614 10100 17620
rect 10060 17066 10088 17614
rect 10140 17536 10192 17542
rect 10140 17478 10192 17484
rect 10048 17060 10100 17066
rect 10048 17002 10100 17008
rect 10060 16250 10088 17002
rect 10048 16244 10100 16250
rect 10048 16186 10100 16192
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 9784 15558 9904 15586
rect 10048 15564 10100 15570
rect 9312 15360 9364 15366
rect 9232 15320 9312 15348
rect 9312 15302 9364 15308
rect 9220 14476 9272 14482
rect 9220 14418 9272 14424
rect 9128 13796 9180 13802
rect 9128 13738 9180 13744
rect 9140 13258 9168 13738
rect 9128 13252 9180 13258
rect 9128 13194 9180 13200
rect 9140 12986 9168 13194
rect 9128 12980 9180 12986
rect 9128 12922 9180 12928
rect 9232 12442 9260 14418
rect 9324 13852 9352 15302
rect 9692 14822 9720 15506
rect 9680 14816 9732 14822
rect 9680 14758 9732 14764
rect 9494 14104 9550 14113
rect 9494 14039 9550 14048
rect 9678 14104 9734 14113
rect 9678 14039 9680 14048
rect 9508 14006 9536 14039
rect 9732 14039 9734 14048
rect 9680 14010 9732 14016
rect 9496 14000 9548 14006
rect 9496 13942 9548 13948
rect 9404 13864 9456 13870
rect 9324 13824 9404 13852
rect 9404 13806 9456 13812
rect 9634 13796 9686 13802
rect 9508 13756 9634 13784
rect 9508 13326 9536 13756
rect 9634 13738 9686 13744
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 9784 12918 9812 15558
rect 10048 15506 10100 15512
rect 9864 15496 9916 15502
rect 10060 15473 10088 15506
rect 9864 15438 9916 15444
rect 10046 15464 10102 15473
rect 9876 14890 9904 15438
rect 10046 15399 10102 15408
rect 9956 15360 10008 15366
rect 9956 15302 10008 15308
rect 9968 14958 9996 15302
rect 10152 15162 10180 17478
rect 10232 16720 10284 16726
rect 10232 16662 10284 16668
rect 10244 15366 10272 16662
rect 10336 16538 10364 17682
rect 10428 17066 10456 19178
rect 10600 18828 10652 18834
rect 10600 18770 10652 18776
rect 10508 17876 10560 17882
rect 10508 17818 10560 17824
rect 10520 17785 10548 17818
rect 10506 17776 10562 17785
rect 10506 17711 10562 17720
rect 10508 17604 10560 17610
rect 10508 17546 10560 17552
rect 10416 17060 10468 17066
rect 10416 17002 10468 17008
rect 10428 16658 10456 17002
rect 10416 16652 10468 16658
rect 10416 16594 10468 16600
rect 10336 16510 10456 16538
rect 10324 16448 10376 16454
rect 10324 16390 10376 16396
rect 10232 15360 10284 15366
rect 10232 15302 10284 15308
rect 10140 15156 10192 15162
rect 10140 15098 10192 15104
rect 9956 14952 10008 14958
rect 9954 14920 9956 14929
rect 10008 14920 10010 14929
rect 9864 14884 9916 14890
rect 9954 14855 10010 14864
rect 9864 14826 9916 14832
rect 9876 14074 9904 14826
rect 10048 14816 10100 14822
rect 10048 14758 10100 14764
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 9864 14068 9916 14074
rect 9864 14010 9916 14016
rect 9968 13530 9996 14418
rect 10060 14346 10088 14758
rect 10048 14340 10100 14346
rect 10048 14282 10100 14288
rect 10140 14272 10192 14278
rect 10140 14214 10192 14220
rect 9956 13524 10008 13530
rect 9956 13466 10008 13472
rect 10152 13258 10180 14214
rect 10244 13394 10272 15302
rect 10336 15026 10364 16390
rect 10428 16046 10456 16510
rect 10416 16040 10468 16046
rect 10416 15982 10468 15988
rect 10416 15156 10468 15162
rect 10416 15098 10468 15104
rect 10324 15020 10376 15026
rect 10324 14962 10376 14968
rect 10428 14346 10456 15098
rect 10416 14340 10468 14346
rect 10416 14282 10468 14288
rect 10232 13388 10284 13394
rect 10232 13330 10284 13336
rect 10140 13252 10192 13258
rect 10140 13194 10192 13200
rect 9772 12912 9824 12918
rect 9772 12854 9824 12860
rect 10048 12912 10100 12918
rect 10048 12854 10100 12860
rect 9220 12436 9272 12442
rect 9220 12378 9272 12384
rect 9956 12232 10008 12238
rect 9956 12174 10008 12180
rect 9968 11694 9996 12174
rect 9680 11688 9732 11694
rect 9126 11656 9182 11665
rect 9680 11630 9732 11636
rect 9956 11688 10008 11694
rect 9956 11630 10008 11636
rect 9126 11591 9182 11600
rect 9140 11558 9168 11591
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 9692 11150 9720 11630
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 9692 10810 9720 11086
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9036 10668 9088 10674
rect 9036 10610 9088 10616
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 8944 10464 8996 10470
rect 8944 10406 8996 10412
rect 8852 9376 8904 9382
rect 8852 9318 8904 9324
rect 8956 9110 8984 10406
rect 9692 10130 9720 10610
rect 10060 10538 10088 12854
rect 10520 11626 10548 17546
rect 10612 17338 10640 18770
rect 10704 17785 10732 19858
rect 10796 18222 10824 22200
rect 10968 20392 11020 20398
rect 10968 20334 11020 20340
rect 10876 19984 10928 19990
rect 10876 19926 10928 19932
rect 10888 19514 10916 19926
rect 10876 19508 10928 19514
rect 10876 19450 10928 19456
rect 10980 19310 11008 20334
rect 11256 20040 11284 22200
rect 11352 20700 11648 20720
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11430 20646 11432 20698
rect 11494 20646 11506 20698
rect 11568 20646 11570 20698
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11352 20624 11648 20644
rect 11336 20528 11388 20534
rect 11612 20528 11664 20534
rect 11388 20488 11612 20516
rect 11336 20470 11388 20476
rect 11612 20470 11664 20476
rect 11256 20012 11468 20040
rect 11060 19984 11112 19990
rect 11060 19926 11112 19932
rect 10968 19304 11020 19310
rect 10968 19246 11020 19252
rect 11072 19174 11100 19926
rect 11336 19916 11388 19922
rect 11164 19876 11336 19904
rect 11164 19446 11192 19876
rect 11336 19858 11388 19864
rect 11440 19802 11468 20012
rect 11256 19774 11468 19802
rect 11152 19440 11204 19446
rect 11152 19382 11204 19388
rect 11060 19168 11112 19174
rect 11060 19110 11112 19116
rect 10968 18624 11020 18630
rect 10968 18566 11020 18572
rect 10784 18216 10836 18222
rect 10784 18158 10836 18164
rect 10784 18080 10836 18086
rect 10784 18022 10836 18028
rect 10690 17776 10746 17785
rect 10690 17711 10746 17720
rect 10600 17332 10652 17338
rect 10600 17274 10652 17280
rect 10612 16590 10640 17274
rect 10692 16652 10744 16658
rect 10692 16594 10744 16600
rect 10600 16584 10652 16590
rect 10600 16526 10652 16532
rect 10600 15904 10652 15910
rect 10600 15846 10652 15852
rect 10612 14618 10640 15846
rect 10704 15570 10732 16594
rect 10692 15564 10744 15570
rect 10692 15506 10744 15512
rect 10600 14612 10652 14618
rect 10600 14554 10652 14560
rect 10704 14482 10732 15506
rect 10692 14476 10744 14482
rect 10692 14418 10744 14424
rect 10600 13796 10652 13802
rect 10600 13738 10652 13744
rect 10612 12918 10640 13738
rect 10796 13462 10824 18022
rect 10876 16108 10928 16114
rect 10876 16050 10928 16056
rect 10888 14890 10916 16050
rect 10980 15706 11008 18566
rect 11072 18290 11100 19110
rect 11152 18964 11204 18970
rect 11152 18906 11204 18912
rect 11060 18284 11112 18290
rect 11060 18226 11112 18232
rect 11060 18080 11112 18086
rect 11060 18022 11112 18028
rect 11072 15994 11100 18022
rect 11164 17134 11192 18906
rect 11256 17746 11284 19774
rect 11352 19612 11648 19632
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11430 19558 11432 19610
rect 11494 19558 11506 19610
rect 11568 19558 11570 19610
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11352 19536 11648 19556
rect 11336 19440 11388 19446
rect 11336 19382 11388 19388
rect 11348 18766 11376 19382
rect 11716 19334 11744 22200
rect 11796 19712 11848 19718
rect 11848 19660 11928 19666
rect 11796 19654 11928 19660
rect 11808 19638 11928 19654
rect 11716 19306 11836 19334
rect 11336 18760 11388 18766
rect 11336 18702 11388 18708
rect 11704 18624 11756 18630
rect 11704 18566 11756 18572
rect 11352 18524 11648 18544
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11430 18470 11432 18522
rect 11494 18470 11506 18522
rect 11568 18470 11570 18522
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11352 18448 11648 18468
rect 11716 18426 11744 18566
rect 11704 18420 11756 18426
rect 11704 18362 11756 18368
rect 11704 18216 11756 18222
rect 11704 18158 11756 18164
rect 11244 17740 11296 17746
rect 11244 17682 11296 17688
rect 11256 17270 11284 17682
rect 11336 17672 11388 17678
rect 11334 17640 11336 17649
rect 11388 17640 11390 17649
rect 11334 17575 11390 17584
rect 11352 17436 11648 17456
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11430 17382 11432 17434
rect 11494 17382 11506 17434
rect 11568 17382 11570 17434
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11352 17360 11648 17380
rect 11716 17338 11744 18158
rect 11808 17649 11836 19306
rect 11794 17640 11850 17649
rect 11794 17575 11850 17584
rect 11704 17332 11756 17338
rect 11704 17274 11756 17280
rect 11244 17264 11296 17270
rect 11244 17206 11296 17212
rect 11900 17202 11928 19638
rect 12072 19304 12124 19310
rect 12072 19246 12124 19252
rect 11980 18760 12032 18766
rect 11980 18702 12032 18708
rect 11888 17196 11940 17202
rect 11888 17138 11940 17144
rect 11152 17128 11204 17134
rect 11152 17070 11204 17076
rect 11164 16250 11192 17070
rect 11888 16992 11940 16998
rect 11888 16934 11940 16940
rect 11244 16720 11296 16726
rect 11244 16662 11296 16668
rect 11794 16688 11850 16697
rect 11152 16244 11204 16250
rect 11152 16186 11204 16192
rect 11256 16114 11284 16662
rect 11794 16623 11850 16632
rect 11352 16348 11648 16368
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11430 16294 11432 16346
rect 11494 16294 11506 16346
rect 11568 16294 11570 16346
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11352 16272 11648 16292
rect 11244 16108 11296 16114
rect 11244 16050 11296 16056
rect 11704 16040 11756 16046
rect 11072 15966 11192 15994
rect 11704 15982 11756 15988
rect 11060 15904 11112 15910
rect 11060 15846 11112 15852
rect 10968 15700 11020 15706
rect 10968 15642 11020 15648
rect 10968 15360 11020 15366
rect 10968 15302 11020 15308
rect 10980 14890 11008 15302
rect 10876 14884 10928 14890
rect 10876 14826 10928 14832
rect 10968 14884 11020 14890
rect 10968 14826 11020 14832
rect 10888 14482 10916 14826
rect 11072 14618 11100 15846
rect 11060 14612 11112 14618
rect 11060 14554 11112 14560
rect 10876 14476 10928 14482
rect 10876 14418 10928 14424
rect 10784 13456 10836 13462
rect 10784 13398 10836 13404
rect 10888 13394 10916 14418
rect 11164 14113 11192 15966
rect 11352 15260 11648 15280
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11430 15206 11432 15258
rect 11494 15206 11506 15258
rect 11568 15206 11570 15258
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11352 15184 11648 15204
rect 11716 15094 11744 15982
rect 11704 15088 11756 15094
rect 11704 15030 11756 15036
rect 11336 14952 11388 14958
rect 11334 14920 11336 14929
rect 11388 14920 11390 14929
rect 11244 14884 11296 14890
rect 11334 14855 11390 14864
rect 11244 14826 11296 14832
rect 11256 14482 11284 14826
rect 11244 14476 11296 14482
rect 11244 14418 11296 14424
rect 11352 14172 11648 14192
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11430 14118 11432 14170
rect 11494 14118 11506 14170
rect 11568 14118 11570 14170
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11150 14104 11206 14113
rect 11352 14096 11648 14116
rect 11150 14039 11206 14048
rect 11808 13394 11836 16623
rect 11900 16454 11928 16934
rect 11992 16522 12020 18702
rect 11980 16516 12032 16522
rect 11980 16458 12032 16464
rect 11888 16448 11940 16454
rect 11888 16390 11940 16396
rect 11888 15972 11940 15978
rect 11888 15914 11940 15920
rect 11900 13530 11928 15914
rect 11992 15638 12020 16458
rect 11980 15632 12032 15638
rect 11980 15574 12032 15580
rect 12084 15162 12112 19246
rect 12176 18970 12204 22200
rect 12256 20256 12308 20262
rect 12256 20198 12308 20204
rect 12164 18964 12216 18970
rect 12164 18906 12216 18912
rect 12164 18828 12216 18834
rect 12164 18770 12216 18776
rect 12176 16250 12204 18770
rect 12268 18698 12296 20198
rect 12348 19916 12400 19922
rect 12400 19876 12480 19904
rect 12348 19858 12400 19864
rect 12452 18970 12480 19876
rect 12636 19530 12664 22200
rect 13096 20534 13124 22200
rect 13556 20534 13584 22200
rect 14016 20534 14044 22200
rect 14476 20602 14504 22200
rect 14464 20596 14516 20602
rect 14464 20538 14516 20544
rect 13084 20528 13136 20534
rect 13084 20470 13136 20476
rect 13544 20528 13596 20534
rect 13544 20470 13596 20476
rect 14004 20528 14056 20534
rect 14004 20470 14056 20476
rect 14936 20466 14964 22200
rect 14924 20460 14976 20466
rect 14924 20402 14976 20408
rect 12808 20392 12860 20398
rect 12808 20334 12860 20340
rect 14280 20392 14332 20398
rect 14280 20334 14332 20340
rect 12820 20058 12848 20334
rect 13268 20324 13320 20330
rect 13268 20266 13320 20272
rect 13820 20324 13872 20330
rect 13820 20266 13872 20272
rect 13912 20324 13964 20330
rect 13912 20266 13964 20272
rect 12808 20052 12860 20058
rect 12808 19994 12860 20000
rect 13176 19712 13228 19718
rect 13176 19654 13228 19660
rect 12636 19502 12940 19530
rect 12532 19440 12584 19446
rect 12808 19440 12860 19446
rect 12584 19388 12808 19394
rect 12532 19382 12860 19388
rect 12544 19366 12848 19382
rect 12532 19304 12584 19310
rect 12532 19246 12584 19252
rect 12440 18964 12492 18970
rect 12440 18906 12492 18912
rect 12256 18692 12308 18698
rect 12256 18634 12308 18640
rect 12440 18080 12492 18086
rect 12440 18022 12492 18028
rect 12452 17338 12480 18022
rect 12256 17332 12308 17338
rect 12256 17274 12308 17280
rect 12440 17332 12492 17338
rect 12440 17274 12492 17280
rect 12164 16244 12216 16250
rect 12164 16186 12216 16192
rect 12268 15910 12296 17274
rect 12440 17196 12492 17202
rect 12440 17138 12492 17144
rect 12348 16992 12400 16998
rect 12348 16934 12400 16940
rect 12360 16046 12388 16934
rect 12348 16040 12400 16046
rect 12348 15982 12400 15988
rect 12256 15904 12308 15910
rect 12256 15846 12308 15852
rect 12452 15638 12480 17138
rect 12440 15632 12492 15638
rect 12440 15574 12492 15580
rect 12254 15464 12310 15473
rect 12254 15399 12256 15408
rect 12308 15399 12310 15408
rect 12256 15370 12308 15376
rect 12072 15156 12124 15162
rect 12072 15098 12124 15104
rect 12452 15042 12480 15574
rect 12544 15162 12572 19246
rect 12716 18760 12768 18766
rect 12716 18702 12768 18708
rect 12728 18426 12756 18702
rect 12716 18420 12768 18426
rect 12716 18362 12768 18368
rect 12808 18352 12860 18358
rect 12808 18294 12860 18300
rect 12716 18284 12768 18290
rect 12716 18226 12768 18232
rect 12728 17542 12756 18226
rect 12820 17746 12848 18294
rect 12912 18222 12940 19502
rect 13084 19508 13136 19514
rect 13084 19450 13136 19456
rect 12992 18828 13044 18834
rect 12992 18770 13044 18776
rect 12900 18216 12952 18222
rect 12900 18158 12952 18164
rect 12808 17740 12860 17746
rect 12808 17682 12860 17688
rect 12716 17536 12768 17542
rect 12716 17478 12768 17484
rect 12624 17332 12676 17338
rect 12624 17274 12676 17280
rect 12532 15156 12584 15162
rect 12532 15098 12584 15104
rect 12360 15014 12480 15042
rect 12164 14544 12216 14550
rect 12162 14512 12164 14521
rect 12216 14512 12218 14521
rect 12162 14447 12218 14456
rect 12256 14476 12308 14482
rect 12256 14418 12308 14424
rect 12164 14408 12216 14414
rect 12164 14350 12216 14356
rect 11980 14272 12032 14278
rect 11980 14214 12032 14220
rect 12072 14272 12124 14278
rect 12072 14214 12124 14220
rect 11888 13524 11940 13530
rect 11888 13466 11940 13472
rect 10876 13388 10928 13394
rect 10876 13330 10928 13336
rect 11796 13388 11848 13394
rect 11796 13330 11848 13336
rect 11808 13274 11836 13330
rect 11808 13246 11928 13274
rect 11352 13084 11648 13104
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11430 13030 11432 13082
rect 11494 13030 11506 13082
rect 11568 13030 11570 13082
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11352 13008 11648 13028
rect 10600 12912 10652 12918
rect 10600 12854 10652 12860
rect 11704 12776 11756 12782
rect 11704 12718 11756 12724
rect 11152 12640 11204 12646
rect 11152 12582 11204 12588
rect 11060 11892 11112 11898
rect 11060 11834 11112 11840
rect 10508 11620 10560 11626
rect 10508 11562 10560 11568
rect 11072 11286 11100 11834
rect 11060 11280 11112 11286
rect 11060 11222 11112 11228
rect 10692 10804 10744 10810
rect 10692 10746 10744 10752
rect 9772 10532 9824 10538
rect 9772 10474 9824 10480
rect 10048 10532 10100 10538
rect 10048 10474 10100 10480
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 9680 10124 9732 10130
rect 9680 10066 9732 10072
rect 9600 9654 9628 10066
rect 9692 9722 9720 10066
rect 9680 9716 9732 9722
rect 9680 9658 9732 9664
rect 9588 9648 9640 9654
rect 9588 9590 9640 9596
rect 9784 9518 9812 10474
rect 10704 10130 10732 10746
rect 10692 10124 10744 10130
rect 10692 10066 10744 10072
rect 11060 10124 11112 10130
rect 11060 10066 11112 10072
rect 11072 9722 11100 10066
rect 11060 9716 11112 9722
rect 11060 9658 11112 9664
rect 9772 9512 9824 9518
rect 9772 9454 9824 9460
rect 9404 9376 9456 9382
rect 9404 9318 9456 9324
rect 8944 9104 8996 9110
rect 8944 9046 8996 9052
rect 9312 9036 9364 9042
rect 9312 8978 9364 8984
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8300 8356 8352 8362
rect 8300 8298 8352 8304
rect 8208 8288 8260 8294
rect 8208 8230 8260 8236
rect 7886 8188 8182 8208
rect 7942 8186 7966 8188
rect 8022 8186 8046 8188
rect 8102 8186 8126 8188
rect 7964 8134 7966 8186
rect 8028 8134 8040 8186
rect 8102 8134 8104 8186
rect 7942 8132 7966 8134
rect 8022 8132 8046 8134
rect 8102 8132 8126 8134
rect 7886 8112 8182 8132
rect 7748 8016 7800 8022
rect 7748 7958 7800 7964
rect 8220 7954 8248 8230
rect 8208 7948 8260 7954
rect 8208 7890 8260 7896
rect 7564 7336 7616 7342
rect 7564 7278 7616 7284
rect 7576 7002 7604 7278
rect 7748 7200 7800 7206
rect 7748 7142 7800 7148
rect 7760 7002 7788 7142
rect 7886 7100 8182 7120
rect 7942 7098 7966 7100
rect 8022 7098 8046 7100
rect 8102 7098 8126 7100
rect 7964 7046 7966 7098
rect 8028 7046 8040 7098
rect 8102 7046 8104 7098
rect 7942 7044 7966 7046
rect 8022 7044 8046 7046
rect 8102 7044 8126 7046
rect 7886 7024 8182 7044
rect 7564 6996 7616 7002
rect 7564 6938 7616 6944
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 8220 6798 8248 7890
rect 8404 7750 8432 8434
rect 9324 8090 9352 8978
rect 9416 8838 9444 9318
rect 9784 9178 9812 9454
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9404 8832 9456 8838
rect 9404 8774 9456 8780
rect 9312 8084 9364 8090
rect 9312 8026 9364 8032
rect 8852 7948 8904 7954
rect 8852 7890 8904 7896
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 8404 7410 8432 7686
rect 8864 7546 8892 7890
rect 8852 7540 8904 7546
rect 8852 7482 8904 7488
rect 8482 7440 8538 7449
rect 8392 7404 8444 7410
rect 8482 7375 8538 7384
rect 8392 7346 8444 7352
rect 8496 7206 8524 7375
rect 9416 7342 9444 8774
rect 9772 8560 9824 8566
rect 9772 8502 9824 8508
rect 9784 8090 9812 8502
rect 9772 8084 9824 8090
rect 9772 8026 9824 8032
rect 9404 7336 9456 7342
rect 9404 7278 9456 7284
rect 8484 7200 8536 7206
rect 8484 7142 8536 7148
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 7288 6724 7340 6730
rect 7288 6666 7340 6672
rect 7886 6012 8182 6032
rect 7942 6010 7966 6012
rect 8022 6010 8046 6012
rect 8102 6010 8126 6012
rect 7964 5958 7966 6010
rect 8028 5958 8040 6010
rect 8102 5958 8104 6010
rect 7942 5956 7966 5958
rect 8022 5956 8046 5958
rect 8102 5956 8126 5958
rect 7886 5936 8182 5956
rect 7886 4924 8182 4944
rect 7942 4922 7966 4924
rect 8022 4922 8046 4924
rect 8102 4922 8126 4924
rect 7964 4870 7966 4922
rect 8028 4870 8040 4922
rect 8102 4870 8104 4922
rect 7942 4868 7966 4870
rect 8022 4868 8046 4870
rect 8102 4868 8126 4870
rect 7886 4848 8182 4868
rect 11164 4622 11192 12582
rect 11352 11996 11648 12016
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11430 11942 11432 11994
rect 11494 11942 11506 11994
rect 11568 11942 11570 11994
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11352 11920 11648 11940
rect 11244 11008 11296 11014
rect 11244 10950 11296 10956
rect 11256 10606 11284 10950
rect 11352 10908 11648 10928
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11430 10854 11432 10906
rect 11494 10854 11506 10906
rect 11568 10854 11570 10906
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11352 10832 11648 10852
rect 11244 10600 11296 10606
rect 11244 10542 11296 10548
rect 11256 10062 11284 10542
rect 11716 10266 11744 12718
rect 11796 12640 11848 12646
rect 11796 12582 11848 12588
rect 11808 12238 11836 12582
rect 11796 12232 11848 12238
rect 11796 12174 11848 12180
rect 11796 10804 11848 10810
rect 11900 10792 11928 13246
rect 11992 12782 12020 14214
rect 12084 14074 12112 14214
rect 12072 14068 12124 14074
rect 12072 14010 12124 14016
rect 12176 13326 12204 14350
rect 12164 13320 12216 13326
rect 12164 13262 12216 13268
rect 12268 12918 12296 14418
rect 12360 13530 12388 15014
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 12452 13530 12480 14894
rect 12532 14884 12584 14890
rect 12532 14826 12584 14832
rect 12544 14521 12572 14826
rect 12530 14512 12586 14521
rect 12530 14447 12586 14456
rect 12532 13728 12584 13734
rect 12532 13670 12584 13676
rect 12348 13524 12400 13530
rect 12348 13466 12400 13472
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12544 12986 12572 13670
rect 12532 12980 12584 12986
rect 12532 12922 12584 12928
rect 12256 12912 12308 12918
rect 12256 12854 12308 12860
rect 11980 12776 12032 12782
rect 11980 12718 12032 12724
rect 12268 11880 12296 12854
rect 12636 12442 12664 17274
rect 12728 16114 12756 17478
rect 12820 17202 12848 17682
rect 12808 17196 12860 17202
rect 12808 17138 12860 17144
rect 12820 16590 12848 17138
rect 12808 16584 12860 16590
rect 12808 16526 12860 16532
rect 12808 16448 12860 16454
rect 12808 16390 12860 16396
rect 12716 16108 12768 16114
rect 12716 16050 12768 16056
rect 12820 14618 12848 16390
rect 12900 15904 12952 15910
rect 12900 15846 12952 15852
rect 12912 15706 12940 15846
rect 12900 15700 12952 15706
rect 12900 15642 12952 15648
rect 12808 14612 12860 14618
rect 12808 14554 12860 14560
rect 12716 14476 12768 14482
rect 12716 14418 12768 14424
rect 12728 13938 12756 14418
rect 12716 13932 12768 13938
rect 12716 13874 12768 13880
rect 12624 12436 12676 12442
rect 12624 12378 12676 12384
rect 12716 12164 12768 12170
rect 12716 12106 12768 12112
rect 12728 11898 12756 12106
rect 13004 11898 13032 18770
rect 13096 17202 13124 19450
rect 13188 17338 13216 19654
rect 13280 19514 13308 20266
rect 13636 20256 13688 20262
rect 13636 20198 13688 20204
rect 13648 19786 13676 20198
rect 13636 19780 13688 19786
rect 13636 19722 13688 19728
rect 13832 19514 13860 20266
rect 13924 20058 13952 20266
rect 14002 20224 14058 20233
rect 14002 20159 14058 20168
rect 13912 20052 13964 20058
rect 13912 19994 13964 20000
rect 14016 19854 14044 20159
rect 14188 19916 14240 19922
rect 14188 19858 14240 19864
rect 14004 19848 14056 19854
rect 14004 19790 14056 19796
rect 13268 19508 13320 19514
rect 13268 19450 13320 19456
rect 13820 19508 13872 19514
rect 13820 19450 13872 19456
rect 13452 19440 13504 19446
rect 13452 19382 13504 19388
rect 13360 19236 13412 19242
rect 13360 19178 13412 19184
rect 13268 19168 13320 19174
rect 13268 19110 13320 19116
rect 13280 18970 13308 19110
rect 13268 18964 13320 18970
rect 13268 18906 13320 18912
rect 13372 18630 13400 19178
rect 13360 18624 13412 18630
rect 13360 18566 13412 18572
rect 13268 18080 13320 18086
rect 13268 18022 13320 18028
rect 13360 18080 13412 18086
rect 13360 18022 13412 18028
rect 13176 17332 13228 17338
rect 13176 17274 13228 17280
rect 13084 17196 13136 17202
rect 13084 17138 13136 17144
rect 13096 15570 13124 17138
rect 13280 16794 13308 18022
rect 13372 17338 13400 18022
rect 13360 17332 13412 17338
rect 13360 17274 13412 17280
rect 13464 16998 13492 19382
rect 14004 19304 14056 19310
rect 14004 19246 14056 19252
rect 14016 18970 14044 19246
rect 14004 18964 14056 18970
rect 14004 18906 14056 18912
rect 13544 18896 13596 18902
rect 13544 18838 13596 18844
rect 13556 17746 13584 18838
rect 13820 18828 13872 18834
rect 13820 18770 13872 18776
rect 13832 18426 13860 18770
rect 13820 18420 13872 18426
rect 13820 18362 13872 18368
rect 14004 18216 14056 18222
rect 14004 18158 14056 18164
rect 14016 17746 14044 18158
rect 13544 17740 13596 17746
rect 13544 17682 13596 17688
rect 14004 17740 14056 17746
rect 14004 17682 14056 17688
rect 13634 17640 13690 17649
rect 13634 17575 13690 17584
rect 13648 17542 13676 17575
rect 13544 17536 13596 17542
rect 13544 17478 13596 17484
rect 13636 17536 13688 17542
rect 13636 17478 13688 17484
rect 13452 16992 13504 16998
rect 13452 16934 13504 16940
rect 13268 16788 13320 16794
rect 13268 16730 13320 16736
rect 13358 16688 13414 16697
rect 13176 16652 13228 16658
rect 13358 16623 13360 16632
rect 13176 16594 13228 16600
rect 13412 16623 13414 16632
rect 13360 16594 13412 16600
rect 13084 15564 13136 15570
rect 13084 15506 13136 15512
rect 13084 15428 13136 15434
rect 13084 15370 13136 15376
rect 12716 11892 12768 11898
rect 12268 11852 12572 11880
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 12084 11150 12112 11698
rect 12348 11620 12400 11626
rect 12348 11562 12400 11568
rect 12256 11348 12308 11354
rect 12256 11290 12308 11296
rect 12072 11144 12124 11150
rect 12072 11086 12124 11092
rect 11848 10764 11928 10792
rect 11796 10746 11848 10752
rect 11704 10260 11756 10266
rect 11704 10202 11756 10208
rect 11244 10056 11296 10062
rect 11244 9998 11296 10004
rect 11352 9820 11648 9840
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11430 9766 11432 9818
rect 11494 9766 11506 9818
rect 11568 9766 11570 9818
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11352 9744 11648 9764
rect 11352 8732 11648 8752
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11430 8678 11432 8730
rect 11494 8678 11506 8730
rect 11568 8678 11570 8730
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11352 8656 11648 8676
rect 11352 7644 11648 7664
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11430 7590 11432 7642
rect 11494 7590 11506 7642
rect 11568 7590 11570 7642
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11352 7568 11648 7588
rect 11352 6556 11648 6576
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11430 6502 11432 6554
rect 11494 6502 11506 6554
rect 11568 6502 11570 6554
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11352 6480 11648 6500
rect 11352 5468 11648 5488
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11430 5414 11432 5466
rect 11494 5414 11506 5466
rect 11568 5414 11570 5466
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11352 5392 11648 5412
rect 11152 4616 11204 4622
rect 11152 4558 11204 4564
rect 11352 4380 11648 4400
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11430 4326 11432 4378
rect 11494 4326 11506 4378
rect 11568 4326 11570 4378
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11352 4304 11648 4324
rect 7886 3836 8182 3856
rect 7942 3834 7966 3836
rect 8022 3834 8046 3836
rect 8102 3834 8126 3836
rect 7964 3782 7966 3834
rect 8028 3782 8040 3834
rect 8102 3782 8104 3834
rect 7942 3780 7966 3782
rect 8022 3780 8046 3782
rect 8102 3780 8126 3782
rect 7886 3760 8182 3780
rect 11352 3292 11648 3312
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11430 3238 11432 3290
rect 11494 3238 11506 3290
rect 11568 3238 11570 3290
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11352 3216 11648 3236
rect 7886 2748 8182 2768
rect 7942 2746 7966 2748
rect 8022 2746 8046 2748
rect 8102 2746 8126 2748
rect 7964 2694 7966 2746
rect 8028 2694 8040 2746
rect 8102 2694 8104 2746
rect 7942 2692 7966 2694
rect 8022 2692 8046 2694
rect 8102 2692 8126 2694
rect 7886 2672 8182 2692
rect 12268 2582 12296 11290
rect 12360 10266 12388 11562
rect 12544 10538 12572 11852
rect 12716 11834 12768 11840
rect 12992 11892 13044 11898
rect 12992 11834 13044 11840
rect 12900 11620 12952 11626
rect 12900 11562 12952 11568
rect 12716 11280 12768 11286
rect 12716 11222 12768 11228
rect 12728 10606 12756 11222
rect 12716 10600 12768 10606
rect 12716 10542 12768 10548
rect 12532 10532 12584 10538
rect 12532 10474 12584 10480
rect 12348 10260 12400 10266
rect 12348 10202 12400 10208
rect 12544 10130 12572 10474
rect 12912 10266 12940 11562
rect 12900 10260 12952 10266
rect 12900 10202 12952 10208
rect 12532 10124 12584 10130
rect 12532 10066 12584 10072
rect 13096 8498 13124 15370
rect 13188 14890 13216 16594
rect 13268 15360 13320 15366
rect 13268 15302 13320 15308
rect 13280 15026 13308 15302
rect 13268 15020 13320 15026
rect 13268 14962 13320 14968
rect 13176 14884 13228 14890
rect 13176 14826 13228 14832
rect 13464 14618 13492 16934
rect 13556 15434 13584 17478
rect 14016 17338 14044 17682
rect 14004 17332 14056 17338
rect 14004 17274 14056 17280
rect 13912 17060 13964 17066
rect 13912 17002 13964 17008
rect 13924 16794 13952 17002
rect 13912 16788 13964 16794
rect 13912 16730 13964 16736
rect 14096 15972 14148 15978
rect 14096 15914 14148 15920
rect 14004 15564 14056 15570
rect 14004 15506 14056 15512
rect 13544 15428 13596 15434
rect 13544 15370 13596 15376
rect 13728 15428 13780 15434
rect 13728 15370 13780 15376
rect 13912 15428 13964 15434
rect 13912 15370 13964 15376
rect 13636 15360 13688 15366
rect 13556 15308 13636 15314
rect 13556 15302 13688 15308
rect 13556 15286 13676 15302
rect 13452 14612 13504 14618
rect 13452 14554 13504 14560
rect 13464 14396 13492 14554
rect 13556 14550 13584 15286
rect 13740 14958 13768 15370
rect 13820 15360 13872 15366
rect 13820 15302 13872 15308
rect 13728 14952 13780 14958
rect 13728 14894 13780 14900
rect 13544 14544 13596 14550
rect 13544 14486 13596 14492
rect 13544 14408 13596 14414
rect 13464 14368 13544 14396
rect 13176 14340 13228 14346
rect 13176 14282 13228 14288
rect 13188 13734 13216 14282
rect 13268 14000 13320 14006
rect 13268 13942 13320 13948
rect 13280 13870 13308 13942
rect 13268 13864 13320 13870
rect 13268 13806 13320 13812
rect 13176 13728 13228 13734
rect 13176 13670 13228 13676
rect 13280 12850 13308 13806
rect 13268 12844 13320 12850
rect 13268 12786 13320 12792
rect 13280 12434 13308 12786
rect 13280 12406 13400 12434
rect 13372 12102 13400 12406
rect 13360 12096 13412 12102
rect 13360 12038 13412 12044
rect 13464 11558 13492 14368
rect 13544 14350 13596 14356
rect 13740 14074 13768 14894
rect 13832 14396 13860 15302
rect 13924 14498 13952 15370
rect 14016 14618 14044 15506
rect 14108 15162 14136 15914
rect 14096 15156 14148 15162
rect 14096 15098 14148 15104
rect 14004 14612 14056 14618
rect 14004 14554 14056 14560
rect 13924 14470 14136 14498
rect 13832 14368 13952 14396
rect 13728 14068 13780 14074
rect 13728 14010 13780 14016
rect 13740 13326 13768 14010
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 13728 13320 13780 13326
rect 13728 13262 13780 13268
rect 13648 12986 13676 13262
rect 13636 12980 13688 12986
rect 13636 12922 13688 12928
rect 13820 12776 13872 12782
rect 13820 12718 13872 12724
rect 13832 12306 13860 12718
rect 13820 12300 13872 12306
rect 13820 12242 13872 12248
rect 13924 12170 13952 14368
rect 14004 13184 14056 13190
rect 14004 13126 14056 13132
rect 14016 12850 14044 13126
rect 14004 12844 14056 12850
rect 14004 12786 14056 12792
rect 14016 12374 14044 12786
rect 14004 12368 14056 12374
rect 14004 12310 14056 12316
rect 13912 12164 13964 12170
rect 13912 12106 13964 12112
rect 13636 12096 13688 12102
rect 13636 12038 13688 12044
rect 13452 11552 13504 11558
rect 13452 11494 13504 11500
rect 13648 11218 13676 12038
rect 13820 11756 13872 11762
rect 13820 11698 13872 11704
rect 13832 11354 13860 11698
rect 13820 11348 13872 11354
rect 13820 11290 13872 11296
rect 13268 11212 13320 11218
rect 13268 11154 13320 11160
rect 13636 11212 13688 11218
rect 13636 11154 13688 11160
rect 13280 10810 13308 11154
rect 13268 10804 13320 10810
rect 13268 10746 13320 10752
rect 13648 10606 13676 11154
rect 13832 10606 13860 11290
rect 13636 10600 13688 10606
rect 13636 10542 13688 10548
rect 13820 10600 13872 10606
rect 13820 10542 13872 10548
rect 14108 9382 14136 14470
rect 14200 11898 14228 19858
rect 14292 19514 14320 20334
rect 14817 20156 15113 20176
rect 14873 20154 14897 20156
rect 14953 20154 14977 20156
rect 15033 20154 15057 20156
rect 14895 20102 14897 20154
rect 14959 20102 14971 20154
rect 15033 20102 15035 20154
rect 14873 20100 14897 20102
rect 14953 20100 14977 20102
rect 15033 20100 15057 20102
rect 14817 20080 15113 20100
rect 15396 19990 15424 22200
rect 15568 20324 15620 20330
rect 15568 20266 15620 20272
rect 15384 19984 15436 19990
rect 15384 19926 15436 19932
rect 15200 19916 15252 19922
rect 15200 19858 15252 19864
rect 14280 19508 14332 19514
rect 14280 19450 14332 19456
rect 15212 19174 15240 19858
rect 15292 19712 15344 19718
rect 15292 19654 15344 19660
rect 15304 19310 15332 19654
rect 15580 19378 15608 20266
rect 15856 19990 15884 22200
rect 16120 20324 16172 20330
rect 16120 20266 16172 20272
rect 16132 20058 16160 20266
rect 16120 20052 16172 20058
rect 16120 19994 16172 20000
rect 16316 19990 16344 22200
rect 16578 20496 16634 20505
rect 16578 20431 16580 20440
rect 16632 20431 16634 20440
rect 16580 20402 16632 20408
rect 16776 19990 16804 22200
rect 17236 20058 17264 22200
rect 17696 20534 17724 22200
rect 18156 20534 18184 22200
rect 18282 20700 18578 20720
rect 18338 20698 18362 20700
rect 18418 20698 18442 20700
rect 18498 20698 18522 20700
rect 18360 20646 18362 20698
rect 18424 20646 18436 20698
rect 18498 20646 18500 20698
rect 18338 20644 18362 20646
rect 18418 20644 18442 20646
rect 18498 20644 18522 20646
rect 18282 20624 18578 20644
rect 18616 20534 18644 22200
rect 19076 20534 19104 22200
rect 19536 20602 19564 22200
rect 19524 20596 19576 20602
rect 19524 20538 19576 20544
rect 17684 20528 17736 20534
rect 17684 20470 17736 20476
rect 18144 20528 18196 20534
rect 18144 20470 18196 20476
rect 18604 20528 18656 20534
rect 18604 20470 18656 20476
rect 19064 20528 19116 20534
rect 19064 20470 19116 20476
rect 19340 20392 19392 20398
rect 19340 20334 19392 20340
rect 18052 20324 18104 20330
rect 18052 20266 18104 20272
rect 18604 20324 18656 20330
rect 18604 20266 18656 20272
rect 18972 20324 19024 20330
rect 18972 20266 19024 20272
rect 17224 20052 17276 20058
rect 17224 19994 17276 20000
rect 15844 19984 15896 19990
rect 15844 19926 15896 19932
rect 16304 19984 16356 19990
rect 16304 19926 16356 19932
rect 16764 19984 16816 19990
rect 16764 19926 16816 19932
rect 16120 19916 16172 19922
rect 16120 19858 16172 19864
rect 16672 19916 16724 19922
rect 16672 19858 16724 19864
rect 17224 19916 17276 19922
rect 17224 19858 17276 19864
rect 17776 19916 17828 19922
rect 17776 19858 17828 19864
rect 16132 19514 16160 19858
rect 16120 19508 16172 19514
rect 16120 19450 16172 19456
rect 16684 19446 16712 19858
rect 17236 19514 17264 19858
rect 17788 19514 17816 19858
rect 18064 19514 18092 20266
rect 18144 19916 18196 19922
rect 18144 19858 18196 19864
rect 17224 19508 17276 19514
rect 17224 19450 17276 19456
rect 17776 19508 17828 19514
rect 17776 19450 17828 19456
rect 18052 19508 18104 19514
rect 18052 19450 18104 19456
rect 16672 19440 16724 19446
rect 16672 19382 16724 19388
rect 15568 19372 15620 19378
rect 15568 19314 15620 19320
rect 15292 19304 15344 19310
rect 15292 19246 15344 19252
rect 16488 19304 16540 19310
rect 16488 19246 16540 19252
rect 17316 19304 17368 19310
rect 17316 19246 17368 19252
rect 17868 19304 17920 19310
rect 17868 19246 17920 19252
rect 17960 19304 18012 19310
rect 17960 19246 18012 19252
rect 15200 19168 15252 19174
rect 15200 19110 15252 19116
rect 14817 19068 15113 19088
rect 14873 19066 14897 19068
rect 14953 19066 14977 19068
rect 15033 19066 15057 19068
rect 14895 19014 14897 19066
rect 14959 19014 14971 19066
rect 15033 19014 15035 19066
rect 14873 19012 14897 19014
rect 14953 19012 14977 19014
rect 15033 19012 15057 19014
rect 14817 18992 15113 19012
rect 14280 18964 14332 18970
rect 14280 18906 14332 18912
rect 14292 14278 14320 18906
rect 16304 18896 16356 18902
rect 16304 18838 16356 18844
rect 14372 18760 14424 18766
rect 14370 18728 14372 18737
rect 14424 18728 14426 18737
rect 14370 18663 14426 18672
rect 14740 18692 14792 18698
rect 14740 18634 14792 18640
rect 14752 17882 14780 18634
rect 15844 18624 15896 18630
rect 15844 18566 15896 18572
rect 16028 18624 16080 18630
rect 16028 18566 16080 18572
rect 15856 18222 15884 18566
rect 16040 18290 16068 18566
rect 16028 18284 16080 18290
rect 16028 18226 16080 18232
rect 15844 18216 15896 18222
rect 15844 18158 15896 18164
rect 16212 18080 16264 18086
rect 16212 18022 16264 18028
rect 14817 17980 15113 18000
rect 14873 17978 14897 17980
rect 14953 17978 14977 17980
rect 15033 17978 15057 17980
rect 14895 17926 14897 17978
rect 14959 17926 14971 17978
rect 15033 17926 15035 17978
rect 14873 17924 14897 17926
rect 14953 17924 14977 17926
rect 15033 17924 15057 17926
rect 14817 17904 15113 17924
rect 14740 17876 14792 17882
rect 14740 17818 14792 17824
rect 15384 17876 15436 17882
rect 15384 17818 15436 17824
rect 15290 17776 15346 17785
rect 15290 17711 15292 17720
rect 15344 17711 15346 17720
rect 15292 17682 15344 17688
rect 14372 17672 14424 17678
rect 14372 17614 14424 17620
rect 14384 17134 14412 17614
rect 15200 17604 15252 17610
rect 15200 17546 15252 17552
rect 14464 17536 14516 17542
rect 14464 17478 14516 17484
rect 14372 17128 14424 17134
rect 14372 17070 14424 17076
rect 14384 16046 14412 17070
rect 14476 16590 14504 17478
rect 15212 17066 15240 17546
rect 15304 17066 15332 17682
rect 15396 17134 15424 17818
rect 15752 17740 15804 17746
rect 15752 17682 15804 17688
rect 15384 17128 15436 17134
rect 15384 17070 15436 17076
rect 15200 17060 15252 17066
rect 15200 17002 15252 17008
rect 15292 17060 15344 17066
rect 15292 17002 15344 17008
rect 14817 16892 15113 16912
rect 14873 16890 14897 16892
rect 14953 16890 14977 16892
rect 15033 16890 15057 16892
rect 14895 16838 14897 16890
rect 14959 16838 14971 16890
rect 15033 16838 15035 16890
rect 14873 16836 14897 16838
rect 14953 16836 14977 16838
rect 15033 16836 15057 16838
rect 14817 16816 15113 16836
rect 15212 16590 15240 17002
rect 14464 16584 14516 16590
rect 14464 16526 14516 16532
rect 15200 16584 15252 16590
rect 15200 16526 15252 16532
rect 15292 16584 15344 16590
rect 15292 16526 15344 16532
rect 14372 16040 14424 16046
rect 14372 15982 14424 15988
rect 14384 14958 14412 15982
rect 14372 14952 14424 14958
rect 14372 14894 14424 14900
rect 14476 14822 14504 16526
rect 15212 16250 15240 16526
rect 15200 16244 15252 16250
rect 15200 16186 15252 16192
rect 14556 15972 14608 15978
rect 14556 15914 14608 15920
rect 14568 15434 14596 15914
rect 15304 15910 15332 16526
rect 15396 16454 15424 17070
rect 15476 17060 15528 17066
rect 15476 17002 15528 17008
rect 15384 16448 15436 16454
rect 15384 16390 15436 16396
rect 15292 15904 15344 15910
rect 15292 15846 15344 15852
rect 14817 15804 15113 15824
rect 14873 15802 14897 15804
rect 14953 15802 14977 15804
rect 15033 15802 15057 15804
rect 14895 15750 14897 15802
rect 14959 15750 14971 15802
rect 15033 15750 15035 15802
rect 14873 15748 14897 15750
rect 14953 15748 14977 15750
rect 15033 15748 15057 15750
rect 14817 15728 15113 15748
rect 15304 15706 15332 15846
rect 15292 15700 15344 15706
rect 15292 15642 15344 15648
rect 14740 15632 14792 15638
rect 14740 15574 14792 15580
rect 14648 15564 14700 15570
rect 14648 15506 14700 15512
rect 14556 15428 14608 15434
rect 14556 15370 14608 15376
rect 14464 14816 14516 14822
rect 14464 14758 14516 14764
rect 14660 14618 14688 15506
rect 14752 15162 14780 15574
rect 15108 15360 15160 15366
rect 15108 15302 15160 15308
rect 14740 15156 14792 15162
rect 14740 15098 14792 15104
rect 14740 15020 14792 15026
rect 14740 14962 14792 14968
rect 14648 14612 14700 14618
rect 14648 14554 14700 14560
rect 14280 14272 14332 14278
rect 14280 14214 14332 14220
rect 14372 14272 14424 14278
rect 14372 14214 14424 14220
rect 14384 14090 14412 14214
rect 14292 14062 14412 14090
rect 14292 13938 14320 14062
rect 14280 13932 14332 13938
rect 14280 13874 14332 13880
rect 14372 12912 14424 12918
rect 14372 12854 14424 12860
rect 14384 12102 14412 12854
rect 14660 12782 14688 14554
rect 14752 14482 14780 14962
rect 15120 14906 15148 15302
rect 15384 15020 15436 15026
rect 15384 14962 15436 14968
rect 15120 14878 15240 14906
rect 14817 14716 15113 14736
rect 14873 14714 14897 14716
rect 14953 14714 14977 14716
rect 15033 14714 15057 14716
rect 14895 14662 14897 14714
rect 14959 14662 14971 14714
rect 15033 14662 15035 14714
rect 14873 14660 14897 14662
rect 14953 14660 14977 14662
rect 15033 14660 15057 14662
rect 14817 14640 15113 14660
rect 15212 14618 15240 14878
rect 15396 14618 15424 14962
rect 15200 14612 15252 14618
rect 15200 14554 15252 14560
rect 15384 14612 15436 14618
rect 15384 14554 15436 14560
rect 14740 14476 14792 14482
rect 14740 14418 14792 14424
rect 14752 13870 14780 14418
rect 15488 14278 15516 17002
rect 15764 16794 15792 17682
rect 16224 17610 16252 18022
rect 16316 17678 16344 18838
rect 16396 18828 16448 18834
rect 16396 18770 16448 18776
rect 16408 17882 16436 18770
rect 16396 17876 16448 17882
rect 16396 17818 16448 17824
rect 16304 17672 16356 17678
rect 16304 17614 16356 17620
rect 16212 17604 16264 17610
rect 16212 17546 16264 17552
rect 16316 17338 16344 17614
rect 16304 17332 16356 17338
rect 16304 17274 16356 17280
rect 15752 16788 15804 16794
rect 15752 16730 15804 16736
rect 15936 16652 15988 16658
rect 15936 16594 15988 16600
rect 15948 16114 15976 16594
rect 15936 16108 15988 16114
rect 15936 16050 15988 16056
rect 15948 15706 15976 16050
rect 15936 15700 15988 15706
rect 15936 15642 15988 15648
rect 16028 15564 16080 15570
rect 16028 15506 16080 15512
rect 16040 15026 16068 15506
rect 16028 15020 16080 15026
rect 16028 14962 16080 14968
rect 15844 14816 15896 14822
rect 15844 14758 15896 14764
rect 16120 14816 16172 14822
rect 16120 14758 16172 14764
rect 16212 14816 16264 14822
rect 16212 14758 16264 14764
rect 15660 14476 15712 14482
rect 15660 14418 15712 14424
rect 15200 14272 15252 14278
rect 15200 14214 15252 14220
rect 15476 14272 15528 14278
rect 15476 14214 15528 14220
rect 14740 13864 14792 13870
rect 14740 13806 14792 13812
rect 14752 12918 14780 13806
rect 14817 13628 15113 13648
rect 14873 13626 14897 13628
rect 14953 13626 14977 13628
rect 15033 13626 15057 13628
rect 14895 13574 14897 13626
rect 14959 13574 14971 13626
rect 15033 13574 15035 13626
rect 14873 13572 14897 13574
rect 14953 13572 14977 13574
rect 15033 13572 15057 13574
rect 14817 13552 15113 13572
rect 14740 12912 14792 12918
rect 14740 12854 14792 12860
rect 14648 12776 14700 12782
rect 14648 12718 14700 12724
rect 14817 12540 15113 12560
rect 14873 12538 14897 12540
rect 14953 12538 14977 12540
rect 15033 12538 15057 12540
rect 14895 12486 14897 12538
rect 14959 12486 14971 12538
rect 15033 12486 15035 12538
rect 14873 12484 14897 12486
rect 14953 12484 14977 12486
rect 15033 12484 15057 12486
rect 14817 12464 15113 12484
rect 14372 12096 14424 12102
rect 14372 12038 14424 12044
rect 14188 11892 14240 11898
rect 14188 11834 14240 11840
rect 14280 11756 14332 11762
rect 14280 11698 14332 11704
rect 14292 11286 14320 11698
rect 15212 11694 15240 14214
rect 15672 13938 15700 14418
rect 15856 13938 15884 14758
rect 16132 14074 16160 14758
rect 16120 14068 16172 14074
rect 16120 14010 16172 14016
rect 15660 13932 15712 13938
rect 15660 13874 15712 13880
rect 15844 13932 15896 13938
rect 15844 13874 15896 13880
rect 15476 13728 15528 13734
rect 15476 13670 15528 13676
rect 15488 13530 15516 13670
rect 15476 13524 15528 13530
rect 15476 13466 15528 13472
rect 15672 12986 15700 13874
rect 16224 13530 16252 14758
rect 16212 13524 16264 13530
rect 16212 13466 16264 13472
rect 15660 12980 15712 12986
rect 15660 12922 15712 12928
rect 16120 12708 16172 12714
rect 16120 12650 16172 12656
rect 15292 12300 15344 12306
rect 15292 12242 15344 12248
rect 15304 11762 15332 12242
rect 15844 12232 15896 12238
rect 15844 12174 15896 12180
rect 15856 11898 15884 12174
rect 16132 12170 16160 12650
rect 16500 12442 16528 19246
rect 16764 18828 16816 18834
rect 16764 18770 16816 18776
rect 16672 18284 16724 18290
rect 16672 18226 16724 18232
rect 16684 16182 16712 18226
rect 16776 18154 16804 18770
rect 17328 18426 17356 19246
rect 17880 18970 17908 19246
rect 17868 18964 17920 18970
rect 17868 18906 17920 18912
rect 17684 18828 17736 18834
rect 17684 18770 17736 18776
rect 17500 18760 17552 18766
rect 17500 18702 17552 18708
rect 17316 18420 17368 18426
rect 17316 18362 17368 18368
rect 17512 18358 17540 18702
rect 17500 18352 17552 18358
rect 17500 18294 17552 18300
rect 17132 18216 17184 18222
rect 17132 18158 17184 18164
rect 16764 18148 16816 18154
rect 16764 18090 16816 18096
rect 16776 16454 16804 18090
rect 16764 16448 16816 16454
rect 16764 16390 16816 16396
rect 16672 16176 16724 16182
rect 16672 16118 16724 16124
rect 16580 15972 16632 15978
rect 16580 15914 16632 15920
rect 16592 13530 16620 15914
rect 16684 15366 16712 16118
rect 16776 15638 16804 16390
rect 16764 15632 16816 15638
rect 16764 15574 16816 15580
rect 16672 15360 16724 15366
rect 16672 15302 16724 15308
rect 16776 14482 16804 15574
rect 17144 15162 17172 18158
rect 17316 16992 17368 16998
rect 17316 16934 17368 16940
rect 17224 16720 17276 16726
rect 17224 16662 17276 16668
rect 17236 16114 17264 16662
rect 17224 16108 17276 16114
rect 17224 16050 17276 16056
rect 17328 16046 17356 16934
rect 17316 16040 17368 16046
rect 17316 15982 17368 15988
rect 17132 15156 17184 15162
rect 17132 15098 17184 15104
rect 17512 14906 17540 18294
rect 17592 16448 17644 16454
rect 17592 16390 17644 16396
rect 17604 15978 17632 16390
rect 17696 16250 17724 18770
rect 17972 18426 18000 19246
rect 18156 18698 18184 19858
rect 18282 19612 18578 19632
rect 18338 19610 18362 19612
rect 18418 19610 18442 19612
rect 18498 19610 18522 19612
rect 18360 19558 18362 19610
rect 18424 19558 18436 19610
rect 18498 19558 18500 19610
rect 18338 19556 18362 19558
rect 18418 19556 18442 19558
rect 18498 19556 18522 19558
rect 18282 19536 18578 19556
rect 18616 19514 18644 20266
rect 18880 20256 18932 20262
rect 18880 20198 18932 20204
rect 18696 19916 18748 19922
rect 18696 19858 18748 19864
rect 18604 19508 18656 19514
rect 18604 19450 18656 19456
rect 18328 19304 18380 19310
rect 18328 19246 18380 19252
rect 18340 18970 18368 19246
rect 18328 18964 18380 18970
rect 18328 18906 18380 18912
rect 18604 18828 18656 18834
rect 18604 18770 18656 18776
rect 18144 18692 18196 18698
rect 18144 18634 18196 18640
rect 18282 18524 18578 18544
rect 18338 18522 18362 18524
rect 18418 18522 18442 18524
rect 18498 18522 18522 18524
rect 18360 18470 18362 18522
rect 18424 18470 18436 18522
rect 18498 18470 18500 18522
rect 18338 18468 18362 18470
rect 18418 18468 18442 18470
rect 18498 18468 18522 18470
rect 18282 18448 18578 18468
rect 17960 18420 18012 18426
rect 17960 18362 18012 18368
rect 18052 18352 18104 18358
rect 18052 18294 18104 18300
rect 17960 17604 18012 17610
rect 17960 17546 18012 17552
rect 17776 17128 17828 17134
rect 17776 17070 17828 17076
rect 17788 16590 17816 17070
rect 17972 17066 18000 17546
rect 17960 17060 18012 17066
rect 17960 17002 18012 17008
rect 18064 16998 18092 18294
rect 18144 18216 18196 18222
rect 18144 18158 18196 18164
rect 18156 17338 18184 18158
rect 18282 17436 18578 17456
rect 18338 17434 18362 17436
rect 18418 17434 18442 17436
rect 18498 17434 18522 17436
rect 18360 17382 18362 17434
rect 18424 17382 18436 17434
rect 18498 17382 18500 17434
rect 18338 17380 18362 17382
rect 18418 17380 18442 17382
rect 18498 17380 18522 17382
rect 18282 17360 18578 17380
rect 18144 17332 18196 17338
rect 18144 17274 18196 17280
rect 18052 16992 18104 16998
rect 18052 16934 18104 16940
rect 18144 16720 18196 16726
rect 18144 16662 18196 16668
rect 17776 16584 17828 16590
rect 17776 16526 17828 16532
rect 17684 16244 17736 16250
rect 17684 16186 17736 16192
rect 17788 15978 17816 16526
rect 17592 15972 17644 15978
rect 17592 15914 17644 15920
rect 17776 15972 17828 15978
rect 17776 15914 17828 15920
rect 17788 15026 17816 15914
rect 18156 15638 18184 16662
rect 18282 16348 18578 16368
rect 18338 16346 18362 16348
rect 18418 16346 18442 16348
rect 18498 16346 18522 16348
rect 18360 16294 18362 16346
rect 18424 16294 18436 16346
rect 18498 16294 18500 16346
rect 18338 16292 18362 16294
rect 18418 16292 18442 16294
rect 18498 16292 18522 16294
rect 18282 16272 18578 16292
rect 18236 15904 18288 15910
rect 18236 15846 18288 15852
rect 17960 15632 18012 15638
rect 17960 15574 18012 15580
rect 18144 15632 18196 15638
rect 18144 15574 18196 15580
rect 17972 15450 18000 15574
rect 17880 15422 18000 15450
rect 18144 15496 18196 15502
rect 18144 15438 18196 15444
rect 18052 15428 18104 15434
rect 17776 15020 17828 15026
rect 17776 14962 17828 14968
rect 17512 14878 17632 14906
rect 16948 14816 17000 14822
rect 16948 14758 17000 14764
rect 17500 14816 17552 14822
rect 17500 14758 17552 14764
rect 16960 14550 16988 14758
rect 17408 14612 17460 14618
rect 17408 14554 17460 14560
rect 16948 14544 17000 14550
rect 16948 14486 17000 14492
rect 16764 14476 16816 14482
rect 16764 14418 16816 14424
rect 17420 14006 17448 14554
rect 17408 14000 17460 14006
rect 17408 13942 17460 13948
rect 16580 13524 16632 13530
rect 16580 13466 16632 13472
rect 17224 13456 17276 13462
rect 17224 13398 17276 13404
rect 16488 12436 16540 12442
rect 16488 12378 16540 12384
rect 16304 12300 16356 12306
rect 16304 12242 16356 12248
rect 16120 12164 16172 12170
rect 16120 12106 16172 12112
rect 15844 11892 15896 11898
rect 15844 11834 15896 11840
rect 16316 11762 16344 12242
rect 16488 11824 16540 11830
rect 16488 11766 16540 11772
rect 15292 11756 15344 11762
rect 15292 11698 15344 11704
rect 16304 11756 16356 11762
rect 16304 11698 16356 11704
rect 15200 11688 15252 11694
rect 15200 11630 15252 11636
rect 14464 11552 14516 11558
rect 14464 11494 14516 11500
rect 14476 11354 14504 11494
rect 14817 11452 15113 11472
rect 14873 11450 14897 11452
rect 14953 11450 14977 11452
rect 15033 11450 15057 11452
rect 14895 11398 14897 11450
rect 14959 11398 14971 11450
rect 15033 11398 15035 11450
rect 14873 11396 14897 11398
rect 14953 11396 14977 11398
rect 15033 11396 15057 11398
rect 14817 11376 15113 11396
rect 15304 11354 15332 11698
rect 14464 11348 14516 11354
rect 14464 11290 14516 11296
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 16500 11286 16528 11766
rect 14280 11280 14332 11286
rect 14280 11222 14332 11228
rect 14924 11280 14976 11286
rect 14924 11222 14976 11228
rect 16488 11280 16540 11286
rect 16488 11222 16540 11228
rect 14936 10810 14964 11222
rect 14924 10804 14976 10810
rect 14924 10746 14976 10752
rect 16500 10674 16528 11222
rect 16488 10668 16540 10674
rect 16488 10610 16540 10616
rect 15200 10532 15252 10538
rect 15200 10474 15252 10480
rect 14817 10364 15113 10384
rect 14873 10362 14897 10364
rect 14953 10362 14977 10364
rect 15033 10362 15057 10364
rect 14895 10310 14897 10362
rect 14959 10310 14971 10362
rect 15033 10310 15035 10362
rect 14873 10308 14897 10310
rect 14953 10308 14977 10310
rect 15033 10308 15057 10310
rect 14817 10288 15113 10308
rect 15212 10266 15240 10474
rect 15752 10464 15804 10470
rect 15752 10406 15804 10412
rect 16120 10464 16172 10470
rect 16120 10406 16172 10412
rect 16948 10464 17000 10470
rect 16948 10406 17000 10412
rect 15200 10260 15252 10266
rect 15200 10202 15252 10208
rect 15764 10198 15792 10406
rect 16132 10198 16160 10406
rect 16960 10266 16988 10406
rect 16948 10260 17000 10266
rect 16948 10202 17000 10208
rect 15752 10192 15804 10198
rect 15752 10134 15804 10140
rect 16120 10192 16172 10198
rect 16120 10134 16172 10140
rect 14096 9376 14148 9382
rect 14096 9318 14148 9324
rect 14817 9276 15113 9296
rect 14873 9274 14897 9276
rect 14953 9274 14977 9276
rect 15033 9274 15057 9276
rect 14895 9222 14897 9274
rect 14959 9222 14971 9274
rect 15033 9222 15035 9274
rect 14873 9220 14897 9222
rect 14953 9220 14977 9222
rect 15033 9220 15057 9222
rect 14817 9200 15113 9220
rect 13084 8492 13136 8498
rect 13084 8434 13136 8440
rect 14817 8188 15113 8208
rect 14873 8186 14897 8188
rect 14953 8186 14977 8188
rect 15033 8186 15057 8188
rect 14895 8134 14897 8186
rect 14959 8134 14971 8186
rect 15033 8134 15035 8186
rect 14873 8132 14897 8134
rect 14953 8132 14977 8134
rect 15033 8132 15057 8134
rect 14817 8112 15113 8132
rect 17236 7478 17264 13398
rect 17316 12844 17368 12850
rect 17316 12786 17368 12792
rect 17328 12646 17356 12786
rect 17316 12640 17368 12646
rect 17316 12582 17368 12588
rect 17328 12306 17356 12582
rect 17316 12300 17368 12306
rect 17316 12242 17368 12248
rect 17328 11218 17356 12242
rect 17316 11212 17368 11218
rect 17316 11154 17368 11160
rect 17512 8906 17540 14758
rect 17604 13190 17632 14878
rect 17880 14822 17908 15422
rect 18052 15370 18104 15376
rect 17960 15360 18012 15366
rect 17960 15302 18012 15308
rect 17868 14816 17920 14822
rect 17868 14758 17920 14764
rect 17972 14618 18000 15302
rect 18064 14958 18092 15370
rect 18052 14952 18104 14958
rect 18052 14894 18104 14900
rect 18156 14618 18184 15438
rect 18248 15434 18276 15846
rect 18236 15428 18288 15434
rect 18236 15370 18288 15376
rect 18282 15260 18578 15280
rect 18338 15258 18362 15260
rect 18418 15258 18442 15260
rect 18498 15258 18522 15260
rect 18360 15206 18362 15258
rect 18424 15206 18436 15258
rect 18498 15206 18500 15258
rect 18338 15204 18362 15206
rect 18418 15204 18442 15206
rect 18498 15204 18522 15206
rect 18282 15184 18578 15204
rect 18616 14618 18644 18770
rect 17960 14612 18012 14618
rect 17960 14554 18012 14560
rect 18144 14612 18196 14618
rect 18144 14554 18196 14560
rect 18604 14612 18656 14618
rect 18604 14554 18656 14560
rect 18282 14172 18578 14192
rect 18338 14170 18362 14172
rect 18418 14170 18442 14172
rect 18498 14170 18522 14172
rect 18360 14118 18362 14170
rect 18424 14118 18436 14170
rect 18498 14118 18500 14170
rect 18338 14116 18362 14118
rect 18418 14116 18442 14118
rect 18498 14116 18522 14118
rect 18282 14096 18578 14116
rect 18052 14000 18104 14006
rect 18052 13942 18104 13948
rect 17776 13728 17828 13734
rect 17776 13670 17828 13676
rect 17788 13326 17816 13670
rect 17960 13388 18012 13394
rect 17960 13330 18012 13336
rect 17776 13320 17828 13326
rect 17776 13262 17828 13268
rect 17592 13184 17644 13190
rect 17592 13126 17644 13132
rect 17604 12782 17632 13126
rect 17788 12850 17816 13262
rect 17776 12844 17828 12850
rect 17776 12786 17828 12792
rect 17592 12776 17644 12782
rect 17592 12718 17644 12724
rect 17788 12374 17816 12786
rect 17972 12442 18000 13330
rect 18064 12850 18092 13942
rect 18282 13084 18578 13104
rect 18338 13082 18362 13084
rect 18418 13082 18442 13084
rect 18498 13082 18522 13084
rect 18360 13030 18362 13082
rect 18424 13030 18436 13082
rect 18498 13030 18500 13082
rect 18338 13028 18362 13030
rect 18418 13028 18442 13030
rect 18498 13028 18522 13030
rect 18282 13008 18578 13028
rect 18052 12844 18104 12850
rect 18052 12786 18104 12792
rect 17960 12436 18012 12442
rect 17960 12378 18012 12384
rect 17776 12368 17828 12374
rect 17776 12310 17828 12316
rect 18282 11996 18578 12016
rect 18338 11994 18362 11996
rect 18418 11994 18442 11996
rect 18498 11994 18522 11996
rect 18360 11942 18362 11994
rect 18424 11942 18436 11994
rect 18498 11942 18500 11994
rect 18338 11940 18362 11942
rect 18418 11940 18442 11942
rect 18498 11940 18522 11942
rect 18282 11920 18578 11940
rect 17592 11008 17644 11014
rect 17592 10950 17644 10956
rect 17604 10538 17632 10950
rect 18282 10908 18578 10928
rect 18338 10906 18362 10908
rect 18418 10906 18442 10908
rect 18498 10906 18522 10908
rect 18360 10854 18362 10906
rect 18424 10854 18436 10906
rect 18498 10854 18500 10906
rect 18338 10852 18362 10854
rect 18418 10852 18442 10854
rect 18498 10852 18522 10854
rect 18282 10832 18578 10852
rect 17592 10532 17644 10538
rect 17592 10474 17644 10480
rect 17604 10062 17632 10474
rect 18708 10266 18736 19858
rect 18788 18828 18840 18834
rect 18788 18770 18840 18776
rect 18800 12986 18828 18770
rect 18788 12980 18840 12986
rect 18788 12922 18840 12928
rect 18788 12164 18840 12170
rect 18788 12106 18840 12112
rect 18800 11694 18828 12106
rect 18788 11688 18840 11694
rect 18788 11630 18840 11636
rect 18696 10260 18748 10266
rect 18696 10202 18748 10208
rect 17592 10056 17644 10062
rect 17592 9998 17644 10004
rect 18282 9820 18578 9840
rect 18338 9818 18362 9820
rect 18418 9818 18442 9820
rect 18498 9818 18522 9820
rect 18360 9766 18362 9818
rect 18424 9766 18436 9818
rect 18498 9766 18500 9818
rect 18338 9764 18362 9766
rect 18418 9764 18442 9766
rect 18498 9764 18522 9766
rect 18282 9744 18578 9764
rect 17500 8900 17552 8906
rect 17500 8842 17552 8848
rect 18282 8732 18578 8752
rect 18338 8730 18362 8732
rect 18418 8730 18442 8732
rect 18498 8730 18522 8732
rect 18360 8678 18362 8730
rect 18424 8678 18436 8730
rect 18498 8678 18500 8730
rect 18338 8676 18362 8678
rect 18418 8676 18442 8678
rect 18498 8676 18522 8678
rect 18282 8656 18578 8676
rect 18282 7644 18578 7664
rect 18338 7642 18362 7644
rect 18418 7642 18442 7644
rect 18498 7642 18522 7644
rect 18360 7590 18362 7642
rect 18424 7590 18436 7642
rect 18498 7590 18500 7642
rect 18338 7588 18362 7590
rect 18418 7588 18442 7590
rect 18498 7588 18522 7590
rect 18282 7568 18578 7588
rect 18892 7546 18920 20198
rect 18984 20058 19012 20266
rect 19248 20256 19300 20262
rect 19248 20198 19300 20204
rect 18972 20052 19024 20058
rect 18972 19994 19024 20000
rect 19156 19984 19208 19990
rect 19156 19926 19208 19932
rect 18972 19712 19024 19718
rect 18972 19654 19024 19660
rect 18984 19310 19012 19654
rect 18972 19304 19024 19310
rect 18972 19246 19024 19252
rect 19168 18630 19196 19926
rect 19260 19786 19288 20198
rect 19248 19780 19300 19786
rect 19248 19722 19300 19728
rect 19352 19174 19380 20334
rect 19996 19990 20024 22200
rect 20456 19990 20484 22200
rect 20916 19990 20944 22200
rect 21376 20466 21404 22200
rect 21364 20460 21416 20466
rect 21364 20402 21416 20408
rect 21836 20330 21864 22200
rect 21824 20324 21876 20330
rect 21824 20266 21876 20272
rect 21180 20256 21232 20262
rect 21180 20198 21232 20204
rect 19984 19984 20036 19990
rect 19984 19926 20036 19932
rect 20444 19984 20496 19990
rect 20444 19926 20496 19932
rect 20904 19984 20956 19990
rect 20904 19926 20956 19932
rect 19708 19916 19760 19922
rect 19708 19858 19760 19864
rect 19432 19848 19484 19854
rect 19432 19790 19484 19796
rect 19444 19514 19472 19790
rect 19432 19508 19484 19514
rect 19432 19450 19484 19456
rect 19340 19168 19392 19174
rect 19340 19110 19392 19116
rect 19156 18624 19208 18630
rect 19156 18566 19208 18572
rect 18972 17536 19024 17542
rect 18972 17478 19024 17484
rect 18984 17202 19012 17478
rect 19340 17264 19392 17270
rect 19340 17206 19392 17212
rect 18972 17196 19024 17202
rect 18972 17138 19024 17144
rect 19156 17060 19208 17066
rect 19156 17002 19208 17008
rect 19168 16794 19196 17002
rect 19156 16788 19208 16794
rect 19156 16730 19208 16736
rect 19352 16046 19380 17206
rect 19340 16040 19392 16046
rect 19340 15982 19392 15988
rect 19064 14816 19116 14822
rect 19064 14758 19116 14764
rect 19076 14414 19104 14758
rect 19064 14408 19116 14414
rect 19064 14350 19116 14356
rect 19076 13870 19104 14350
rect 19064 13864 19116 13870
rect 19064 13806 19116 13812
rect 19248 13864 19300 13870
rect 19248 13806 19300 13812
rect 18972 13184 19024 13190
rect 18972 13126 19024 13132
rect 18984 12782 19012 13126
rect 19156 12844 19208 12850
rect 19156 12786 19208 12792
rect 18972 12776 19024 12782
rect 18972 12718 19024 12724
rect 19168 12170 19196 12786
rect 19260 12374 19288 13806
rect 19248 12368 19300 12374
rect 19248 12310 19300 12316
rect 19156 12164 19208 12170
rect 19156 12106 19208 12112
rect 19260 11762 19288 12310
rect 19248 11756 19300 11762
rect 19248 11698 19300 11704
rect 19260 10674 19288 11698
rect 19248 10668 19300 10674
rect 19248 10610 19300 10616
rect 19720 7546 19748 19858
rect 19984 19848 20036 19854
rect 19984 19790 20036 19796
rect 19800 19780 19852 19786
rect 19800 19722 19852 19728
rect 19812 12434 19840 19722
rect 19892 17672 19944 17678
rect 19892 17614 19944 17620
rect 19904 17134 19932 17614
rect 19892 17128 19944 17134
rect 19892 17070 19944 17076
rect 19892 16448 19944 16454
rect 19892 16390 19944 16396
rect 19904 16250 19932 16390
rect 19892 16244 19944 16250
rect 19892 16186 19944 16192
rect 19812 12406 19932 12434
rect 18880 7540 18932 7546
rect 18880 7482 18932 7488
rect 19708 7540 19760 7546
rect 19708 7482 19760 7488
rect 17224 7472 17276 7478
rect 17224 7414 17276 7420
rect 18788 7336 18840 7342
rect 18786 7304 18788 7313
rect 19064 7336 19116 7342
rect 18840 7304 18842 7313
rect 19064 7278 19116 7284
rect 18786 7239 18842 7248
rect 14817 7100 15113 7120
rect 14873 7098 14897 7100
rect 14953 7098 14977 7100
rect 15033 7098 15057 7100
rect 14895 7046 14897 7098
rect 14959 7046 14971 7098
rect 15033 7046 15035 7098
rect 14873 7044 14897 7046
rect 14953 7044 14977 7046
rect 15033 7044 15057 7046
rect 14817 7024 15113 7044
rect 19076 6662 19104 7278
rect 19800 6860 19852 6866
rect 19800 6802 19852 6808
rect 19064 6656 19116 6662
rect 19064 6598 19116 6604
rect 18282 6556 18578 6576
rect 18338 6554 18362 6556
rect 18418 6554 18442 6556
rect 18498 6554 18522 6556
rect 18360 6502 18362 6554
rect 18424 6502 18436 6554
rect 18498 6502 18500 6554
rect 18338 6500 18362 6502
rect 18418 6500 18442 6502
rect 18498 6500 18522 6502
rect 18282 6480 18578 6500
rect 14817 6012 15113 6032
rect 14873 6010 14897 6012
rect 14953 6010 14977 6012
rect 15033 6010 15057 6012
rect 14895 5958 14897 6010
rect 14959 5958 14971 6010
rect 15033 5958 15035 6010
rect 14873 5956 14897 5958
rect 14953 5956 14977 5958
rect 15033 5956 15057 5958
rect 14817 5936 15113 5956
rect 19812 5914 19840 6802
rect 19904 6458 19932 12406
rect 19996 6730 20024 19790
rect 20720 19236 20772 19242
rect 20720 19178 20772 19184
rect 20536 18624 20588 18630
rect 20536 18566 20588 18572
rect 19984 6724 20036 6730
rect 19984 6666 20036 6672
rect 19892 6452 19944 6458
rect 19892 6394 19944 6400
rect 20076 6248 20128 6254
rect 20076 6190 20128 6196
rect 19800 5908 19852 5914
rect 19800 5850 19852 5856
rect 20088 5642 20116 6190
rect 20548 5914 20576 18566
rect 20732 14074 20760 19178
rect 20812 19168 20864 19174
rect 20812 19110 20864 19116
rect 20720 14068 20772 14074
rect 20720 14010 20772 14016
rect 20536 5908 20588 5914
rect 20536 5850 20588 5856
rect 20076 5636 20128 5642
rect 20076 5578 20128 5584
rect 18282 5468 18578 5488
rect 18338 5466 18362 5468
rect 18418 5466 18442 5468
rect 18498 5466 18522 5468
rect 18360 5414 18362 5466
rect 18424 5414 18436 5466
rect 18498 5414 18500 5466
rect 18338 5412 18362 5414
rect 18418 5412 18442 5414
rect 18498 5412 18522 5414
rect 18282 5392 18578 5412
rect 20824 5370 20852 19110
rect 21192 18766 21220 20198
rect 22296 19310 22324 22200
rect 22756 20398 22784 22200
rect 22744 20392 22796 20398
rect 22744 20334 22796 20340
rect 21364 19304 21416 19310
rect 21364 19246 21416 19252
rect 22284 19304 22336 19310
rect 22284 19246 22336 19252
rect 21376 18970 21404 19246
rect 21364 18964 21416 18970
rect 21364 18906 21416 18912
rect 21180 18760 21232 18766
rect 21180 18702 21232 18708
rect 21088 12300 21140 12306
rect 21088 12242 21140 12248
rect 21100 11898 21128 12242
rect 21088 11892 21140 11898
rect 21088 11834 21140 11840
rect 21364 11688 21416 11694
rect 21364 11630 21416 11636
rect 21376 11529 21404 11630
rect 21362 11520 21418 11529
rect 21362 11455 21418 11464
rect 20812 5364 20864 5370
rect 20812 5306 20864 5312
rect 20996 5160 21048 5166
rect 20996 5102 21048 5108
rect 14817 4924 15113 4944
rect 14873 4922 14897 4924
rect 14953 4922 14977 4924
rect 15033 4922 15057 4924
rect 14895 4870 14897 4922
rect 14959 4870 14971 4922
rect 15033 4870 15035 4922
rect 14873 4868 14897 4870
rect 14953 4868 14977 4870
rect 15033 4868 15057 4870
rect 14817 4848 15113 4868
rect 21008 4486 21036 5102
rect 20996 4480 21048 4486
rect 20996 4422 21048 4428
rect 18282 4380 18578 4400
rect 18338 4378 18362 4380
rect 18418 4378 18442 4380
rect 18498 4378 18522 4380
rect 18360 4326 18362 4378
rect 18424 4326 18436 4378
rect 18498 4326 18500 4378
rect 18338 4324 18362 4326
rect 18418 4324 18442 4326
rect 18498 4324 18522 4326
rect 18282 4304 18578 4324
rect 14817 3836 15113 3856
rect 14873 3834 14897 3836
rect 14953 3834 14977 3836
rect 15033 3834 15057 3836
rect 14895 3782 14897 3834
rect 14959 3782 14971 3834
rect 15033 3782 15035 3834
rect 14873 3780 14897 3782
rect 14953 3780 14977 3782
rect 15033 3780 15057 3782
rect 14817 3760 15113 3780
rect 18282 3292 18578 3312
rect 18338 3290 18362 3292
rect 18418 3290 18442 3292
rect 18498 3290 18522 3292
rect 18360 3238 18362 3290
rect 18424 3238 18436 3290
rect 18498 3238 18500 3290
rect 18338 3236 18362 3238
rect 18418 3236 18442 3238
rect 18498 3236 18522 3238
rect 18282 3216 18578 3236
rect 14817 2748 15113 2768
rect 14873 2746 14897 2748
rect 14953 2746 14977 2748
rect 15033 2746 15057 2748
rect 14895 2694 14897 2746
rect 14959 2694 14971 2746
rect 15033 2694 15035 2746
rect 14873 2692 14897 2694
rect 14953 2692 14977 2694
rect 15033 2692 15057 2694
rect 14817 2672 15113 2692
rect 5448 2576 5500 2582
rect 5448 2518 5500 2524
rect 12256 2576 12308 2582
rect 12256 2518 12308 2524
rect 3976 2372 4028 2378
rect 3976 2314 4028 2320
rect 11704 2372 11756 2378
rect 11704 2314 11756 2320
rect 4421 2204 4717 2224
rect 4477 2202 4501 2204
rect 4557 2202 4581 2204
rect 4637 2202 4661 2204
rect 4499 2150 4501 2202
rect 4563 2150 4575 2202
rect 4637 2150 4639 2202
rect 4477 2148 4501 2150
rect 4557 2148 4581 2150
rect 4637 2148 4661 2150
rect 4421 2128 4717 2148
rect 11352 2204 11648 2224
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11430 2150 11432 2202
rect 11494 2150 11506 2202
rect 11568 2150 11570 2202
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11352 2128 11648 2148
rect 3882 2000 3938 2009
rect 3882 1935 3938 1944
rect 3146 1592 3202 1601
rect 3146 1527 3202 1536
rect 11716 1170 11744 2314
rect 18282 2204 18578 2224
rect 18338 2202 18362 2204
rect 18418 2202 18442 2204
rect 18498 2202 18522 2204
rect 18360 2150 18362 2202
rect 18424 2150 18436 2202
rect 18498 2150 18500 2202
rect 18338 2148 18362 2150
rect 18418 2148 18442 2150
rect 18498 2148 18522 2150
rect 18282 2128 18578 2148
rect 11532 1142 11744 1170
rect 2778 1048 2834 1057
rect 2778 983 2834 992
rect 11532 800 11560 1142
rect 2226 640 2282 649
rect 2226 575 2282 584
rect 2134 232 2190 241
rect 2134 167 2190 176
rect 11518 0 11574 800
<< via2 >>
rect 3974 22616 4030 22672
rect 1582 19780 1638 19816
rect 1582 19760 1584 19780
rect 1584 19760 1636 19780
rect 1636 19760 1638 19780
rect 1582 19352 1638 19408
rect 1582 18828 1638 18864
rect 1582 18808 1584 18828
rect 1584 18808 1636 18828
rect 1636 18808 1638 18828
rect 1674 18420 1730 18456
rect 1674 18400 1676 18420
rect 1676 18400 1728 18420
rect 1728 18400 1730 18420
rect 1582 17060 1638 17096
rect 1582 17040 1584 17060
rect 1584 17040 1636 17060
rect 1636 17040 1638 17060
rect 1582 16496 1638 16552
rect 1582 16108 1638 16144
rect 1582 16088 1584 16108
rect 1584 16088 1636 16108
rect 1636 16088 1638 16108
rect 1582 15564 1638 15600
rect 1582 15544 1584 15564
rect 1584 15544 1636 15564
rect 1636 15544 1638 15564
rect 1674 15156 1730 15192
rect 1674 15136 1676 15156
rect 1676 15136 1728 15156
rect 1728 15136 1730 15156
rect 1674 14220 1676 14240
rect 1676 14220 1728 14240
rect 1728 14220 1730 14240
rect 1674 14184 1730 14220
rect 1582 13812 1584 13832
rect 1584 13812 1636 13832
rect 1636 13812 1638 13832
rect 1582 13776 1638 13812
rect 1490 11328 1546 11384
rect 1398 10512 1454 10568
rect 1398 9968 1454 10024
rect 1398 9052 1400 9072
rect 1400 9052 1452 9072
rect 1452 9052 1454 9072
rect 1398 9016 1454 9052
rect 1858 9460 1860 9480
rect 1860 9460 1912 9480
rect 1912 9460 1914 9480
rect 1858 9424 1914 9460
rect 2962 21664 3018 21720
rect 2870 20712 2926 20768
rect 2778 20476 2780 20496
rect 2780 20476 2832 20496
rect 2832 20476 2834 20496
rect 2778 20440 2834 20476
rect 2778 20304 2834 20360
rect 2226 17484 2228 17504
rect 2228 17484 2280 17504
rect 2280 17484 2282 17504
rect 2226 17448 2282 17484
rect 2226 14612 2282 14648
rect 2226 14592 2228 14612
rect 2228 14592 2280 14612
rect 2280 14592 2282 14612
rect 2502 18672 2558 18728
rect 3054 21256 3110 21312
rect 2778 17992 2834 18048
rect 4066 22208 4122 22264
rect 4421 20698 4477 20700
rect 4501 20698 4557 20700
rect 4581 20698 4637 20700
rect 4661 20698 4717 20700
rect 4421 20646 4447 20698
rect 4447 20646 4477 20698
rect 4501 20646 4511 20698
rect 4511 20646 4557 20698
rect 4581 20646 4627 20698
rect 4627 20646 4637 20698
rect 4661 20646 4691 20698
rect 4691 20646 4717 20698
rect 4421 20644 4477 20646
rect 4501 20644 4557 20646
rect 4581 20644 4637 20646
rect 4661 20644 4717 20646
rect 4158 20460 4214 20496
rect 4158 20440 4160 20460
rect 4160 20440 4212 20460
rect 4212 20440 4214 20460
rect 4066 19252 4068 19272
rect 4068 19252 4120 19272
rect 4120 19252 4122 19272
rect 4066 19216 4122 19252
rect 4618 20032 4674 20088
rect 4421 19610 4477 19612
rect 4501 19610 4557 19612
rect 4581 19610 4637 19612
rect 4661 19610 4717 19612
rect 4421 19558 4447 19610
rect 4447 19558 4477 19610
rect 4501 19558 4511 19610
rect 4511 19558 4557 19610
rect 4581 19558 4627 19610
rect 4627 19558 4637 19610
rect 4661 19558 4691 19610
rect 4691 19558 4717 19610
rect 4421 19556 4477 19558
rect 4501 19556 4557 19558
rect 4581 19556 4637 19558
rect 4661 19556 4717 19558
rect 3330 18128 3386 18184
rect 1858 8064 1914 8120
rect 2870 12280 2926 12336
rect 4421 18522 4477 18524
rect 4501 18522 4557 18524
rect 4581 18522 4637 18524
rect 4661 18522 4717 18524
rect 4421 18470 4447 18522
rect 4447 18470 4477 18522
rect 4501 18470 4511 18522
rect 4511 18470 4557 18522
rect 4581 18470 4627 18522
rect 4627 18470 4637 18522
rect 4661 18470 4691 18522
rect 4691 18470 4717 18522
rect 4421 18468 4477 18470
rect 4501 18468 4557 18470
rect 4581 18468 4637 18470
rect 4661 18468 4717 18470
rect 5078 19216 5134 19272
rect 5354 19780 5410 19816
rect 5354 19760 5356 19780
rect 5356 19760 5408 19780
rect 5408 19760 5410 19780
rect 5078 18536 5134 18592
rect 5814 20576 5870 20632
rect 4421 17434 4477 17436
rect 4501 17434 4557 17436
rect 4581 17434 4637 17436
rect 4661 17434 4717 17436
rect 4421 17382 4447 17434
rect 4447 17382 4477 17434
rect 4501 17382 4511 17434
rect 4511 17382 4557 17434
rect 4581 17382 4627 17434
rect 4627 17382 4637 17434
rect 4661 17382 4691 17434
rect 4691 17382 4717 17434
rect 4421 17380 4477 17382
rect 4501 17380 4557 17382
rect 4581 17380 4637 17382
rect 4661 17380 4717 17382
rect 4421 16346 4477 16348
rect 4501 16346 4557 16348
rect 4581 16346 4637 16348
rect 4661 16346 4717 16348
rect 4421 16294 4447 16346
rect 4447 16294 4477 16346
rect 4501 16294 4511 16346
rect 4511 16294 4557 16346
rect 4581 16294 4627 16346
rect 4627 16294 4637 16346
rect 4661 16294 4691 16346
rect 4691 16294 4717 16346
rect 4421 16292 4477 16294
rect 4501 16292 4557 16294
rect 4581 16292 4637 16294
rect 4661 16292 4717 16294
rect 4066 15952 4122 16008
rect 4618 15988 4620 16008
rect 4620 15988 4672 16008
rect 4672 15988 4674 16008
rect 4618 15952 4674 15988
rect 4421 15258 4477 15260
rect 4501 15258 4557 15260
rect 4581 15258 4637 15260
rect 4661 15258 4717 15260
rect 4421 15206 4447 15258
rect 4447 15206 4477 15258
rect 4501 15206 4511 15258
rect 4511 15206 4557 15258
rect 4581 15206 4627 15258
rect 4627 15206 4637 15258
rect 4661 15206 4691 15258
rect 4691 15206 4717 15258
rect 4421 15204 4477 15206
rect 4501 15204 4557 15206
rect 4581 15204 4637 15206
rect 4661 15204 4717 15206
rect 4421 14170 4477 14172
rect 4501 14170 4557 14172
rect 4581 14170 4637 14172
rect 4661 14170 4717 14172
rect 4421 14118 4447 14170
rect 4447 14118 4477 14170
rect 4501 14118 4511 14170
rect 4511 14118 4557 14170
rect 4581 14118 4627 14170
rect 4627 14118 4637 14170
rect 4661 14118 4691 14170
rect 4691 14118 4717 14170
rect 4421 14116 4477 14118
rect 4501 14116 4557 14118
rect 4581 14116 4637 14118
rect 4661 14116 4717 14118
rect 5078 14048 5134 14104
rect 4342 13912 4398 13968
rect 4066 13232 4122 13288
rect 3606 12824 3662 12880
rect 3146 11872 3202 11928
rect 2870 11600 2926 11656
rect 4421 13082 4477 13084
rect 4501 13082 4557 13084
rect 4581 13082 4637 13084
rect 4661 13082 4717 13084
rect 4421 13030 4447 13082
rect 4447 13030 4477 13082
rect 4501 13030 4511 13082
rect 4511 13030 4557 13082
rect 4581 13030 4627 13082
rect 4627 13030 4637 13082
rect 4661 13030 4691 13082
rect 4691 13030 4717 13082
rect 4421 13028 4477 13030
rect 4501 13028 4557 13030
rect 4581 13028 4637 13030
rect 4661 13028 4717 13030
rect 3422 10920 3478 10976
rect 1398 7656 1454 7712
rect 1582 7248 1638 7304
rect 1398 7112 1454 7168
rect 1398 6704 1454 6760
rect 1398 6196 1400 6216
rect 1400 6196 1452 6216
rect 1452 6196 1454 6216
rect 1398 6160 1454 6196
rect 1398 5772 1454 5808
rect 1398 5752 1400 5772
rect 1400 5752 1452 5772
rect 1452 5752 1454 5772
rect 1398 5208 1454 5264
rect 1858 4800 1914 4856
rect 1398 4392 1454 4448
rect 1674 3848 1730 3904
rect 1674 3440 1730 3496
rect 2778 8608 2834 8664
rect 1766 2932 1768 2952
rect 1768 2932 1820 2952
rect 1820 2932 1822 2952
rect 1766 2896 1822 2932
rect 1674 2508 1730 2544
rect 1674 2488 1676 2508
rect 1676 2488 1728 2508
rect 1728 2488 1730 2508
rect 3882 7384 3938 7440
rect 4421 11994 4477 11996
rect 4501 11994 4557 11996
rect 4581 11994 4637 11996
rect 4661 11994 4717 11996
rect 4421 11942 4447 11994
rect 4447 11942 4477 11994
rect 4501 11942 4511 11994
rect 4511 11942 4557 11994
rect 4581 11942 4627 11994
rect 4627 11942 4637 11994
rect 4661 11942 4691 11994
rect 4691 11942 4717 11994
rect 4421 11940 4477 11942
rect 4501 11940 4557 11942
rect 4581 11940 4637 11942
rect 4661 11940 4717 11942
rect 4421 10906 4477 10908
rect 4501 10906 4557 10908
rect 4581 10906 4637 10908
rect 4661 10906 4717 10908
rect 4421 10854 4447 10906
rect 4447 10854 4477 10906
rect 4501 10854 4511 10906
rect 4511 10854 4557 10906
rect 4581 10854 4627 10906
rect 4627 10854 4637 10906
rect 4661 10854 4691 10906
rect 4691 10854 4717 10906
rect 4421 10852 4477 10854
rect 4501 10852 4557 10854
rect 4581 10852 4637 10854
rect 4661 10852 4717 10854
rect 4421 9818 4477 9820
rect 4501 9818 4557 9820
rect 4581 9818 4637 9820
rect 4661 9818 4717 9820
rect 4421 9766 4447 9818
rect 4447 9766 4477 9818
rect 4501 9766 4511 9818
rect 4511 9766 4557 9818
rect 4581 9766 4627 9818
rect 4627 9766 4637 9818
rect 4661 9766 4691 9818
rect 4691 9766 4717 9818
rect 4421 9764 4477 9766
rect 4501 9764 4557 9766
rect 4581 9764 4637 9766
rect 4661 9764 4717 9766
rect 4421 8730 4477 8732
rect 4501 8730 4557 8732
rect 4581 8730 4637 8732
rect 4661 8730 4717 8732
rect 4421 8678 4447 8730
rect 4447 8678 4477 8730
rect 4501 8678 4511 8730
rect 4511 8678 4557 8730
rect 4581 8678 4627 8730
rect 4627 8678 4637 8730
rect 4661 8678 4691 8730
rect 4691 8678 4717 8730
rect 4421 8676 4477 8678
rect 4501 8676 4557 8678
rect 4581 8676 4637 8678
rect 4661 8676 4717 8678
rect 4421 7642 4477 7644
rect 4501 7642 4557 7644
rect 4581 7642 4637 7644
rect 4661 7642 4717 7644
rect 4421 7590 4447 7642
rect 4447 7590 4477 7642
rect 4501 7590 4511 7642
rect 4511 7590 4557 7642
rect 4581 7590 4627 7642
rect 4627 7590 4637 7642
rect 4661 7590 4691 7642
rect 4691 7590 4717 7642
rect 4421 7588 4477 7590
rect 4501 7588 4557 7590
rect 4581 7588 4637 7590
rect 4661 7588 4717 7590
rect 5630 16632 5686 16688
rect 6550 20460 6606 20496
rect 6550 20440 6552 20460
rect 6552 20440 6604 20460
rect 6604 20440 6606 20460
rect 6090 18536 6146 18592
rect 5998 15952 6054 16008
rect 4421 6554 4477 6556
rect 4501 6554 4557 6556
rect 4581 6554 4637 6556
rect 4661 6554 4717 6556
rect 4421 6502 4447 6554
rect 4447 6502 4477 6554
rect 4501 6502 4511 6554
rect 4511 6502 4557 6554
rect 4581 6502 4627 6554
rect 4627 6502 4637 6554
rect 4661 6502 4691 6554
rect 4691 6502 4717 6554
rect 4421 6500 4477 6502
rect 4501 6500 4557 6502
rect 4581 6500 4637 6502
rect 4661 6500 4717 6502
rect 4421 5466 4477 5468
rect 4501 5466 4557 5468
rect 4581 5466 4637 5468
rect 4661 5466 4717 5468
rect 4421 5414 4447 5466
rect 4447 5414 4477 5466
rect 4501 5414 4511 5466
rect 4511 5414 4557 5466
rect 4581 5414 4627 5466
rect 4627 5414 4637 5466
rect 4661 5414 4691 5466
rect 4691 5414 4717 5466
rect 4421 5412 4477 5414
rect 4501 5412 4557 5414
rect 4581 5412 4637 5414
rect 4661 5412 4717 5414
rect 4421 4378 4477 4380
rect 4501 4378 4557 4380
rect 4581 4378 4637 4380
rect 4661 4378 4717 4380
rect 4421 4326 4447 4378
rect 4447 4326 4477 4378
rect 4501 4326 4511 4378
rect 4511 4326 4557 4378
rect 4581 4326 4627 4378
rect 4627 4326 4637 4378
rect 4661 4326 4691 4378
rect 4691 4326 4717 4378
rect 4421 4324 4477 4326
rect 4501 4324 4557 4326
rect 4581 4324 4637 4326
rect 4661 4324 4717 4326
rect 4421 3290 4477 3292
rect 4501 3290 4557 3292
rect 4581 3290 4637 3292
rect 4661 3290 4717 3292
rect 4421 3238 4447 3290
rect 4447 3238 4477 3290
rect 4501 3238 4511 3290
rect 4511 3238 4557 3290
rect 4581 3238 4627 3290
rect 4627 3238 4637 3290
rect 4661 3238 4691 3290
rect 4691 3238 4717 3290
rect 4421 3236 4477 3238
rect 4501 3236 4557 3238
rect 4581 3236 4637 3238
rect 4661 3236 4717 3238
rect 6090 13948 6092 13968
rect 6092 13948 6144 13968
rect 6144 13948 6146 13968
rect 6090 13912 6146 13948
rect 5906 11736 5962 11792
rect 6826 20440 6882 20496
rect 6642 16652 6698 16688
rect 6642 16632 6644 16652
rect 6644 16632 6696 16652
rect 6696 16632 6698 16652
rect 7286 20052 7342 20088
rect 7286 20032 7288 20052
rect 7288 20032 7340 20052
rect 7340 20032 7342 20052
rect 7654 20596 7710 20632
rect 7654 20576 7656 20596
rect 7656 20576 7708 20596
rect 7708 20576 7710 20596
rect 7886 20154 7942 20156
rect 7966 20154 8022 20156
rect 8046 20154 8102 20156
rect 8126 20154 8182 20156
rect 7886 20102 7912 20154
rect 7912 20102 7942 20154
rect 7966 20102 7976 20154
rect 7976 20102 8022 20154
rect 8046 20102 8092 20154
rect 8092 20102 8102 20154
rect 8126 20102 8156 20154
rect 8156 20102 8182 20154
rect 7886 20100 7942 20102
rect 7966 20100 8022 20102
rect 8046 20100 8102 20102
rect 8126 20100 8182 20102
rect 8390 20052 8446 20088
rect 8390 20032 8392 20052
rect 8392 20032 8444 20052
rect 8444 20032 8446 20052
rect 7886 19066 7942 19068
rect 7966 19066 8022 19068
rect 8046 19066 8102 19068
rect 8126 19066 8182 19068
rect 7886 19014 7912 19066
rect 7912 19014 7942 19066
rect 7966 19014 7976 19066
rect 7976 19014 8022 19066
rect 8046 19014 8092 19066
rect 8092 19014 8102 19066
rect 8126 19014 8156 19066
rect 8156 19014 8182 19066
rect 7886 19012 7942 19014
rect 7966 19012 8022 19014
rect 8046 19012 8102 19014
rect 8126 19012 8182 19014
rect 7886 17978 7942 17980
rect 7966 17978 8022 17980
rect 8046 17978 8102 17980
rect 8126 17978 8182 17980
rect 7886 17926 7912 17978
rect 7912 17926 7942 17978
rect 7966 17926 7976 17978
rect 7976 17926 8022 17978
rect 8046 17926 8092 17978
rect 8092 17926 8102 17978
rect 8126 17926 8156 17978
rect 8156 17926 8182 17978
rect 7886 17924 7942 17926
rect 7966 17924 8022 17926
rect 8046 17924 8102 17926
rect 8126 17924 8182 17926
rect 6642 13096 6698 13152
rect 7886 16890 7942 16892
rect 7966 16890 8022 16892
rect 8046 16890 8102 16892
rect 8126 16890 8182 16892
rect 7886 16838 7912 16890
rect 7912 16838 7942 16890
rect 7966 16838 7976 16890
rect 7976 16838 8022 16890
rect 8046 16838 8092 16890
rect 8092 16838 8102 16890
rect 8126 16838 8156 16890
rect 8156 16838 8182 16890
rect 7886 16836 7942 16838
rect 7966 16836 8022 16838
rect 8046 16836 8102 16838
rect 8126 16836 8182 16838
rect 7886 15802 7942 15804
rect 7966 15802 8022 15804
rect 8046 15802 8102 15804
rect 8126 15802 8182 15804
rect 7886 15750 7912 15802
rect 7912 15750 7942 15802
rect 7966 15750 7976 15802
rect 7976 15750 8022 15802
rect 8046 15750 8092 15802
rect 8092 15750 8102 15802
rect 8126 15750 8156 15802
rect 8156 15750 8182 15802
rect 7886 15748 7942 15750
rect 7966 15748 8022 15750
rect 8046 15748 8102 15750
rect 8126 15748 8182 15750
rect 7886 14714 7942 14716
rect 7966 14714 8022 14716
rect 8046 14714 8102 14716
rect 8126 14714 8182 14716
rect 7886 14662 7912 14714
rect 7912 14662 7942 14714
rect 7966 14662 7976 14714
rect 7976 14662 8022 14714
rect 8046 14662 8092 14714
rect 8092 14662 8102 14714
rect 8126 14662 8156 14714
rect 8156 14662 8182 14714
rect 7886 14660 7942 14662
rect 7966 14660 8022 14662
rect 8046 14660 8102 14662
rect 8126 14660 8182 14662
rect 7886 13626 7942 13628
rect 7966 13626 8022 13628
rect 8046 13626 8102 13628
rect 8126 13626 8182 13628
rect 7886 13574 7912 13626
rect 7912 13574 7942 13626
rect 7966 13574 7976 13626
rect 7976 13574 8022 13626
rect 8046 13574 8092 13626
rect 8092 13574 8102 13626
rect 8126 13574 8156 13626
rect 8156 13574 8182 13626
rect 7886 13572 7942 13574
rect 7966 13572 8022 13574
rect 8046 13572 8102 13574
rect 8126 13572 8182 13574
rect 8114 13132 8116 13152
rect 8116 13132 8168 13152
rect 8168 13132 8170 13152
rect 8114 13096 8170 13132
rect 7886 12538 7942 12540
rect 7966 12538 8022 12540
rect 8046 12538 8102 12540
rect 8126 12538 8182 12540
rect 7886 12486 7912 12538
rect 7912 12486 7942 12538
rect 7966 12486 7976 12538
rect 7976 12486 8022 12538
rect 8046 12486 8092 12538
rect 8092 12486 8102 12538
rect 8126 12486 8156 12538
rect 8156 12486 8182 12538
rect 7886 12484 7942 12486
rect 7966 12484 8022 12486
rect 8046 12484 8102 12486
rect 8126 12484 8182 12486
rect 7470 11756 7526 11792
rect 7470 11736 7472 11756
rect 7472 11736 7524 11756
rect 7524 11736 7526 11756
rect 8942 20032 8998 20088
rect 8850 19796 8852 19816
rect 8852 19796 8904 19816
rect 8904 19796 8906 19816
rect 8850 19760 8906 19796
rect 8850 18128 8906 18184
rect 9126 17720 9182 17776
rect 7886 11450 7942 11452
rect 7966 11450 8022 11452
rect 8046 11450 8102 11452
rect 8126 11450 8182 11452
rect 7886 11398 7912 11450
rect 7912 11398 7942 11450
rect 7966 11398 7976 11450
rect 7976 11398 8022 11450
rect 8046 11398 8092 11450
rect 8092 11398 8102 11450
rect 8126 11398 8156 11450
rect 8156 11398 8182 11450
rect 7886 11396 7942 11398
rect 7966 11396 8022 11398
rect 8046 11396 8102 11398
rect 8126 11396 8182 11398
rect 7886 10362 7942 10364
rect 7966 10362 8022 10364
rect 8046 10362 8102 10364
rect 8126 10362 8182 10364
rect 7886 10310 7912 10362
rect 7912 10310 7942 10362
rect 7966 10310 7976 10362
rect 7976 10310 8022 10362
rect 8046 10310 8092 10362
rect 8092 10310 8102 10362
rect 8126 10310 8156 10362
rect 8156 10310 8182 10362
rect 7886 10308 7942 10310
rect 7966 10308 8022 10310
rect 8046 10308 8102 10310
rect 8126 10308 8182 10310
rect 7886 9274 7942 9276
rect 7966 9274 8022 9276
rect 8046 9274 8102 9276
rect 8126 9274 8182 9276
rect 7886 9222 7912 9274
rect 7912 9222 7942 9274
rect 7966 9222 7976 9274
rect 7976 9222 8022 9274
rect 8046 9222 8092 9274
rect 8092 9222 8102 9274
rect 8126 9222 8156 9274
rect 8156 9222 8182 9274
rect 7886 9220 7942 9222
rect 7966 9220 8022 9222
rect 8046 9220 8102 9222
rect 8126 9220 8182 9222
rect 10046 20204 10048 20224
rect 10048 20204 10100 20224
rect 10100 20204 10102 20224
rect 10046 20168 10102 20204
rect 10506 20304 10562 20360
rect 10506 20052 10562 20088
rect 10506 20032 10508 20052
rect 10508 20032 10560 20052
rect 10560 20032 10562 20052
rect 9402 16632 9458 16688
rect 9494 14048 9550 14104
rect 9678 14068 9734 14104
rect 9678 14048 9680 14068
rect 9680 14048 9732 14068
rect 9732 14048 9734 14068
rect 10046 15408 10102 15464
rect 10506 17720 10562 17776
rect 9954 14900 9956 14920
rect 9956 14900 10008 14920
rect 10008 14900 10010 14920
rect 9954 14864 10010 14900
rect 9126 11600 9182 11656
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11378 20698
rect 11378 20646 11408 20698
rect 11432 20646 11442 20698
rect 11442 20646 11488 20698
rect 11512 20646 11558 20698
rect 11558 20646 11568 20698
rect 11592 20646 11622 20698
rect 11622 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 10690 17720 10746 17776
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11378 19610
rect 11378 19558 11408 19610
rect 11432 19558 11442 19610
rect 11442 19558 11488 19610
rect 11512 19558 11558 19610
rect 11558 19558 11568 19610
rect 11592 19558 11622 19610
rect 11622 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11378 18522
rect 11378 18470 11408 18522
rect 11432 18470 11442 18522
rect 11442 18470 11488 18522
rect 11512 18470 11558 18522
rect 11558 18470 11568 18522
rect 11592 18470 11622 18522
rect 11622 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 11334 17620 11336 17640
rect 11336 17620 11388 17640
rect 11388 17620 11390 17640
rect 11334 17584 11390 17620
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11378 17434
rect 11378 17382 11408 17434
rect 11432 17382 11442 17434
rect 11442 17382 11488 17434
rect 11512 17382 11558 17434
rect 11558 17382 11568 17434
rect 11592 17382 11622 17434
rect 11622 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11794 17584 11850 17640
rect 11794 16632 11850 16688
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11378 16346
rect 11378 16294 11408 16346
rect 11432 16294 11442 16346
rect 11442 16294 11488 16346
rect 11512 16294 11558 16346
rect 11558 16294 11568 16346
rect 11592 16294 11622 16346
rect 11622 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11378 15258
rect 11378 15206 11408 15258
rect 11432 15206 11442 15258
rect 11442 15206 11488 15258
rect 11512 15206 11558 15258
rect 11558 15206 11568 15258
rect 11592 15206 11622 15258
rect 11622 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11334 14900 11336 14920
rect 11336 14900 11388 14920
rect 11388 14900 11390 14920
rect 11334 14864 11390 14900
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11378 14170
rect 11378 14118 11408 14170
rect 11432 14118 11442 14170
rect 11442 14118 11488 14170
rect 11512 14118 11558 14170
rect 11558 14118 11568 14170
rect 11592 14118 11622 14170
rect 11622 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11150 14048 11206 14104
rect 12254 15428 12310 15464
rect 12254 15408 12256 15428
rect 12256 15408 12308 15428
rect 12308 15408 12310 15428
rect 12162 14492 12164 14512
rect 12164 14492 12216 14512
rect 12216 14492 12218 14512
rect 12162 14456 12218 14492
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11378 13082
rect 11378 13030 11408 13082
rect 11432 13030 11442 13082
rect 11442 13030 11488 13082
rect 11512 13030 11558 13082
rect 11558 13030 11568 13082
rect 11592 13030 11622 13082
rect 11622 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 7886 8186 7942 8188
rect 7966 8186 8022 8188
rect 8046 8186 8102 8188
rect 8126 8186 8182 8188
rect 7886 8134 7912 8186
rect 7912 8134 7942 8186
rect 7966 8134 7976 8186
rect 7976 8134 8022 8186
rect 8046 8134 8092 8186
rect 8092 8134 8102 8186
rect 8126 8134 8156 8186
rect 8156 8134 8182 8186
rect 7886 8132 7942 8134
rect 7966 8132 8022 8134
rect 8046 8132 8102 8134
rect 8126 8132 8182 8134
rect 7886 7098 7942 7100
rect 7966 7098 8022 7100
rect 8046 7098 8102 7100
rect 8126 7098 8182 7100
rect 7886 7046 7912 7098
rect 7912 7046 7942 7098
rect 7966 7046 7976 7098
rect 7976 7046 8022 7098
rect 8046 7046 8092 7098
rect 8092 7046 8102 7098
rect 8126 7046 8156 7098
rect 8156 7046 8182 7098
rect 7886 7044 7942 7046
rect 7966 7044 8022 7046
rect 8046 7044 8102 7046
rect 8126 7044 8182 7046
rect 8482 7384 8538 7440
rect 7886 6010 7942 6012
rect 7966 6010 8022 6012
rect 8046 6010 8102 6012
rect 8126 6010 8182 6012
rect 7886 5958 7912 6010
rect 7912 5958 7942 6010
rect 7966 5958 7976 6010
rect 7976 5958 8022 6010
rect 8046 5958 8092 6010
rect 8092 5958 8102 6010
rect 8126 5958 8156 6010
rect 8156 5958 8182 6010
rect 7886 5956 7942 5958
rect 7966 5956 8022 5958
rect 8046 5956 8102 5958
rect 8126 5956 8182 5958
rect 7886 4922 7942 4924
rect 7966 4922 8022 4924
rect 8046 4922 8102 4924
rect 8126 4922 8182 4924
rect 7886 4870 7912 4922
rect 7912 4870 7942 4922
rect 7966 4870 7976 4922
rect 7976 4870 8022 4922
rect 8046 4870 8092 4922
rect 8092 4870 8102 4922
rect 8126 4870 8156 4922
rect 8156 4870 8182 4922
rect 7886 4868 7942 4870
rect 7966 4868 8022 4870
rect 8046 4868 8102 4870
rect 8126 4868 8182 4870
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11378 11994
rect 11378 11942 11408 11994
rect 11432 11942 11442 11994
rect 11442 11942 11488 11994
rect 11512 11942 11558 11994
rect 11558 11942 11568 11994
rect 11592 11942 11622 11994
rect 11622 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11378 10906
rect 11378 10854 11408 10906
rect 11432 10854 11442 10906
rect 11442 10854 11488 10906
rect 11512 10854 11558 10906
rect 11558 10854 11568 10906
rect 11592 10854 11622 10906
rect 11622 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 12530 14456 12586 14512
rect 14002 20168 14058 20224
rect 13634 17584 13690 17640
rect 13358 16652 13414 16688
rect 13358 16632 13360 16652
rect 13360 16632 13412 16652
rect 13412 16632 13414 16652
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11378 9818
rect 11378 9766 11408 9818
rect 11432 9766 11442 9818
rect 11442 9766 11488 9818
rect 11512 9766 11558 9818
rect 11558 9766 11568 9818
rect 11592 9766 11622 9818
rect 11622 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11378 8730
rect 11378 8678 11408 8730
rect 11432 8678 11442 8730
rect 11442 8678 11488 8730
rect 11512 8678 11558 8730
rect 11558 8678 11568 8730
rect 11592 8678 11622 8730
rect 11622 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11378 7642
rect 11378 7590 11408 7642
rect 11432 7590 11442 7642
rect 11442 7590 11488 7642
rect 11512 7590 11558 7642
rect 11558 7590 11568 7642
rect 11592 7590 11622 7642
rect 11622 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11378 6554
rect 11378 6502 11408 6554
rect 11432 6502 11442 6554
rect 11442 6502 11488 6554
rect 11512 6502 11558 6554
rect 11558 6502 11568 6554
rect 11592 6502 11622 6554
rect 11622 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11378 5466
rect 11378 5414 11408 5466
rect 11432 5414 11442 5466
rect 11442 5414 11488 5466
rect 11512 5414 11558 5466
rect 11558 5414 11568 5466
rect 11592 5414 11622 5466
rect 11622 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11378 4378
rect 11378 4326 11408 4378
rect 11432 4326 11442 4378
rect 11442 4326 11488 4378
rect 11512 4326 11558 4378
rect 11558 4326 11568 4378
rect 11592 4326 11622 4378
rect 11622 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 7886 3834 7942 3836
rect 7966 3834 8022 3836
rect 8046 3834 8102 3836
rect 8126 3834 8182 3836
rect 7886 3782 7912 3834
rect 7912 3782 7942 3834
rect 7966 3782 7976 3834
rect 7976 3782 8022 3834
rect 8046 3782 8092 3834
rect 8092 3782 8102 3834
rect 8126 3782 8156 3834
rect 8156 3782 8182 3834
rect 7886 3780 7942 3782
rect 7966 3780 8022 3782
rect 8046 3780 8102 3782
rect 8126 3780 8182 3782
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11378 3290
rect 11378 3238 11408 3290
rect 11432 3238 11442 3290
rect 11442 3238 11488 3290
rect 11512 3238 11558 3290
rect 11558 3238 11568 3290
rect 11592 3238 11622 3290
rect 11622 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 7886 2746 7942 2748
rect 7966 2746 8022 2748
rect 8046 2746 8102 2748
rect 8126 2746 8182 2748
rect 7886 2694 7912 2746
rect 7912 2694 7942 2746
rect 7966 2694 7976 2746
rect 7976 2694 8022 2746
rect 8046 2694 8092 2746
rect 8092 2694 8102 2746
rect 8126 2694 8156 2746
rect 8156 2694 8182 2746
rect 7886 2692 7942 2694
rect 7966 2692 8022 2694
rect 8046 2692 8102 2694
rect 8126 2692 8182 2694
rect 14817 20154 14873 20156
rect 14897 20154 14953 20156
rect 14977 20154 15033 20156
rect 15057 20154 15113 20156
rect 14817 20102 14843 20154
rect 14843 20102 14873 20154
rect 14897 20102 14907 20154
rect 14907 20102 14953 20154
rect 14977 20102 15023 20154
rect 15023 20102 15033 20154
rect 15057 20102 15087 20154
rect 15087 20102 15113 20154
rect 14817 20100 14873 20102
rect 14897 20100 14953 20102
rect 14977 20100 15033 20102
rect 15057 20100 15113 20102
rect 16578 20460 16634 20496
rect 16578 20440 16580 20460
rect 16580 20440 16632 20460
rect 16632 20440 16634 20460
rect 18282 20698 18338 20700
rect 18362 20698 18418 20700
rect 18442 20698 18498 20700
rect 18522 20698 18578 20700
rect 18282 20646 18308 20698
rect 18308 20646 18338 20698
rect 18362 20646 18372 20698
rect 18372 20646 18418 20698
rect 18442 20646 18488 20698
rect 18488 20646 18498 20698
rect 18522 20646 18552 20698
rect 18552 20646 18578 20698
rect 18282 20644 18338 20646
rect 18362 20644 18418 20646
rect 18442 20644 18498 20646
rect 18522 20644 18578 20646
rect 14817 19066 14873 19068
rect 14897 19066 14953 19068
rect 14977 19066 15033 19068
rect 15057 19066 15113 19068
rect 14817 19014 14843 19066
rect 14843 19014 14873 19066
rect 14897 19014 14907 19066
rect 14907 19014 14953 19066
rect 14977 19014 15023 19066
rect 15023 19014 15033 19066
rect 15057 19014 15087 19066
rect 15087 19014 15113 19066
rect 14817 19012 14873 19014
rect 14897 19012 14953 19014
rect 14977 19012 15033 19014
rect 15057 19012 15113 19014
rect 14370 18708 14372 18728
rect 14372 18708 14424 18728
rect 14424 18708 14426 18728
rect 14370 18672 14426 18708
rect 14817 17978 14873 17980
rect 14897 17978 14953 17980
rect 14977 17978 15033 17980
rect 15057 17978 15113 17980
rect 14817 17926 14843 17978
rect 14843 17926 14873 17978
rect 14897 17926 14907 17978
rect 14907 17926 14953 17978
rect 14977 17926 15023 17978
rect 15023 17926 15033 17978
rect 15057 17926 15087 17978
rect 15087 17926 15113 17978
rect 14817 17924 14873 17926
rect 14897 17924 14953 17926
rect 14977 17924 15033 17926
rect 15057 17924 15113 17926
rect 15290 17740 15346 17776
rect 15290 17720 15292 17740
rect 15292 17720 15344 17740
rect 15344 17720 15346 17740
rect 14817 16890 14873 16892
rect 14897 16890 14953 16892
rect 14977 16890 15033 16892
rect 15057 16890 15113 16892
rect 14817 16838 14843 16890
rect 14843 16838 14873 16890
rect 14897 16838 14907 16890
rect 14907 16838 14953 16890
rect 14977 16838 15023 16890
rect 15023 16838 15033 16890
rect 15057 16838 15087 16890
rect 15087 16838 15113 16890
rect 14817 16836 14873 16838
rect 14897 16836 14953 16838
rect 14977 16836 15033 16838
rect 15057 16836 15113 16838
rect 14817 15802 14873 15804
rect 14897 15802 14953 15804
rect 14977 15802 15033 15804
rect 15057 15802 15113 15804
rect 14817 15750 14843 15802
rect 14843 15750 14873 15802
rect 14897 15750 14907 15802
rect 14907 15750 14953 15802
rect 14977 15750 15023 15802
rect 15023 15750 15033 15802
rect 15057 15750 15087 15802
rect 15087 15750 15113 15802
rect 14817 15748 14873 15750
rect 14897 15748 14953 15750
rect 14977 15748 15033 15750
rect 15057 15748 15113 15750
rect 14817 14714 14873 14716
rect 14897 14714 14953 14716
rect 14977 14714 15033 14716
rect 15057 14714 15113 14716
rect 14817 14662 14843 14714
rect 14843 14662 14873 14714
rect 14897 14662 14907 14714
rect 14907 14662 14953 14714
rect 14977 14662 15023 14714
rect 15023 14662 15033 14714
rect 15057 14662 15087 14714
rect 15087 14662 15113 14714
rect 14817 14660 14873 14662
rect 14897 14660 14953 14662
rect 14977 14660 15033 14662
rect 15057 14660 15113 14662
rect 14817 13626 14873 13628
rect 14897 13626 14953 13628
rect 14977 13626 15033 13628
rect 15057 13626 15113 13628
rect 14817 13574 14843 13626
rect 14843 13574 14873 13626
rect 14897 13574 14907 13626
rect 14907 13574 14953 13626
rect 14977 13574 15023 13626
rect 15023 13574 15033 13626
rect 15057 13574 15087 13626
rect 15087 13574 15113 13626
rect 14817 13572 14873 13574
rect 14897 13572 14953 13574
rect 14977 13572 15033 13574
rect 15057 13572 15113 13574
rect 14817 12538 14873 12540
rect 14897 12538 14953 12540
rect 14977 12538 15033 12540
rect 15057 12538 15113 12540
rect 14817 12486 14843 12538
rect 14843 12486 14873 12538
rect 14897 12486 14907 12538
rect 14907 12486 14953 12538
rect 14977 12486 15023 12538
rect 15023 12486 15033 12538
rect 15057 12486 15087 12538
rect 15087 12486 15113 12538
rect 14817 12484 14873 12486
rect 14897 12484 14953 12486
rect 14977 12484 15033 12486
rect 15057 12484 15113 12486
rect 18282 19610 18338 19612
rect 18362 19610 18418 19612
rect 18442 19610 18498 19612
rect 18522 19610 18578 19612
rect 18282 19558 18308 19610
rect 18308 19558 18338 19610
rect 18362 19558 18372 19610
rect 18372 19558 18418 19610
rect 18442 19558 18488 19610
rect 18488 19558 18498 19610
rect 18522 19558 18552 19610
rect 18552 19558 18578 19610
rect 18282 19556 18338 19558
rect 18362 19556 18418 19558
rect 18442 19556 18498 19558
rect 18522 19556 18578 19558
rect 18282 18522 18338 18524
rect 18362 18522 18418 18524
rect 18442 18522 18498 18524
rect 18522 18522 18578 18524
rect 18282 18470 18308 18522
rect 18308 18470 18338 18522
rect 18362 18470 18372 18522
rect 18372 18470 18418 18522
rect 18442 18470 18488 18522
rect 18488 18470 18498 18522
rect 18522 18470 18552 18522
rect 18552 18470 18578 18522
rect 18282 18468 18338 18470
rect 18362 18468 18418 18470
rect 18442 18468 18498 18470
rect 18522 18468 18578 18470
rect 18282 17434 18338 17436
rect 18362 17434 18418 17436
rect 18442 17434 18498 17436
rect 18522 17434 18578 17436
rect 18282 17382 18308 17434
rect 18308 17382 18338 17434
rect 18362 17382 18372 17434
rect 18372 17382 18418 17434
rect 18442 17382 18488 17434
rect 18488 17382 18498 17434
rect 18522 17382 18552 17434
rect 18552 17382 18578 17434
rect 18282 17380 18338 17382
rect 18362 17380 18418 17382
rect 18442 17380 18498 17382
rect 18522 17380 18578 17382
rect 18282 16346 18338 16348
rect 18362 16346 18418 16348
rect 18442 16346 18498 16348
rect 18522 16346 18578 16348
rect 18282 16294 18308 16346
rect 18308 16294 18338 16346
rect 18362 16294 18372 16346
rect 18372 16294 18418 16346
rect 18442 16294 18488 16346
rect 18488 16294 18498 16346
rect 18522 16294 18552 16346
rect 18552 16294 18578 16346
rect 18282 16292 18338 16294
rect 18362 16292 18418 16294
rect 18442 16292 18498 16294
rect 18522 16292 18578 16294
rect 14817 11450 14873 11452
rect 14897 11450 14953 11452
rect 14977 11450 15033 11452
rect 15057 11450 15113 11452
rect 14817 11398 14843 11450
rect 14843 11398 14873 11450
rect 14897 11398 14907 11450
rect 14907 11398 14953 11450
rect 14977 11398 15023 11450
rect 15023 11398 15033 11450
rect 15057 11398 15087 11450
rect 15087 11398 15113 11450
rect 14817 11396 14873 11398
rect 14897 11396 14953 11398
rect 14977 11396 15033 11398
rect 15057 11396 15113 11398
rect 14817 10362 14873 10364
rect 14897 10362 14953 10364
rect 14977 10362 15033 10364
rect 15057 10362 15113 10364
rect 14817 10310 14843 10362
rect 14843 10310 14873 10362
rect 14897 10310 14907 10362
rect 14907 10310 14953 10362
rect 14977 10310 15023 10362
rect 15023 10310 15033 10362
rect 15057 10310 15087 10362
rect 15087 10310 15113 10362
rect 14817 10308 14873 10310
rect 14897 10308 14953 10310
rect 14977 10308 15033 10310
rect 15057 10308 15113 10310
rect 14817 9274 14873 9276
rect 14897 9274 14953 9276
rect 14977 9274 15033 9276
rect 15057 9274 15113 9276
rect 14817 9222 14843 9274
rect 14843 9222 14873 9274
rect 14897 9222 14907 9274
rect 14907 9222 14953 9274
rect 14977 9222 15023 9274
rect 15023 9222 15033 9274
rect 15057 9222 15087 9274
rect 15087 9222 15113 9274
rect 14817 9220 14873 9222
rect 14897 9220 14953 9222
rect 14977 9220 15033 9222
rect 15057 9220 15113 9222
rect 14817 8186 14873 8188
rect 14897 8186 14953 8188
rect 14977 8186 15033 8188
rect 15057 8186 15113 8188
rect 14817 8134 14843 8186
rect 14843 8134 14873 8186
rect 14897 8134 14907 8186
rect 14907 8134 14953 8186
rect 14977 8134 15023 8186
rect 15023 8134 15033 8186
rect 15057 8134 15087 8186
rect 15087 8134 15113 8186
rect 14817 8132 14873 8134
rect 14897 8132 14953 8134
rect 14977 8132 15033 8134
rect 15057 8132 15113 8134
rect 18282 15258 18338 15260
rect 18362 15258 18418 15260
rect 18442 15258 18498 15260
rect 18522 15258 18578 15260
rect 18282 15206 18308 15258
rect 18308 15206 18338 15258
rect 18362 15206 18372 15258
rect 18372 15206 18418 15258
rect 18442 15206 18488 15258
rect 18488 15206 18498 15258
rect 18522 15206 18552 15258
rect 18552 15206 18578 15258
rect 18282 15204 18338 15206
rect 18362 15204 18418 15206
rect 18442 15204 18498 15206
rect 18522 15204 18578 15206
rect 18282 14170 18338 14172
rect 18362 14170 18418 14172
rect 18442 14170 18498 14172
rect 18522 14170 18578 14172
rect 18282 14118 18308 14170
rect 18308 14118 18338 14170
rect 18362 14118 18372 14170
rect 18372 14118 18418 14170
rect 18442 14118 18488 14170
rect 18488 14118 18498 14170
rect 18522 14118 18552 14170
rect 18552 14118 18578 14170
rect 18282 14116 18338 14118
rect 18362 14116 18418 14118
rect 18442 14116 18498 14118
rect 18522 14116 18578 14118
rect 18282 13082 18338 13084
rect 18362 13082 18418 13084
rect 18442 13082 18498 13084
rect 18522 13082 18578 13084
rect 18282 13030 18308 13082
rect 18308 13030 18338 13082
rect 18362 13030 18372 13082
rect 18372 13030 18418 13082
rect 18442 13030 18488 13082
rect 18488 13030 18498 13082
rect 18522 13030 18552 13082
rect 18552 13030 18578 13082
rect 18282 13028 18338 13030
rect 18362 13028 18418 13030
rect 18442 13028 18498 13030
rect 18522 13028 18578 13030
rect 18282 11994 18338 11996
rect 18362 11994 18418 11996
rect 18442 11994 18498 11996
rect 18522 11994 18578 11996
rect 18282 11942 18308 11994
rect 18308 11942 18338 11994
rect 18362 11942 18372 11994
rect 18372 11942 18418 11994
rect 18442 11942 18488 11994
rect 18488 11942 18498 11994
rect 18522 11942 18552 11994
rect 18552 11942 18578 11994
rect 18282 11940 18338 11942
rect 18362 11940 18418 11942
rect 18442 11940 18498 11942
rect 18522 11940 18578 11942
rect 18282 10906 18338 10908
rect 18362 10906 18418 10908
rect 18442 10906 18498 10908
rect 18522 10906 18578 10908
rect 18282 10854 18308 10906
rect 18308 10854 18338 10906
rect 18362 10854 18372 10906
rect 18372 10854 18418 10906
rect 18442 10854 18488 10906
rect 18488 10854 18498 10906
rect 18522 10854 18552 10906
rect 18552 10854 18578 10906
rect 18282 10852 18338 10854
rect 18362 10852 18418 10854
rect 18442 10852 18498 10854
rect 18522 10852 18578 10854
rect 18282 9818 18338 9820
rect 18362 9818 18418 9820
rect 18442 9818 18498 9820
rect 18522 9818 18578 9820
rect 18282 9766 18308 9818
rect 18308 9766 18338 9818
rect 18362 9766 18372 9818
rect 18372 9766 18418 9818
rect 18442 9766 18488 9818
rect 18488 9766 18498 9818
rect 18522 9766 18552 9818
rect 18552 9766 18578 9818
rect 18282 9764 18338 9766
rect 18362 9764 18418 9766
rect 18442 9764 18498 9766
rect 18522 9764 18578 9766
rect 18282 8730 18338 8732
rect 18362 8730 18418 8732
rect 18442 8730 18498 8732
rect 18522 8730 18578 8732
rect 18282 8678 18308 8730
rect 18308 8678 18338 8730
rect 18362 8678 18372 8730
rect 18372 8678 18418 8730
rect 18442 8678 18488 8730
rect 18488 8678 18498 8730
rect 18522 8678 18552 8730
rect 18552 8678 18578 8730
rect 18282 8676 18338 8678
rect 18362 8676 18418 8678
rect 18442 8676 18498 8678
rect 18522 8676 18578 8678
rect 18282 7642 18338 7644
rect 18362 7642 18418 7644
rect 18442 7642 18498 7644
rect 18522 7642 18578 7644
rect 18282 7590 18308 7642
rect 18308 7590 18338 7642
rect 18362 7590 18372 7642
rect 18372 7590 18418 7642
rect 18442 7590 18488 7642
rect 18488 7590 18498 7642
rect 18522 7590 18552 7642
rect 18552 7590 18578 7642
rect 18282 7588 18338 7590
rect 18362 7588 18418 7590
rect 18442 7588 18498 7590
rect 18522 7588 18578 7590
rect 18786 7284 18788 7304
rect 18788 7284 18840 7304
rect 18840 7284 18842 7304
rect 18786 7248 18842 7284
rect 14817 7098 14873 7100
rect 14897 7098 14953 7100
rect 14977 7098 15033 7100
rect 15057 7098 15113 7100
rect 14817 7046 14843 7098
rect 14843 7046 14873 7098
rect 14897 7046 14907 7098
rect 14907 7046 14953 7098
rect 14977 7046 15023 7098
rect 15023 7046 15033 7098
rect 15057 7046 15087 7098
rect 15087 7046 15113 7098
rect 14817 7044 14873 7046
rect 14897 7044 14953 7046
rect 14977 7044 15033 7046
rect 15057 7044 15113 7046
rect 18282 6554 18338 6556
rect 18362 6554 18418 6556
rect 18442 6554 18498 6556
rect 18522 6554 18578 6556
rect 18282 6502 18308 6554
rect 18308 6502 18338 6554
rect 18362 6502 18372 6554
rect 18372 6502 18418 6554
rect 18442 6502 18488 6554
rect 18488 6502 18498 6554
rect 18522 6502 18552 6554
rect 18552 6502 18578 6554
rect 18282 6500 18338 6502
rect 18362 6500 18418 6502
rect 18442 6500 18498 6502
rect 18522 6500 18578 6502
rect 14817 6010 14873 6012
rect 14897 6010 14953 6012
rect 14977 6010 15033 6012
rect 15057 6010 15113 6012
rect 14817 5958 14843 6010
rect 14843 5958 14873 6010
rect 14897 5958 14907 6010
rect 14907 5958 14953 6010
rect 14977 5958 15023 6010
rect 15023 5958 15033 6010
rect 15057 5958 15087 6010
rect 15087 5958 15113 6010
rect 14817 5956 14873 5958
rect 14897 5956 14953 5958
rect 14977 5956 15033 5958
rect 15057 5956 15113 5958
rect 18282 5466 18338 5468
rect 18362 5466 18418 5468
rect 18442 5466 18498 5468
rect 18522 5466 18578 5468
rect 18282 5414 18308 5466
rect 18308 5414 18338 5466
rect 18362 5414 18372 5466
rect 18372 5414 18418 5466
rect 18442 5414 18488 5466
rect 18488 5414 18498 5466
rect 18522 5414 18552 5466
rect 18552 5414 18578 5466
rect 18282 5412 18338 5414
rect 18362 5412 18418 5414
rect 18442 5412 18498 5414
rect 18522 5412 18578 5414
rect 21362 11464 21418 11520
rect 14817 4922 14873 4924
rect 14897 4922 14953 4924
rect 14977 4922 15033 4924
rect 15057 4922 15113 4924
rect 14817 4870 14843 4922
rect 14843 4870 14873 4922
rect 14897 4870 14907 4922
rect 14907 4870 14953 4922
rect 14977 4870 15023 4922
rect 15023 4870 15033 4922
rect 15057 4870 15087 4922
rect 15087 4870 15113 4922
rect 14817 4868 14873 4870
rect 14897 4868 14953 4870
rect 14977 4868 15033 4870
rect 15057 4868 15113 4870
rect 18282 4378 18338 4380
rect 18362 4378 18418 4380
rect 18442 4378 18498 4380
rect 18522 4378 18578 4380
rect 18282 4326 18308 4378
rect 18308 4326 18338 4378
rect 18362 4326 18372 4378
rect 18372 4326 18418 4378
rect 18442 4326 18488 4378
rect 18488 4326 18498 4378
rect 18522 4326 18552 4378
rect 18552 4326 18578 4378
rect 18282 4324 18338 4326
rect 18362 4324 18418 4326
rect 18442 4324 18498 4326
rect 18522 4324 18578 4326
rect 14817 3834 14873 3836
rect 14897 3834 14953 3836
rect 14977 3834 15033 3836
rect 15057 3834 15113 3836
rect 14817 3782 14843 3834
rect 14843 3782 14873 3834
rect 14897 3782 14907 3834
rect 14907 3782 14953 3834
rect 14977 3782 15023 3834
rect 15023 3782 15033 3834
rect 15057 3782 15087 3834
rect 15087 3782 15113 3834
rect 14817 3780 14873 3782
rect 14897 3780 14953 3782
rect 14977 3780 15033 3782
rect 15057 3780 15113 3782
rect 18282 3290 18338 3292
rect 18362 3290 18418 3292
rect 18442 3290 18498 3292
rect 18522 3290 18578 3292
rect 18282 3238 18308 3290
rect 18308 3238 18338 3290
rect 18362 3238 18372 3290
rect 18372 3238 18418 3290
rect 18442 3238 18488 3290
rect 18488 3238 18498 3290
rect 18522 3238 18552 3290
rect 18552 3238 18578 3290
rect 18282 3236 18338 3238
rect 18362 3236 18418 3238
rect 18442 3236 18498 3238
rect 18522 3236 18578 3238
rect 14817 2746 14873 2748
rect 14897 2746 14953 2748
rect 14977 2746 15033 2748
rect 15057 2746 15113 2748
rect 14817 2694 14843 2746
rect 14843 2694 14873 2746
rect 14897 2694 14907 2746
rect 14907 2694 14953 2746
rect 14977 2694 15023 2746
rect 15023 2694 15033 2746
rect 15057 2694 15087 2746
rect 15087 2694 15113 2746
rect 14817 2692 14873 2694
rect 14897 2692 14953 2694
rect 14977 2692 15033 2694
rect 15057 2692 15113 2694
rect 4421 2202 4477 2204
rect 4501 2202 4557 2204
rect 4581 2202 4637 2204
rect 4661 2202 4717 2204
rect 4421 2150 4447 2202
rect 4447 2150 4477 2202
rect 4501 2150 4511 2202
rect 4511 2150 4557 2202
rect 4581 2150 4627 2202
rect 4627 2150 4637 2202
rect 4661 2150 4691 2202
rect 4691 2150 4717 2202
rect 4421 2148 4477 2150
rect 4501 2148 4557 2150
rect 4581 2148 4637 2150
rect 4661 2148 4717 2150
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11378 2202
rect 11378 2150 11408 2202
rect 11432 2150 11442 2202
rect 11442 2150 11488 2202
rect 11512 2150 11558 2202
rect 11558 2150 11568 2202
rect 11592 2150 11622 2202
rect 11622 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 3882 1944 3938 2000
rect 3146 1536 3202 1592
rect 18282 2202 18338 2204
rect 18362 2202 18418 2204
rect 18442 2202 18498 2204
rect 18522 2202 18578 2204
rect 18282 2150 18308 2202
rect 18308 2150 18338 2202
rect 18362 2150 18372 2202
rect 18372 2150 18418 2202
rect 18442 2150 18488 2202
rect 18488 2150 18498 2202
rect 18522 2150 18552 2202
rect 18552 2150 18578 2202
rect 18282 2148 18338 2150
rect 18362 2148 18418 2150
rect 18442 2148 18498 2150
rect 18522 2148 18578 2150
rect 2778 992 2834 1048
rect 2226 584 2282 640
rect 2134 176 2190 232
<< metal3 >>
rect 0 22674 800 22704
rect 3969 22674 4035 22677
rect 0 22672 4035 22674
rect 0 22616 3974 22672
rect 4030 22616 4035 22672
rect 0 22614 4035 22616
rect 0 22584 800 22614
rect 3969 22611 4035 22614
rect 0 22266 800 22296
rect 4061 22266 4127 22269
rect 0 22264 4127 22266
rect 0 22208 4066 22264
rect 4122 22208 4127 22264
rect 0 22206 4127 22208
rect 0 22176 800 22206
rect 4061 22203 4127 22206
rect 0 21722 800 21752
rect 2957 21722 3023 21725
rect 0 21720 3023 21722
rect 0 21664 2962 21720
rect 3018 21664 3023 21720
rect 0 21662 3023 21664
rect 0 21632 800 21662
rect 2957 21659 3023 21662
rect 0 21314 800 21344
rect 3049 21314 3115 21317
rect 0 21312 3115 21314
rect 0 21256 3054 21312
rect 3110 21256 3115 21312
rect 0 21254 3115 21256
rect 0 21224 800 21254
rect 3049 21251 3115 21254
rect 0 20770 800 20800
rect 2865 20770 2931 20773
rect 0 20768 2931 20770
rect 0 20712 2870 20768
rect 2926 20712 2931 20768
rect 0 20710 2931 20712
rect 0 20680 800 20710
rect 2865 20707 2931 20710
rect 4409 20704 4729 20705
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 20639 4729 20640
rect 11340 20704 11660 20705
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 20639 11660 20640
rect 18270 20704 18590 20705
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18590 20704
rect 18270 20639 18590 20640
rect 5809 20634 5875 20637
rect 7649 20634 7715 20637
rect 5809 20632 7715 20634
rect 5809 20576 5814 20632
rect 5870 20576 7654 20632
rect 7710 20576 7715 20632
rect 5809 20574 7715 20576
rect 5809 20571 5875 20574
rect 7649 20571 7715 20574
rect 2773 20498 2839 20501
rect 4153 20498 4219 20501
rect 6545 20498 6611 20501
rect 2773 20496 3618 20498
rect 2773 20440 2778 20496
rect 2834 20440 3618 20496
rect 2773 20438 3618 20440
rect 2773 20435 2839 20438
rect 0 20362 800 20392
rect 2773 20362 2839 20365
rect 0 20360 2839 20362
rect 0 20304 2778 20360
rect 2834 20304 2839 20360
rect 0 20302 2839 20304
rect 3558 20362 3618 20438
rect 4153 20496 6611 20498
rect 4153 20440 4158 20496
rect 4214 20440 6550 20496
rect 6606 20440 6611 20496
rect 4153 20438 6611 20440
rect 4153 20435 4219 20438
rect 6545 20435 6611 20438
rect 6821 20498 6887 20501
rect 16573 20498 16639 20501
rect 6821 20496 16639 20498
rect 6821 20440 6826 20496
rect 6882 20440 16578 20496
rect 16634 20440 16639 20496
rect 6821 20438 16639 20440
rect 6821 20435 6887 20438
rect 16573 20435 16639 20438
rect 10501 20362 10567 20365
rect 3558 20360 10567 20362
rect 3558 20304 10506 20360
rect 10562 20304 10567 20360
rect 3558 20302 10567 20304
rect 0 20272 800 20302
rect 2773 20299 2839 20302
rect 10501 20299 10567 20302
rect 10041 20226 10107 20229
rect 13997 20226 14063 20229
rect 10041 20224 14063 20226
rect 10041 20168 10046 20224
rect 10102 20168 14002 20224
rect 14058 20168 14063 20224
rect 10041 20166 14063 20168
rect 10041 20163 10107 20166
rect 13997 20163 14063 20166
rect 7874 20160 8194 20161
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8194 20160
rect 7874 20095 8194 20096
rect 14805 20160 15125 20161
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 20095 15125 20096
rect 4613 20090 4679 20093
rect 7281 20090 7347 20093
rect 4613 20088 7347 20090
rect 4613 20032 4618 20088
rect 4674 20032 7286 20088
rect 7342 20032 7347 20088
rect 4613 20030 7347 20032
rect 4613 20027 4679 20030
rect 7281 20027 7347 20030
rect 8385 20090 8451 20093
rect 8937 20090 9003 20093
rect 10501 20090 10567 20093
rect 8385 20088 10567 20090
rect 8385 20032 8390 20088
rect 8446 20032 8942 20088
rect 8998 20032 10506 20088
rect 10562 20032 10567 20088
rect 8385 20030 10567 20032
rect 8385 20027 8451 20030
rect 8937 20027 9003 20030
rect 10501 20027 10567 20030
rect 0 19818 800 19848
rect 1577 19818 1643 19821
rect 0 19816 1643 19818
rect 0 19760 1582 19816
rect 1638 19760 1643 19816
rect 0 19758 1643 19760
rect 0 19728 800 19758
rect 1577 19755 1643 19758
rect 5349 19818 5415 19821
rect 8845 19818 8911 19821
rect 5349 19816 8911 19818
rect 5349 19760 5354 19816
rect 5410 19760 8850 19816
rect 8906 19760 8911 19816
rect 5349 19758 8911 19760
rect 5349 19755 5415 19758
rect 8845 19755 8911 19758
rect 4409 19616 4729 19617
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 19551 4729 19552
rect 11340 19616 11660 19617
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 19551 11660 19552
rect 18270 19616 18590 19617
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18590 19616
rect 18270 19551 18590 19552
rect 0 19410 800 19440
rect 1577 19410 1643 19413
rect 0 19408 1643 19410
rect 0 19352 1582 19408
rect 1638 19352 1643 19408
rect 0 19350 1643 19352
rect 0 19320 800 19350
rect 1577 19347 1643 19350
rect 4061 19274 4127 19277
rect 5073 19274 5139 19277
rect 4061 19272 5139 19274
rect 4061 19216 4066 19272
rect 4122 19216 5078 19272
rect 5134 19216 5139 19272
rect 4061 19214 5139 19216
rect 4061 19211 4127 19214
rect 5073 19211 5139 19214
rect 7874 19072 8194 19073
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8194 19072
rect 7874 19007 8194 19008
rect 14805 19072 15125 19073
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 19007 15125 19008
rect 0 18866 800 18896
rect 1577 18866 1643 18869
rect 0 18864 1643 18866
rect 0 18808 1582 18864
rect 1638 18808 1643 18864
rect 0 18806 1643 18808
rect 0 18776 800 18806
rect 1577 18803 1643 18806
rect 2497 18730 2563 18733
rect 14365 18730 14431 18733
rect 2497 18728 14431 18730
rect 2497 18672 2502 18728
rect 2558 18672 14370 18728
rect 14426 18672 14431 18728
rect 2497 18670 14431 18672
rect 2497 18667 2563 18670
rect 14365 18667 14431 18670
rect 5073 18594 5139 18597
rect 6085 18594 6151 18597
rect 5073 18592 6151 18594
rect 5073 18536 5078 18592
rect 5134 18536 6090 18592
rect 6146 18536 6151 18592
rect 5073 18534 6151 18536
rect 5073 18531 5139 18534
rect 6085 18531 6151 18534
rect 4409 18528 4729 18529
rect 0 18458 800 18488
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 18463 4729 18464
rect 11340 18528 11660 18529
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 18463 11660 18464
rect 18270 18528 18590 18529
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18590 18528
rect 18270 18463 18590 18464
rect 1669 18458 1735 18461
rect 0 18456 1735 18458
rect 0 18400 1674 18456
rect 1730 18400 1735 18456
rect 0 18398 1735 18400
rect 0 18368 800 18398
rect 1669 18395 1735 18398
rect 3325 18186 3391 18189
rect 8845 18186 8911 18189
rect 3325 18184 8911 18186
rect 3325 18128 3330 18184
rect 3386 18128 8850 18184
rect 8906 18128 8911 18184
rect 3325 18126 8911 18128
rect 3325 18123 3391 18126
rect 8845 18123 8911 18126
rect 0 18050 800 18080
rect 2773 18050 2839 18053
rect 0 18048 2839 18050
rect 0 17992 2778 18048
rect 2834 17992 2839 18048
rect 0 17990 2839 17992
rect 0 17960 800 17990
rect 2773 17987 2839 17990
rect 7874 17984 8194 17985
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8194 17984
rect 7874 17919 8194 17920
rect 14805 17984 15125 17985
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 14805 17919 15125 17920
rect 9121 17778 9187 17781
rect 10501 17778 10567 17781
rect 9121 17776 10567 17778
rect 9121 17720 9126 17776
rect 9182 17720 10506 17776
rect 10562 17720 10567 17776
rect 9121 17718 10567 17720
rect 9121 17715 9187 17718
rect 10501 17715 10567 17718
rect 10685 17778 10751 17781
rect 15285 17778 15351 17781
rect 10685 17776 15351 17778
rect 10685 17720 10690 17776
rect 10746 17720 15290 17776
rect 15346 17720 15351 17776
rect 10685 17718 15351 17720
rect 10685 17715 10751 17718
rect 15285 17715 15351 17718
rect 11329 17642 11395 17645
rect 11789 17642 11855 17645
rect 13629 17642 13695 17645
rect 11329 17640 13695 17642
rect 11329 17584 11334 17640
rect 11390 17584 11794 17640
rect 11850 17584 13634 17640
rect 13690 17584 13695 17640
rect 11329 17582 13695 17584
rect 11329 17579 11395 17582
rect 11789 17579 11855 17582
rect 13629 17579 13695 17582
rect 0 17506 800 17536
rect 2221 17506 2287 17509
rect 0 17504 2287 17506
rect 0 17448 2226 17504
rect 2282 17448 2287 17504
rect 0 17446 2287 17448
rect 0 17416 800 17446
rect 2221 17443 2287 17446
rect 4409 17440 4729 17441
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 17375 4729 17376
rect 11340 17440 11660 17441
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 17375 11660 17376
rect 18270 17440 18590 17441
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18590 17440
rect 18270 17375 18590 17376
rect 0 17098 800 17128
rect 1577 17098 1643 17101
rect 0 17096 1643 17098
rect 0 17040 1582 17096
rect 1638 17040 1643 17096
rect 0 17038 1643 17040
rect 0 17008 800 17038
rect 1577 17035 1643 17038
rect 7874 16896 8194 16897
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8194 16896
rect 7874 16831 8194 16832
rect 14805 16896 15125 16897
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 16831 15125 16832
rect 5625 16690 5691 16693
rect 6637 16690 6703 16693
rect 5625 16688 6703 16690
rect 5625 16632 5630 16688
rect 5686 16632 6642 16688
rect 6698 16632 6703 16688
rect 5625 16630 6703 16632
rect 5625 16627 5691 16630
rect 6637 16627 6703 16630
rect 9397 16690 9463 16693
rect 11789 16690 11855 16693
rect 13353 16690 13419 16693
rect 9397 16688 13419 16690
rect 9397 16632 9402 16688
rect 9458 16632 11794 16688
rect 11850 16632 13358 16688
rect 13414 16632 13419 16688
rect 9397 16630 13419 16632
rect 9397 16627 9463 16630
rect 11789 16627 11855 16630
rect 13353 16627 13419 16630
rect 0 16554 800 16584
rect 1577 16554 1643 16557
rect 0 16552 1643 16554
rect 0 16496 1582 16552
rect 1638 16496 1643 16552
rect 0 16494 1643 16496
rect 0 16464 800 16494
rect 1577 16491 1643 16494
rect 4409 16352 4729 16353
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 16287 4729 16288
rect 11340 16352 11660 16353
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 16287 11660 16288
rect 18270 16352 18590 16353
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18590 16352
rect 18270 16287 18590 16288
rect 0 16146 800 16176
rect 1577 16146 1643 16149
rect 0 16144 1643 16146
rect 0 16088 1582 16144
rect 1638 16088 1643 16144
rect 0 16086 1643 16088
rect 0 16056 800 16086
rect 1577 16083 1643 16086
rect 4061 16010 4127 16013
rect 4613 16010 4679 16013
rect 5993 16010 6059 16013
rect 4061 16008 6059 16010
rect 4061 15952 4066 16008
rect 4122 15952 4618 16008
rect 4674 15952 5998 16008
rect 6054 15952 6059 16008
rect 4061 15950 6059 15952
rect 4061 15947 4127 15950
rect 4613 15947 4679 15950
rect 5993 15947 6059 15950
rect 7874 15808 8194 15809
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8194 15808
rect 7874 15743 8194 15744
rect 14805 15808 15125 15809
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 15743 15125 15744
rect 0 15602 800 15632
rect 1577 15602 1643 15605
rect 0 15600 1643 15602
rect 0 15544 1582 15600
rect 1638 15544 1643 15600
rect 0 15542 1643 15544
rect 0 15512 800 15542
rect 1577 15539 1643 15542
rect 10041 15466 10107 15469
rect 12249 15466 12315 15469
rect 10041 15464 12315 15466
rect 10041 15408 10046 15464
rect 10102 15408 12254 15464
rect 12310 15408 12315 15464
rect 10041 15406 12315 15408
rect 10041 15403 10107 15406
rect 12249 15403 12315 15406
rect 4409 15264 4729 15265
rect 0 15194 800 15224
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 15199 4729 15200
rect 11340 15264 11660 15265
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 15199 11660 15200
rect 18270 15264 18590 15265
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18590 15264
rect 18270 15199 18590 15200
rect 1669 15194 1735 15197
rect 0 15192 1735 15194
rect 0 15136 1674 15192
rect 1730 15136 1735 15192
rect 0 15134 1735 15136
rect 0 15104 800 15134
rect 1669 15131 1735 15134
rect 9949 14922 10015 14925
rect 11329 14922 11395 14925
rect 9949 14920 11395 14922
rect 9949 14864 9954 14920
rect 10010 14864 11334 14920
rect 11390 14864 11395 14920
rect 9949 14862 11395 14864
rect 9949 14859 10015 14862
rect 11329 14859 11395 14862
rect 7874 14720 8194 14721
rect 0 14650 800 14680
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8194 14720
rect 7874 14655 8194 14656
rect 14805 14720 15125 14721
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 14655 15125 14656
rect 2221 14650 2287 14653
rect 0 14648 2287 14650
rect 0 14592 2226 14648
rect 2282 14592 2287 14648
rect 0 14590 2287 14592
rect 0 14560 800 14590
rect 2221 14587 2287 14590
rect 12157 14514 12223 14517
rect 12525 14514 12591 14517
rect 12157 14512 12591 14514
rect 12157 14456 12162 14512
rect 12218 14456 12530 14512
rect 12586 14456 12591 14512
rect 12157 14454 12591 14456
rect 12157 14451 12223 14454
rect 12525 14451 12591 14454
rect 0 14242 800 14272
rect 1669 14242 1735 14245
rect 0 14240 1735 14242
rect 0 14184 1674 14240
rect 1730 14184 1735 14240
rect 0 14182 1735 14184
rect 0 14152 800 14182
rect 1669 14179 1735 14182
rect 4409 14176 4729 14177
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 14111 4729 14112
rect 11340 14176 11660 14177
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 14111 11660 14112
rect 18270 14176 18590 14177
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18590 14176
rect 18270 14111 18590 14112
rect 5073 14106 5139 14109
rect 9489 14106 9555 14109
rect 5073 14104 9555 14106
rect 5073 14048 5078 14104
rect 5134 14048 9494 14104
rect 9550 14048 9555 14104
rect 5073 14046 9555 14048
rect 5073 14043 5139 14046
rect 9489 14043 9555 14046
rect 9673 14106 9739 14109
rect 11145 14106 11211 14109
rect 9673 14104 11211 14106
rect 9673 14048 9678 14104
rect 9734 14048 11150 14104
rect 11206 14048 11211 14104
rect 9673 14046 11211 14048
rect 9673 14043 9739 14046
rect 11145 14043 11211 14046
rect 4337 13970 4403 13973
rect 6085 13970 6151 13973
rect 4337 13968 6151 13970
rect 4337 13912 4342 13968
rect 4398 13912 6090 13968
rect 6146 13912 6151 13968
rect 4337 13910 6151 13912
rect 4337 13907 4403 13910
rect 6085 13907 6151 13910
rect 0 13834 800 13864
rect 1577 13834 1643 13837
rect 0 13832 1643 13834
rect 0 13776 1582 13832
rect 1638 13776 1643 13832
rect 0 13774 1643 13776
rect 0 13744 800 13774
rect 1577 13771 1643 13774
rect 7874 13632 8194 13633
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8194 13632
rect 7874 13567 8194 13568
rect 14805 13632 15125 13633
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 13567 15125 13568
rect 0 13290 800 13320
rect 4061 13290 4127 13293
rect 0 13288 4127 13290
rect 0 13232 4066 13288
rect 4122 13232 4127 13288
rect 0 13230 4127 13232
rect 0 13200 800 13230
rect 4061 13227 4127 13230
rect 6637 13154 6703 13157
rect 8109 13154 8175 13157
rect 6637 13152 8175 13154
rect 6637 13096 6642 13152
rect 6698 13096 8114 13152
rect 8170 13096 8175 13152
rect 6637 13094 8175 13096
rect 6637 13091 6703 13094
rect 8109 13091 8175 13094
rect 4409 13088 4729 13089
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 13023 4729 13024
rect 11340 13088 11660 13089
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 13023 11660 13024
rect 18270 13088 18590 13089
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18590 13088
rect 18270 13023 18590 13024
rect 0 12882 800 12912
rect 3601 12882 3667 12885
rect 0 12880 3667 12882
rect 0 12824 3606 12880
rect 3662 12824 3667 12880
rect 0 12822 3667 12824
rect 0 12792 800 12822
rect 3601 12819 3667 12822
rect 7874 12544 8194 12545
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8194 12544
rect 7874 12479 8194 12480
rect 14805 12544 15125 12545
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 12479 15125 12480
rect 0 12338 800 12368
rect 2865 12338 2931 12341
rect 0 12336 2931 12338
rect 0 12280 2870 12336
rect 2926 12280 2931 12336
rect 0 12278 2931 12280
rect 0 12248 800 12278
rect 2865 12275 2931 12278
rect 4409 12000 4729 12001
rect 0 11930 800 11960
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 11935 4729 11936
rect 11340 12000 11660 12001
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 11935 11660 11936
rect 18270 12000 18590 12001
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18590 12000
rect 18270 11935 18590 11936
rect 3141 11930 3207 11933
rect 0 11928 3207 11930
rect 0 11872 3146 11928
rect 3202 11872 3207 11928
rect 0 11870 3207 11872
rect 0 11840 800 11870
rect 3141 11867 3207 11870
rect 5901 11794 5967 11797
rect 7465 11794 7531 11797
rect 5901 11792 7531 11794
rect 5901 11736 5906 11792
rect 5962 11736 7470 11792
rect 7526 11736 7531 11792
rect 5901 11734 7531 11736
rect 5901 11731 5967 11734
rect 7465 11731 7531 11734
rect 2865 11658 2931 11661
rect 9121 11658 9187 11661
rect 2865 11656 9187 11658
rect 2865 11600 2870 11656
rect 2926 11600 9126 11656
rect 9182 11600 9187 11656
rect 2865 11598 9187 11600
rect 2865 11595 2931 11598
rect 9121 11595 9187 11598
rect 21357 11522 21423 11525
rect 22200 11522 23000 11552
rect 21357 11520 23000 11522
rect 21357 11464 21362 11520
rect 21418 11464 23000 11520
rect 21357 11462 23000 11464
rect 21357 11459 21423 11462
rect 7874 11456 8194 11457
rect 0 11386 800 11416
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8194 11456
rect 7874 11391 8194 11392
rect 14805 11456 15125 11457
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 22200 11432 23000 11462
rect 14805 11391 15125 11392
rect 1485 11386 1551 11389
rect 0 11384 1551 11386
rect 0 11328 1490 11384
rect 1546 11328 1551 11384
rect 0 11326 1551 11328
rect 0 11296 800 11326
rect 1485 11323 1551 11326
rect 0 10978 800 11008
rect 3417 10978 3483 10981
rect 0 10976 3483 10978
rect 0 10920 3422 10976
rect 3478 10920 3483 10976
rect 0 10918 3483 10920
rect 0 10888 800 10918
rect 3417 10915 3483 10918
rect 4409 10912 4729 10913
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 10847 4729 10848
rect 11340 10912 11660 10913
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 10847 11660 10848
rect 18270 10912 18590 10913
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18590 10912
rect 18270 10847 18590 10848
rect 1393 10570 1459 10573
rect 1350 10568 1459 10570
rect 1350 10512 1398 10568
rect 1454 10512 1459 10568
rect 1350 10507 1459 10512
rect 0 10434 800 10464
rect 1350 10434 1410 10507
rect 0 10374 1410 10434
rect 0 10344 800 10374
rect 7874 10368 8194 10369
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8194 10368
rect 7874 10303 8194 10304
rect 14805 10368 15125 10369
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14805 10303 15125 10304
rect 0 10026 800 10056
rect 1393 10026 1459 10029
rect 0 10024 1459 10026
rect 0 9968 1398 10024
rect 1454 9968 1459 10024
rect 0 9966 1459 9968
rect 0 9936 800 9966
rect 1393 9963 1459 9966
rect 4409 9824 4729 9825
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 9759 4729 9760
rect 11340 9824 11660 9825
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 9759 11660 9760
rect 18270 9824 18590 9825
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18590 9824
rect 18270 9759 18590 9760
rect 0 9482 800 9512
rect 1853 9482 1919 9485
rect 0 9480 1919 9482
rect 0 9424 1858 9480
rect 1914 9424 1919 9480
rect 0 9422 1919 9424
rect 0 9392 800 9422
rect 1853 9419 1919 9422
rect 7874 9280 8194 9281
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8194 9280
rect 7874 9215 8194 9216
rect 14805 9280 15125 9281
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 9215 15125 9216
rect 0 9074 800 9104
rect 1393 9074 1459 9077
rect 0 9072 1459 9074
rect 0 9016 1398 9072
rect 1454 9016 1459 9072
rect 0 9014 1459 9016
rect 0 8984 800 9014
rect 1393 9011 1459 9014
rect 4409 8736 4729 8737
rect 0 8666 800 8696
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 8671 4729 8672
rect 11340 8736 11660 8737
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 8671 11660 8672
rect 18270 8736 18590 8737
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18590 8736
rect 18270 8671 18590 8672
rect 2773 8666 2839 8669
rect 0 8664 2839 8666
rect 0 8608 2778 8664
rect 2834 8608 2839 8664
rect 0 8606 2839 8608
rect 0 8576 800 8606
rect 2773 8603 2839 8606
rect 7874 8192 8194 8193
rect 0 8122 800 8152
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8194 8192
rect 7874 8127 8194 8128
rect 14805 8192 15125 8193
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 8127 15125 8128
rect 1853 8122 1919 8125
rect 0 8120 1919 8122
rect 0 8064 1858 8120
rect 1914 8064 1919 8120
rect 0 8062 1919 8064
rect 0 8032 800 8062
rect 1853 8059 1919 8062
rect 0 7714 800 7744
rect 1393 7714 1459 7717
rect 0 7712 1459 7714
rect 0 7656 1398 7712
rect 1454 7656 1459 7712
rect 0 7654 1459 7656
rect 0 7624 800 7654
rect 1393 7651 1459 7654
rect 4409 7648 4729 7649
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 7583 4729 7584
rect 11340 7648 11660 7649
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 7583 11660 7584
rect 18270 7648 18590 7649
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18590 7648
rect 18270 7583 18590 7584
rect 3877 7442 3943 7445
rect 8477 7442 8543 7445
rect 3877 7440 8543 7442
rect 3877 7384 3882 7440
rect 3938 7384 8482 7440
rect 8538 7384 8543 7440
rect 3877 7382 8543 7384
rect 3877 7379 3943 7382
rect 8477 7379 8543 7382
rect 1577 7306 1643 7309
rect 18781 7306 18847 7309
rect 1577 7304 18847 7306
rect 1577 7248 1582 7304
rect 1638 7248 18786 7304
rect 18842 7248 18847 7304
rect 1577 7246 18847 7248
rect 1577 7243 1643 7246
rect 18781 7243 18847 7246
rect 0 7170 800 7200
rect 1393 7170 1459 7173
rect 0 7168 1459 7170
rect 0 7112 1398 7168
rect 1454 7112 1459 7168
rect 0 7110 1459 7112
rect 0 7080 800 7110
rect 1393 7107 1459 7110
rect 7874 7104 8194 7105
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8194 7104
rect 7874 7039 8194 7040
rect 14805 7104 15125 7105
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 7039 15125 7040
rect 0 6762 800 6792
rect 1393 6762 1459 6765
rect 0 6760 1459 6762
rect 0 6704 1398 6760
rect 1454 6704 1459 6760
rect 0 6702 1459 6704
rect 0 6672 800 6702
rect 1393 6699 1459 6702
rect 4409 6560 4729 6561
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 6495 4729 6496
rect 11340 6560 11660 6561
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 6495 11660 6496
rect 18270 6560 18590 6561
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18590 6560
rect 18270 6495 18590 6496
rect 0 6218 800 6248
rect 1393 6218 1459 6221
rect 0 6216 1459 6218
rect 0 6160 1398 6216
rect 1454 6160 1459 6216
rect 0 6158 1459 6160
rect 0 6128 800 6158
rect 1393 6155 1459 6158
rect 7874 6016 8194 6017
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8194 6016
rect 7874 5951 8194 5952
rect 14805 6016 15125 6017
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 5951 15125 5952
rect 0 5810 800 5840
rect 1393 5810 1459 5813
rect 0 5808 1459 5810
rect 0 5752 1398 5808
rect 1454 5752 1459 5808
rect 0 5750 1459 5752
rect 0 5720 800 5750
rect 1393 5747 1459 5750
rect 4409 5472 4729 5473
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 5407 4729 5408
rect 11340 5472 11660 5473
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 5407 11660 5408
rect 18270 5472 18590 5473
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18590 5472
rect 18270 5407 18590 5408
rect 0 5266 800 5296
rect 1393 5266 1459 5269
rect 0 5264 1459 5266
rect 0 5208 1398 5264
rect 1454 5208 1459 5264
rect 0 5206 1459 5208
rect 0 5176 800 5206
rect 1393 5203 1459 5206
rect 7874 4928 8194 4929
rect 0 4858 800 4888
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8194 4928
rect 7874 4863 8194 4864
rect 14805 4928 15125 4929
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 4863 15125 4864
rect 1853 4858 1919 4861
rect 0 4856 1919 4858
rect 0 4800 1858 4856
rect 1914 4800 1919 4856
rect 0 4798 1919 4800
rect 0 4768 800 4798
rect 1853 4795 1919 4798
rect 0 4450 800 4480
rect 1393 4450 1459 4453
rect 0 4448 1459 4450
rect 0 4392 1398 4448
rect 1454 4392 1459 4448
rect 0 4390 1459 4392
rect 0 4360 800 4390
rect 1393 4387 1459 4390
rect 4409 4384 4729 4385
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 4319 4729 4320
rect 11340 4384 11660 4385
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 4319 11660 4320
rect 18270 4384 18590 4385
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18590 4384
rect 18270 4319 18590 4320
rect 0 3906 800 3936
rect 1669 3906 1735 3909
rect 0 3904 1735 3906
rect 0 3848 1674 3904
rect 1730 3848 1735 3904
rect 0 3846 1735 3848
rect 0 3816 800 3846
rect 1669 3843 1735 3846
rect 7874 3840 8194 3841
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8194 3840
rect 7874 3775 8194 3776
rect 14805 3840 15125 3841
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 14805 3775 15125 3776
rect 0 3498 800 3528
rect 1669 3498 1735 3501
rect 0 3496 1735 3498
rect 0 3440 1674 3496
rect 1730 3440 1735 3496
rect 0 3438 1735 3440
rect 0 3408 800 3438
rect 1669 3435 1735 3438
rect 4409 3296 4729 3297
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 3231 4729 3232
rect 11340 3296 11660 3297
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 3231 11660 3232
rect 18270 3296 18590 3297
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18590 3296
rect 18270 3231 18590 3232
rect 0 2954 800 2984
rect 1761 2954 1827 2957
rect 0 2952 1827 2954
rect 0 2896 1766 2952
rect 1822 2896 1827 2952
rect 0 2894 1827 2896
rect 0 2864 800 2894
rect 1761 2891 1827 2894
rect 7874 2752 8194 2753
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8194 2752
rect 7874 2687 8194 2688
rect 14805 2752 15125 2753
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2687 15125 2688
rect 0 2546 800 2576
rect 1669 2546 1735 2549
rect 0 2544 1735 2546
rect 0 2488 1674 2544
rect 1730 2488 1735 2544
rect 0 2486 1735 2488
rect 0 2456 800 2486
rect 1669 2483 1735 2486
rect 4409 2208 4729 2209
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2143 4729 2144
rect 11340 2208 11660 2209
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2143 11660 2144
rect 18270 2208 18590 2209
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18590 2208
rect 18270 2143 18590 2144
rect 0 2002 800 2032
rect 3877 2002 3943 2005
rect 0 2000 3943 2002
rect 0 1944 3882 2000
rect 3938 1944 3943 2000
rect 0 1942 3943 1944
rect 0 1912 800 1942
rect 3877 1939 3943 1942
rect 0 1594 800 1624
rect 3141 1594 3207 1597
rect 0 1592 3207 1594
rect 0 1536 3146 1592
rect 3202 1536 3207 1592
rect 0 1534 3207 1536
rect 0 1504 800 1534
rect 3141 1531 3207 1534
rect 0 1050 800 1080
rect 2773 1050 2839 1053
rect 0 1048 2839 1050
rect 0 992 2778 1048
rect 2834 992 2839 1048
rect 0 990 2839 992
rect 0 960 800 990
rect 2773 987 2839 990
rect 0 642 800 672
rect 2221 642 2287 645
rect 0 640 2287 642
rect 0 584 2226 640
rect 2282 584 2287 640
rect 0 582 2287 584
rect 0 552 800 582
rect 2221 579 2287 582
rect 0 234 800 264
rect 2129 234 2195 237
rect 0 232 2195 234
rect 0 176 2134 232
rect 2190 176 2195 232
rect 0 174 2195 176
rect 0 144 800 174
rect 2129 171 2195 174
<< via3 >>
rect 4417 20700 4481 20704
rect 4417 20644 4421 20700
rect 4421 20644 4477 20700
rect 4477 20644 4481 20700
rect 4417 20640 4481 20644
rect 4497 20700 4561 20704
rect 4497 20644 4501 20700
rect 4501 20644 4557 20700
rect 4557 20644 4561 20700
rect 4497 20640 4561 20644
rect 4577 20700 4641 20704
rect 4577 20644 4581 20700
rect 4581 20644 4637 20700
rect 4637 20644 4641 20700
rect 4577 20640 4641 20644
rect 4657 20700 4721 20704
rect 4657 20644 4661 20700
rect 4661 20644 4717 20700
rect 4717 20644 4721 20700
rect 4657 20640 4721 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 18278 20700 18342 20704
rect 18278 20644 18282 20700
rect 18282 20644 18338 20700
rect 18338 20644 18342 20700
rect 18278 20640 18342 20644
rect 18358 20700 18422 20704
rect 18358 20644 18362 20700
rect 18362 20644 18418 20700
rect 18418 20644 18422 20700
rect 18358 20640 18422 20644
rect 18438 20700 18502 20704
rect 18438 20644 18442 20700
rect 18442 20644 18498 20700
rect 18498 20644 18502 20700
rect 18438 20640 18502 20644
rect 18518 20700 18582 20704
rect 18518 20644 18522 20700
rect 18522 20644 18578 20700
rect 18578 20644 18582 20700
rect 18518 20640 18582 20644
rect 7882 20156 7946 20160
rect 7882 20100 7886 20156
rect 7886 20100 7942 20156
rect 7942 20100 7946 20156
rect 7882 20096 7946 20100
rect 7962 20156 8026 20160
rect 7962 20100 7966 20156
rect 7966 20100 8022 20156
rect 8022 20100 8026 20156
rect 7962 20096 8026 20100
rect 8042 20156 8106 20160
rect 8042 20100 8046 20156
rect 8046 20100 8102 20156
rect 8102 20100 8106 20156
rect 8042 20096 8106 20100
rect 8122 20156 8186 20160
rect 8122 20100 8126 20156
rect 8126 20100 8182 20156
rect 8182 20100 8186 20156
rect 8122 20096 8186 20100
rect 14813 20156 14877 20160
rect 14813 20100 14817 20156
rect 14817 20100 14873 20156
rect 14873 20100 14877 20156
rect 14813 20096 14877 20100
rect 14893 20156 14957 20160
rect 14893 20100 14897 20156
rect 14897 20100 14953 20156
rect 14953 20100 14957 20156
rect 14893 20096 14957 20100
rect 14973 20156 15037 20160
rect 14973 20100 14977 20156
rect 14977 20100 15033 20156
rect 15033 20100 15037 20156
rect 14973 20096 15037 20100
rect 15053 20156 15117 20160
rect 15053 20100 15057 20156
rect 15057 20100 15113 20156
rect 15113 20100 15117 20156
rect 15053 20096 15117 20100
rect 4417 19612 4481 19616
rect 4417 19556 4421 19612
rect 4421 19556 4477 19612
rect 4477 19556 4481 19612
rect 4417 19552 4481 19556
rect 4497 19612 4561 19616
rect 4497 19556 4501 19612
rect 4501 19556 4557 19612
rect 4557 19556 4561 19612
rect 4497 19552 4561 19556
rect 4577 19612 4641 19616
rect 4577 19556 4581 19612
rect 4581 19556 4637 19612
rect 4637 19556 4641 19612
rect 4577 19552 4641 19556
rect 4657 19612 4721 19616
rect 4657 19556 4661 19612
rect 4661 19556 4717 19612
rect 4717 19556 4721 19612
rect 4657 19552 4721 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 18278 19612 18342 19616
rect 18278 19556 18282 19612
rect 18282 19556 18338 19612
rect 18338 19556 18342 19612
rect 18278 19552 18342 19556
rect 18358 19612 18422 19616
rect 18358 19556 18362 19612
rect 18362 19556 18418 19612
rect 18418 19556 18422 19612
rect 18358 19552 18422 19556
rect 18438 19612 18502 19616
rect 18438 19556 18442 19612
rect 18442 19556 18498 19612
rect 18498 19556 18502 19612
rect 18438 19552 18502 19556
rect 18518 19612 18582 19616
rect 18518 19556 18522 19612
rect 18522 19556 18578 19612
rect 18578 19556 18582 19612
rect 18518 19552 18582 19556
rect 7882 19068 7946 19072
rect 7882 19012 7886 19068
rect 7886 19012 7942 19068
rect 7942 19012 7946 19068
rect 7882 19008 7946 19012
rect 7962 19068 8026 19072
rect 7962 19012 7966 19068
rect 7966 19012 8022 19068
rect 8022 19012 8026 19068
rect 7962 19008 8026 19012
rect 8042 19068 8106 19072
rect 8042 19012 8046 19068
rect 8046 19012 8102 19068
rect 8102 19012 8106 19068
rect 8042 19008 8106 19012
rect 8122 19068 8186 19072
rect 8122 19012 8126 19068
rect 8126 19012 8182 19068
rect 8182 19012 8186 19068
rect 8122 19008 8186 19012
rect 14813 19068 14877 19072
rect 14813 19012 14817 19068
rect 14817 19012 14873 19068
rect 14873 19012 14877 19068
rect 14813 19008 14877 19012
rect 14893 19068 14957 19072
rect 14893 19012 14897 19068
rect 14897 19012 14953 19068
rect 14953 19012 14957 19068
rect 14893 19008 14957 19012
rect 14973 19068 15037 19072
rect 14973 19012 14977 19068
rect 14977 19012 15033 19068
rect 15033 19012 15037 19068
rect 14973 19008 15037 19012
rect 15053 19068 15117 19072
rect 15053 19012 15057 19068
rect 15057 19012 15113 19068
rect 15113 19012 15117 19068
rect 15053 19008 15117 19012
rect 4417 18524 4481 18528
rect 4417 18468 4421 18524
rect 4421 18468 4477 18524
rect 4477 18468 4481 18524
rect 4417 18464 4481 18468
rect 4497 18524 4561 18528
rect 4497 18468 4501 18524
rect 4501 18468 4557 18524
rect 4557 18468 4561 18524
rect 4497 18464 4561 18468
rect 4577 18524 4641 18528
rect 4577 18468 4581 18524
rect 4581 18468 4637 18524
rect 4637 18468 4641 18524
rect 4577 18464 4641 18468
rect 4657 18524 4721 18528
rect 4657 18468 4661 18524
rect 4661 18468 4717 18524
rect 4717 18468 4721 18524
rect 4657 18464 4721 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 18278 18524 18342 18528
rect 18278 18468 18282 18524
rect 18282 18468 18338 18524
rect 18338 18468 18342 18524
rect 18278 18464 18342 18468
rect 18358 18524 18422 18528
rect 18358 18468 18362 18524
rect 18362 18468 18418 18524
rect 18418 18468 18422 18524
rect 18358 18464 18422 18468
rect 18438 18524 18502 18528
rect 18438 18468 18442 18524
rect 18442 18468 18498 18524
rect 18498 18468 18502 18524
rect 18438 18464 18502 18468
rect 18518 18524 18582 18528
rect 18518 18468 18522 18524
rect 18522 18468 18578 18524
rect 18578 18468 18582 18524
rect 18518 18464 18582 18468
rect 7882 17980 7946 17984
rect 7882 17924 7886 17980
rect 7886 17924 7942 17980
rect 7942 17924 7946 17980
rect 7882 17920 7946 17924
rect 7962 17980 8026 17984
rect 7962 17924 7966 17980
rect 7966 17924 8022 17980
rect 8022 17924 8026 17980
rect 7962 17920 8026 17924
rect 8042 17980 8106 17984
rect 8042 17924 8046 17980
rect 8046 17924 8102 17980
rect 8102 17924 8106 17980
rect 8042 17920 8106 17924
rect 8122 17980 8186 17984
rect 8122 17924 8126 17980
rect 8126 17924 8182 17980
rect 8182 17924 8186 17980
rect 8122 17920 8186 17924
rect 14813 17980 14877 17984
rect 14813 17924 14817 17980
rect 14817 17924 14873 17980
rect 14873 17924 14877 17980
rect 14813 17920 14877 17924
rect 14893 17980 14957 17984
rect 14893 17924 14897 17980
rect 14897 17924 14953 17980
rect 14953 17924 14957 17980
rect 14893 17920 14957 17924
rect 14973 17980 15037 17984
rect 14973 17924 14977 17980
rect 14977 17924 15033 17980
rect 15033 17924 15037 17980
rect 14973 17920 15037 17924
rect 15053 17980 15117 17984
rect 15053 17924 15057 17980
rect 15057 17924 15113 17980
rect 15113 17924 15117 17980
rect 15053 17920 15117 17924
rect 4417 17436 4481 17440
rect 4417 17380 4421 17436
rect 4421 17380 4477 17436
rect 4477 17380 4481 17436
rect 4417 17376 4481 17380
rect 4497 17436 4561 17440
rect 4497 17380 4501 17436
rect 4501 17380 4557 17436
rect 4557 17380 4561 17436
rect 4497 17376 4561 17380
rect 4577 17436 4641 17440
rect 4577 17380 4581 17436
rect 4581 17380 4637 17436
rect 4637 17380 4641 17436
rect 4577 17376 4641 17380
rect 4657 17436 4721 17440
rect 4657 17380 4661 17436
rect 4661 17380 4717 17436
rect 4717 17380 4721 17436
rect 4657 17376 4721 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 18278 17436 18342 17440
rect 18278 17380 18282 17436
rect 18282 17380 18338 17436
rect 18338 17380 18342 17436
rect 18278 17376 18342 17380
rect 18358 17436 18422 17440
rect 18358 17380 18362 17436
rect 18362 17380 18418 17436
rect 18418 17380 18422 17436
rect 18358 17376 18422 17380
rect 18438 17436 18502 17440
rect 18438 17380 18442 17436
rect 18442 17380 18498 17436
rect 18498 17380 18502 17436
rect 18438 17376 18502 17380
rect 18518 17436 18582 17440
rect 18518 17380 18522 17436
rect 18522 17380 18578 17436
rect 18578 17380 18582 17436
rect 18518 17376 18582 17380
rect 7882 16892 7946 16896
rect 7882 16836 7886 16892
rect 7886 16836 7942 16892
rect 7942 16836 7946 16892
rect 7882 16832 7946 16836
rect 7962 16892 8026 16896
rect 7962 16836 7966 16892
rect 7966 16836 8022 16892
rect 8022 16836 8026 16892
rect 7962 16832 8026 16836
rect 8042 16892 8106 16896
rect 8042 16836 8046 16892
rect 8046 16836 8102 16892
rect 8102 16836 8106 16892
rect 8042 16832 8106 16836
rect 8122 16892 8186 16896
rect 8122 16836 8126 16892
rect 8126 16836 8182 16892
rect 8182 16836 8186 16892
rect 8122 16832 8186 16836
rect 14813 16892 14877 16896
rect 14813 16836 14817 16892
rect 14817 16836 14873 16892
rect 14873 16836 14877 16892
rect 14813 16832 14877 16836
rect 14893 16892 14957 16896
rect 14893 16836 14897 16892
rect 14897 16836 14953 16892
rect 14953 16836 14957 16892
rect 14893 16832 14957 16836
rect 14973 16892 15037 16896
rect 14973 16836 14977 16892
rect 14977 16836 15033 16892
rect 15033 16836 15037 16892
rect 14973 16832 15037 16836
rect 15053 16892 15117 16896
rect 15053 16836 15057 16892
rect 15057 16836 15113 16892
rect 15113 16836 15117 16892
rect 15053 16832 15117 16836
rect 4417 16348 4481 16352
rect 4417 16292 4421 16348
rect 4421 16292 4477 16348
rect 4477 16292 4481 16348
rect 4417 16288 4481 16292
rect 4497 16348 4561 16352
rect 4497 16292 4501 16348
rect 4501 16292 4557 16348
rect 4557 16292 4561 16348
rect 4497 16288 4561 16292
rect 4577 16348 4641 16352
rect 4577 16292 4581 16348
rect 4581 16292 4637 16348
rect 4637 16292 4641 16348
rect 4577 16288 4641 16292
rect 4657 16348 4721 16352
rect 4657 16292 4661 16348
rect 4661 16292 4717 16348
rect 4717 16292 4721 16348
rect 4657 16288 4721 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 18278 16348 18342 16352
rect 18278 16292 18282 16348
rect 18282 16292 18338 16348
rect 18338 16292 18342 16348
rect 18278 16288 18342 16292
rect 18358 16348 18422 16352
rect 18358 16292 18362 16348
rect 18362 16292 18418 16348
rect 18418 16292 18422 16348
rect 18358 16288 18422 16292
rect 18438 16348 18502 16352
rect 18438 16292 18442 16348
rect 18442 16292 18498 16348
rect 18498 16292 18502 16348
rect 18438 16288 18502 16292
rect 18518 16348 18582 16352
rect 18518 16292 18522 16348
rect 18522 16292 18578 16348
rect 18578 16292 18582 16348
rect 18518 16288 18582 16292
rect 7882 15804 7946 15808
rect 7882 15748 7886 15804
rect 7886 15748 7942 15804
rect 7942 15748 7946 15804
rect 7882 15744 7946 15748
rect 7962 15804 8026 15808
rect 7962 15748 7966 15804
rect 7966 15748 8022 15804
rect 8022 15748 8026 15804
rect 7962 15744 8026 15748
rect 8042 15804 8106 15808
rect 8042 15748 8046 15804
rect 8046 15748 8102 15804
rect 8102 15748 8106 15804
rect 8042 15744 8106 15748
rect 8122 15804 8186 15808
rect 8122 15748 8126 15804
rect 8126 15748 8182 15804
rect 8182 15748 8186 15804
rect 8122 15744 8186 15748
rect 14813 15804 14877 15808
rect 14813 15748 14817 15804
rect 14817 15748 14873 15804
rect 14873 15748 14877 15804
rect 14813 15744 14877 15748
rect 14893 15804 14957 15808
rect 14893 15748 14897 15804
rect 14897 15748 14953 15804
rect 14953 15748 14957 15804
rect 14893 15744 14957 15748
rect 14973 15804 15037 15808
rect 14973 15748 14977 15804
rect 14977 15748 15033 15804
rect 15033 15748 15037 15804
rect 14973 15744 15037 15748
rect 15053 15804 15117 15808
rect 15053 15748 15057 15804
rect 15057 15748 15113 15804
rect 15113 15748 15117 15804
rect 15053 15744 15117 15748
rect 4417 15260 4481 15264
rect 4417 15204 4421 15260
rect 4421 15204 4477 15260
rect 4477 15204 4481 15260
rect 4417 15200 4481 15204
rect 4497 15260 4561 15264
rect 4497 15204 4501 15260
rect 4501 15204 4557 15260
rect 4557 15204 4561 15260
rect 4497 15200 4561 15204
rect 4577 15260 4641 15264
rect 4577 15204 4581 15260
rect 4581 15204 4637 15260
rect 4637 15204 4641 15260
rect 4577 15200 4641 15204
rect 4657 15260 4721 15264
rect 4657 15204 4661 15260
rect 4661 15204 4717 15260
rect 4717 15204 4721 15260
rect 4657 15200 4721 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 18278 15260 18342 15264
rect 18278 15204 18282 15260
rect 18282 15204 18338 15260
rect 18338 15204 18342 15260
rect 18278 15200 18342 15204
rect 18358 15260 18422 15264
rect 18358 15204 18362 15260
rect 18362 15204 18418 15260
rect 18418 15204 18422 15260
rect 18358 15200 18422 15204
rect 18438 15260 18502 15264
rect 18438 15204 18442 15260
rect 18442 15204 18498 15260
rect 18498 15204 18502 15260
rect 18438 15200 18502 15204
rect 18518 15260 18582 15264
rect 18518 15204 18522 15260
rect 18522 15204 18578 15260
rect 18578 15204 18582 15260
rect 18518 15200 18582 15204
rect 7882 14716 7946 14720
rect 7882 14660 7886 14716
rect 7886 14660 7942 14716
rect 7942 14660 7946 14716
rect 7882 14656 7946 14660
rect 7962 14716 8026 14720
rect 7962 14660 7966 14716
rect 7966 14660 8022 14716
rect 8022 14660 8026 14716
rect 7962 14656 8026 14660
rect 8042 14716 8106 14720
rect 8042 14660 8046 14716
rect 8046 14660 8102 14716
rect 8102 14660 8106 14716
rect 8042 14656 8106 14660
rect 8122 14716 8186 14720
rect 8122 14660 8126 14716
rect 8126 14660 8182 14716
rect 8182 14660 8186 14716
rect 8122 14656 8186 14660
rect 14813 14716 14877 14720
rect 14813 14660 14817 14716
rect 14817 14660 14873 14716
rect 14873 14660 14877 14716
rect 14813 14656 14877 14660
rect 14893 14716 14957 14720
rect 14893 14660 14897 14716
rect 14897 14660 14953 14716
rect 14953 14660 14957 14716
rect 14893 14656 14957 14660
rect 14973 14716 15037 14720
rect 14973 14660 14977 14716
rect 14977 14660 15033 14716
rect 15033 14660 15037 14716
rect 14973 14656 15037 14660
rect 15053 14716 15117 14720
rect 15053 14660 15057 14716
rect 15057 14660 15113 14716
rect 15113 14660 15117 14716
rect 15053 14656 15117 14660
rect 4417 14172 4481 14176
rect 4417 14116 4421 14172
rect 4421 14116 4477 14172
rect 4477 14116 4481 14172
rect 4417 14112 4481 14116
rect 4497 14172 4561 14176
rect 4497 14116 4501 14172
rect 4501 14116 4557 14172
rect 4557 14116 4561 14172
rect 4497 14112 4561 14116
rect 4577 14172 4641 14176
rect 4577 14116 4581 14172
rect 4581 14116 4637 14172
rect 4637 14116 4641 14172
rect 4577 14112 4641 14116
rect 4657 14172 4721 14176
rect 4657 14116 4661 14172
rect 4661 14116 4717 14172
rect 4717 14116 4721 14172
rect 4657 14112 4721 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 18278 14172 18342 14176
rect 18278 14116 18282 14172
rect 18282 14116 18338 14172
rect 18338 14116 18342 14172
rect 18278 14112 18342 14116
rect 18358 14172 18422 14176
rect 18358 14116 18362 14172
rect 18362 14116 18418 14172
rect 18418 14116 18422 14172
rect 18358 14112 18422 14116
rect 18438 14172 18502 14176
rect 18438 14116 18442 14172
rect 18442 14116 18498 14172
rect 18498 14116 18502 14172
rect 18438 14112 18502 14116
rect 18518 14172 18582 14176
rect 18518 14116 18522 14172
rect 18522 14116 18578 14172
rect 18578 14116 18582 14172
rect 18518 14112 18582 14116
rect 7882 13628 7946 13632
rect 7882 13572 7886 13628
rect 7886 13572 7942 13628
rect 7942 13572 7946 13628
rect 7882 13568 7946 13572
rect 7962 13628 8026 13632
rect 7962 13572 7966 13628
rect 7966 13572 8022 13628
rect 8022 13572 8026 13628
rect 7962 13568 8026 13572
rect 8042 13628 8106 13632
rect 8042 13572 8046 13628
rect 8046 13572 8102 13628
rect 8102 13572 8106 13628
rect 8042 13568 8106 13572
rect 8122 13628 8186 13632
rect 8122 13572 8126 13628
rect 8126 13572 8182 13628
rect 8182 13572 8186 13628
rect 8122 13568 8186 13572
rect 14813 13628 14877 13632
rect 14813 13572 14817 13628
rect 14817 13572 14873 13628
rect 14873 13572 14877 13628
rect 14813 13568 14877 13572
rect 14893 13628 14957 13632
rect 14893 13572 14897 13628
rect 14897 13572 14953 13628
rect 14953 13572 14957 13628
rect 14893 13568 14957 13572
rect 14973 13628 15037 13632
rect 14973 13572 14977 13628
rect 14977 13572 15033 13628
rect 15033 13572 15037 13628
rect 14973 13568 15037 13572
rect 15053 13628 15117 13632
rect 15053 13572 15057 13628
rect 15057 13572 15113 13628
rect 15113 13572 15117 13628
rect 15053 13568 15117 13572
rect 4417 13084 4481 13088
rect 4417 13028 4421 13084
rect 4421 13028 4477 13084
rect 4477 13028 4481 13084
rect 4417 13024 4481 13028
rect 4497 13084 4561 13088
rect 4497 13028 4501 13084
rect 4501 13028 4557 13084
rect 4557 13028 4561 13084
rect 4497 13024 4561 13028
rect 4577 13084 4641 13088
rect 4577 13028 4581 13084
rect 4581 13028 4637 13084
rect 4637 13028 4641 13084
rect 4577 13024 4641 13028
rect 4657 13084 4721 13088
rect 4657 13028 4661 13084
rect 4661 13028 4717 13084
rect 4717 13028 4721 13084
rect 4657 13024 4721 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 18278 13084 18342 13088
rect 18278 13028 18282 13084
rect 18282 13028 18338 13084
rect 18338 13028 18342 13084
rect 18278 13024 18342 13028
rect 18358 13084 18422 13088
rect 18358 13028 18362 13084
rect 18362 13028 18418 13084
rect 18418 13028 18422 13084
rect 18358 13024 18422 13028
rect 18438 13084 18502 13088
rect 18438 13028 18442 13084
rect 18442 13028 18498 13084
rect 18498 13028 18502 13084
rect 18438 13024 18502 13028
rect 18518 13084 18582 13088
rect 18518 13028 18522 13084
rect 18522 13028 18578 13084
rect 18578 13028 18582 13084
rect 18518 13024 18582 13028
rect 7882 12540 7946 12544
rect 7882 12484 7886 12540
rect 7886 12484 7942 12540
rect 7942 12484 7946 12540
rect 7882 12480 7946 12484
rect 7962 12540 8026 12544
rect 7962 12484 7966 12540
rect 7966 12484 8022 12540
rect 8022 12484 8026 12540
rect 7962 12480 8026 12484
rect 8042 12540 8106 12544
rect 8042 12484 8046 12540
rect 8046 12484 8102 12540
rect 8102 12484 8106 12540
rect 8042 12480 8106 12484
rect 8122 12540 8186 12544
rect 8122 12484 8126 12540
rect 8126 12484 8182 12540
rect 8182 12484 8186 12540
rect 8122 12480 8186 12484
rect 14813 12540 14877 12544
rect 14813 12484 14817 12540
rect 14817 12484 14873 12540
rect 14873 12484 14877 12540
rect 14813 12480 14877 12484
rect 14893 12540 14957 12544
rect 14893 12484 14897 12540
rect 14897 12484 14953 12540
rect 14953 12484 14957 12540
rect 14893 12480 14957 12484
rect 14973 12540 15037 12544
rect 14973 12484 14977 12540
rect 14977 12484 15033 12540
rect 15033 12484 15037 12540
rect 14973 12480 15037 12484
rect 15053 12540 15117 12544
rect 15053 12484 15057 12540
rect 15057 12484 15113 12540
rect 15113 12484 15117 12540
rect 15053 12480 15117 12484
rect 4417 11996 4481 12000
rect 4417 11940 4421 11996
rect 4421 11940 4477 11996
rect 4477 11940 4481 11996
rect 4417 11936 4481 11940
rect 4497 11996 4561 12000
rect 4497 11940 4501 11996
rect 4501 11940 4557 11996
rect 4557 11940 4561 11996
rect 4497 11936 4561 11940
rect 4577 11996 4641 12000
rect 4577 11940 4581 11996
rect 4581 11940 4637 11996
rect 4637 11940 4641 11996
rect 4577 11936 4641 11940
rect 4657 11996 4721 12000
rect 4657 11940 4661 11996
rect 4661 11940 4717 11996
rect 4717 11940 4721 11996
rect 4657 11936 4721 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 18278 11996 18342 12000
rect 18278 11940 18282 11996
rect 18282 11940 18338 11996
rect 18338 11940 18342 11996
rect 18278 11936 18342 11940
rect 18358 11996 18422 12000
rect 18358 11940 18362 11996
rect 18362 11940 18418 11996
rect 18418 11940 18422 11996
rect 18358 11936 18422 11940
rect 18438 11996 18502 12000
rect 18438 11940 18442 11996
rect 18442 11940 18498 11996
rect 18498 11940 18502 11996
rect 18438 11936 18502 11940
rect 18518 11996 18582 12000
rect 18518 11940 18522 11996
rect 18522 11940 18578 11996
rect 18578 11940 18582 11996
rect 18518 11936 18582 11940
rect 7882 11452 7946 11456
rect 7882 11396 7886 11452
rect 7886 11396 7942 11452
rect 7942 11396 7946 11452
rect 7882 11392 7946 11396
rect 7962 11452 8026 11456
rect 7962 11396 7966 11452
rect 7966 11396 8022 11452
rect 8022 11396 8026 11452
rect 7962 11392 8026 11396
rect 8042 11452 8106 11456
rect 8042 11396 8046 11452
rect 8046 11396 8102 11452
rect 8102 11396 8106 11452
rect 8042 11392 8106 11396
rect 8122 11452 8186 11456
rect 8122 11396 8126 11452
rect 8126 11396 8182 11452
rect 8182 11396 8186 11452
rect 8122 11392 8186 11396
rect 14813 11452 14877 11456
rect 14813 11396 14817 11452
rect 14817 11396 14873 11452
rect 14873 11396 14877 11452
rect 14813 11392 14877 11396
rect 14893 11452 14957 11456
rect 14893 11396 14897 11452
rect 14897 11396 14953 11452
rect 14953 11396 14957 11452
rect 14893 11392 14957 11396
rect 14973 11452 15037 11456
rect 14973 11396 14977 11452
rect 14977 11396 15033 11452
rect 15033 11396 15037 11452
rect 14973 11392 15037 11396
rect 15053 11452 15117 11456
rect 15053 11396 15057 11452
rect 15057 11396 15113 11452
rect 15113 11396 15117 11452
rect 15053 11392 15117 11396
rect 4417 10908 4481 10912
rect 4417 10852 4421 10908
rect 4421 10852 4477 10908
rect 4477 10852 4481 10908
rect 4417 10848 4481 10852
rect 4497 10908 4561 10912
rect 4497 10852 4501 10908
rect 4501 10852 4557 10908
rect 4557 10852 4561 10908
rect 4497 10848 4561 10852
rect 4577 10908 4641 10912
rect 4577 10852 4581 10908
rect 4581 10852 4637 10908
rect 4637 10852 4641 10908
rect 4577 10848 4641 10852
rect 4657 10908 4721 10912
rect 4657 10852 4661 10908
rect 4661 10852 4717 10908
rect 4717 10852 4721 10908
rect 4657 10848 4721 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 18278 10908 18342 10912
rect 18278 10852 18282 10908
rect 18282 10852 18338 10908
rect 18338 10852 18342 10908
rect 18278 10848 18342 10852
rect 18358 10908 18422 10912
rect 18358 10852 18362 10908
rect 18362 10852 18418 10908
rect 18418 10852 18422 10908
rect 18358 10848 18422 10852
rect 18438 10908 18502 10912
rect 18438 10852 18442 10908
rect 18442 10852 18498 10908
rect 18498 10852 18502 10908
rect 18438 10848 18502 10852
rect 18518 10908 18582 10912
rect 18518 10852 18522 10908
rect 18522 10852 18578 10908
rect 18578 10852 18582 10908
rect 18518 10848 18582 10852
rect 7882 10364 7946 10368
rect 7882 10308 7886 10364
rect 7886 10308 7942 10364
rect 7942 10308 7946 10364
rect 7882 10304 7946 10308
rect 7962 10364 8026 10368
rect 7962 10308 7966 10364
rect 7966 10308 8022 10364
rect 8022 10308 8026 10364
rect 7962 10304 8026 10308
rect 8042 10364 8106 10368
rect 8042 10308 8046 10364
rect 8046 10308 8102 10364
rect 8102 10308 8106 10364
rect 8042 10304 8106 10308
rect 8122 10364 8186 10368
rect 8122 10308 8126 10364
rect 8126 10308 8182 10364
rect 8182 10308 8186 10364
rect 8122 10304 8186 10308
rect 14813 10364 14877 10368
rect 14813 10308 14817 10364
rect 14817 10308 14873 10364
rect 14873 10308 14877 10364
rect 14813 10304 14877 10308
rect 14893 10364 14957 10368
rect 14893 10308 14897 10364
rect 14897 10308 14953 10364
rect 14953 10308 14957 10364
rect 14893 10304 14957 10308
rect 14973 10364 15037 10368
rect 14973 10308 14977 10364
rect 14977 10308 15033 10364
rect 15033 10308 15037 10364
rect 14973 10304 15037 10308
rect 15053 10364 15117 10368
rect 15053 10308 15057 10364
rect 15057 10308 15113 10364
rect 15113 10308 15117 10364
rect 15053 10304 15117 10308
rect 4417 9820 4481 9824
rect 4417 9764 4421 9820
rect 4421 9764 4477 9820
rect 4477 9764 4481 9820
rect 4417 9760 4481 9764
rect 4497 9820 4561 9824
rect 4497 9764 4501 9820
rect 4501 9764 4557 9820
rect 4557 9764 4561 9820
rect 4497 9760 4561 9764
rect 4577 9820 4641 9824
rect 4577 9764 4581 9820
rect 4581 9764 4637 9820
rect 4637 9764 4641 9820
rect 4577 9760 4641 9764
rect 4657 9820 4721 9824
rect 4657 9764 4661 9820
rect 4661 9764 4717 9820
rect 4717 9764 4721 9820
rect 4657 9760 4721 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 18278 9820 18342 9824
rect 18278 9764 18282 9820
rect 18282 9764 18338 9820
rect 18338 9764 18342 9820
rect 18278 9760 18342 9764
rect 18358 9820 18422 9824
rect 18358 9764 18362 9820
rect 18362 9764 18418 9820
rect 18418 9764 18422 9820
rect 18358 9760 18422 9764
rect 18438 9820 18502 9824
rect 18438 9764 18442 9820
rect 18442 9764 18498 9820
rect 18498 9764 18502 9820
rect 18438 9760 18502 9764
rect 18518 9820 18582 9824
rect 18518 9764 18522 9820
rect 18522 9764 18578 9820
rect 18578 9764 18582 9820
rect 18518 9760 18582 9764
rect 7882 9276 7946 9280
rect 7882 9220 7886 9276
rect 7886 9220 7942 9276
rect 7942 9220 7946 9276
rect 7882 9216 7946 9220
rect 7962 9276 8026 9280
rect 7962 9220 7966 9276
rect 7966 9220 8022 9276
rect 8022 9220 8026 9276
rect 7962 9216 8026 9220
rect 8042 9276 8106 9280
rect 8042 9220 8046 9276
rect 8046 9220 8102 9276
rect 8102 9220 8106 9276
rect 8042 9216 8106 9220
rect 8122 9276 8186 9280
rect 8122 9220 8126 9276
rect 8126 9220 8182 9276
rect 8182 9220 8186 9276
rect 8122 9216 8186 9220
rect 14813 9276 14877 9280
rect 14813 9220 14817 9276
rect 14817 9220 14873 9276
rect 14873 9220 14877 9276
rect 14813 9216 14877 9220
rect 14893 9276 14957 9280
rect 14893 9220 14897 9276
rect 14897 9220 14953 9276
rect 14953 9220 14957 9276
rect 14893 9216 14957 9220
rect 14973 9276 15037 9280
rect 14973 9220 14977 9276
rect 14977 9220 15033 9276
rect 15033 9220 15037 9276
rect 14973 9216 15037 9220
rect 15053 9276 15117 9280
rect 15053 9220 15057 9276
rect 15057 9220 15113 9276
rect 15113 9220 15117 9276
rect 15053 9216 15117 9220
rect 4417 8732 4481 8736
rect 4417 8676 4421 8732
rect 4421 8676 4477 8732
rect 4477 8676 4481 8732
rect 4417 8672 4481 8676
rect 4497 8732 4561 8736
rect 4497 8676 4501 8732
rect 4501 8676 4557 8732
rect 4557 8676 4561 8732
rect 4497 8672 4561 8676
rect 4577 8732 4641 8736
rect 4577 8676 4581 8732
rect 4581 8676 4637 8732
rect 4637 8676 4641 8732
rect 4577 8672 4641 8676
rect 4657 8732 4721 8736
rect 4657 8676 4661 8732
rect 4661 8676 4717 8732
rect 4717 8676 4721 8732
rect 4657 8672 4721 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 18278 8732 18342 8736
rect 18278 8676 18282 8732
rect 18282 8676 18338 8732
rect 18338 8676 18342 8732
rect 18278 8672 18342 8676
rect 18358 8732 18422 8736
rect 18358 8676 18362 8732
rect 18362 8676 18418 8732
rect 18418 8676 18422 8732
rect 18358 8672 18422 8676
rect 18438 8732 18502 8736
rect 18438 8676 18442 8732
rect 18442 8676 18498 8732
rect 18498 8676 18502 8732
rect 18438 8672 18502 8676
rect 18518 8732 18582 8736
rect 18518 8676 18522 8732
rect 18522 8676 18578 8732
rect 18578 8676 18582 8732
rect 18518 8672 18582 8676
rect 7882 8188 7946 8192
rect 7882 8132 7886 8188
rect 7886 8132 7942 8188
rect 7942 8132 7946 8188
rect 7882 8128 7946 8132
rect 7962 8188 8026 8192
rect 7962 8132 7966 8188
rect 7966 8132 8022 8188
rect 8022 8132 8026 8188
rect 7962 8128 8026 8132
rect 8042 8188 8106 8192
rect 8042 8132 8046 8188
rect 8046 8132 8102 8188
rect 8102 8132 8106 8188
rect 8042 8128 8106 8132
rect 8122 8188 8186 8192
rect 8122 8132 8126 8188
rect 8126 8132 8182 8188
rect 8182 8132 8186 8188
rect 8122 8128 8186 8132
rect 14813 8188 14877 8192
rect 14813 8132 14817 8188
rect 14817 8132 14873 8188
rect 14873 8132 14877 8188
rect 14813 8128 14877 8132
rect 14893 8188 14957 8192
rect 14893 8132 14897 8188
rect 14897 8132 14953 8188
rect 14953 8132 14957 8188
rect 14893 8128 14957 8132
rect 14973 8188 15037 8192
rect 14973 8132 14977 8188
rect 14977 8132 15033 8188
rect 15033 8132 15037 8188
rect 14973 8128 15037 8132
rect 15053 8188 15117 8192
rect 15053 8132 15057 8188
rect 15057 8132 15113 8188
rect 15113 8132 15117 8188
rect 15053 8128 15117 8132
rect 4417 7644 4481 7648
rect 4417 7588 4421 7644
rect 4421 7588 4477 7644
rect 4477 7588 4481 7644
rect 4417 7584 4481 7588
rect 4497 7644 4561 7648
rect 4497 7588 4501 7644
rect 4501 7588 4557 7644
rect 4557 7588 4561 7644
rect 4497 7584 4561 7588
rect 4577 7644 4641 7648
rect 4577 7588 4581 7644
rect 4581 7588 4637 7644
rect 4637 7588 4641 7644
rect 4577 7584 4641 7588
rect 4657 7644 4721 7648
rect 4657 7588 4661 7644
rect 4661 7588 4717 7644
rect 4717 7588 4721 7644
rect 4657 7584 4721 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 18278 7644 18342 7648
rect 18278 7588 18282 7644
rect 18282 7588 18338 7644
rect 18338 7588 18342 7644
rect 18278 7584 18342 7588
rect 18358 7644 18422 7648
rect 18358 7588 18362 7644
rect 18362 7588 18418 7644
rect 18418 7588 18422 7644
rect 18358 7584 18422 7588
rect 18438 7644 18502 7648
rect 18438 7588 18442 7644
rect 18442 7588 18498 7644
rect 18498 7588 18502 7644
rect 18438 7584 18502 7588
rect 18518 7644 18582 7648
rect 18518 7588 18522 7644
rect 18522 7588 18578 7644
rect 18578 7588 18582 7644
rect 18518 7584 18582 7588
rect 7882 7100 7946 7104
rect 7882 7044 7886 7100
rect 7886 7044 7942 7100
rect 7942 7044 7946 7100
rect 7882 7040 7946 7044
rect 7962 7100 8026 7104
rect 7962 7044 7966 7100
rect 7966 7044 8022 7100
rect 8022 7044 8026 7100
rect 7962 7040 8026 7044
rect 8042 7100 8106 7104
rect 8042 7044 8046 7100
rect 8046 7044 8102 7100
rect 8102 7044 8106 7100
rect 8042 7040 8106 7044
rect 8122 7100 8186 7104
rect 8122 7044 8126 7100
rect 8126 7044 8182 7100
rect 8182 7044 8186 7100
rect 8122 7040 8186 7044
rect 14813 7100 14877 7104
rect 14813 7044 14817 7100
rect 14817 7044 14873 7100
rect 14873 7044 14877 7100
rect 14813 7040 14877 7044
rect 14893 7100 14957 7104
rect 14893 7044 14897 7100
rect 14897 7044 14953 7100
rect 14953 7044 14957 7100
rect 14893 7040 14957 7044
rect 14973 7100 15037 7104
rect 14973 7044 14977 7100
rect 14977 7044 15033 7100
rect 15033 7044 15037 7100
rect 14973 7040 15037 7044
rect 15053 7100 15117 7104
rect 15053 7044 15057 7100
rect 15057 7044 15113 7100
rect 15113 7044 15117 7100
rect 15053 7040 15117 7044
rect 4417 6556 4481 6560
rect 4417 6500 4421 6556
rect 4421 6500 4477 6556
rect 4477 6500 4481 6556
rect 4417 6496 4481 6500
rect 4497 6556 4561 6560
rect 4497 6500 4501 6556
rect 4501 6500 4557 6556
rect 4557 6500 4561 6556
rect 4497 6496 4561 6500
rect 4577 6556 4641 6560
rect 4577 6500 4581 6556
rect 4581 6500 4637 6556
rect 4637 6500 4641 6556
rect 4577 6496 4641 6500
rect 4657 6556 4721 6560
rect 4657 6500 4661 6556
rect 4661 6500 4717 6556
rect 4717 6500 4721 6556
rect 4657 6496 4721 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 18278 6556 18342 6560
rect 18278 6500 18282 6556
rect 18282 6500 18338 6556
rect 18338 6500 18342 6556
rect 18278 6496 18342 6500
rect 18358 6556 18422 6560
rect 18358 6500 18362 6556
rect 18362 6500 18418 6556
rect 18418 6500 18422 6556
rect 18358 6496 18422 6500
rect 18438 6556 18502 6560
rect 18438 6500 18442 6556
rect 18442 6500 18498 6556
rect 18498 6500 18502 6556
rect 18438 6496 18502 6500
rect 18518 6556 18582 6560
rect 18518 6500 18522 6556
rect 18522 6500 18578 6556
rect 18578 6500 18582 6556
rect 18518 6496 18582 6500
rect 7882 6012 7946 6016
rect 7882 5956 7886 6012
rect 7886 5956 7942 6012
rect 7942 5956 7946 6012
rect 7882 5952 7946 5956
rect 7962 6012 8026 6016
rect 7962 5956 7966 6012
rect 7966 5956 8022 6012
rect 8022 5956 8026 6012
rect 7962 5952 8026 5956
rect 8042 6012 8106 6016
rect 8042 5956 8046 6012
rect 8046 5956 8102 6012
rect 8102 5956 8106 6012
rect 8042 5952 8106 5956
rect 8122 6012 8186 6016
rect 8122 5956 8126 6012
rect 8126 5956 8182 6012
rect 8182 5956 8186 6012
rect 8122 5952 8186 5956
rect 14813 6012 14877 6016
rect 14813 5956 14817 6012
rect 14817 5956 14873 6012
rect 14873 5956 14877 6012
rect 14813 5952 14877 5956
rect 14893 6012 14957 6016
rect 14893 5956 14897 6012
rect 14897 5956 14953 6012
rect 14953 5956 14957 6012
rect 14893 5952 14957 5956
rect 14973 6012 15037 6016
rect 14973 5956 14977 6012
rect 14977 5956 15033 6012
rect 15033 5956 15037 6012
rect 14973 5952 15037 5956
rect 15053 6012 15117 6016
rect 15053 5956 15057 6012
rect 15057 5956 15113 6012
rect 15113 5956 15117 6012
rect 15053 5952 15117 5956
rect 4417 5468 4481 5472
rect 4417 5412 4421 5468
rect 4421 5412 4477 5468
rect 4477 5412 4481 5468
rect 4417 5408 4481 5412
rect 4497 5468 4561 5472
rect 4497 5412 4501 5468
rect 4501 5412 4557 5468
rect 4557 5412 4561 5468
rect 4497 5408 4561 5412
rect 4577 5468 4641 5472
rect 4577 5412 4581 5468
rect 4581 5412 4637 5468
rect 4637 5412 4641 5468
rect 4577 5408 4641 5412
rect 4657 5468 4721 5472
rect 4657 5412 4661 5468
rect 4661 5412 4717 5468
rect 4717 5412 4721 5468
rect 4657 5408 4721 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 18278 5468 18342 5472
rect 18278 5412 18282 5468
rect 18282 5412 18338 5468
rect 18338 5412 18342 5468
rect 18278 5408 18342 5412
rect 18358 5468 18422 5472
rect 18358 5412 18362 5468
rect 18362 5412 18418 5468
rect 18418 5412 18422 5468
rect 18358 5408 18422 5412
rect 18438 5468 18502 5472
rect 18438 5412 18442 5468
rect 18442 5412 18498 5468
rect 18498 5412 18502 5468
rect 18438 5408 18502 5412
rect 18518 5468 18582 5472
rect 18518 5412 18522 5468
rect 18522 5412 18578 5468
rect 18578 5412 18582 5468
rect 18518 5408 18582 5412
rect 7882 4924 7946 4928
rect 7882 4868 7886 4924
rect 7886 4868 7942 4924
rect 7942 4868 7946 4924
rect 7882 4864 7946 4868
rect 7962 4924 8026 4928
rect 7962 4868 7966 4924
rect 7966 4868 8022 4924
rect 8022 4868 8026 4924
rect 7962 4864 8026 4868
rect 8042 4924 8106 4928
rect 8042 4868 8046 4924
rect 8046 4868 8102 4924
rect 8102 4868 8106 4924
rect 8042 4864 8106 4868
rect 8122 4924 8186 4928
rect 8122 4868 8126 4924
rect 8126 4868 8182 4924
rect 8182 4868 8186 4924
rect 8122 4864 8186 4868
rect 14813 4924 14877 4928
rect 14813 4868 14817 4924
rect 14817 4868 14873 4924
rect 14873 4868 14877 4924
rect 14813 4864 14877 4868
rect 14893 4924 14957 4928
rect 14893 4868 14897 4924
rect 14897 4868 14953 4924
rect 14953 4868 14957 4924
rect 14893 4864 14957 4868
rect 14973 4924 15037 4928
rect 14973 4868 14977 4924
rect 14977 4868 15033 4924
rect 15033 4868 15037 4924
rect 14973 4864 15037 4868
rect 15053 4924 15117 4928
rect 15053 4868 15057 4924
rect 15057 4868 15113 4924
rect 15113 4868 15117 4924
rect 15053 4864 15117 4868
rect 4417 4380 4481 4384
rect 4417 4324 4421 4380
rect 4421 4324 4477 4380
rect 4477 4324 4481 4380
rect 4417 4320 4481 4324
rect 4497 4380 4561 4384
rect 4497 4324 4501 4380
rect 4501 4324 4557 4380
rect 4557 4324 4561 4380
rect 4497 4320 4561 4324
rect 4577 4380 4641 4384
rect 4577 4324 4581 4380
rect 4581 4324 4637 4380
rect 4637 4324 4641 4380
rect 4577 4320 4641 4324
rect 4657 4380 4721 4384
rect 4657 4324 4661 4380
rect 4661 4324 4717 4380
rect 4717 4324 4721 4380
rect 4657 4320 4721 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 18278 4380 18342 4384
rect 18278 4324 18282 4380
rect 18282 4324 18338 4380
rect 18338 4324 18342 4380
rect 18278 4320 18342 4324
rect 18358 4380 18422 4384
rect 18358 4324 18362 4380
rect 18362 4324 18418 4380
rect 18418 4324 18422 4380
rect 18358 4320 18422 4324
rect 18438 4380 18502 4384
rect 18438 4324 18442 4380
rect 18442 4324 18498 4380
rect 18498 4324 18502 4380
rect 18438 4320 18502 4324
rect 18518 4380 18582 4384
rect 18518 4324 18522 4380
rect 18522 4324 18578 4380
rect 18578 4324 18582 4380
rect 18518 4320 18582 4324
rect 7882 3836 7946 3840
rect 7882 3780 7886 3836
rect 7886 3780 7942 3836
rect 7942 3780 7946 3836
rect 7882 3776 7946 3780
rect 7962 3836 8026 3840
rect 7962 3780 7966 3836
rect 7966 3780 8022 3836
rect 8022 3780 8026 3836
rect 7962 3776 8026 3780
rect 8042 3836 8106 3840
rect 8042 3780 8046 3836
rect 8046 3780 8102 3836
rect 8102 3780 8106 3836
rect 8042 3776 8106 3780
rect 8122 3836 8186 3840
rect 8122 3780 8126 3836
rect 8126 3780 8182 3836
rect 8182 3780 8186 3836
rect 8122 3776 8186 3780
rect 14813 3836 14877 3840
rect 14813 3780 14817 3836
rect 14817 3780 14873 3836
rect 14873 3780 14877 3836
rect 14813 3776 14877 3780
rect 14893 3836 14957 3840
rect 14893 3780 14897 3836
rect 14897 3780 14953 3836
rect 14953 3780 14957 3836
rect 14893 3776 14957 3780
rect 14973 3836 15037 3840
rect 14973 3780 14977 3836
rect 14977 3780 15033 3836
rect 15033 3780 15037 3836
rect 14973 3776 15037 3780
rect 15053 3836 15117 3840
rect 15053 3780 15057 3836
rect 15057 3780 15113 3836
rect 15113 3780 15117 3836
rect 15053 3776 15117 3780
rect 4417 3292 4481 3296
rect 4417 3236 4421 3292
rect 4421 3236 4477 3292
rect 4477 3236 4481 3292
rect 4417 3232 4481 3236
rect 4497 3292 4561 3296
rect 4497 3236 4501 3292
rect 4501 3236 4557 3292
rect 4557 3236 4561 3292
rect 4497 3232 4561 3236
rect 4577 3292 4641 3296
rect 4577 3236 4581 3292
rect 4581 3236 4637 3292
rect 4637 3236 4641 3292
rect 4577 3232 4641 3236
rect 4657 3292 4721 3296
rect 4657 3236 4661 3292
rect 4661 3236 4717 3292
rect 4717 3236 4721 3292
rect 4657 3232 4721 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 18278 3292 18342 3296
rect 18278 3236 18282 3292
rect 18282 3236 18338 3292
rect 18338 3236 18342 3292
rect 18278 3232 18342 3236
rect 18358 3292 18422 3296
rect 18358 3236 18362 3292
rect 18362 3236 18418 3292
rect 18418 3236 18422 3292
rect 18358 3232 18422 3236
rect 18438 3292 18502 3296
rect 18438 3236 18442 3292
rect 18442 3236 18498 3292
rect 18498 3236 18502 3292
rect 18438 3232 18502 3236
rect 18518 3292 18582 3296
rect 18518 3236 18522 3292
rect 18522 3236 18578 3292
rect 18578 3236 18582 3292
rect 18518 3232 18582 3236
rect 7882 2748 7946 2752
rect 7882 2692 7886 2748
rect 7886 2692 7942 2748
rect 7942 2692 7946 2748
rect 7882 2688 7946 2692
rect 7962 2748 8026 2752
rect 7962 2692 7966 2748
rect 7966 2692 8022 2748
rect 8022 2692 8026 2748
rect 7962 2688 8026 2692
rect 8042 2748 8106 2752
rect 8042 2692 8046 2748
rect 8046 2692 8102 2748
rect 8102 2692 8106 2748
rect 8042 2688 8106 2692
rect 8122 2748 8186 2752
rect 8122 2692 8126 2748
rect 8126 2692 8182 2748
rect 8182 2692 8186 2748
rect 8122 2688 8186 2692
rect 14813 2748 14877 2752
rect 14813 2692 14817 2748
rect 14817 2692 14873 2748
rect 14873 2692 14877 2748
rect 14813 2688 14877 2692
rect 14893 2748 14957 2752
rect 14893 2692 14897 2748
rect 14897 2692 14953 2748
rect 14953 2692 14957 2748
rect 14893 2688 14957 2692
rect 14973 2748 15037 2752
rect 14973 2692 14977 2748
rect 14977 2692 15033 2748
rect 15033 2692 15037 2748
rect 14973 2688 15037 2692
rect 15053 2748 15117 2752
rect 15053 2692 15057 2748
rect 15057 2692 15113 2748
rect 15113 2692 15117 2748
rect 15053 2688 15117 2692
rect 4417 2204 4481 2208
rect 4417 2148 4421 2204
rect 4421 2148 4477 2204
rect 4477 2148 4481 2204
rect 4417 2144 4481 2148
rect 4497 2204 4561 2208
rect 4497 2148 4501 2204
rect 4501 2148 4557 2204
rect 4557 2148 4561 2204
rect 4497 2144 4561 2148
rect 4577 2204 4641 2208
rect 4577 2148 4581 2204
rect 4581 2148 4637 2204
rect 4637 2148 4641 2204
rect 4577 2144 4641 2148
rect 4657 2204 4721 2208
rect 4657 2148 4661 2204
rect 4661 2148 4717 2204
rect 4717 2148 4721 2204
rect 4657 2144 4721 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 18278 2204 18342 2208
rect 18278 2148 18282 2204
rect 18282 2148 18338 2204
rect 18338 2148 18342 2204
rect 18278 2144 18342 2148
rect 18358 2204 18422 2208
rect 18358 2148 18362 2204
rect 18362 2148 18418 2204
rect 18418 2148 18422 2204
rect 18358 2144 18422 2148
rect 18438 2204 18502 2208
rect 18438 2148 18442 2204
rect 18442 2148 18498 2204
rect 18498 2148 18502 2204
rect 18438 2144 18502 2148
rect 18518 2204 18582 2208
rect 18518 2148 18522 2204
rect 18522 2148 18578 2204
rect 18578 2148 18582 2204
rect 18518 2144 18582 2148
<< metal4 >>
rect 4409 20704 4729 20720
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 19616 4729 20640
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 18528 4729 19552
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 17440 4729 18464
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 16352 4729 17376
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 15264 4729 16288
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 14176 4729 15200
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 13088 4729 14112
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 12000 4729 13024
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 10912 4729 11936
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 9824 4729 10848
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 8736 4729 9760
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 7648 4729 8672
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 6560 4729 7584
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 5472 4729 6496
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 4384 4729 5408
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 3296 4729 4320
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 2208 4729 3232
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2128 4729 2144
rect 7874 20160 8195 20720
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8195 20160
rect 7874 19072 8195 20096
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8195 19072
rect 7874 17984 8195 19008
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8195 17984
rect 7874 16896 8195 17920
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8195 16896
rect 7874 15808 8195 16832
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8195 15808
rect 7874 14720 8195 15744
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8195 14720
rect 7874 13632 8195 14656
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8195 13632
rect 7874 12544 8195 13568
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8195 12544
rect 7874 11456 8195 12480
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8195 11456
rect 7874 10368 8195 11392
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8195 10368
rect 7874 9280 8195 10304
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8195 9280
rect 7874 8192 8195 9216
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8195 8192
rect 7874 7104 8195 8128
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8195 7104
rect 7874 6016 8195 7040
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8195 6016
rect 7874 4928 8195 5952
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8195 4928
rect 7874 3840 8195 4864
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8195 3840
rect 7874 2752 8195 3776
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8195 2752
rect 7874 2128 8195 2688
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 14805 20160 15125 20720
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 19072 15125 20096
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 17984 15125 19008
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 14805 16896 15125 17920
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 15808 15125 16832
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 14720 15125 15744
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 13632 15125 14656
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 12544 15125 13568
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 11456 15125 12480
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 10368 15125 11392
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14805 9280 15125 10304
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 8192 15125 9216
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 7104 15125 8128
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 6016 15125 7040
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 4928 15125 5952
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 3840 15125 4864
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 14805 2752 15125 3776
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2128 15125 2688
rect 18270 20704 18591 20720
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18591 20704
rect 18270 19616 18591 20640
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18591 19616
rect 18270 18528 18591 19552
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18591 18528
rect 18270 17440 18591 18464
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18591 17440
rect 18270 16352 18591 17376
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18591 16352
rect 18270 15264 18591 16288
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18591 15264
rect 18270 14176 18591 15200
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18591 14176
rect 18270 13088 18591 14112
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18591 13088
rect 18270 12000 18591 13024
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18591 12000
rect 18270 10912 18591 11936
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18591 10912
rect 18270 9824 18591 10848
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18591 9824
rect 18270 8736 18591 9760
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18591 8736
rect 18270 7648 18591 8672
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18591 7648
rect 18270 6560 18591 7584
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18591 6560
rect 18270 5472 18591 6496
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18591 5472
rect 18270 4384 18591 5408
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18591 4384
rect 18270 3296 18591 4320
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18591 3296
rect 18270 2208 18591 3232
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18591 2208
rect 18270 2128 18591 2144
use sky130_fd_sc_hd__fill_2  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3
timestamp 1624635492
transform 1 0 1380 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1624635492
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_9
timestamp 1624635492
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9
timestamp 1624635492
transform 1 0 1932 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input43 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 1932 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1624635492
transform 1 0 1564 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1624635492
transform 1 0 2116 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1624635492
transform 1 0 2116 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_15
timestamp 1624635492
transform 1 0 2484 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15
timestamp 1624635492
transform 1 0 2484 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1624635492
transform 1 0 2668 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1624635492
transform 1 0 2668 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 3404 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1624635492
transform -1 0 3404 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21
timestamp 1624635492
transform 1 0 3036 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3404 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_21
timestamp 1624635492
transform 1 0 3036 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_25
timestamp 1624635492
transform 1 0 3404 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1624635492
transform -1 0 3772 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1624635492
transform -1 0 4048 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_29
timestamp 1624635492
transform 1 0 3772 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1624635492
transform -1 0 4140 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_33 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 4140 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1624635492
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1624635492
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1624635492
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1624635492
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56
timestamp 1624635492
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_59
timestamp 1624635492
transform 1 0 6532 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_45
timestamp 1624635492
transform 1 0 5244 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_58
timestamp 1624635492
transform 1 0 6440 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_71
timestamp 1624635492
transform 1 0 7636 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83
timestamp 1624635492
transform 1 0 8740 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_70
timestamp 1624635492
transform 1 0 7544 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_82
timestamp 1624635492
transform 1 0 8648 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1624635492
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_88
timestamp 1624635492
transform 1 0 9200 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_100
timestamp 1624635492
transform 1 0 10304 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_94
timestamp 1624635492
transform 1 0 9752 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1624635492
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1624635492
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output60
timestamp 1624635492
transform -1 0 12420 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output60_A
timestamp 1624635492
transform -1 0 12788 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_112
timestamp 1624635492
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_117
timestamp 1624635492
transform 1 0 11868 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_123
timestamp 1624635492
transform 1 0 12420 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_106 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 10856 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_115
timestamp 1624635492
transform 1 0 11684 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1624635492
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_127
timestamp 1624635492
transform 1 0 12788 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_139 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 13892 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_127
timestamp 1624635492
transform 1 0 12788 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_139
timestamp 1624635492
transform 1 0 13892 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_146
timestamp 1624635492
transform 1 0 14536 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_158
timestamp 1624635492
transform 1 0 15640 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_151
timestamp 1624635492
transform 1 0 14996 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_163
timestamp 1624635492
transform 1 0 16100 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1624635492
transform 1 0 17112 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1624635492
transform 1 0 16836 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_170
timestamp 1624635492
transform 1 0 16744 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_175
timestamp 1624635492
transform 1 0 17204 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1624635492
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_172
timestamp 1624635492
transform 1 0 16928 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1624635492
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1624635492
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_199
timestamp 1624635492
transform 1 0 19412 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_204
timestamp 1624635492
transform 1 0 19872 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1624635492
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_208
timestamp 1624635492
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1624635492
transform -1 0 21896 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1624635492
transform -1 0 21896 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_216
timestamp 1624635492
transform 1 0 20976 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_222 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 21528 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_220
timestamp 1624635492
transform 1 0 21344 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1624635492
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1624635492
transform 1 0 1564 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1624635492
transform 1 0 2116 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1624635492
transform -1 0 2852 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1624635492
transform 1 0 1380 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_9
timestamp 1624635492
transform 1 0 1932 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_15
timestamp 1624635492
transform 1 0 2484 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_19
timestamp 1624635492
transform 1 0 2852 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1624635492
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1624635492
transform -1 0 3220 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_23
timestamp 1624635492
transform 1 0 3220 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_30
timestamp 1624635492
transform 1 0 3864 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_42
timestamp 1624635492
transform 1 0 4968 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_54
timestamp 1624635492
transform 1 0 6072 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_66
timestamp 1624635492
transform 1 0 7176 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_78
timestamp 1624635492
transform 1 0 8280 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1624635492
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_87
timestamp 1624635492
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_99
timestamp 1624635492
transform 1 0 10212 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_111
timestamp 1624635492
transform 1 0 11316 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_123
timestamp 1624635492
transform 1 0 12420 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1624635492
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_135
timestamp 1624635492
transform 1 0 13524 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_144
timestamp 1624635492
transform 1 0 14352 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_156
timestamp 1624635492
transform 1 0 15456 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_168
timestamp 1624635492
transform 1 0 16560 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_180
timestamp 1624635492
transform 1 0 17664 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1624635492
transform 1 0 19504 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_192
timestamp 1624635492
transform 1 0 18768 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_201
timestamp 1624635492
transform 1 0 19596 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1624635492
transform -1 0 21896 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_213
timestamp 1624635492
transform 1 0 20700 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_221
timestamp 1624635492
transform 1 0 21436 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1624635492
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1624635492
transform 1 0 1564 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1624635492
transform -1 0 2300 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1624635492
transform -1 0 2668 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1624635492
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_9
timestamp 1624635492
transform 1 0 1932 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_13
timestamp 1624635492
transform 1 0 2300 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_17
timestamp 1624635492
transform 1 0 2668 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_29
timestamp 1624635492
transform 1 0 3772 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_41
timestamp 1624635492
transform 1 0 4876 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1624635492
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_53
timestamp 1624635492
transform 1 0 5980 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_58
timestamp 1624635492
transform 1 0 6440 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_70
timestamp 1624635492
transform 1 0 7544 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_82
timestamp 1624635492
transform 1 0 8648 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_94
timestamp 1624635492
transform 1 0 9752 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1624635492
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_106
timestamp 1624635492
transform 1 0 10856 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_115
timestamp 1624635492
transform 1 0 11684 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_127
timestamp 1624635492
transform 1 0 12788 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_139
timestamp 1624635492
transform 1 0 13892 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_151
timestamp 1624635492
transform 1 0 14996 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_163
timestamp 1624635492
transform 1 0 16100 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1624635492
transform 1 0 16836 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_172
timestamp 1624635492
transform 1 0 16928 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1624635492
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1624635492
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1624635492
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1624635492
transform -1 0 21896 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_220
timestamp 1624635492
transform 1 0 21344 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1624635492
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1624635492
transform 1 0 1840 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1624635492
transform -1 0 2484 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_6
timestamp 1624635492
transform 1 0 1656 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_11
timestamp 1624635492
transform 1 0 2116 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1624635492
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1624635492
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_27
timestamp 1624635492
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_30
timestamp 1624635492
transform 1 0 3864 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_42
timestamp 1624635492
transform 1 0 4968 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_54
timestamp 1624635492
transform 1 0 6072 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_66
timestamp 1624635492
transform 1 0 7176 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_78
timestamp 1624635492
transform 1 0 8280 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1624635492
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_87
timestamp 1624635492
transform 1 0 9108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_99
timestamp 1624635492
transform 1 0 10212 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_111
timestamp 1624635492
transform 1 0 11316 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_123
timestamp 1624635492
transform 1 0 12420 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1624635492
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_135
timestamp 1624635492
transform 1 0 13524 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_144
timestamp 1624635492
transform 1 0 14352 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_156
timestamp 1624635492
transform 1 0 15456 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_168
timestamp 1624635492
transform 1 0 16560 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_180
timestamp 1624635492
transform 1 0 17664 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1624635492
transform 1 0 19504 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_192
timestamp 1624635492
transform 1 0 18768 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_201
timestamp 1624635492
transform 1 0 19596 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1624635492
transform -1 0 21896 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_213
timestamp 1624635492
transform 1 0 20700 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_221
timestamp 1624635492
transform 1 0 21436 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1624635492
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1624635492
transform 1 0 1380 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1624635492
transform -1 0 2024 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1624635492
transform -1 0 2392 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_6
timestamp 1624635492
transform 1 0 1656 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_10
timestamp 1624635492
transform 1 0 2024 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_14
timestamp 1624635492
transform 1 0 2392 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_26
timestamp 1624635492
transform 1 0 3496 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_38
timestamp 1624635492
transform 1 0 4600 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1624635492
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_50
timestamp 1624635492
transform 1 0 5704 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_56
timestamp 1624635492
transform 1 0 6256 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_58
timestamp 1624635492
transform 1 0 6440 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_70
timestamp 1624635492
transform 1 0 7544 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_82
timestamp 1624635492
transform 1 0 8648 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_94
timestamp 1624635492
transform 1 0 9752 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1624635492
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_106
timestamp 1624635492
transform 1 0 10856 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_115
timestamp 1624635492
transform 1 0 11684 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_127
timestamp 1624635492
transform 1 0 12788 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_139
timestamp 1624635492
transform 1 0 13892 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_151
timestamp 1624635492
transform 1 0 14996 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_163
timestamp 1624635492
transform 1 0 16100 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1624635492
transform 1 0 16836 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_172
timestamp 1624635492
transform 1 0 16928 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1624635492
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1624635492
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_208
timestamp 1624635492
transform 1 0 20240 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _107_
timestamp 1624635492
transform -1 0 21068 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1624635492
transform -1 0 21896 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1624635492
transform -1 0 21436 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_217
timestamp 1624635492
transform 1 0 21068 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_221
timestamp 1624635492
transform 1 0 21436 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_6
timestamp 1624635492
transform 1 0 1656 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_6
timestamp 1624635492
transform 1 0 1656 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1624635492
transform -1 0 2024 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1624635492
transform -1 0 2024 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1624635492
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1624635492
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1624635492
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1624635492
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_10
timestamp 1624635492
transform 1 0 2024 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_10
timestamp 1624635492
transform 1 0 2024 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1624635492
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_22
timestamp 1624635492
transform 1 0 3128 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_28
timestamp 1624635492
transform 1 0 3680 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_30
timestamp 1624635492
transform 1 0 3864 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_22
timestamp 1624635492
transform 1 0 3128 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_34
timestamp 1624635492
transform 1 0 4232 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1624635492
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_42
timestamp 1624635492
transform 1 0 4968 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_54
timestamp 1624635492
transform 1 0 6072 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_46
timestamp 1624635492
transform 1 0 5336 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_54
timestamp 1624635492
transform 1 0 6072 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_58
timestamp 1624635492
transform 1 0 6440 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_66
timestamp 1624635492
transform 1 0 7176 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_78
timestamp 1624635492
transform 1 0 8280 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_70
timestamp 1624635492
transform 1 0 7544 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_82
timestamp 1624635492
transform 1 0 8648 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1624635492
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_87
timestamp 1624635492
transform 1 0 9108 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_99
timestamp 1624635492
transform 1 0 10212 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_94
timestamp 1624635492
transform 1 0 9752 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1624635492
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_111
timestamp 1624635492
transform 1 0 11316 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_123
timestamp 1624635492
transform 1 0 12420 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_106
timestamp 1624635492
transform 1 0 10856 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_115
timestamp 1624635492
transform 1 0 11684 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1624635492
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_135
timestamp 1624635492
transform 1 0 13524 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_144
timestamp 1624635492
transform 1 0 14352 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_127
timestamp 1624635492
transform 1 0 12788 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_139
timestamp 1624635492
transform 1 0 13892 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_156
timestamp 1624635492
transform 1 0 15456 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_151
timestamp 1624635492
transform 1 0 14996 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_163
timestamp 1624635492
transform 1 0 16100 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1624635492
transform 1 0 16836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_168
timestamp 1624635492
transform 1 0 16560 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_180
timestamp 1624635492
transform 1 0 17664 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_172
timestamp 1624635492
transform 1 0 16928 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1624635492
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _105_
timestamp 1624635492
transform 1 0 20056 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1624635492
transform 1 0 19504 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_192
timestamp 1624635492
transform 1 0 18768 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_201
timestamp 1624635492
transform 1 0 19596 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_196
timestamp 1624635492
transform 1 0 19136 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_204
timestamp 1624635492
transform 1 0 19872 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_213
timestamp 1624635492
transform 1 0 20700 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_209
timestamp 1624635492
transform 1 0 20332 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_214
timestamp 1624635492
transform 1 0 20792 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_209
timestamp 1624635492
transform 1 0 20332 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1624635492
transform -1 0 20700 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1624635492
transform -1 0 21160 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _106_
timestamp 1624635492
transform -1 0 20792 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_221
timestamp 1624635492
transform 1 0 21436 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_222
timestamp 1624635492
transform 1 0 21528 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_218
timestamp 1624635492
transform 1 0 21160 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1624635492
transform -1 0 21896 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1624635492
transform -1 0 21896 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1624635492
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1624635492
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1624635492
transform -1 0 2024 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_6
timestamp 1624635492
transform 1 0 1656 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_10
timestamp 1624635492
transform 1 0 2024 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 4324 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1624635492
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 3956 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_22
timestamp 1624635492
transform 1 0 3128 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_28
timestamp 1624635492
transform 1 0 3680 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_30
timestamp 1624635492
transform 1 0 3864 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_33
timestamp 1624635492
transform 1 0 4140 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1624635492
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_56
timestamp 1624635492
transform 1 0 6256 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _039_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 8280 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1624635492
transform 1 0 7268 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_8_64
timestamp 1624635492
transform 1 0 6992 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_76
timestamp 1624635492
transform 1 0 8096 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_81
timestamp 1624635492
transform 1 0 8556 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1624635492
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_85
timestamp 1624635492
transform 1 0 8924 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_87
timestamp 1624635492
transform 1 0 9108 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_99
timestamp 1624635492
transform 1 0 10212 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_111
timestamp 1624635492
transform 1 0 11316 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_123
timestamp 1624635492
transform 1 0 12420 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1624635492
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_135
timestamp 1624635492
transform 1 0 13524 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_144
timestamp 1624635492
transform 1 0 14352 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_156
timestamp 1624635492
transform 1 0 15456 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_168
timestamp 1624635492
transform 1 0 16560 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_180
timestamp 1624635492
transform 1 0 17664 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _104_
timestamp 1624635492
transform 1 0 19780 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1624635492
transform 1 0 19504 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1624635492
transform -1 0 20424 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_192
timestamp 1624635492
transform 1 0 18768 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_201
timestamp 1624635492
transform 1 0 19596 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_206
timestamp 1624635492
transform 1 0 20056 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1624635492
transform -1 0 21896 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_210
timestamp 1624635492
transform 1 0 20424 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_222
timestamp 1624635492
transform 1 0 21528 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1624635492
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1624635492
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1624635492
transform 1 0 1840 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1624635492
transform -1 0 2484 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1624635492
transform -1 0 2852 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_6
timestamp 1624635492
transform 1 0 1656 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_11
timestamp 1624635492
transform 1 0 2116 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_15
timestamp 1624635492
transform 1 0 2484 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_19
timestamp 1624635492
transform 1 0 2852 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1624635492
transform 1 0 4600 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1624635492
transform 1 0 3588 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 3220 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_25
timestamp 1624635492
transform 1 0 3404 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_36
timestamp 1624635492
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _067_
timestamp 1624635492
transform 1 0 5612 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1624635492
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 6716 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_47
timestamp 1624635492
transform 1 0 5428 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1624635492
transform 1 0 5888 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_56
timestamp 1624635492
transform 1 0 6256 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_58
timestamp 1624635492
transform 1 0 6440 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1624635492
transform -1 0 8924 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1624635492
transform -1 0 7912 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_63
timestamp 1624635492
transform 1 0 6900 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_74
timestamp 1624635492
transform 1 0 7912 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 9108 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 9476 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_85
timestamp 1624635492
transform 1 0 8924 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_89
timestamp 1624635492
transform 1 0 9292 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1624635492
transform 1 0 9660 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1624635492
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_105
timestamp 1624635492
transform 1 0 10764 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_113
timestamp 1624635492
transform 1 0 11500 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_115
timestamp 1624635492
transform 1 0 11684 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_127
timestamp 1624635492
transform 1 0 12788 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_139
timestamp 1624635492
transform 1 0 13892 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_151
timestamp 1624635492
transform 1 0 14996 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_163
timestamp 1624635492
transform 1 0 16100 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1624635492
transform 1 0 16836 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_172
timestamp 1624635492
transform 1 0 16928 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_184
timestamp 1624635492
transform 1 0 18032 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _102_
timestamp 1624635492
transform -1 0 18860 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _103_
timestamp 1624635492
transform 1 0 19044 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_193
timestamp 1624635492
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_198
timestamp 1624635492
transform 1 0 19320 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1624635492
transform -1 0 21896 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_210
timestamp 1624635492
transform 1 0 20424 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_222
timestamp 1624635492
transform 1 0 21528 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1624635492
transform 1 0 2760 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 2024 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1624635492
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1624635492
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_6
timestamp 1624635492
transform 1 0 1656 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_13
timestamp 1624635492
transform 1 0 2300 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_17
timestamp 1624635492
transform 1 0 2668 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 5520 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1624635492
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_27
timestamp 1624635492
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_30
timestamp 1624635492
transform 1 0 3864 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 5704 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_48
timestamp 1624635492
transform 1 0 5520 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 8832 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_66
timestamp 1624635492
transform 1 0 7176 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1624635492
transform 1 0 9292 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1624635492
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_84
timestamp 1624635492
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_87
timestamp 1624635492
transform 1 0 9108 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_98
timestamp 1624635492
transform 1 0 10120 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_110
timestamp 1624635492
transform 1 0 11224 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_122
timestamp 1624635492
transform 1 0 12328 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1624635492
transform 1 0 14260 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_134
timestamp 1624635492
transform 1 0 13432 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_142
timestamp 1624635492
transform 1 0 14168 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_144
timestamp 1624635492
transform 1 0 14352 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_156
timestamp 1624635492
transform 1 0 15456 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_168
timestamp 1624635492
transform 1 0 16560 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_180
timestamp 1624635492
transform 1 0 17664 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1624635492
transform 1 0 19504 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_192
timestamp 1624635492
transform 1 0 18768 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_201
timestamp 1624635492
transform 1 0 19596 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1624635492
transform -1 0 21896 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_213
timestamp 1624635492
transform 1 0 20700 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_221
timestamp 1624635492
transform 1 0 21436 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _069_
timestamp 1624635492
transform 1 0 1748 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 2300 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1624635492
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1624635492
transform -1 0 1564 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_5
timestamp 1624635492
transform 1 0 1564 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_10
timestamp 1624635492
transform 1 0 2024 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 4048 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_11_29
timestamp 1624635492
transform 1 0 3772 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 6624 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1624635492
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_48
timestamp 1624635492
transform 1 0 5520 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_56
timestamp 1624635492
transform 1 0 6256 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_58
timestamp 1624635492
transform 1 0 6440 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1624635492
transform -1 0 9108 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_76
timestamp 1624635492
transform 1 0 8096 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_87
timestamp 1624635492
transform 1 0 9108 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_99
timestamp 1624635492
transform 1 0 10212 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1624635492
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_111
timestamp 1624635492
transform 1 0 11316 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_115
timestamp 1624635492
transform 1 0 11684 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_127
timestamp 1624635492
transform 1 0 12788 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_139
timestamp 1624635492
transform 1 0 13892 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_151
timestamp 1624635492
transform 1 0 14996 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_163
timestamp 1624635492
transform 1 0 16100 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1624635492
transform 1 0 16836 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_172
timestamp 1624635492
transform 1 0 16928 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1624635492
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1624635492
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1624635492
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1624635492
transform -1 0 21896 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_220
timestamp 1624635492
transform 1 0 21344 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _070_
timestamp 1624635492
transform -1 0 2024 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 2208 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1624635492
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 1624635492
transform 1 0 2668 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1624635492
transform -1 0 1564 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_5
timestamp 1624635492
transform 1 0 1564 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_10
timestamp 1624635492
transform 1 0 2024 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_15
timestamp 1624635492
transform 1 0 2484 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_20
timestamp 1624635492
transform 1 0 2944 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1624635492
transform 1 0 4876 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1624635492
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1624635492
transform -1 0 3312 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1624635492
transform -1 0 4048 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1624635492
transform 1 0 3312 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_28
timestamp 1624635492
transform 1 0 3680 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_32
timestamp 1624635492
transform 1 0 4048 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_40
timestamp 1624635492
transform 1 0 4784 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_50
timestamp 1624635492
transform 1 0 5704 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_62
timestamp 1624635492
transform 1 0 6808 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1624635492
transform 1 0 7084 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_12_74
timestamp 1624635492
transform 1 0 7912 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1624635492
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 9752 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_87
timestamp 1624635492
transform 1 0 9108 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_92
timestamp 1624635492
transform 1 0 9568 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_96
timestamp 1624635492
transform 1 0 9936 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_108
timestamp 1624635492
transform 1 0 11040 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_120
timestamp 1624635492
transform 1 0 12144 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1624635492
transform 1 0 14260 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_132
timestamp 1624635492
transform 1 0 13248 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_140
timestamp 1624635492
transform 1 0 13984 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_144
timestamp 1624635492
transform 1 0 14352 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_156
timestamp 1624635492
transform 1 0 15456 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_168
timestamp 1624635492
transform 1 0 16560 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_180
timestamp 1624635492
transform 1 0 17664 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1624635492
transform 1 0 19504 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_192
timestamp 1624635492
transform 1 0 18768 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_201
timestamp 1624635492
transform 1 0 19596 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1624635492
transform -1 0 21896 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_213
timestamp 1624635492
transform 1 0 20700 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_221
timestamp 1624635492
transform 1 0 21436 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_6
timestamp 1624635492
transform 1 0 1656 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_6
timestamp 1624635492
transform 1 0 1656 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1624635492
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1624635492
transform 1 0 1840 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1624635492
transform 1 0 1380 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1624635492
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1624635492
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_18
timestamp 1624635492
transform 1 0 2760 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_11
timestamp 1624635492
transform 1 0 2116 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1624635492
transform 1 0 2944 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1624635492
transform -1 0 2760 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 3312 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_14_30
timestamp 1624635492
transform 1 0 3864 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_28
timestamp 1624635492
transform 1 0 3680 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_24
timestamp 1624635492
transform 1 0 3312 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_29
timestamp 1624635492
transform 1 0 3772 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 3956 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1624635492
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_41
timestamp 1624635492
transform 1 0 4876 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_37
timestamp 1624635492
transform 1 0 4508 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_33
timestamp 1624635492
transform 1 0 4140 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 4692 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 4324 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1624635492
transform -1 0 4876 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_13_41
timestamp 1624635492
transform 1 0 4876 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 5244 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1624635492
transform 1 0 6624 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1624635492
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_53
timestamp 1624635492
transform 1 0 5980 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_58
timestamp 1624635492
transform 1 0 6440 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_61
timestamp 1624635492
transform 1 0 6716 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1624635492
transform -1 0 7176 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 7912 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1624635492
transform 1 0 7728 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_13_69
timestamp 1624635492
transform 1 0 7452 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_73
timestamp 1624635492
transform 1 0 7820 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_66
timestamp 1624635492
transform 1 0 7176 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_81
timestamp 1624635492
transform 1 0 8556 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 10764 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1624635492
transform 1 0 9568 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1624635492
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_90
timestamp 1624635492
transform 1 0 9384 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_101
timestamp 1624635492
transform 1 0 10396 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_85
timestamp 1624635492
transform 1 0 8924 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_87
timestamp 1624635492
transform 1 0 9108 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_105
timestamp 1624635492
transform 1 0 10764 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_113
timestamp 1624635492
transform 1 0 11500 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_109
timestamp 1624635492
transform 1 0 11132 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 11132 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1624635492
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l1_in_0_
timestamp 1624635492
transform -1 0 11960 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_122
timestamp 1624635492
transform 1 0 12328 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_118
timestamp 1624635492
transform 1 0 11960 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1624635492
transform 1 0 12420 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_115
timestamp 1624635492
transform 1 0 11684 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1624635492
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_127
timestamp 1624635492
transform 1 0 12788 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_139
timestamp 1624635492
transform 1 0 13892 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_126
timestamp 1624635492
transform 1 0 12696 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_138
timestamp 1624635492
transform 1 0 13800 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_142
timestamp 1624635492
transform 1 0 14168 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_144
timestamp 1624635492
transform 1 0 14352 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 15180 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_151
timestamp 1624635492
transform 1 0 14996 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_163
timestamp 1624635492
transform 1 0 16100 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_152
timestamp 1624635492
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_155
timestamp 1624635492
transform 1 0 15364 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_26.mux_l2_in_0_
timestamp 1624635492
transform -1 0 17388 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1624635492
transform 1 0 16836 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_172
timestamp 1624635492
transform 1 0 16928 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1624635492
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_167
timestamp 1624635492
transform 1 0 16468 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_177
timestamp 1624635492
transform 1 0 17388 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1624635492
transform 1 0 19504 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1624635492
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1624635492
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_189
timestamp 1624635492
transform 1 0 18492 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_197
timestamp 1624635492
transform 1 0 19228 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_201
timestamp 1624635492
transform 1 0 19596 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1624635492
transform -1 0 21896 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1624635492
transform -1 0 21896 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_220
timestamp 1624635492
transform 1 0 21344 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_213
timestamp 1624635492
transform 1 0 20700 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_221
timestamp 1624635492
transform 1 0 21436 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 4232 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1624635492
transform -1 0 2576 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1624635492
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1624635492
transform -1 0 1564 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_5
timestamp 1624635492
transform 1 0 1564 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_16
timestamp 1624635492
transform 1 0 2576 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1624635492
transform 1 0 4416 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_34
timestamp 1624635492
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 6624 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1624635492
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 5428 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 5796 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_45
timestamp 1624635492
transform 1 0 5244 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_49
timestamp 1624635492
transform 1 0 5612 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_53
timestamp 1624635492
transform 1 0 5980 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_58
timestamp 1624635492
transform 1 0 6440 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1624635492
transform 1 0 8556 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_76
timestamp 1624635492
transform 1 0 8096 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_80
timestamp 1624635492
transform 1 0 8464 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_left_track_1.prog_clk
timestamp 1624635492
transform -1 0 9844 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_90
timestamp 1624635492
transform 1 0 9384 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_95
timestamp 1624635492
transform 1 0 9844 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 11868 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1624635492
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A0
timestamp 1624635492
transform -1 0 11408 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_107
timestamp 1624635492
transform 1 0 10948 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_112
timestamp 1624635492
transform 1 0 11408 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_115
timestamp 1624635492
transform 1 0 11684 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 13524 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_133
timestamp 1624635492
transform 1 0 13340 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1624635492
transform -1 0 16652 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_26.mux_l1_in_0_
timestamp 1624635492
transform -1 0 16192 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_151
timestamp 1624635492
transform 1 0 14996 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_164
timestamp 1624635492
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 18584 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1624635492
transform 1 0 16836 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1624635492
transform 1 0 16652 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_172
timestamp 1624635492
transform 1 0 16928 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_190
timestamp 1624635492
transform 1 0 18584 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_202
timestamp 1624635492
transform 1 0 19688 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1624635492
transform -1 0 21896 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_214
timestamp 1624635492
transform 1 0 20792 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_222
timestamp 1624635492
transform 1 0 21528 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1624635492
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 1840 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1624635492
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1624635492
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_6
timestamp 1624635492
transform 1 0 1656 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_11
timestamp 1624635492
transform 1 0 2116 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1624635492
transform -1 0 4876 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1624635492
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1624635492
transform -1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_23
timestamp 1624635492
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1624635492
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_30
timestamp 1624635492
transform 1 0 3864 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_41
timestamp 1624635492
transform 1 0 4876 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1624635492
transform 1 0 5060 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1624635492
transform 1 0 5796 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l2_in_0__S
timestamp 1624635492
transform 1 0 6808 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_46
timestamp 1624635492
transform 1 0 5336 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_50
timestamp 1624635492
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_60
timestamp 1624635492
transform 1 0 6624 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 8648 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_64
timestamp 1624635492
transform 1 0 6992 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_82
timestamp 1624635492
transform 1 0 8648 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1624635492
transform 1 0 9292 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 10212 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1624635492
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_87
timestamp 1624635492
transform 1 0 9108 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_92
timestamp 1624635492
transform 1 0 9568 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_98
timestamp 1624635492
transform 1 0 10120 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 12144 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_115
timestamp 1624635492
transform 1 0 11684 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_119
timestamp 1624635492
transform 1 0 12052 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1624635492
transform -1 0 14076 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1624635492
transform 1 0 14260 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_136
timestamp 1624635492
transform 1 0 13616 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1624635492
transform 1 0 14076 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_144
timestamp 1624635492
transform 1 0 14352 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 14536 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 16192 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_162
timestamp 1624635492
transform 1 0 16008 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_180
timestamp 1624635492
transform 1 0 17664 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1624635492
transform 1 0 19504 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_192
timestamp 1624635492
transform 1 0 18768 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_201
timestamp 1624635492
transform 1 0 19596 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1624635492
transform -1 0 21896 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_213
timestamp 1624635492
transform 1 0 20700 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_221
timestamp 1624635492
transform 1 0 21436 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp 1624635492
transform 1 0 1748 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 2208 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1624635492
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1624635492
transform 1 0 2668 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1624635492
transform -1 0 1564 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_5
timestamp 1624635492
transform 1 0 1564 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_10
timestamp 1624635492
transform 1 0 2024 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_15
timestamp 1624635492
transform 1 0 2484 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_20
timestamp 1624635492
transform 1 0 2944 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1624635492
transform 1 0 4324 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1624635492
transform 1 0 3312 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_33
timestamp 1624635492
transform 1 0 4140 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1624635492
transform 1 0 6624 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1624635492
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_left_track_1.prog_clk
timestamp 1624635492
transform 1 0 5888 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1624635492
transform -1 0 5520 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_44
timestamp 1624635492
transform 1 0 5152 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_48
timestamp 1624635492
transform 1 0 5520 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_55
timestamp 1624635492
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_58
timestamp 1624635492
transform 1 0 6440 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1624635492
transform 1 0 7912 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_69
timestamp 1624635492
transform 1 0 7452 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_73
timestamp 1624635492
transform 1 0 7820 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_83
timestamp 1624635492
transform 1 0 8740 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 9660 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_91
timestamp 1624635492
transform 1 0 9476 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_0_
timestamp 1624635492
transform -1 0 12880 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1624635492
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 11684 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_109
timestamp 1624635492
transform 1 0 11132 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_113
timestamp 1624635492
transform 1 0 11500 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_117
timestamp 1624635492
transform 1 0 11868 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_0_
timestamp 1624635492
transform -1 0 13892 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l2_in_0_
timestamp 1624635492
transform -1 0 14904 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_128
timestamp 1624635492
transform 1 0 12880 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_139
timestamp 1624635492
transform 1 0 13892 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1624635492
transform -1 0 16376 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_0_
timestamp 1624635492
transform -1 0 15916 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_150
timestamp 1624635492
transform 1 0 14904 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_161
timestamp 1624635492
transform 1 0 15916 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_166
timestamp 1624635492
transform 1 0 16376 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 19136 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1624635492
transform 1 0 16836 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 16928 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_170
timestamp 1624635492
transform 1 0 16744 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_174
timestamp 1624635492
transform 1 0 17112 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_196
timestamp 1624635492
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_208
timestamp 1624635492
transform 1 0 20240 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1624635492
transform -1 0 21896 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1624635492
transform 1 0 21160 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1624635492
transform -1 0 20976 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_216
timestamp 1624635492
transform 1 0 20976 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_221
timestamp 1624635492
transform 1 0 21436 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _068_
timestamp 1624635492
transform 1 0 1748 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 2484 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 2668 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1624635492
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 1564 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_5
timestamp 1624635492
transform 1 0 1564 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_10
timestamp 1624635492
transform 1 0 2024 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_15
timestamp 1624635492
transform 1 0 2484 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_20
timestamp 1624635492
transform 1 0 2944 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 4048 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1624635492
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1624635492
transform -1 0 3404 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_25
timestamp 1624635492
transform 1 0 3404 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_30
timestamp 1624635492
transform 1 0 3864 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 7360 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_48
timestamp 1624635492
transform 1 0 5520 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1624635492
transform 1 0 7544 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_left_track_1.prog_clk
timestamp 1624635492
transform 1 0 8556 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_68
timestamp 1624635492
transform 1 0 7360 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_79
timestamp 1624635492
transform 1 0 8372 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1624635492
transform -1 0 10580 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1624635492
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1624635492
transform -1 0 9292 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_84
timestamp 1624635492
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_89
timestamp 1624635492
transform 1 0 9292 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_93
timestamp 1624635492
transform 1 0 9660 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_103
timestamp 1624635492
transform 1 0 10580 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1624635492
transform 1 0 10764 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1624635492
transform -1 0 12420 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1624635492
transform 1 0 12604 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 11408 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_108
timestamp 1624635492
transform 1 0 11040 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_112
timestamp 1624635492
transform 1 0 11408 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_123
timestamp 1624635492
transform 1 0 12420 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1624635492
transform 1 0 14260 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_left_track_1.prog_clk
timestamp 1624635492
transform 1 0 13616 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_134
timestamp 1624635492
transform 1 0 13432 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_139
timestamp 1624635492
transform 1 0 13892 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_144
timestamp 1624635492
transform 1 0 14352 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 14536 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l2_in_0_
timestamp 1624635492
transform 1 0 16192 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_162
timestamp 1624635492
transform 1 0 16008 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 17296 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_18_173
timestamp 1624635492
transform 1 0 17020 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1624635492
transform 1 0 18952 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 21436 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1624635492
transform 1 0 19504 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_192
timestamp 1624635492
transform 1 0 18768 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_197
timestamp 1624635492
transform 1 0 19228 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_201
timestamp 1624635492
transform 1 0 19596 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1624635492
transform -1 0 21896 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_221
timestamp 1624635492
transform 1 0 21436 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1624635492
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1624635492
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1624635492
transform 1 0 1380 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1624635492
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp 1624635492
transform 1 0 1748 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1624635492
transform -1 0 1840 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_5
timestamp 1624635492
transform 1 0 1564 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 2300 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_10
timestamp 1624635492
transform 1 0 2024 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_8
timestamp 1624635492
transform 1 0 1840 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_18
timestamp 1624635492
transform 1 0 2760 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_13
timestamp 1624635492
transform 1 0 2300 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_19
timestamp 1624635492
transform 1 0 2852 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_15
timestamp 1624635492
transform 1 0 2484 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1624635492
transform -1 0 3220 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_39.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 2484 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1624635492
transform 1 0 2208 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 4416 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 6072 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l2_in_0_
timestamp 1624635492
transform 1 0 4324 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1624635492
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1624635492
transform -1 0 3588 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1624635492
transform -1 0 4048 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_36
timestamp 1624635492
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_23
timestamp 1624635492
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_27
timestamp 1624635492
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_32
timestamp 1624635492
transform 1 0 4048 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_44
timestamp 1624635492
transform 1 0 5152 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l1_in_0_
timestamp 1624635492
transform 1 0 5336 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_60
timestamp 1624635492
transform 1 0 6624 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_55
timestamp 1624635492
transform 1 0 6164 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_58
timestamp 1624635492
transform 1 0 6440 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_54
timestamp 1624635492
transform 1 0 6072 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1624635492
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1624635492
transform 1 0 6716 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1624635492
transform 1 0 6348 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_left_track_1.prog_clk
timestamp 1624635492
transform 1 0 6808 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1624635492
transform -1 0 7820 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 7728 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1624635492
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_70
timestamp 1624635492
transform 1 0 7544 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_65
timestamp 1624635492
transform 1 0 7084 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_69
timestamp 1624635492
transform 1 0 7452 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_73
timestamp 1624635492
transform 1 0 7820 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_87
timestamp 1624635492
transform 1 0 9108 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_84
timestamp 1624635492
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_93
timestamp 1624635492
transform 1 0 9660 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_88
timestamp 1624635492
transform 1 0 9200 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_left_track_1.prog_clk
timestamp 1624635492
transform 1 0 9384 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1624635492
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1624635492
transform 1 0 9292 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_102
timestamp 1624635492
transform 1 0 10488 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_98
timestamp 1624635492
transform 1 0 10120 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_101
timestamp 1624635492
transform 1 0 10396 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_97
timestamp 1624635492
transform 1 0 10028 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 10488 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 9844 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1624635492
transform -1 0 10488 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_104
timestamp 1624635492
transform 1 0 10672 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_112
timestamp 1624635492
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_108
timestamp 1624635492
transform 1 0 11040 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 10856 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1624635492
transform -1 0 11408 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1624635492
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_1_
timestamp 1624635492
transform 1 0 10856 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_115
timestamp 1624635492
transform 1 0 11684 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_115
timestamp 1624635492
transform 1 0 11684 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_1_
timestamp 1624635492
transform 1 0 11868 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 13340 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1624635492
transform 1 0 13524 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1624635492
transform 1 0 13156 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1624635492
transform 1 0 14260 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_133
timestamp 1624635492
transform 1 0 13340 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_144
timestamp 1624635492
transform 1 0 14352 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_126
timestamp 1624635492
transform 1 0 12696 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_130
timestamp 1624635492
transform 1 0 13064 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_140
timestamp 1624635492
transform 1 0 13984 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_144
timestamp 1624635492
transform 1 0 14352 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_154
timestamp 1624635492
transform 1 0 15272 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_149
timestamp 1624635492
transform 1 0 14812 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_149
timestamp 1624635492
transform 1 0 14812 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 15456 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_left_track_1.prog_clk
timestamp 1624635492
transform 1 0 14536 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1624635492
transform 1 0 14996 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1624635492
transform 1 0 14536 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_166
timestamp 1624635492
transform 1 0 16376 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_162
timestamp 1624635492
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_158
timestamp 1624635492
transform 1 0 15640 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1624635492
transform 1 0 16100 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 16468 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_20_174
timestamp 1624635492
transform 1 0 17112 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_170
timestamp 1624635492
transform 1 0 16744 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_172
timestamp 1624635492
transform 1 0 16928 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_167
timestamp 1624635492
transform 1 0 16468 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A1
timestamp 1624635492
transform -1 0 16744 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 17204 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_left_track_1.prog_clk
timestamp 1624635492
transform -1 0 17388 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1624635492
transform 1 0 16836 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_177
timestamp 1624635492
transform 1 0 17388 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_177
timestamp 1624635492
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1624635492
transform -1 0 18400 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1624635492
transform -1 0 18400 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1624635492
transform 1 0 18584 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1624635492
transform 1 0 19504 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_188
timestamp 1624635492
transform 1 0 18400 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_199
timestamp 1624635492
transform 1 0 19412 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_188
timestamp 1624635492
transform 1 0 18400 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_201
timestamp 1624635492
transform 1 0 19596 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1624635492
transform -1 0 21896 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1624635492
transform -1 0 21896 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_211
timestamp 1624635492
transform 1 0 20516 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_213
timestamp 1624635492
transform 1 0 20700 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_221
timestamp 1624635492
transform 1 0 21436 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp 1624635492
transform 1 0 2116 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 2576 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1624635492
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output61
timestamp 1624635492
transform -1 0 1932 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1624635492
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_9
timestamp 1624635492
transform 1 0 1932 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_14
timestamp 1624635492
transform 1 0 2392 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_19
timestamp 1624635492
transform 1 0 2852 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1624635492
transform 1 0 3128 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 6164 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1624635492
transform 1 0 3588 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1624635492
transform 1 0 4048 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_25
timestamp 1624635492
transform 1 0 3404 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_30
timestamp 1624635492
transform 1 0 3864 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_35
timestamp 1624635492
transform 1 0 4324 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1624635492
transform 1 0 6624 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1624635492
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_55
timestamp 1624635492
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_58
timestamp 1624635492
transform 1 0 6440 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 9568 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1624635492
transform -1 0 7820 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_69
timestamp 1624635492
transform 1 0 7452 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_73
timestamp 1624635492
transform 1 0 7820 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 11224 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_92
timestamp 1624635492
transform 1 0 9568 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1624635492
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_left_track_1.prog_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 13708 0 1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_21_110
timestamp 1624635492
transform 1 0 11224 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_115
timestamp 1624635492
transform 1 0 11684 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 15364 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_137
timestamp 1624635492
transform 1 0 13708 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1624635492
transform -1 0 16376 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_155
timestamp 1624635492
transform 1 0 15364 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_166
timestamp 1624635492
transform 1 0 16376 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 19228 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1624635492
transform 1 0 16836 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_170
timestamp 1624635492
transform 1 0 16744 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_172
timestamp 1624635492
transform 1 0 16928 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_176
timestamp 1624635492
transform 1 0 17296 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_179
timestamp 1624635492
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_197
timestamp 1624635492
transform 1 0 19228 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1624635492
transform -1 0 21896 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_209
timestamp 1624635492
transform 1 0 20332 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_221
timestamp 1624635492
transform 1 0 21436 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l2_in_0_
timestamp 1624635492
transform 1 0 2760 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1624635492
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output72
timestamp 1624635492
transform -1 0 1932 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output73
timestamp 1624635492
transform -1 0 2484 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1624635492
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_9
timestamp 1624635492
transform 1 0 1932 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_15
timestamp 1624635492
transform 1 0 2484 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 4048 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1624635492
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1624635492
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_30
timestamp 1624635492
transform 1 0 3864 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1624635492
transform -1 0 6164 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 6348 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_22_48
timestamp 1624635492
transform 1 0 5520 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_55
timestamp 1624635492
transform 1 0 6164 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input55
timestamp 1624635492
transform 1 0 8004 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input57
timestamp 1624635492
transform 1 0 8464 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_73
timestamp 1624635492
transform 1 0 7820 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_78
timestamp 1624635492
transform 1 0 8280 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_83
timestamp 1624635492
transform 1 0 8740 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 10580 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l3_in_0_
timestamp 1624635492
transform -1 0 10396 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1624635492
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1624635492
transform -1 0 9292 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_89
timestamp 1624635492
transform 1 0 9292 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_101
timestamp 1624635492
transform 1 0 10396 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_0_
timestamp 1624635492
transform 1 0 12236 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_119
timestamp 1624635492
transform 1 0 12052 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1624635492
transform -1 0 14076 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1624635492
transform 1 0 14260 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_130
timestamp 1624635492
transform 1 0 13064 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1624635492
transform 1 0 14076 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_144
timestamp 1624635492
transform 1 0 14352 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 16836 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_left_track_1.prog_clk
timestamp 1624635492
transform -1 0 14812 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_149
timestamp 1624635492
transform 1 0 14812 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_153
timestamp 1624635492
transform 1 0 15180 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l2_in_0_
timestamp 1624635492
transform -1 0 18492 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 17204 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_171
timestamp 1624635492
transform 1 0 16836 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_175
timestamp 1624635492
transform 1 0 17204 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_179
timestamp 1624635492
transform 1 0 17572 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1624635492
transform 1 0 19504 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_189
timestamp 1624635492
transform 1 0 18492 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_197
timestamp 1624635492
transform 1 0 19228 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_201
timestamp 1624635492
transform 1 0 19596 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1624635492
transform -1 0 21896 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_213
timestamp 1624635492
transform 1 0 20700 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_221
timestamp 1624635492
transform 1 0 21436 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp 1624635492
transform 1 0 2116 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 2576 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1624635492
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output74
timestamp 1624635492
transform -1 0 1932 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1624635492
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_9
timestamp 1624635492
transform 1 0 1932 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_14
timestamp 1624635492
transform 1 0 2392 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l1_in_0_
timestamp 1624635492
transform 1 0 4232 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_32
timestamp 1624635492
transform 1 0 4048 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1624635492
transform -1 0 7452 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1624635492
transform 1 0 5336 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1624635492
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_43
timestamp 1624635492
transform 1 0 5060 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_55
timestamp 1624635492
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_58
timestamp 1624635492
transform 1 0 6440 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1624635492
transform -1 0 8096 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 9752 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_23_69
timestamp 1624635492
transform 1 0 7452 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_76
timestamp 1624635492
transform 1 0 8096 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 11408 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_94
timestamp 1624635492
transform 1 0 9752 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1624635492
transform -1 0 12880 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1624635492
transform 1 0 11592 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1624635492
transform -1 0 11868 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_112
timestamp 1624635492
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_117
timestamp 1624635492
transform 1 0 11868 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 14536 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_128
timestamp 1624635492
transform 1 0 12880 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1624635492
transform 1 0 14720 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1624635492
transform -1 0 16652 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_146
timestamp 1624635492
transform 1 0 14536 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_157
timestamp 1624635492
transform 1 0 15548 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 17940 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1624635492
transform 1 0 16836 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 17480 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 16928 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1624635492
transform 1 0 16652 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_174
timestamp 1624635492
transform 1 0 17112 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_180
timestamp 1624635492
transform 1 0 17664 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_199
timestamp 1624635492
transform 1 0 19412 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1624635492
transform -1 0 21896 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_211
timestamp 1624635492
transform 1 0 20516 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp 1624635492
transform 1 0 2116 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1624635492
transform -1 0 2852 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1624635492
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output75
timestamp 1624635492
transform -1 0 1932 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1624635492
transform 1 0 1380 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_9
timestamp 1624635492
transform 1 0 1932 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_14
timestamp 1624635492
transform 1 0 2392 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_19
timestamp 1624635492
transform 1 0 2852 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 5980 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 3036 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 4048 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1624635492
transform 1 0 3772 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_24
timestamp 1624635492
transform 1 0 3312 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_28
timestamp 1624635492
transform 1 0 3680 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_30
timestamp 1624635492
transform 1 0 3864 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_35
timestamp 1624635492
transform 1 0 4324 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _066_
timestamp 1624635492
transform 1 0 6164 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 6624 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_24_53
timestamp 1624635492
transform 1 0 5980 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_58
timestamp 1624635492
transform 1 0 6440 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1624635492
transform 1 0 8280 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_76
timestamp 1624635492
transform 1 0 8096 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_81
timestamp 1624635492
transform 1 0 8556 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1624635492
transform 1 0 9292 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1624635492
transform 1 0 9016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_left_track_1.prog_clk
timestamp 1624635492
transform -1 0 10580 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_85
timestamp 1624635492
transform 1 0 8924 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_87
timestamp 1624635492
transform 1 0 9108 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_98
timestamp 1624635492
transform 1 0 10120 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_103
timestamp 1624635492
transform 1 0 10580 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 12328 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1624635492
transform -1 0 12696 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_122
timestamp 1624635492
transform 1 0 12328 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1624635492
transform 1 0 13248 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1624635492
transform 1 0 14260 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 13064 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 14352 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_126
timestamp 1624635492
transform 1 0 12696 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_130
timestamp 1624635492
transform 1 0 13064 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1624635492
transform 1 0 14076 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 15732 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_left_track_1.prog_clk
timestamp 1624635492
transform -1 0 15548 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 14904 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_146
timestamp 1624635492
transform 1 0 14536 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_152
timestamp 1624635492
transform 1 0 15088 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_157
timestamp 1624635492
transform 1 0 15548 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_0_
timestamp 1624635492
transform -1 0 18492 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_175
timestamp 1624635492
transform 1 0 17204 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_179
timestamp 1624635492
transform 1 0 17572 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1624635492
transform 1 0 18676 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1624635492
transform 1 0 19504 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 19136 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_189
timestamp 1624635492
transform 1 0 18492 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1624635492
transform 1 0 18952 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_198
timestamp 1624635492
transform 1 0 19320 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_201
timestamp 1624635492
transform 1 0 19596 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1624635492
transform -1 0 21896 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_213
timestamp 1624635492
transform 1 0 20700 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_221
timestamp 1624635492
transform 1 0 21436 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp 1624635492
transform 1 0 2116 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp 1624635492
transform 1 0 2576 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1624635492
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output76
timestamp 1624635492
transform -1 0 1932 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1624635492
transform 1 0 1380 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_9
timestamp 1624635492
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_14
timestamp 1624635492
transform 1 0 2392 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_19
timestamp 1624635492
transform 1 0 2852 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 4600 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 3036 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 3496 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 3956 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_24
timestamp 1624635492
transform 1 0 3312 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_29
timestamp 1624635492
transform 1 0 3772 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_34
timestamp 1624635492
transform 1 0 4232 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1624635492
transform 1 0 6348 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1624635492
transform 1 0 6624 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_54
timestamp 1624635492
transform 1 0 6072 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_58
timestamp 1624635492
transform 1 0 6440 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 8648 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1624635492
transform 1 0 7636 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1624635492
transform 1 0 7084 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_63
timestamp 1624635492
transform 1 0 6900 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_68
timestamp 1624635492
transform 1 0 7360 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_80
timestamp 1624635492
transform 1 0 8464 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_0_
timestamp 1624635492
transform 1 0 10580 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_25_98
timestamp 1624635492
transform 1 0 10120 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_102
timestamp 1624635492
transform 1 0 10488 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1624635492
transform 1 0 11868 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1624635492
transform 1 0 11592 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_112
timestamp 1624635492
transform 1 0 11408 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_115
timestamp 1624635492
transform 1 0 11684 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 13800 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_left_track_1.prog_clk
timestamp 1624635492
transform 1 0 12880 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1624635492
transform -1 0 13524 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_126
timestamp 1624635492
transform 1 0 12696 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_131
timestamp 1624635492
transform 1 0 13156 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_135
timestamp 1624635492
transform 1 0 13524 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_0_
timestamp 1624635492
transform -1 0 16560 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_25_154
timestamp 1624635492
transform 1 0 15272 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_158
timestamp 1624635492
transform 1 0 15640 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 19688 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l2_in_0_
timestamp 1624635492
transform -1 0 17940 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1624635492
transform 1 0 16836 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_168
timestamp 1624635492
transform 1 0 16560 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_172
timestamp 1624635492
transform 1 0 16928 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_183
timestamp 1624635492
transform 1 0 17940 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 20056 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_202
timestamp 1624635492
transform 1 0 19688 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_206
timestamp 1624635492
transform 1 0 20056 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1624635492
transform -1 0 21896 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_218
timestamp 1624635492
transform 1 0 21160 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_222
timestamp 1624635492
transform 1 0 21528 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_9
timestamp 1624635492
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1624635492
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_9
timestamp 1624635492
transform 1 0 1932 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1624635492
transform 1 0 1380 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output78
timestamp 1624635492
transform -1 0 1932 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output77
timestamp 1624635492
transform -1 0 1932 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1624635492
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1624635492
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_15
timestamp 1624635492
transform 1 0 2484 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_19
timestamp 1624635492
transform 1 0 2852 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_14
timestamp 1624635492
transform 1 0 2392 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output80
timestamp 1624635492
transform -1 0 2484 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1624635492
transform 1 0 2576 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp 1624635492
transform 1 0 2116 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 4140 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1624635492
transform 1 0 3128 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1624635492
transform 1 0 4692 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 4324 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l1_in_0_
timestamp 1624635492
transform 1 0 4324 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1624635492
transform 1 0 3772 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_25
timestamp 1624635492
transform 1 0 3404 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_30
timestamp 1624635492
transform 1 0 3864 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_35
timestamp 1624635492
transform 1 0 4324 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_33
timestamp 1624635492
transform 1 0 4140 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_44
timestamp 1624635492
transform 1 0 5152 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_48
timestamp 1624635492
transform 1 0 5520 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1624635492
transform 1 0 5704 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1624635492
transform 1 0 5336 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_27_60
timestamp 1624635492
transform 1 0 6624 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_55
timestamp 1624635492
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_58
timestamp 1624635492
transform 1 0 6440 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_53
timestamp 1624635492
transform 1 0 5980 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1624635492
transform -1 0 6624 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1624635492
transform -1 0 6808 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1624635492
transform 1 0 6164 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1624635492
transform 1 0 6348 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_62
timestamp 1624635492
transform 1 0 6808 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1624635492
transform -1 0 9016 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1624635492
transform -1 0 7268 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 8464 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1624635492
transform 1 0 7452 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1624635492
transform 1 0 8464 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_67
timestamp 1624635492
transform 1 0 7268 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_78
timestamp 1624635492
transform 1 0 8280 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_83
timestamp 1624635492
transform 1 0 8740 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_80
timestamp 1624635492
transform 1 0 8464 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 9200 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1624635492
transform 1 0 9292 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1624635492
transform 1 0 9016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1624635492
transform 1 0 10304 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_87
timestamp 1624635492
transform 1 0 9108 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_98
timestamp 1624635492
transform 1 0 10120 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_103
timestamp 1624635492
transform 1 0 10580 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_86
timestamp 1624635492
transform 1 0 9016 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_104
timestamp 1624635492
transform 1 0 10672 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_113
timestamp 1624635492
transform 1 0 11500 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_109
timestamp 1624635492
transform 1 0 11132 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1624635492
transform 1 0 10856 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1624635492
transform 1 0 11592 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_123
timestamp 1624635492
transform 1 0 12420 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_117
timestamp 1624635492
transform 1 0 11868 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_121
timestamp 1624635492
transform 1 0 12236 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1624635492
transform -1 0 11868 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_left_track_1.prog_clk
timestamp 1624635492
transform 1 0 12420 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1624635492
transform -1 0 12420 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 10764 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_26_126
timestamp 1624635492
transform 1 0 12696 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1624635492
transform -1 0 13708 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1624635492
transform -1 0 13616 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1624635492
transform -1 0 13984 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1624635492
transform -1 0 14076 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_137
timestamp 1624635492
transform 1 0 13708 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_136
timestamp 1624635492
transform 1 0 13616 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1624635492
transform 1 0 14260 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1624635492
transform -1 0 14352 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 14536 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1624635492
transform 1 0 14076 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_140
timestamp 1624635492
transform 1 0 13984 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_144
timestamp 1624635492
transform 1 0 14352 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 16100 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 14812 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1624635492
transform -1 0 15824 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_26_146
timestamp 1624635492
transform 1 0 14536 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_150
timestamp 1624635492
transform 1 0 14904 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_160
timestamp 1624635492
transform 1 0 15824 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_148
timestamp 1624635492
transform 1 0 14720 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_165
timestamp 1624635492
transform 1 0 16284 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_177
timestamp 1624635492
transform 1 0 17388 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_172
timestamp 1624635492
transform 1 0 16928 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1624635492
transform 1 0 16652 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 16652 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1624635492
transform 1 0 16836 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1624635492
transform -1 0 17388 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_181
timestamp 1624635492
transform 1 0 17756 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_179
timestamp 1624635492
transform 1 0 17572 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 17848 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 17756 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l2_in_0_
timestamp 1624635492
transform 1 0 19504 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1624635492
transform 1 0 19504 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 19596 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A0
timestamp 1624635492
transform -1 0 20148 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_197
timestamp 1624635492
transform 1 0 19228 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_203
timestamp 1624635492
transform 1 0 19780 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_207
timestamp 1624635492
transform 1 0 20148 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_198
timestamp 1624635492
transform 1 0 19320 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1624635492
transform -1 0 21896 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1624635492
transform -1 0 21896 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_219
timestamp 1624635492
transform 1 0 21252 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_209
timestamp 1624635492
transform 1 0 20332 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_221
timestamp 1624635492
transform 1 0 21436 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l2_in_0_
timestamp 1624635492
transform -1 0 3588 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1624635492
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output69
timestamp 1624635492
transform -1 0 1932 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output79
timestamp 1624635492
transform -1 0 2484 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1624635492
transform 1 0 1380 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_9
timestamp 1624635492
transform 1 0 1932 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_15
timestamp 1624635492
transform 1 0 2484 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1624635492
transform 1 0 4048 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 6256 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1624635492
transform 1 0 3772 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_27
timestamp 1624635492
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_30
timestamp 1624635492
transform 1 0 3864 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_35
timestamp 1624635492
transform 1 0 4324 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_39
timestamp 1624635492
transform 1 0 4692 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 6440 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_56
timestamp 1624635492
transform 1 0 6256 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_61
timestamp 1624635492
transform 1 0 6716 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 7176 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_28_65
timestamp 1624635492
transform 1 0 7084 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_82
timestamp 1624635492
transform 1 0 8648 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1624635492
transform -1 0 10120 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1624635492
transform 1 0 9016 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1624635492
transform 1 0 10304 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_87
timestamp 1624635492
transform 1 0 9108 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_98
timestamp 1624635492
transform 1 0 10120 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_103
timestamp 1624635492
transform 1 0 10580 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 13156 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 1624635492
transform -1 0 11500 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input30
timestamp 1624635492
transform -1 0 11040 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_108
timestamp 1624635492
transform 1 0 11040 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_113
timestamp 1624635492
transform 1 0 11500 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1624635492
transform 1 0 14260 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input31
timestamp 1624635492
transform -1 0 13616 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 1624635492
transform -1 0 14076 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1624635492
transform -1 0 14536 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_131
timestamp 1624635492
transform 1 0 13156 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_136
timestamp 1624635492
transform 1 0 13616 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1624635492
transform 1 0 14076 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1624635492
transform -1 0 15640 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1624635492
transform 1 0 15824 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_28_146
timestamp 1624635492
transform 1 0 14536 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_158
timestamp 1624635492
transform 1 0 15640 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1624635492
transform 1 0 16836 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_0_
timestamp 1624635492
transform -1 0 18400 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_169
timestamp 1624635492
transform 1 0 16652 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_174
timestamp 1624635492
transform 1 0 17112 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_178
timestamp 1624635492
transform 1 0 17480 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1624635492
transform -1 0 18860 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1624635492
transform 1 0 19504 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 19228 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_188
timestamp 1624635492
transform 1 0 18400 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_193
timestamp 1624635492
transform 1 0 18860 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_197
timestamp 1624635492
transform 1 0 19228 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_201
timestamp 1624635492
transform 1 0 19596 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1624635492
transform -1 0 21896 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_213
timestamp 1624635492
transform 1 0 20700 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_221
timestamp 1624635492
transform 1 0 21436 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 2852 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1624635492
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output62
timestamp 1624635492
transform -1 0 1932 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output68
timestamp 1624635492
transform -1 0 2484 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1624635492
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_9
timestamp 1624635492
transform 1 0 1932 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_15
timestamp 1624635492
transform 1 0 2484 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1624635492
transform 1 0 4784 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_29_35
timestamp 1624635492
transform 1 0 4324 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_39
timestamp 1624635492
transform 1 0 4692 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1624635492
transform 1 0 5796 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1624635492
transform 1 0 6808 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1624635492
transform 1 0 6348 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1624635492
transform 1 0 6440 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_49
timestamp 1624635492
transform 1 0 5612 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_54
timestamp 1624635492
transform 1 0 6072 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_60
timestamp 1624635492
transform 1 0 6624 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 7820 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 8280 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_71
timestamp 1624635492
transform 1 0 7636 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_76
timestamp 1624635492
transform 1 0 8096 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_81
timestamp 1624635492
transform 1 0 8556 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1624635492
transform 1 0 9292 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 8832 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1624635492
transform 1 0 10304 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_87
timestamp 1624635492
transform 1 0 9108 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_98
timestamp 1624635492
transform 1 0 10120 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_103
timestamp 1624635492
transform 1 0 10580 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1624635492
transform -1 0 12696 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1624635492
transform 1 0 11592 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1624635492
transform 1 0 10764 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1624635492
transform -1 0 11408 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_108
timestamp 1624635492
transform 1 0 11040 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_112
timestamp 1624635492
transform 1 0 11408 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_115
timestamp 1624635492
transform 1 0 11684 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 15548 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1624635492
transform 1 0 12880 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_126
timestamp 1624635492
transform 1 0 12696 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_137
timestamp 1624635492
transform 1 0 13708 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1624635492
transform 1 0 15732 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_157
timestamp 1624635492
transform 1 0 15548 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 17388 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 18032 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1624635492
transform 1 0 16836 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_left_track_1.prog_clk
timestamp 1624635492
transform -1 0 18492 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_168
timestamp 1624635492
transform 1 0 16560 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_172
timestamp 1624635492
transform 1 0 16928 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_177
timestamp 1624635492
transform 1 0 17388 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_184
timestamp 1624635492
transform 1 0 18032 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 18860 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_189
timestamp 1624635492
transform 1 0 18492 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_193
timestamp 1624635492
transform 1 0 18860 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_205
timestamp 1624635492
transform 1 0 19964 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1624635492
transform -1 0 21896 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1624635492
transform 1 0 21068 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp 1624635492
transform 1 0 2668 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1624635492
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output63
timestamp 1624635492
transform -1 0 1932 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output67
timestamp 1624635492
transform -1 0 2484 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1624635492
transform 1 0 1380 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_9
timestamp 1624635492
transform 1 0 1932 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_15
timestamp 1624635492
transform 1 0 2484 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_20
timestamp 1624635492
transform 1 0 2944 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1624635492
transform 1 0 3128 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp 1624635492
transform 1 0 4048 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1624635492
transform 1 0 4508 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1624635492
transform 1 0 3772 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_25
timestamp 1624635492
transform 1 0 3404 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_30
timestamp 1624635492
transform 1 0 3864 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_35
timestamp 1624635492
transform 1 0 4324 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_40
timestamp 1624635492
transform 1 0 4784 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp 1624635492
transform -1 0 6900 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 4968 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_58
timestamp 1624635492
transform 1 0 6440 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1624635492
transform 1 0 8464 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1624635492
transform -1 0 8280 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1624635492
transform 1 0 7084 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_63
timestamp 1624635492
transform 1 0 6900 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_67
timestamp 1624635492
transform 1 0 7268 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_78
timestamp 1624635492
transform 1 0 8280 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_83
timestamp 1624635492
transform 1 0 8740 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 10764 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1624635492
transform 1 0 9016 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_87
timestamp 1624635492
transform 1 0 9108 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1624635492
transform -1 0 12604 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1624635492
transform 1 0 10948 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1624635492
transform -1 0 11592 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_105
timestamp 1624635492
transform 1 0 10764 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_110
timestamp 1624635492
transform 1 0 11224 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_114
timestamp 1624635492
transform 1 0 11592 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_125
timestamp 1624635492
transform 1 0 12604 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 13248 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 14076 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1624635492
transform 1 0 14260 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1624635492
transform -1 0 13616 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1624635492
transform -1 0 14536 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_132
timestamp 1624635492
transform 1 0 13248 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_136
timestamp 1624635492
transform 1 0 13616 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1624635492
transform 1 0 14076 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 17480 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1624635492
transform -1 0 15548 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_30_146
timestamp 1624635492
transform 1 0 14536 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_157
timestamp 1624635492
transform 1 0 15548 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_161
timestamp 1624635492
transform 1 0 15916 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 17940 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 18400 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_178
timestamp 1624635492
transform 1 0 17480 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_183
timestamp 1624635492
transform 1 0 17940 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 18584 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1624635492
transform 1 0 19504 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output90_A
timestamp 1624635492
transform 1 0 19044 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_188
timestamp 1624635492
transform 1 0 18400 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_193
timestamp 1624635492
transform 1 0 18860 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_197
timestamp 1624635492
transform 1 0 19228 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_201
timestamp 1624635492
transform 1 0 19596 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1624635492
transform -1 0 21896 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1624635492
transform -1 0 21436 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_213
timestamp 1624635492
transform 1 0 20700 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_221
timestamp 1624635492
transform 1 0 21436 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 4140 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1624635492
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output64
timestamp 1624635492
transform -1 0 1932 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output66
timestamp 1624635492
transform -1 0 2484 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1624635492
transform 1 0 1380 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_9
timestamp 1624635492
transform 1 0 1932 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_15
timestamp 1624635492
transform 1 0 2484 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 6164 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1624635492
transform -1 0 4508 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_33
timestamp 1624635492
transform 1 0 4140 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_37
timestamp 1624635492
transform 1 0 4508 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1624635492
transform 1 0 6624 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1624635492
transform 1 0 6348 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_55
timestamp 1624635492
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_58
timestamp 1624635492
transform 1 0 6440 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 8924 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1624635492
transform -1 0 7268 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_63
timestamp 1624635492
transform 1 0 6900 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_67
timestamp 1624635492
transform 1 0 7268 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1624635492
transform -1 0 9476 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 9660 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_31_85
timestamp 1624635492
transform 1 0 8924 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_91
timestamp 1624635492
transform 1 0 9476 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 12788 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 12328 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1624635492
transform 1 0 11592 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1624635492
transform -1 0 11868 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_109
timestamp 1624635492
transform 1 0 11132 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_113
timestamp 1624635492
transform 1 0 11500 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_117
timestamp 1624635492
transform 1 0 11868 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_122
timestamp 1624635492
transform 1 0 12328 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp 1624635492
transform -1 0 13248 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp 1624635492
transform 1 0 13800 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp 1624635492
transform 1 0 14260 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1624635492
transform -1 0 13616 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_127
timestamp 1624635492
transform 1 0 12788 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_132
timestamp 1624635492
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_136
timestamp 1624635492
transform 1 0 13616 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_141
timestamp 1624635492
transform 1 0 14076 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1624635492
transform -1 0 14996 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp 1624635492
transform -1 0 15548 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 1624635492
transform -1 0 16100 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 16284 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_146
timestamp 1624635492
transform 1 0 14536 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_151
timestamp 1624635492
transform 1 0 14996 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_157
timestamp 1624635492
transform 1 0 15548 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_163
timestamp 1624635492
transform 1 0 16100 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp 1624635492
transform 1 0 17112 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 1624635492
transform -1 0 17848 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 1624635492
transform 1 0 18032 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1624635492
transform 1 0 16836 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_168
timestamp 1624635492
transform 1 0 16560 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_172
timestamp 1624635492
transform 1 0 16928 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_177
timestamp 1624635492
transform 1 0 17388 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_182
timestamp 1624635492
transform 1 0 17848 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_187
timestamp 1624635492
transform 1 0 18308 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp 1624635492
transform 1 0 18492 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp 1624635492
transform -1 0 19228 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 19412 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output91_A
timestamp 1624635492
transform 1 0 19780 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_192
timestamp 1624635492
transform 1 0 18768 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_197
timestamp 1624635492
transform 1 0 19228 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_201
timestamp 1624635492
transform 1 0 19596 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_205
timestamp 1624635492
transform 1 0 19964 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 21436 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1624635492
transform -1 0 21896 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_221
timestamp 1624635492
transform 1 0 21436 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1624635492
transform -1 0 3588 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1624635492
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input56
timestamp 1624635492
transform 1 0 2208 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output65
timestamp 1624635492
transform -1 0 1932 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1624635492
transform 1 0 1380 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_9
timestamp 1624635492
transform 1 0 1932 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_16
timestamp 1624635492
transform 1 0 2576 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1624635492
transform 1 0 4048 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1624635492
transform -1 0 5336 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1624635492
transform 1 0 3772 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_27
timestamp 1624635492
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_30
timestamp 1624635492
transform 1 0 3864 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_35
timestamp 1624635492
transform 1 0 4324 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 6992 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_32_46
timestamp 1624635492
transform 1 0 5336 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1624635492
transform 1 0 8004 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 7176 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1624635492
transform -1 0 7820 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_64
timestamp 1624635492
transform 1 0 6992 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_69
timestamp 1624635492
transform 1 0 7452 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_73
timestamp 1624635492
transform 1 0 7820 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 11500 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1624635492
transform 1 0 9016 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1624635492
transform 1 0 9292 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_84
timestamp 1624635492
transform 1 0 8832 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_87
timestamp 1624635492
transform 1 0 9108 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_92
timestamp 1624635492
transform 1 0 9568 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_96
timestamp 1624635492
transform 1 0 9936 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 12604 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 12144 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_113
timestamp 1624635492
transform 1 0 11500 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_120
timestamp 1624635492
transform 1 0 12144 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_125
timestamp 1624635492
transform 1 0 12604 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp 1624635492
transform -1 0 13432 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1624635492
transform 1 0 13616 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1624635492
transform 1 0 14260 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1624635492
transform -1 0 12972 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_129
timestamp 1624635492
transform 1 0 12972 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_134
timestamp 1624635492
transform 1 0 13432 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_139
timestamp 1624635492
transform 1 0 13892 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_144
timestamp 1624635492
transform 1 0 14352 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 14904 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output96
timestamp 1624635492
transform -1 0 15732 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output97
timestamp 1624635492
transform -1 0 16284 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_150
timestamp 1624635492
transform 1 0 14904 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_154
timestamp 1624635492
transform 1 0 15272 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_159
timestamp 1624635492
transform 1 0 15732 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_165
timestamp 1624635492
transform 1 0 16284 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp 1624635492
transform -1 0 18400 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output98
timestamp 1624635492
transform -1 0 16836 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output99
timestamp 1624635492
transform -1 0 17388 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output100
timestamp 1624635492
transform -1 0 17940 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_171
timestamp 1624635492
transform 1 0 16836 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_177
timestamp 1624635492
transform 1 0 17388 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_183
timestamp 1624635492
transform 1 0 17940 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 18860 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1624635492
transform 1 0 19504 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output87
timestamp 1624635492
transform -1 0 20332 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 19044 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 19780 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_188
timestamp 1624635492
transform 1 0 18400 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_193
timestamp 1624635492
transform 1 0 18860 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_197
timestamp 1624635492
transform 1 0 19228 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_203
timestamp 1624635492
transform 1 0 19780 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1624635492
transform -1 0 21896 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output88
timestamp 1624635492
transform -1 0 20884 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output89
timestamp 1624635492
transform -1 0 21436 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_209
timestamp 1624635492
transform 1 0 20332 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_215
timestamp 1624635492
transform 1 0 20884 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_221
timestamp 1624635492
transform 1 0 21436 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1624635492
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1624635492
transform 1 0 1564 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input52
timestamp 1624635492
transform 1 0 2116 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input53
timestamp 1624635492
transform 1 0 2668 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1624635492
transform 1 0 1380 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_9
timestamp 1624635492
transform 1 0 1932 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_15
timestamp 1624635492
transform 1 0 2484 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1624635492
transform 1 0 4048 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1624635492
transform 1 0 3772 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input54
timestamp 1624635492
transform 1 0 3220 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_21
timestamp 1624635492
transform 1 0 3036 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_27
timestamp 1624635492
transform 1 0 3588 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_30
timestamp 1624635492
transform 1 0 3864 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_41
timestamp 1624635492
transform 1 0 4876 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1624635492
transform 1 0 5428 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1624635492
transform 1 0 6440 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input58
timestamp 1624635492
transform 1 0 6716 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1624635492
transform -1 0 5244 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_45
timestamp 1624635492
transform 1 0 5244 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_56
timestamp 1624635492
transform 1 0 6256 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1624635492
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1624635492
transform 1 0 8372 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output70
timestamp 1624635492
transform -1 0 7636 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output71
timestamp 1624635492
transform -1 0 8188 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_65
timestamp 1624635492
transform 1 0 7084 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_71
timestamp 1624635492
transform 1 0 7636 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_77
timestamp 1624635492
transform 1 0 8188 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_82
timestamp 1624635492
transform 1 0 8648 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1624635492
transform 1 0 9384 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1624635492
transform 1 0 9108 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1624635492
transform 1 0 10396 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_86
timestamp 1624635492
transform 1 0 9016 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_88
timestamp 1624635492
transform 1 0 9200 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_99
timestamp 1624635492
transform 1 0 10212 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_104
timestamp 1624635492
transform 1 0 10672 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1624635492
transform 1 0 11776 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1624635492
transform 1 0 12052 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output94
timestamp 1624635492
transform 1 0 12512 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output95
timestamp 1624635492
transform 1 0 11224 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1624635492
transform -1 0 11040 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_108
timestamp 1624635492
transform 1 0 11040 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_114
timestamp 1624635492
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_117
timestamp 1624635492
transform 1 0 11868 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_122
timestamp 1624635492
transform 1 0 12328 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1624635492
transform 1 0 14444 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output81
timestamp 1624635492
transform -1 0 13432 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output92
timestamp 1624635492
transform -1 0 13984 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_128
timestamp 1624635492
transform 1 0 12880 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_134
timestamp 1624635492
transform 1 0 13432 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_140
timestamp 1624635492
transform 1 0 13984 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_144
timestamp 1624635492
transform 1 0 14352 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output90
timestamp 1624635492
transform 1 0 16008 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output91
timestamp 1624635492
transform 1 0 15456 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output93
timestamp 1624635492
transform -1 0 15088 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_146
timestamp 1624635492
transform 1 0 14536 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_152
timestamp 1624635492
transform 1 0 15088 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_160
timestamp 1624635492
transform 1 0 15824 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1624635492
transform 1 0 16376 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1624635492
transform 1 0 17112 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output82
timestamp 1624635492
transform -1 0 18032 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output83
timestamp 1624635492
transform -1 0 18584 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output86
timestamp 1624635492
transform 1 0 16560 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1624635492
transform -1 0 17388 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_172
timestamp 1624635492
transform 1 0 16928 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_177
timestamp 1624635492
transform 1 0 17388 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_184
timestamp 1624635492
transform 1 0 18032 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1624635492
transform 1 0 19780 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output84
timestamp 1624635492
transform -1 0 19136 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output85
timestamp 1624635492
transform -1 0 20424 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 19504 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_190
timestamp 1624635492
transform 1 0 18584 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_196
timestamp 1624635492
transform 1 0 19136 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_200
timestamp 1624635492
transform 1 0 19504 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_204
timestamp 1624635492
transform 1 0 19872 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1624635492
transform -1 0 21896 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input59
timestamp 1624635492
transform -1 0 21436 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1624635492
transform -1 0 20884 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_210
timestamp 1624635492
transform 1 0 20424 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_215
timestamp 1624635492
transform 1 0 20884 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_221
timestamp 1624635492
transform 1 0 21436 0 1 20128
box -38 -48 222 592
<< labels >>
rlabel metal3 s 22200 11432 23000 11552 6 ccff_head
port 0 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 ccff_tail
port 1 nsew signal tristate
rlabel metal3 s 0 4360 800 4480 6 chanx_left_in[0]
port 2 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 chanx_left_in[10]
port 3 nsew signal input
rlabel metal3 s 0 9392 800 9512 6 chanx_left_in[11]
port 4 nsew signal input
rlabel metal3 s 0 9936 800 10056 6 chanx_left_in[12]
port 5 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 chanx_left_in[13]
port 6 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 chanx_left_in[14]
port 7 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 chanx_left_in[15]
port 8 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 chanx_left_in[16]
port 9 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 chanx_left_in[17]
port 10 nsew signal input
rlabel metal3 s 0 12792 800 12912 6 chanx_left_in[18]
port 11 nsew signal input
rlabel metal3 s 0 13200 800 13320 6 chanx_left_in[19]
port 12 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 chanx_left_in[1]
port 13 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 chanx_left_in[2]
port 14 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 chanx_left_in[3]
port 15 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 chanx_left_in[4]
port 16 nsew signal input
rlabel metal3 s 0 6672 800 6792 6 chanx_left_in[5]
port 17 nsew signal input
rlabel metal3 s 0 7080 800 7200 6 chanx_left_in[6]
port 18 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 chanx_left_in[7]
port 19 nsew signal input
rlabel metal3 s 0 8032 800 8152 6 chanx_left_in[8]
port 20 nsew signal input
rlabel metal3 s 0 8576 800 8696 6 chanx_left_in[9]
port 21 nsew signal input
rlabel metal3 s 0 13744 800 13864 6 chanx_left_out[0]
port 22 nsew signal tristate
rlabel metal3 s 0 18368 800 18488 6 chanx_left_out[10]
port 23 nsew signal tristate
rlabel metal3 s 0 18776 800 18896 6 chanx_left_out[11]
port 24 nsew signal tristate
rlabel metal3 s 0 19320 800 19440 6 chanx_left_out[12]
port 25 nsew signal tristate
rlabel metal3 s 0 19728 800 19848 6 chanx_left_out[13]
port 26 nsew signal tristate
rlabel metal3 s 0 20272 800 20392 6 chanx_left_out[14]
port 27 nsew signal tristate
rlabel metal3 s 0 20680 800 20800 6 chanx_left_out[15]
port 28 nsew signal tristate
rlabel metal3 s 0 21224 800 21344 6 chanx_left_out[16]
port 29 nsew signal tristate
rlabel metal3 s 0 21632 800 21752 6 chanx_left_out[17]
port 30 nsew signal tristate
rlabel metal3 s 0 22176 800 22296 6 chanx_left_out[18]
port 31 nsew signal tristate
rlabel metal3 s 0 22584 800 22704 6 chanx_left_out[19]
port 32 nsew signal tristate
rlabel metal3 s 0 14152 800 14272 6 chanx_left_out[1]
port 33 nsew signal tristate
rlabel metal3 s 0 14560 800 14680 6 chanx_left_out[2]
port 34 nsew signal tristate
rlabel metal3 s 0 15104 800 15224 6 chanx_left_out[3]
port 35 nsew signal tristate
rlabel metal3 s 0 15512 800 15632 6 chanx_left_out[4]
port 36 nsew signal tristate
rlabel metal3 s 0 16056 800 16176 6 chanx_left_out[5]
port 37 nsew signal tristate
rlabel metal3 s 0 16464 800 16584 6 chanx_left_out[6]
port 38 nsew signal tristate
rlabel metal3 s 0 17008 800 17128 6 chanx_left_out[7]
port 39 nsew signal tristate
rlabel metal3 s 0 17416 800 17536 6 chanx_left_out[8]
port 40 nsew signal tristate
rlabel metal3 s 0 17960 800 18080 6 chanx_left_out[9]
port 41 nsew signal tristate
rlabel metal2 s 3882 22200 3938 23000 6 chany_top_in[0]
port 42 nsew signal input
rlabel metal2 s 8482 22200 8538 23000 6 chany_top_in[10]
port 43 nsew signal input
rlabel metal2 s 8942 22200 8998 23000 6 chany_top_in[11]
port 44 nsew signal input
rlabel metal2 s 9402 22200 9458 23000 6 chany_top_in[12]
port 45 nsew signal input
rlabel metal2 s 9862 22200 9918 23000 6 chany_top_in[13]
port 46 nsew signal input
rlabel metal2 s 10322 22200 10378 23000 6 chany_top_in[14]
port 47 nsew signal input
rlabel metal2 s 10782 22200 10838 23000 6 chany_top_in[15]
port 48 nsew signal input
rlabel metal2 s 11242 22200 11298 23000 6 chany_top_in[16]
port 49 nsew signal input
rlabel metal2 s 11702 22200 11758 23000 6 chany_top_in[17]
port 50 nsew signal input
rlabel metal2 s 12162 22200 12218 23000 6 chany_top_in[18]
port 51 nsew signal input
rlabel metal2 s 12622 22200 12678 23000 6 chany_top_in[19]
port 52 nsew signal input
rlabel metal2 s 4342 22200 4398 23000 6 chany_top_in[1]
port 53 nsew signal input
rlabel metal2 s 4802 22200 4858 23000 6 chany_top_in[2]
port 54 nsew signal input
rlabel metal2 s 5262 22200 5318 23000 6 chany_top_in[3]
port 55 nsew signal input
rlabel metal2 s 5722 22200 5778 23000 6 chany_top_in[4]
port 56 nsew signal input
rlabel metal2 s 6182 22200 6238 23000 6 chany_top_in[5]
port 57 nsew signal input
rlabel metal2 s 6642 22200 6698 23000 6 chany_top_in[6]
port 58 nsew signal input
rlabel metal2 s 7102 22200 7158 23000 6 chany_top_in[7]
port 59 nsew signal input
rlabel metal2 s 7562 22200 7618 23000 6 chany_top_in[8]
port 60 nsew signal input
rlabel metal2 s 8022 22200 8078 23000 6 chany_top_in[9]
port 61 nsew signal input
rlabel metal2 s 13082 22200 13138 23000 6 chany_top_out[0]
port 62 nsew signal tristate
rlabel metal2 s 17682 22200 17738 23000 6 chany_top_out[10]
port 63 nsew signal tristate
rlabel metal2 s 18142 22200 18198 23000 6 chany_top_out[11]
port 64 nsew signal tristate
rlabel metal2 s 18602 22200 18658 23000 6 chany_top_out[12]
port 65 nsew signal tristate
rlabel metal2 s 19062 22200 19118 23000 6 chany_top_out[13]
port 66 nsew signal tristate
rlabel metal2 s 19522 22200 19578 23000 6 chany_top_out[14]
port 67 nsew signal tristate
rlabel metal2 s 19982 22200 20038 23000 6 chany_top_out[15]
port 68 nsew signal tristate
rlabel metal2 s 20442 22200 20498 23000 6 chany_top_out[16]
port 69 nsew signal tristate
rlabel metal2 s 20902 22200 20958 23000 6 chany_top_out[17]
port 70 nsew signal tristate
rlabel metal2 s 21362 22200 21418 23000 6 chany_top_out[18]
port 71 nsew signal tristate
rlabel metal2 s 21822 22200 21878 23000 6 chany_top_out[19]
port 72 nsew signal tristate
rlabel metal2 s 13542 22200 13598 23000 6 chany_top_out[1]
port 73 nsew signal tristate
rlabel metal2 s 14002 22200 14058 23000 6 chany_top_out[2]
port 74 nsew signal tristate
rlabel metal2 s 14462 22200 14518 23000 6 chany_top_out[3]
port 75 nsew signal tristate
rlabel metal2 s 14922 22200 14978 23000 6 chany_top_out[4]
port 76 nsew signal tristate
rlabel metal2 s 15382 22200 15438 23000 6 chany_top_out[5]
port 77 nsew signal tristate
rlabel metal2 s 15842 22200 15898 23000 6 chany_top_out[6]
port 78 nsew signal tristate
rlabel metal2 s 16302 22200 16358 23000 6 chany_top_out[7]
port 79 nsew signal tristate
rlabel metal2 s 16762 22200 16818 23000 6 chany_top_out[8]
port 80 nsew signal tristate
rlabel metal2 s 17222 22200 17278 23000 6 chany_top_out[9]
port 81 nsew signal tristate
rlabel metal3 s 0 2456 800 2576 6 left_bottom_grid_pin_11_
port 82 nsew signal input
rlabel metal3 s 0 2864 800 2984 6 left_bottom_grid_pin_13_
port 83 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 left_bottom_grid_pin_15_
port 84 nsew signal input
rlabel metal3 s 0 3816 800 3936 6 left_bottom_grid_pin_17_
port 85 nsew signal input
rlabel metal3 s 0 144 800 264 6 left_bottom_grid_pin_1_
port 86 nsew signal input
rlabel metal3 s 0 552 800 672 6 left_bottom_grid_pin_3_
port 87 nsew signal input
rlabel metal3 s 0 960 800 1080 6 left_bottom_grid_pin_5_
port 88 nsew signal input
rlabel metal3 s 0 1504 800 1624 6 left_bottom_grid_pin_7_
port 89 nsew signal input
rlabel metal3 s 0 1912 800 2032 6 left_bottom_grid_pin_9_
port 90 nsew signal input
rlabel metal2 s 22282 22200 22338 23000 6 prog_clk_0_N_in
port 91 nsew signal input
rlabel metal2 s 202 22200 258 23000 6 top_left_grid_pin_42_
port 92 nsew signal input
rlabel metal2 s 662 22200 718 23000 6 top_left_grid_pin_43_
port 93 nsew signal input
rlabel metal2 s 1122 22200 1178 23000 6 top_left_grid_pin_44_
port 94 nsew signal input
rlabel metal2 s 1582 22200 1638 23000 6 top_left_grid_pin_45_
port 95 nsew signal input
rlabel metal2 s 2042 22200 2098 23000 6 top_left_grid_pin_46_
port 96 nsew signal input
rlabel metal2 s 2502 22200 2558 23000 6 top_left_grid_pin_47_
port 97 nsew signal input
rlabel metal2 s 2962 22200 3018 23000 6 top_left_grid_pin_48_
port 98 nsew signal input
rlabel metal2 s 3422 22200 3478 23000 6 top_left_grid_pin_49_
port 99 nsew signal input
rlabel metal2 s 22742 22200 22798 23000 6 top_right_grid_pin_1_
port 100 nsew signal input
rlabel metal4 s 18271 2128 18591 20720 6 VPWR
port 101 nsew power bidirectional
rlabel metal4 s 11340 2128 11660 20720 6 VPWR
port 102 nsew power bidirectional
rlabel metal4 s 4409 2128 4729 20720 6 VPWR
port 103 nsew power bidirectional
rlabel metal4 s 14805 2128 15125 20720 6 VGND
port 104 nsew ground bidirectional
rlabel metal4 s 7875 2128 8195 20720 6 VGND
port 105 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
